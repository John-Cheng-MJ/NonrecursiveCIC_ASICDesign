module add_signed_116_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [27:0] A, B;
  output [28:0] Z;
  wire [27:0] A, B;
  wire [28:0] Z;
  wire n_89, n_90, n_93, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_103, n_104, n_105, n_106, n_107, n_109, n_110;
  wire n_111, n_112, n_113, n_115, n_116, n_117, n_118, n_119;
  wire n_121, n_122, n_123, n_124, n_125, n_127, n_128, n_129;
  wire n_130, n_131, n_133, n_134, n_135, n_136, n_137, n_139;
  wire n_140, n_141, n_142, n_143, n_145, n_146, n_147, n_148;
  wire n_149, n_151, n_152, n_153, n_154, n_155, n_157, n_158;
  wire n_159, n_160, n_161, n_163, n_164, n_165, n_166, n_167;
  wire n_169, n_170, n_171, n_172, n_173, n_175, n_176, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_185, n_187, n_189;
  wire n_190, n_192, n_193, n_195, n_197, n_199, n_200, n_202;
  wire n_203, n_205, n_207, n_209, n_210, n_212, n_213, n_215;
  wire n_217, n_219, n_220, n_222, n_223, n_225, n_227, n_229;
  wire n_230, n_232, n_233, n_235, n_237, n_239, n_240, n_242;
  wire n_244, n_245, n_246, n_248, n_249, n_250, n_252, n_253;
  wire n_254, n_255, n_257, n_259, n_261, n_262, n_263, n_265;
  wire n_266, n_267, n_269, n_270, n_272, n_274, n_276, n_277;
  wire n_278, n_280, n_281, n_282, n_284, n_286, n_287, n_288;
  wire n_290, n_291, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_309, n_312, n_314, n_315, n_316, n_319, n_320;
  wire n_321, n_324, n_326, n_327, n_328, n_330, n_331, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_346, n_347, n_348, n_350, n_351;
  wire n_352, n_354, n_355, n_356, n_358, n_359, n_360, n_361;
  wire n_363, n_364, n_365, n_367, n_368, n_369, n_370, n_372;
  wire n_373, n_374, n_376, n_377, n_378, n_379, n_381, n_382;
  wire n_384, n_385, n_387, n_388, n_389, n_390, n_392, n_393;
  wire n_394, n_396, n_397, n_398, n_399, n_401, n_402, n_404;
  wire n_405, n_407, n_408, n_409, n_410, n_412, n_413, n_414;
  wire n_415, n_417, n_418, n_419, n_420, n_422, n_423;
  not g3 (Z[28], n_89);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_90, A[0], B[0]);
  nor g9 (n_93, A[1], B[1]);
  nand g10 (n_96, A[1], B[1]);
  nor g11 (n_103, A[2], B[2]);
  nand g12 (n_98, A[2], B[2]);
  nor g13 (n_99, A[3], B[3]);
  nand g14 (n_100, A[3], B[3]);
  nor g15 (n_109, A[4], B[4]);
  nand g16 (n_104, A[4], B[4]);
  nor g17 (n_105, A[5], B[5]);
  nand g18 (n_106, A[5], B[5]);
  nor g19 (n_115, A[6], B[6]);
  nand g20 (n_110, A[6], B[6]);
  nor g21 (n_111, A[7], B[7]);
  nand g22 (n_112, A[7], B[7]);
  nor g23 (n_121, A[8], B[8]);
  nand g24 (n_116, A[8], B[8]);
  nor g25 (n_117, A[9], B[9]);
  nand g26 (n_118, A[9], B[9]);
  nor g27 (n_127, A[10], B[10]);
  nand g28 (n_122, A[10], B[10]);
  nor g29 (n_123, A[11], B[11]);
  nand g30 (n_124, A[11], B[11]);
  nor g31 (n_133, A[12], B[12]);
  nand g32 (n_128, A[12], B[12]);
  nor g33 (n_129, A[13], B[13]);
  nand g34 (n_130, A[13], B[13]);
  nor g35 (n_139, A[14], B[14]);
  nand g36 (n_134, A[14], B[14]);
  nor g37 (n_135, A[15], B[15]);
  nand g38 (n_136, A[15], B[15]);
  nor g39 (n_145, A[16], B[16]);
  nand g40 (n_140, A[16], B[16]);
  nor g41 (n_141, A[17], B[17]);
  nand g42 (n_142, A[17], B[17]);
  nor g43 (n_151, A[18], B[18]);
  nand g44 (n_146, A[18], B[18]);
  nor g45 (n_147, A[19], B[19]);
  nand g46 (n_148, A[19], B[19]);
  nor g47 (n_157, A[20], B[20]);
  nand g48 (n_152, A[20], B[20]);
  nor g49 (n_153, A[21], B[21]);
  nand g50 (n_154, A[21], B[21]);
  nor g51 (n_163, A[22], B[22]);
  nand g52 (n_158, A[22], B[22]);
  nor g53 (n_159, A[23], B[23]);
  nand g54 (n_160, A[23], B[23]);
  nor g55 (n_169, A[24], B[24]);
  nand g56 (n_164, A[24], B[24]);
  nor g57 (n_165, A[25], B[25]);
  nand g58 (n_166, A[25], B[25]);
  nor g59 (n_175, A[26], B[26]);
  nand g60 (n_170, A[26], B[26]);
  nand g65 (n_176, n_96, n_97);
  nor g66 (n_101, n_98, n_99);
  nor g69 (n_179, n_103, n_99);
  nor g70 (n_107, n_104, n_105);
  nor g73 (n_185, n_109, n_105);
  nor g74 (n_113, n_110, n_111);
  nor g77 (n_187, n_115, n_111);
  nor g78 (n_119, n_116, n_117);
  nor g81 (n_195, n_121, n_117);
  nor g82 (n_125, n_122, n_123);
  nor g85 (n_197, n_127, n_123);
  nor g86 (n_131, n_128, n_129);
  nor g89 (n_205, n_133, n_129);
  nor g90 (n_137, n_134, n_135);
  nor g93 (n_207, n_139, n_135);
  nor g94 (n_143, n_140, n_141);
  nor g97 (n_215, n_145, n_141);
  nor g98 (n_149, n_146, n_147);
  nor g101 (n_217, n_151, n_147);
  nor g102 (n_155, n_152, n_153);
  nor g105 (n_225, n_157, n_153);
  nor g106 (n_161, n_158, n_159);
  nor g109 (n_227, n_163, n_159);
  nor g110 (n_167, n_164, n_165);
  nor g113 (n_235, n_169, n_165);
  nor g114 (n_173, n_170, n_171);
  nor g117 (n_237, n_175, n_171);
  nand g120 (n_363, n_98, n_178);
  nand g121 (n_181, n_179, n_176);
  nand g122 (n_242, n_180, n_181);
  nor g123 (n_183, n_115, n_182);
  nand g132 (n_250, n_185, n_187);
  nor g133 (n_193, n_127, n_192);
  nand g142 (n_257, n_195, n_197);
  nor g143 (n_203, n_139, n_202);
  nand g152 (n_265, n_205, n_207);
  nor g153 (n_213, n_151, n_212);
  nand g162 (n_272, n_215, n_217);
  nor g163 (n_223, n_163, n_222);
  nand g172 (n_280, n_225, n_227);
  nor g173 (n_233, n_175, n_232);
  nand g182 (n_319, n_235, n_237);
  nand g185 (n_367, n_104, n_244);
  nand g186 (n_245, n_185, n_242);
  nand g187 (n_369, n_182, n_245);
  nand g190 (n_372, n_248, n_249);
  nand g193 (n_284, n_252, n_253);
  nor g194 (n_255, n_133, n_254);
  nor g197 (n_294, n_133, n_257);
  nor g203 (n_263, n_261, n_254);
  nor g206 (n_300, n_257, n_261);
  nor g207 (n_267, n_265, n_254);
  nor g210 (n_303, n_257, n_265);
  nor g211 (n_270, n_157, n_269);
  nor g214 (n_334, n_157, n_272);
  nor g220 (n_278, n_276, n_269);
  nor g223 (n_340, n_272, n_276);
  nor g224 (n_282, n_280, n_269);
  nor g227 (n_309, n_272, n_280);
  nand g230 (n_376, n_116, n_286);
  nand g231 (n_287, n_195, n_284);
  nand g232 (n_378, n_192, n_287);
  nand g235 (n_381, n_290, n_291);
  nand g238 (n_384, n_254, n_293);
  nand g239 (n_296, n_294, n_284);
  nand g240 (n_387, n_295, n_296);
  nand g241 (n_299, n_297, n_284);
  nand g242 (n_389, n_298, n_299);
  nand g243 (n_302, n_300, n_284);
  nand g244 (n_392, n_301, n_302);
  nand g245 (n_305, n_303, n_284);
  nand g246 (n_324, n_304, n_305);
  nor g247 (n_307, n_169, n_306);
  nand g256 (n_348, n_235, n_309);
  nor g257 (n_316, n_314, n_306);
  nor g262 (n_321, n_319, n_306);
  nand g269 (n_396, n_140, n_326);
  nand g270 (n_327, n_215, n_324);
  nand g271 (n_398, n_212, n_327);
  nand g274 (n_401, n_330, n_331);
  nand g277 (n_404, n_269, n_333);
  nand g278 (n_336, n_334, n_324);
  nand g279 (n_407, n_335, n_336);
  nand g280 (n_339, n_337, n_324);
  nand g281 (n_409, n_338, n_339);
  nand g282 (n_342, n_340, n_324);
  nand g283 (n_412, n_341, n_342);
  nand g284 (n_343, n_309, n_324);
  nand g285 (n_414, n_306, n_343);
  nand g288 (n_417, n_346, n_347);
  nand g291 (n_419, n_350, n_351);
  nand g294 (n_422, n_354, n_355);
  nand g297 (n_89, n_358, n_359);
  xnor g301 (Z[2], n_176, n_361);
  xnor g304 (Z[3], n_363, n_364);
  xnor g306 (Z[4], n_242, n_365);
  xnor g309 (Z[5], n_367, n_368);
  xnor g311 (Z[6], n_369, n_370);
  xnor g314 (Z[7], n_372, n_373);
  xnor g316 (Z[8], n_284, n_374);
  xnor g319 (Z[9], n_376, n_377);
  xnor g321 (Z[10], n_378, n_379);
  xnor g324 (Z[11], n_381, n_382);
  xnor g327 (Z[12], n_384, n_385);
  xnor g330 (Z[13], n_387, n_388);
  xnor g332 (Z[14], n_389, n_390);
  xnor g335 (Z[15], n_392, n_393);
  xnor g337 (Z[16], n_324, n_394);
  xnor g340 (Z[17], n_396, n_397);
  xnor g342 (Z[18], n_398, n_399);
  xnor g345 (Z[19], n_401, n_402);
  xnor g348 (Z[20], n_404, n_405);
  xnor g351 (Z[21], n_407, n_408);
  xnor g353 (Z[22], n_409, n_410);
  xnor g356 (Z[23], n_412, n_413);
  xnor g358 (Z[24], n_414, n_415);
  xnor g361 (Z[25], n_417, n_418);
  xnor g363 (Z[26], n_419, n_420);
  xnor g366 (Z[27], n_422, n_423);
  and g369 (n_171, A[27], B[27]);
  or g370 (n_172, A[27], B[27]);
  and g371 (n_212, wc, n_142);
  not gc (wc, n_143);
  and g372 (n_219, wc0, n_148);
  not gc0 (wc0, n_149);
  and g373 (n_222, wc1, n_154);
  not gc1 (wc1, n_155);
  and g374 (n_229, wc2, n_160);
  not gc2 (wc2, n_161);
  and g375 (n_232, wc3, n_166);
  not gc3 (wc3, n_167);
  and g376 (n_192, wc4, n_118);
  not gc4 (wc4, n_119);
  and g377 (n_199, wc5, n_124);
  not gc5 (wc5, n_125);
  and g378 (n_202, wc6, n_130);
  not gc6 (wc6, n_131);
  and g379 (n_209, wc7, n_136);
  not gc7 (wc7, n_137);
  and g380 (n_182, wc8, n_106);
  not gc8 (wc8, n_107);
  and g381 (n_189, wc9, n_112);
  not gc9 (wc9, n_113);
  and g382 (n_180, wc10, n_100);
  not gc10 (wc10, n_101);
  or g383 (n_97, n_90, n_93);
  or g384 (n_246, wc11, n_115);
  not gc11 (wc11, n_185);
  or g385 (n_288, wc12, n_127);
  not gc12 (wc12, n_195);
  or g386 (n_261, wc13, n_139);
  not gc13 (wc13, n_205);
  or g387 (n_328, wc14, n_151);
  not gc14 (wc14, n_215);
  or g388 (n_276, wc15, n_163);
  not gc15 (wc15, n_225);
  or g389 (n_314, wc16, n_175);
  not gc16 (wc16, n_235);
  or g390 (n_360, wc17, n_93);
  not gc17 (wc17, n_96);
  or g391 (n_361, wc18, n_103);
  not gc18 (wc18, n_98);
  or g392 (n_364, wc19, n_99);
  not gc19 (wc19, n_100);
  or g393 (n_365, wc20, n_109);
  not gc20 (wc20, n_104);
  or g394 (n_368, wc21, n_105);
  not gc21 (wc21, n_106);
  or g395 (n_370, wc22, n_115);
  not gc22 (wc22, n_110);
  or g396 (n_373, wc23, n_111);
  not gc23 (wc23, n_112);
  or g397 (n_374, wc24, n_121);
  not gc24 (wc24, n_116);
  or g398 (n_377, wc25, n_117);
  not gc25 (wc25, n_118);
  or g399 (n_379, wc26, n_127);
  not gc26 (wc26, n_122);
  or g400 (n_382, wc27, n_123);
  not gc27 (wc27, n_124);
  or g401 (n_385, wc28, n_133);
  not gc28 (wc28, n_128);
  or g402 (n_388, wc29, n_129);
  not gc29 (wc29, n_130);
  or g403 (n_390, wc30, n_139);
  not gc30 (wc30, n_134);
  or g404 (n_393, wc31, n_135);
  not gc31 (wc31, n_136);
  or g405 (n_394, wc32, n_145);
  not gc32 (wc32, n_140);
  or g406 (n_397, wc33, n_141);
  not gc33 (wc33, n_142);
  or g407 (n_399, wc34, n_151);
  not gc34 (wc34, n_146);
  or g408 (n_402, wc35, n_147);
  not gc35 (wc35, n_148);
  or g409 (n_405, wc36, n_157);
  not gc36 (wc36, n_152);
  or g410 (n_408, wc37, n_153);
  not gc37 (wc37, n_154);
  or g411 (n_410, wc38, n_163);
  not gc38 (wc38, n_158);
  or g412 (n_413, wc39, n_159);
  not gc39 (wc39, n_160);
  or g413 (n_415, wc40, n_169);
  not gc40 (wc40, n_164);
  or g414 (n_418, wc41, n_165);
  not gc41 (wc41, n_166);
  or g415 (n_420, wc42, n_175);
  not gc42 (wc42, n_170);
  and g416 (n_220, wc43, n_217);
  not gc43 (wc43, n_212);
  and g417 (n_230, wc44, n_227);
  not gc44 (wc44, n_222);
  and g418 (n_239, n_172, wc45);
  not gc45 (wc45, n_173);
  and g419 (n_200, wc46, n_197);
  not gc46 (wc46, n_192);
  and g420 (n_210, wc47, n_207);
  not gc47 (wc47, n_202);
  and g421 (n_190, wc48, n_187);
  not gc48 (wc48, n_182);
  and g422 (n_297, wc49, n_205);
  not gc49 (wc49, n_257);
  and g423 (n_337, wc50, n_225);
  not gc50 (wc50, n_272);
  xor g424 (Z[1], n_90, n_360);
  or g425 (n_423, wc51, n_171);
  not gc51 (wc51, n_172);
  and g426 (n_269, wc52, n_219);
  not gc52 (wc52, n_220);
  and g427 (n_281, wc53, n_229);
  not gc53 (wc53, n_230);
  and g428 (n_240, wc54, n_237);
  not gc54 (wc54, n_232);
  and g429 (n_254, wc55, n_199);
  not gc55 (wc55, n_200);
  and g430 (n_266, wc56, n_209);
  not gc56 (wc56, n_210);
  and g431 (n_252, wc57, n_189);
  not gc57 (wc57, n_190);
  or g432 (n_178, wc58, n_103);
  not gc58 (wc58, n_176);
  and g433 (n_248, wc59, n_110);
  not gc59 (wc59, n_183);
  and g434 (n_290, wc60, n_122);
  not gc60 (wc60, n_193);
  and g435 (n_262, wc61, n_134);
  not gc61 (wc61, n_203);
  and g436 (n_330, wc62, n_146);
  not gc62 (wc62, n_213);
  and g437 (n_277, wc63, n_158);
  not gc63 (wc63, n_223);
  and g438 (n_315, wc64, n_170);
  not gc64 (wc64, n_233);
  or g439 (n_344, wc65, n_169);
  not gc65 (wc65, n_309);
  or g440 (n_352, n_314, wc66);
  not gc66 (wc66, n_309);
  and g441 (n_320, wc67, n_239);
  not gc67 (wc67, n_240);
  or g442 (n_356, wc68, n_319);
  not gc68 (wc68, n_309);
  and g443 (n_259, wc69, n_205);
  not gc69 (wc69, n_254);
  and g444 (n_274, wc70, n_225);
  not gc70 (wc70, n_269);
  and g445 (n_306, n_281, wc71);
  not gc71 (wc71, n_282);
  and g446 (n_304, n_266, wc72);
  not gc72 (wc72, n_267);
  or g447 (n_253, n_250, wc73);
  not gc73 (wc73, n_242);
  or g448 (n_244, wc74, n_109);
  not gc74 (wc74, n_242);
  or g449 (n_249, n_246, wc75);
  not gc75 (wc75, n_242);
  and g450 (n_295, wc76, n_128);
  not gc76 (wc76, n_255);
  and g451 (n_298, wc77, n_202);
  not gc77 (wc77, n_259);
  and g452 (n_301, n_262, wc78);
  not gc78 (wc78, n_263);
  and g453 (n_335, wc79, n_152);
  not gc79 (wc79, n_270);
  and g454 (n_338, wc80, n_222);
  not gc80 (wc80, n_274);
  and g455 (n_341, n_277, wc81);
  not gc81 (wc81, n_278);
  and g456 (n_312, wc82, n_235);
  not gc82 (wc82, n_306);
  and g457 (n_358, n_320, wc83);
  not gc83 (wc83, n_321);
  or g458 (n_286, wc84, n_121);
  not gc84 (wc84, n_284);
  or g459 (n_291, n_288, wc85);
  not gc85 (wc85, n_284);
  or g460 (n_293, wc86, n_257);
  not gc86 (wc86, n_284);
  and g461 (n_346, wc87, n_164);
  not gc87 (wc87, n_307);
  and g462 (n_350, wc88, n_232);
  not gc88 (wc88, n_312);
  and g463 (n_354, n_315, wc89);
  not gc89 (wc89, n_316);
  or g464 (n_359, n_356, wc90);
  not gc90 (wc90, n_324);
  or g465 (n_326, wc91, n_145);
  not gc91 (wc91, n_324);
  or g466 (n_331, n_328, wc92);
  not gc92 (wc92, n_324);
  or g467 (n_333, wc93, n_272);
  not gc93 (wc93, n_324);
  or g468 (n_347, n_344, wc94);
  not gc94 (wc94, n_324);
  or g469 (n_351, n_348, wc95);
  not gc95 (wc95, n_324);
  or g470 (n_355, n_352, wc96);
  not gc96 (wc96, n_324);
endmodule

module add_signed_116_GENERIC(A, B, Z);
  input [27:0] A, B;
  output [28:0] Z;
  wire [27:0] A, B;
  wire [28:0] Z;
  add_signed_116_GENERIC_REAL g1(.A ({A[26], A[26:0]}), .B ({B[26],
       B[26:0]}), .Z (Z));
endmodule

module add_signed_1220_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [66:0] A, B;
  output [67:0] Z;
  wire [66:0] A, B;
  wire [67:0] Z;
  wire n_206, n_207, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540;
  not g3 (Z[67], n_206);
  nand g4 (n_207, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_212, A[1], B[1]);
  nand g13 (n_216, n_212, n_213, n_214);
  xor g14 (n_215, A[1], B[1]);
  nand g16 (n_217, A[2], B[2]);
  nand g17 (n_218, A[2], n_216);
  nand g18 (n_219, B[2], n_216);
  nand g19 (n_221, n_217, n_218, n_219);
  xor g20 (n_220, A[2], B[2]);
  xor g21 (Z[2], n_216, n_220);
  nand g22 (n_222, A[3], B[3]);
  nand g23 (n_223, A[3], n_221);
  nand g24 (n_224, B[3], n_221);
  nand g25 (n_226, n_222, n_223, n_224);
  xor g26 (n_225, A[3], B[3]);
  xor g27 (Z[3], n_221, n_225);
  nand g28 (n_227, A[4], B[4]);
  nand g29 (n_228, A[4], n_226);
  nand g30 (n_229, B[4], n_226);
  nand g31 (n_231, n_227, n_228, n_229);
  xor g32 (n_230, A[4], B[4]);
  xor g33 (Z[4], n_226, n_230);
  nand g34 (n_232, A[5], B[5]);
  nand g35 (n_233, A[5], n_231);
  nand g36 (n_234, B[5], n_231);
  nand g37 (n_236, n_232, n_233, n_234);
  xor g38 (n_235, A[5], B[5]);
  xor g39 (Z[5], n_231, n_235);
  nand g40 (n_237, A[6], B[6]);
  nand g41 (n_238, A[6], n_236);
  nand g42 (n_239, B[6], n_236);
  nand g43 (n_241, n_237, n_238, n_239);
  xor g44 (n_240, A[6], B[6]);
  xor g45 (Z[6], n_236, n_240);
  nand g46 (n_242, A[7], B[7]);
  nand g47 (n_243, A[7], n_241);
  nand g48 (n_244, B[7], n_241);
  nand g49 (n_246, n_242, n_243, n_244);
  xor g50 (n_245, A[7], B[7]);
  xor g51 (Z[7], n_241, n_245);
  nand g52 (n_247, A[8], B[8]);
  nand g53 (n_248, A[8], n_246);
  nand g54 (n_249, B[8], n_246);
  nand g55 (n_251, n_247, n_248, n_249);
  xor g56 (n_250, A[8], B[8]);
  xor g57 (Z[8], n_246, n_250);
  nand g58 (n_252, A[9], B[9]);
  nand g59 (n_253, A[9], n_251);
  nand g60 (n_254, B[9], n_251);
  nand g61 (n_256, n_252, n_253, n_254);
  xor g62 (n_255, A[9], B[9]);
  xor g63 (Z[9], n_251, n_255);
  nand g64 (n_257, A[10], B[10]);
  nand g65 (n_258, A[10], n_256);
  nand g66 (n_259, B[10], n_256);
  nand g67 (n_261, n_257, n_258, n_259);
  xor g68 (n_260, A[10], B[10]);
  xor g69 (Z[10], n_256, n_260);
  nand g70 (n_262, A[11], B[11]);
  nand g71 (n_263, A[11], n_261);
  nand g72 (n_264, B[11], n_261);
  nand g73 (n_266, n_262, n_263, n_264);
  xor g74 (n_265, A[11], B[11]);
  xor g75 (Z[11], n_261, n_265);
  nand g76 (n_267, A[12], B[12]);
  nand g77 (n_268, A[12], n_266);
  nand g78 (n_269, B[12], n_266);
  nand g79 (n_271, n_267, n_268, n_269);
  xor g80 (n_270, A[12], B[12]);
  xor g81 (Z[12], n_266, n_270);
  nand g82 (n_272, A[13], B[13]);
  nand g83 (n_273, A[13], n_271);
  nand g84 (n_274, B[13], n_271);
  nand g85 (n_276, n_272, n_273, n_274);
  xor g86 (n_275, A[13], B[13]);
  xor g87 (Z[13], n_271, n_275);
  nand g88 (n_277, A[14], B[14]);
  nand g89 (n_278, A[14], n_276);
  nand g90 (n_279, B[14], n_276);
  nand g91 (n_281, n_277, n_278, n_279);
  xor g92 (n_280, A[14], B[14]);
  xor g93 (Z[14], n_276, n_280);
  nand g94 (n_282, A[15], B[15]);
  nand g95 (n_283, A[15], n_281);
  nand g96 (n_284, B[15], n_281);
  nand g97 (n_286, n_282, n_283, n_284);
  xor g98 (n_285, A[15], B[15]);
  xor g99 (Z[15], n_281, n_285);
  nand g100 (n_287, A[16], B[16]);
  nand g101 (n_288, A[16], n_286);
  nand g102 (n_289, B[16], n_286);
  nand g103 (n_291, n_287, n_288, n_289);
  xor g104 (n_290, A[16], B[16]);
  xor g105 (Z[16], n_286, n_290);
  nand g106 (n_292, A[17], B[17]);
  nand g107 (n_293, A[17], n_291);
  nand g108 (n_294, B[17], n_291);
  nand g109 (n_296, n_292, n_293, n_294);
  xor g110 (n_295, A[17], B[17]);
  xor g111 (Z[17], n_291, n_295);
  nand g112 (n_297, A[18], B[18]);
  nand g113 (n_298, A[18], n_296);
  nand g114 (n_299, B[18], n_296);
  nand g115 (n_301, n_297, n_298, n_299);
  xor g116 (n_300, A[18], B[18]);
  xor g117 (Z[18], n_296, n_300);
  nand g118 (n_302, A[19], B[19]);
  nand g119 (n_303, A[19], n_301);
  nand g120 (n_304, B[19], n_301);
  nand g121 (n_306, n_302, n_303, n_304);
  xor g122 (n_305, A[19], B[19]);
  xor g123 (Z[19], n_301, n_305);
  nand g124 (n_307, A[20], B[20]);
  nand g125 (n_308, A[20], n_306);
  nand g126 (n_309, B[20], n_306);
  nand g127 (n_311, n_307, n_308, n_309);
  xor g128 (n_310, A[20], B[20]);
  xor g129 (Z[20], n_306, n_310);
  nand g130 (n_312, A[21], B[21]);
  nand g131 (n_313, A[21], n_311);
  nand g132 (n_314, B[21], n_311);
  nand g133 (n_316, n_312, n_313, n_314);
  xor g134 (n_315, A[21], B[21]);
  xor g135 (Z[21], n_311, n_315);
  nand g136 (n_317, A[22], B[22]);
  nand g137 (n_318, A[22], n_316);
  nand g138 (n_319, B[22], n_316);
  nand g139 (n_321, n_317, n_318, n_319);
  xor g140 (n_320, A[22], B[22]);
  xor g141 (Z[22], n_316, n_320);
  nand g142 (n_322, A[23], B[23]);
  nand g143 (n_323, A[23], n_321);
  nand g144 (n_324, B[23], n_321);
  nand g145 (n_326, n_322, n_323, n_324);
  xor g146 (n_325, A[23], B[23]);
  xor g147 (Z[23], n_321, n_325);
  nand g148 (n_327, A[24], B[24]);
  nand g149 (n_328, A[24], n_326);
  nand g150 (n_329, B[24], n_326);
  nand g151 (n_331, n_327, n_328, n_329);
  xor g152 (n_330, A[24], B[24]);
  xor g153 (Z[24], n_326, n_330);
  nand g154 (n_332, A[25], B[25]);
  nand g155 (n_333, A[25], n_331);
  nand g156 (n_334, B[25], n_331);
  nand g157 (n_336, n_332, n_333, n_334);
  xor g158 (n_335, A[25], B[25]);
  xor g159 (Z[25], n_331, n_335);
  nand g160 (n_337, A[26], B[26]);
  nand g161 (n_338, A[26], n_336);
  nand g162 (n_339, B[26], n_336);
  nand g163 (n_341, n_337, n_338, n_339);
  xor g164 (n_340, A[26], B[26]);
  xor g165 (Z[26], n_336, n_340);
  nand g166 (n_342, A[27], B[27]);
  nand g167 (n_343, A[27], n_341);
  nand g168 (n_344, B[27], n_341);
  nand g169 (n_346, n_342, n_343, n_344);
  xor g170 (n_345, A[27], B[27]);
  xor g171 (Z[27], n_341, n_345);
  nand g172 (n_347, A[28], B[28]);
  nand g173 (n_348, A[28], n_346);
  nand g174 (n_349, B[28], n_346);
  nand g175 (n_351, n_347, n_348, n_349);
  xor g176 (n_350, A[28], B[28]);
  xor g177 (Z[28], n_346, n_350);
  nand g178 (n_352, A[29], B[29]);
  nand g179 (n_353, A[29], n_351);
  nand g180 (n_354, B[29], n_351);
  nand g181 (n_356, n_352, n_353, n_354);
  xor g182 (n_355, A[29], B[29]);
  xor g183 (Z[29], n_351, n_355);
  nand g184 (n_357, A[30], B[30]);
  nand g185 (n_358, A[30], n_356);
  nand g186 (n_359, B[30], n_356);
  nand g187 (n_361, n_357, n_358, n_359);
  xor g188 (n_360, A[30], B[30]);
  xor g189 (Z[30], n_356, n_360);
  nand g190 (n_362, A[31], B[31]);
  nand g191 (n_363, A[31], n_361);
  nand g192 (n_364, B[31], n_361);
  nand g193 (n_366, n_362, n_363, n_364);
  xor g194 (n_365, A[31], B[31]);
  xor g195 (Z[31], n_361, n_365);
  nand g196 (n_367, A[32], B[32]);
  nand g197 (n_368, A[32], n_366);
  nand g198 (n_369, B[32], n_366);
  nand g199 (n_371, n_367, n_368, n_369);
  xor g200 (n_370, A[32], B[32]);
  xor g201 (Z[32], n_366, n_370);
  nand g202 (n_372, A[33], B[33]);
  nand g203 (n_373, A[33], n_371);
  nand g204 (n_374, B[33], n_371);
  nand g205 (n_376, n_372, n_373, n_374);
  xor g206 (n_375, A[33], B[33]);
  xor g207 (Z[33], n_371, n_375);
  nand g208 (n_377, A[34], B[34]);
  nand g209 (n_378, A[34], n_376);
  nand g210 (n_379, B[34], n_376);
  nand g211 (n_381, n_377, n_378, n_379);
  xor g212 (n_380, A[34], B[34]);
  xor g213 (Z[34], n_376, n_380);
  nand g214 (n_382, A[35], B[35]);
  nand g215 (n_383, A[35], n_381);
  nand g216 (n_384, B[35], n_381);
  nand g217 (n_386, n_382, n_383, n_384);
  xor g218 (n_385, A[35], B[35]);
  xor g219 (Z[35], n_381, n_385);
  nand g220 (n_387, A[36], B[36]);
  nand g221 (n_388, A[36], n_386);
  nand g222 (n_389, B[36], n_386);
  nand g223 (n_391, n_387, n_388, n_389);
  xor g224 (n_390, A[36], B[36]);
  xor g225 (Z[36], n_386, n_390);
  nand g226 (n_392, A[37], B[37]);
  nand g227 (n_393, A[37], n_391);
  nand g228 (n_394, B[37], n_391);
  nand g229 (n_396, n_392, n_393, n_394);
  xor g230 (n_395, A[37], B[37]);
  xor g231 (Z[37], n_391, n_395);
  nand g232 (n_397, A[38], B[38]);
  nand g233 (n_398, A[38], n_396);
  nand g234 (n_399, B[38], n_396);
  nand g235 (n_401, n_397, n_398, n_399);
  xor g236 (n_400, A[38], B[38]);
  xor g237 (Z[38], n_396, n_400);
  nand g238 (n_402, A[39], B[39]);
  nand g239 (n_403, A[39], n_401);
  nand g240 (n_404, B[39], n_401);
  nand g241 (n_406, n_402, n_403, n_404);
  xor g242 (n_405, A[39], B[39]);
  xor g243 (Z[39], n_401, n_405);
  nand g244 (n_407, A[40], B[40]);
  nand g245 (n_408, A[40], n_406);
  nand g246 (n_409, B[40], n_406);
  nand g247 (n_411, n_407, n_408, n_409);
  xor g248 (n_410, A[40], B[40]);
  xor g249 (Z[40], n_406, n_410);
  nand g250 (n_412, A[41], B[41]);
  nand g251 (n_413, A[41], n_411);
  nand g252 (n_414, B[41], n_411);
  nand g253 (n_416, n_412, n_413, n_414);
  xor g254 (n_415, A[41], B[41]);
  xor g255 (Z[41], n_411, n_415);
  nand g256 (n_417, A[42], B[42]);
  nand g257 (n_418, A[42], n_416);
  nand g258 (n_419, B[42], n_416);
  nand g259 (n_421, n_417, n_418, n_419);
  xor g260 (n_420, A[42], B[42]);
  xor g261 (Z[42], n_416, n_420);
  nand g262 (n_422, A[43], B[43]);
  nand g263 (n_423, A[43], n_421);
  nand g264 (n_424, B[43], n_421);
  nand g265 (n_426, n_422, n_423, n_424);
  xor g266 (n_425, A[43], B[43]);
  xor g267 (Z[43], n_421, n_425);
  nand g268 (n_427, A[44], B[44]);
  nand g269 (n_428, A[44], n_426);
  nand g270 (n_429, B[44], n_426);
  nand g271 (n_431, n_427, n_428, n_429);
  xor g272 (n_430, A[44], B[44]);
  xor g273 (Z[44], n_426, n_430);
  nand g274 (n_432, A[45], B[45]);
  nand g275 (n_433, A[45], n_431);
  nand g276 (n_434, B[45], n_431);
  nand g277 (n_436, n_432, n_433, n_434);
  xor g278 (n_435, A[45], B[45]);
  xor g279 (Z[45], n_431, n_435);
  nand g280 (n_437, A[46], B[46]);
  nand g281 (n_438, A[46], n_436);
  nand g282 (n_439, B[46], n_436);
  nand g283 (n_441, n_437, n_438, n_439);
  xor g284 (n_440, A[46], B[46]);
  xor g285 (Z[46], n_436, n_440);
  nand g286 (n_442, A[47], B[47]);
  nand g287 (n_443, A[47], n_441);
  nand g288 (n_444, B[47], n_441);
  nand g289 (n_446, n_442, n_443, n_444);
  xor g290 (n_445, A[47], B[47]);
  xor g291 (Z[47], n_441, n_445);
  nand g292 (n_447, A[48], B[48]);
  nand g293 (n_448, A[48], n_446);
  nand g294 (n_449, B[48], n_446);
  nand g295 (n_451, n_447, n_448, n_449);
  xor g296 (n_450, A[48], B[48]);
  xor g297 (Z[48], n_446, n_450);
  nand g298 (n_452, A[49], B[49]);
  nand g299 (n_453, A[49], n_451);
  nand g300 (n_454, B[49], n_451);
  nand g301 (n_456, n_452, n_453, n_454);
  xor g302 (n_455, A[49], B[49]);
  xor g303 (Z[49], n_451, n_455);
  nand g304 (n_457, A[50], B[50]);
  nand g305 (n_458, A[50], n_456);
  nand g306 (n_459, B[50], n_456);
  nand g307 (n_461, n_457, n_458, n_459);
  xor g308 (n_460, A[50], B[50]);
  xor g309 (Z[50], n_456, n_460);
  nand g310 (n_462, A[51], B[51]);
  nand g311 (n_463, A[51], n_461);
  nand g312 (n_464, B[51], n_461);
  nand g313 (n_466, n_462, n_463, n_464);
  xor g314 (n_465, A[51], B[51]);
  xor g315 (Z[51], n_461, n_465);
  nand g316 (n_467, A[52], B[52]);
  nand g317 (n_468, A[52], n_466);
  nand g318 (n_469, B[52], n_466);
  nand g319 (n_471, n_467, n_468, n_469);
  xor g320 (n_470, A[52], B[52]);
  xor g321 (Z[52], n_466, n_470);
  nand g322 (n_472, A[53], B[53]);
  nand g323 (n_473, A[53], n_471);
  nand g324 (n_474, B[53], n_471);
  nand g325 (n_476, n_472, n_473, n_474);
  xor g326 (n_475, A[53], B[53]);
  xor g327 (Z[53], n_471, n_475);
  nand g328 (n_477, A[54], B[54]);
  nand g329 (n_478, A[54], n_476);
  nand g330 (n_479, B[54], n_476);
  nand g331 (n_481, n_477, n_478, n_479);
  xor g332 (n_480, A[54], B[54]);
  xor g333 (Z[54], n_476, n_480);
  nand g334 (n_482, A[55], B[55]);
  nand g335 (n_483, A[55], n_481);
  nand g336 (n_484, B[55], n_481);
  nand g337 (n_486, n_482, n_483, n_484);
  xor g338 (n_485, A[55], B[55]);
  xor g339 (Z[55], n_481, n_485);
  nand g340 (n_487, A[56], B[56]);
  nand g341 (n_488, A[56], n_486);
  nand g342 (n_489, B[56], n_486);
  nand g343 (n_491, n_487, n_488, n_489);
  xor g344 (n_490, A[56], B[56]);
  xor g345 (Z[56], n_486, n_490);
  nand g346 (n_492, A[57], B[57]);
  nand g347 (n_493, A[57], n_491);
  nand g348 (n_494, B[57], n_491);
  nand g349 (n_496, n_492, n_493, n_494);
  xor g350 (n_495, A[57], B[57]);
  xor g351 (Z[57], n_491, n_495);
  nand g352 (n_497, A[58], B[58]);
  nand g353 (n_498, A[58], n_496);
  nand g354 (n_499, B[58], n_496);
  nand g355 (n_501, n_497, n_498, n_499);
  xor g356 (n_500, A[58], B[58]);
  xor g357 (Z[58], n_496, n_500);
  nand g358 (n_502, A[59], B[59]);
  nand g359 (n_503, A[59], n_501);
  nand g360 (n_504, B[59], n_501);
  nand g361 (n_506, n_502, n_503, n_504);
  xor g362 (n_505, A[59], B[59]);
  xor g363 (Z[59], n_501, n_505);
  nand g364 (n_507, A[60], B[60]);
  nand g365 (n_508, A[60], n_506);
  nand g366 (n_509, B[60], n_506);
  nand g367 (n_511, n_507, n_508, n_509);
  xor g368 (n_510, A[60], B[60]);
  xor g369 (Z[60], n_506, n_510);
  nand g370 (n_512, A[61], B[61]);
  nand g371 (n_513, A[61], n_511);
  nand g372 (n_514, B[61], n_511);
  nand g373 (n_516, n_512, n_513, n_514);
  xor g374 (n_515, A[61], B[61]);
  xor g375 (Z[61], n_511, n_515);
  nand g376 (n_517, A[62], B[62]);
  nand g377 (n_518, A[62], n_516);
  nand g378 (n_519, B[62], n_516);
  nand g379 (n_521, n_517, n_518, n_519);
  xor g380 (n_520, A[62], B[62]);
  xor g381 (Z[62], n_516, n_520);
  nand g382 (n_522, A[63], B[63]);
  nand g383 (n_523, A[63], n_521);
  nand g384 (n_524, B[63], n_521);
  nand g385 (n_526, n_522, n_523, n_524);
  xor g386 (n_525, A[63], B[63]);
  xor g387 (Z[63], n_521, n_525);
  nand g388 (n_527, A[64], B[64]);
  nand g389 (n_528, A[64], n_526);
  nand g390 (n_529, B[64], n_526);
  nand g391 (n_531, n_527, n_528, n_529);
  xor g392 (n_530, A[64], B[64]);
  xor g393 (Z[64], n_526, n_530);
  nand g394 (n_532, A[65], B[65]);
  nand g395 (n_533, A[65], n_531);
  nand g396 (n_534, B[65], n_531);
  nand g397 (n_536, n_532, n_533, n_534);
  xor g398 (n_535, A[65], B[65]);
  xor g399 (Z[65], n_531, n_535);
  nand g403 (n_206, n_537, n_538, n_539);
  xor g405 (Z[66], n_536, n_540);
  or g407 (n_537, A[66], B[66]);
  xor g408 (n_540, A[66], B[66]);
  or g409 (n_213, wc, n_207);
  not gc (wc, A[1]);
  or g410 (n_214, wc0, n_207);
  not gc0 (wc0, B[1]);
  xnor g411 (Z[1], n_207, n_215);
  or g412 (n_538, A[66], wc1);
  not gc1 (wc1, n_536);
  or g413 (n_539, B[66], wc2);
  not gc2 (wc2, n_536);
endmodule

module add_signed_1220_GENERIC(A, B, Z);
  input [66:0] A, B;
  output [67:0] Z;
  wire [66:0] A, B;
  wire [67:0] Z;
  add_signed_1220_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_1220_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [66:0] A, B;
  output [67:0] Z;
  wire [66:0] A, B;
  wire [67:0] Z;
  wire n_206, n_207, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540;
  not g3 (Z[67], n_206);
  nand g4 (n_207, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_212, A[1], B[1]);
  nand g13 (n_216, n_212, n_213, n_214);
  xor g14 (n_215, A[1], B[1]);
  nand g16 (n_217, A[2], B[2]);
  nand g17 (n_218, A[2], n_216);
  nand g18 (n_219, B[2], n_216);
  nand g19 (n_221, n_217, n_218, n_219);
  xor g20 (n_220, A[2], B[2]);
  xor g21 (Z[2], n_216, n_220);
  nand g22 (n_222, A[3], B[3]);
  nand g23 (n_223, A[3], n_221);
  nand g24 (n_224, B[3], n_221);
  nand g25 (n_226, n_222, n_223, n_224);
  xor g26 (n_225, A[3], B[3]);
  xor g27 (Z[3], n_221, n_225);
  nand g28 (n_227, A[4], B[4]);
  nand g29 (n_228, A[4], n_226);
  nand g30 (n_229, B[4], n_226);
  nand g31 (n_231, n_227, n_228, n_229);
  xor g32 (n_230, A[4], B[4]);
  xor g33 (Z[4], n_226, n_230);
  nand g34 (n_232, A[5], B[5]);
  nand g35 (n_233, A[5], n_231);
  nand g36 (n_234, B[5], n_231);
  nand g37 (n_236, n_232, n_233, n_234);
  xor g38 (n_235, A[5], B[5]);
  xor g39 (Z[5], n_231, n_235);
  nand g40 (n_237, A[6], B[6]);
  nand g41 (n_238, A[6], n_236);
  nand g42 (n_239, B[6], n_236);
  nand g43 (n_241, n_237, n_238, n_239);
  xor g44 (n_240, A[6], B[6]);
  xor g45 (Z[6], n_236, n_240);
  nand g46 (n_242, A[7], B[7]);
  nand g47 (n_243, A[7], n_241);
  nand g48 (n_244, B[7], n_241);
  nand g49 (n_246, n_242, n_243, n_244);
  xor g50 (n_245, A[7], B[7]);
  xor g51 (Z[7], n_241, n_245);
  nand g52 (n_247, A[8], B[8]);
  nand g53 (n_248, A[8], n_246);
  nand g54 (n_249, B[8], n_246);
  nand g55 (n_251, n_247, n_248, n_249);
  xor g56 (n_250, A[8], B[8]);
  xor g57 (Z[8], n_246, n_250);
  nand g58 (n_252, A[9], B[9]);
  nand g59 (n_253, A[9], n_251);
  nand g60 (n_254, B[9], n_251);
  nand g61 (n_256, n_252, n_253, n_254);
  xor g62 (n_255, A[9], B[9]);
  xor g63 (Z[9], n_251, n_255);
  nand g64 (n_257, A[10], B[10]);
  nand g65 (n_258, A[10], n_256);
  nand g66 (n_259, B[10], n_256);
  nand g67 (n_261, n_257, n_258, n_259);
  xor g68 (n_260, A[10], B[10]);
  xor g69 (Z[10], n_256, n_260);
  nand g70 (n_262, A[11], B[11]);
  nand g71 (n_263, A[11], n_261);
  nand g72 (n_264, B[11], n_261);
  nand g73 (n_266, n_262, n_263, n_264);
  xor g74 (n_265, A[11], B[11]);
  xor g75 (Z[11], n_261, n_265);
  nand g76 (n_267, A[12], B[12]);
  nand g77 (n_268, A[12], n_266);
  nand g78 (n_269, B[12], n_266);
  nand g79 (n_271, n_267, n_268, n_269);
  xor g80 (n_270, A[12], B[12]);
  xor g81 (Z[12], n_266, n_270);
  nand g82 (n_272, A[13], B[13]);
  nand g83 (n_273, A[13], n_271);
  nand g84 (n_274, B[13], n_271);
  nand g85 (n_276, n_272, n_273, n_274);
  xor g86 (n_275, A[13], B[13]);
  xor g87 (Z[13], n_271, n_275);
  nand g88 (n_277, A[14], B[14]);
  nand g89 (n_278, A[14], n_276);
  nand g90 (n_279, B[14], n_276);
  nand g91 (n_281, n_277, n_278, n_279);
  xor g92 (n_280, A[14], B[14]);
  xor g93 (Z[14], n_276, n_280);
  nand g94 (n_282, A[15], B[15]);
  nand g95 (n_283, A[15], n_281);
  nand g96 (n_284, B[15], n_281);
  nand g97 (n_286, n_282, n_283, n_284);
  xor g98 (n_285, A[15], B[15]);
  xor g99 (Z[15], n_281, n_285);
  nand g100 (n_287, A[16], B[16]);
  nand g101 (n_288, A[16], n_286);
  nand g102 (n_289, B[16], n_286);
  nand g103 (n_291, n_287, n_288, n_289);
  xor g104 (n_290, A[16], B[16]);
  xor g105 (Z[16], n_286, n_290);
  nand g106 (n_292, A[17], B[17]);
  nand g107 (n_293, A[17], n_291);
  nand g108 (n_294, B[17], n_291);
  nand g109 (n_296, n_292, n_293, n_294);
  xor g110 (n_295, A[17], B[17]);
  xor g111 (Z[17], n_291, n_295);
  nand g112 (n_297, A[18], B[18]);
  nand g113 (n_298, A[18], n_296);
  nand g114 (n_299, B[18], n_296);
  nand g115 (n_301, n_297, n_298, n_299);
  xor g116 (n_300, A[18], B[18]);
  xor g117 (Z[18], n_296, n_300);
  nand g118 (n_302, A[19], B[19]);
  nand g119 (n_303, A[19], n_301);
  nand g120 (n_304, B[19], n_301);
  nand g121 (n_306, n_302, n_303, n_304);
  xor g122 (n_305, A[19], B[19]);
  xor g123 (Z[19], n_301, n_305);
  nand g124 (n_307, A[20], B[20]);
  nand g125 (n_308, A[20], n_306);
  nand g126 (n_309, B[20], n_306);
  nand g127 (n_311, n_307, n_308, n_309);
  xor g128 (n_310, A[20], B[20]);
  xor g129 (Z[20], n_306, n_310);
  nand g130 (n_312, A[21], B[21]);
  nand g131 (n_313, A[21], n_311);
  nand g132 (n_314, B[21], n_311);
  nand g133 (n_316, n_312, n_313, n_314);
  xor g134 (n_315, A[21], B[21]);
  xor g135 (Z[21], n_311, n_315);
  nand g136 (n_317, A[22], B[22]);
  nand g137 (n_318, A[22], n_316);
  nand g138 (n_319, B[22], n_316);
  nand g139 (n_321, n_317, n_318, n_319);
  xor g140 (n_320, A[22], B[22]);
  xor g141 (Z[22], n_316, n_320);
  nand g142 (n_322, A[23], B[23]);
  nand g143 (n_323, A[23], n_321);
  nand g144 (n_324, B[23], n_321);
  nand g145 (n_326, n_322, n_323, n_324);
  xor g146 (n_325, A[23], B[23]);
  xor g147 (Z[23], n_321, n_325);
  nand g148 (n_327, A[24], B[24]);
  nand g149 (n_328, A[24], n_326);
  nand g150 (n_329, B[24], n_326);
  nand g151 (n_331, n_327, n_328, n_329);
  xor g152 (n_330, A[24], B[24]);
  xor g153 (Z[24], n_326, n_330);
  nand g154 (n_332, A[25], B[25]);
  nand g155 (n_333, A[25], n_331);
  nand g156 (n_334, B[25], n_331);
  nand g157 (n_336, n_332, n_333, n_334);
  xor g158 (n_335, A[25], B[25]);
  xor g159 (Z[25], n_331, n_335);
  nand g160 (n_337, A[26], B[26]);
  nand g161 (n_338, A[26], n_336);
  nand g162 (n_339, B[26], n_336);
  nand g163 (n_341, n_337, n_338, n_339);
  xor g164 (n_340, A[26], B[26]);
  xor g165 (Z[26], n_336, n_340);
  nand g166 (n_342, A[27], B[27]);
  nand g167 (n_343, A[27], n_341);
  nand g168 (n_344, B[27], n_341);
  nand g169 (n_346, n_342, n_343, n_344);
  xor g170 (n_345, A[27], B[27]);
  xor g171 (Z[27], n_341, n_345);
  nand g172 (n_347, A[28], B[28]);
  nand g173 (n_348, A[28], n_346);
  nand g174 (n_349, B[28], n_346);
  nand g175 (n_351, n_347, n_348, n_349);
  xor g176 (n_350, A[28], B[28]);
  xor g177 (Z[28], n_346, n_350);
  nand g178 (n_352, A[29], B[29]);
  nand g179 (n_353, A[29], n_351);
  nand g180 (n_354, B[29], n_351);
  nand g181 (n_356, n_352, n_353, n_354);
  xor g182 (n_355, A[29], B[29]);
  xor g183 (Z[29], n_351, n_355);
  nand g184 (n_357, A[30], B[30]);
  nand g185 (n_358, A[30], n_356);
  nand g186 (n_359, B[30], n_356);
  nand g187 (n_361, n_357, n_358, n_359);
  xor g188 (n_360, A[30], B[30]);
  xor g189 (Z[30], n_356, n_360);
  nand g190 (n_362, A[31], B[31]);
  nand g191 (n_363, A[31], n_361);
  nand g192 (n_364, B[31], n_361);
  nand g193 (n_366, n_362, n_363, n_364);
  xor g194 (n_365, A[31], B[31]);
  xor g195 (Z[31], n_361, n_365);
  nand g196 (n_367, A[32], B[32]);
  nand g197 (n_368, A[32], n_366);
  nand g198 (n_369, B[32], n_366);
  nand g199 (n_371, n_367, n_368, n_369);
  xor g200 (n_370, A[32], B[32]);
  xor g201 (Z[32], n_366, n_370);
  nand g202 (n_372, A[33], B[33]);
  nand g203 (n_373, A[33], n_371);
  nand g204 (n_374, B[33], n_371);
  nand g205 (n_376, n_372, n_373, n_374);
  xor g206 (n_375, A[33], B[33]);
  xor g207 (Z[33], n_371, n_375);
  nand g208 (n_377, A[34], B[34]);
  nand g209 (n_378, A[34], n_376);
  nand g210 (n_379, B[34], n_376);
  nand g211 (n_381, n_377, n_378, n_379);
  xor g212 (n_380, A[34], B[34]);
  xor g213 (Z[34], n_376, n_380);
  nand g214 (n_382, A[35], B[35]);
  nand g215 (n_383, A[35], n_381);
  nand g216 (n_384, B[35], n_381);
  nand g217 (n_386, n_382, n_383, n_384);
  xor g218 (n_385, A[35], B[35]);
  xor g219 (Z[35], n_381, n_385);
  nand g220 (n_387, A[36], B[36]);
  nand g221 (n_388, A[36], n_386);
  nand g222 (n_389, B[36], n_386);
  nand g223 (n_391, n_387, n_388, n_389);
  xor g224 (n_390, A[36], B[36]);
  xor g225 (Z[36], n_386, n_390);
  nand g226 (n_392, A[37], B[37]);
  nand g227 (n_393, A[37], n_391);
  nand g228 (n_394, B[37], n_391);
  nand g229 (n_396, n_392, n_393, n_394);
  xor g230 (n_395, A[37], B[37]);
  xor g231 (Z[37], n_391, n_395);
  nand g232 (n_397, A[38], B[38]);
  nand g233 (n_398, A[38], n_396);
  nand g234 (n_399, B[38], n_396);
  nand g235 (n_401, n_397, n_398, n_399);
  xor g236 (n_400, A[38], B[38]);
  xor g237 (Z[38], n_396, n_400);
  nand g238 (n_402, A[39], B[39]);
  nand g239 (n_403, A[39], n_401);
  nand g240 (n_404, B[39], n_401);
  nand g241 (n_406, n_402, n_403, n_404);
  xor g242 (n_405, A[39], B[39]);
  xor g243 (Z[39], n_401, n_405);
  nand g244 (n_407, A[40], B[40]);
  nand g245 (n_408, A[40], n_406);
  nand g246 (n_409, B[40], n_406);
  nand g247 (n_411, n_407, n_408, n_409);
  xor g248 (n_410, A[40], B[40]);
  xor g249 (Z[40], n_406, n_410);
  nand g250 (n_412, A[41], B[41]);
  nand g251 (n_413, A[41], n_411);
  nand g252 (n_414, B[41], n_411);
  nand g253 (n_416, n_412, n_413, n_414);
  xor g254 (n_415, A[41], B[41]);
  xor g255 (Z[41], n_411, n_415);
  nand g256 (n_417, A[42], B[42]);
  nand g257 (n_418, A[42], n_416);
  nand g258 (n_419, B[42], n_416);
  nand g259 (n_421, n_417, n_418, n_419);
  xor g260 (n_420, A[42], B[42]);
  xor g261 (Z[42], n_416, n_420);
  nand g262 (n_422, A[43], B[43]);
  nand g263 (n_423, A[43], n_421);
  nand g264 (n_424, B[43], n_421);
  nand g265 (n_426, n_422, n_423, n_424);
  xor g266 (n_425, A[43], B[43]);
  xor g267 (Z[43], n_421, n_425);
  nand g268 (n_427, A[44], B[44]);
  nand g269 (n_428, A[44], n_426);
  nand g270 (n_429, B[44], n_426);
  nand g271 (n_431, n_427, n_428, n_429);
  xor g272 (n_430, A[44], B[44]);
  xor g273 (Z[44], n_426, n_430);
  nand g274 (n_432, A[45], B[45]);
  nand g275 (n_433, A[45], n_431);
  nand g276 (n_434, B[45], n_431);
  nand g277 (n_436, n_432, n_433, n_434);
  xor g278 (n_435, A[45], B[45]);
  xor g279 (Z[45], n_431, n_435);
  nand g280 (n_437, A[46], B[46]);
  nand g281 (n_438, A[46], n_436);
  nand g282 (n_439, B[46], n_436);
  nand g283 (n_441, n_437, n_438, n_439);
  xor g284 (n_440, A[46], B[46]);
  xor g285 (Z[46], n_436, n_440);
  nand g286 (n_442, A[47], B[47]);
  nand g287 (n_443, A[47], n_441);
  nand g288 (n_444, B[47], n_441);
  nand g289 (n_446, n_442, n_443, n_444);
  xor g290 (n_445, A[47], B[47]);
  xor g291 (Z[47], n_441, n_445);
  nand g292 (n_447, A[48], B[48]);
  nand g293 (n_448, A[48], n_446);
  nand g294 (n_449, B[48], n_446);
  nand g295 (n_451, n_447, n_448, n_449);
  xor g296 (n_450, A[48], B[48]);
  xor g297 (Z[48], n_446, n_450);
  nand g298 (n_452, A[49], B[49]);
  nand g299 (n_453, A[49], n_451);
  nand g300 (n_454, B[49], n_451);
  nand g301 (n_456, n_452, n_453, n_454);
  xor g302 (n_455, A[49], B[49]);
  xor g303 (Z[49], n_451, n_455);
  nand g304 (n_457, A[50], B[50]);
  nand g305 (n_458, A[50], n_456);
  nand g306 (n_459, B[50], n_456);
  nand g307 (n_461, n_457, n_458, n_459);
  xor g308 (n_460, A[50], B[50]);
  xor g309 (Z[50], n_456, n_460);
  nand g310 (n_462, A[51], B[51]);
  nand g311 (n_463, A[51], n_461);
  nand g312 (n_464, B[51], n_461);
  nand g313 (n_466, n_462, n_463, n_464);
  xor g314 (n_465, A[51], B[51]);
  xor g315 (Z[51], n_461, n_465);
  nand g316 (n_467, A[52], B[52]);
  nand g317 (n_468, A[52], n_466);
  nand g318 (n_469, B[52], n_466);
  nand g319 (n_471, n_467, n_468, n_469);
  xor g320 (n_470, A[52], B[52]);
  xor g321 (Z[52], n_466, n_470);
  nand g322 (n_472, A[53], B[53]);
  nand g323 (n_473, A[53], n_471);
  nand g324 (n_474, B[53], n_471);
  nand g325 (n_476, n_472, n_473, n_474);
  xor g326 (n_475, A[53], B[53]);
  xor g327 (Z[53], n_471, n_475);
  nand g328 (n_477, A[54], B[54]);
  nand g329 (n_478, A[54], n_476);
  nand g330 (n_479, B[54], n_476);
  nand g331 (n_481, n_477, n_478, n_479);
  xor g332 (n_480, A[54], B[54]);
  xor g333 (Z[54], n_476, n_480);
  nand g334 (n_482, A[55], B[55]);
  nand g335 (n_483, A[55], n_481);
  nand g336 (n_484, B[55], n_481);
  nand g337 (n_486, n_482, n_483, n_484);
  xor g338 (n_485, A[55], B[55]);
  xor g339 (Z[55], n_481, n_485);
  nand g340 (n_487, A[56], B[56]);
  nand g341 (n_488, A[56], n_486);
  nand g342 (n_489, B[56], n_486);
  nand g343 (n_491, n_487, n_488, n_489);
  xor g344 (n_490, A[56], B[56]);
  xor g345 (Z[56], n_486, n_490);
  nand g346 (n_492, A[57], B[57]);
  nand g347 (n_493, A[57], n_491);
  nand g348 (n_494, B[57], n_491);
  nand g349 (n_496, n_492, n_493, n_494);
  xor g350 (n_495, A[57], B[57]);
  xor g351 (Z[57], n_491, n_495);
  nand g352 (n_497, A[58], B[58]);
  nand g353 (n_498, A[58], n_496);
  nand g354 (n_499, B[58], n_496);
  nand g355 (n_501, n_497, n_498, n_499);
  xor g356 (n_500, A[58], B[58]);
  xor g357 (Z[58], n_496, n_500);
  nand g358 (n_502, A[59], B[59]);
  nand g359 (n_503, A[59], n_501);
  nand g360 (n_504, B[59], n_501);
  nand g361 (n_506, n_502, n_503, n_504);
  xor g362 (n_505, A[59], B[59]);
  xor g363 (Z[59], n_501, n_505);
  nand g364 (n_507, A[60], B[60]);
  nand g365 (n_508, A[60], n_506);
  nand g366 (n_509, B[60], n_506);
  nand g367 (n_511, n_507, n_508, n_509);
  xor g368 (n_510, A[60], B[60]);
  xor g369 (Z[60], n_506, n_510);
  nand g370 (n_512, A[61], B[61]);
  nand g371 (n_513, A[61], n_511);
  nand g372 (n_514, B[61], n_511);
  nand g373 (n_516, n_512, n_513, n_514);
  xor g374 (n_515, A[61], B[61]);
  xor g375 (Z[61], n_511, n_515);
  nand g376 (n_517, A[62], B[62]);
  nand g377 (n_518, A[62], n_516);
  nand g378 (n_519, B[62], n_516);
  nand g379 (n_521, n_517, n_518, n_519);
  xor g380 (n_520, A[62], B[62]);
  xor g381 (Z[62], n_516, n_520);
  nand g382 (n_522, A[63], B[63]);
  nand g383 (n_523, A[63], n_521);
  nand g384 (n_524, B[63], n_521);
  nand g385 (n_526, n_522, n_523, n_524);
  xor g386 (n_525, A[63], B[63]);
  xor g387 (Z[63], n_521, n_525);
  nand g388 (n_527, A[64], B[64]);
  nand g389 (n_528, A[64], n_526);
  nand g390 (n_529, B[64], n_526);
  nand g391 (n_531, n_527, n_528, n_529);
  xor g392 (n_530, A[64], B[64]);
  xor g393 (Z[64], n_526, n_530);
  nand g394 (n_532, A[65], B[65]);
  nand g395 (n_533, A[65], n_531);
  nand g396 (n_534, B[65], n_531);
  nand g397 (n_536, n_532, n_533, n_534);
  xor g398 (n_535, A[65], B[65]);
  xor g399 (Z[65], n_531, n_535);
  nand g403 (n_206, n_537, n_538, n_539);
  xor g405 (Z[66], n_536, n_540);
  or g407 (n_537, A[66], B[66]);
  xor g408 (n_540, A[66], B[66]);
  or g409 (n_213, wc, n_207);
  not gc (wc, A[1]);
  or g410 (n_214, wc0, n_207);
  not gc0 (wc0, B[1]);
  xnor g411 (Z[1], n_207, n_215);
  or g412 (n_538, A[66], wc1);
  not gc1 (wc1, n_536);
  or g413 (n_539, B[66], wc2);
  not gc2 (wc2, n_536);
endmodule

module add_signed_1220_1_GENERIC(A, B, Z);
  input [66:0] A, B;
  output [67:0] Z;
  wire [66:0] A, B;
  wire [67:0] Z;
  add_signed_1220_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_1220_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [66:0] A, B;
  output [67:0] Z;
  wire [66:0] A, B;
  wire [67:0] Z;
  wire n_206, n_207, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540;
  not g3 (Z[67], n_206);
  nand g4 (n_207, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_212, A[1], B[1]);
  nand g13 (n_216, n_212, n_213, n_214);
  xor g14 (n_215, A[1], B[1]);
  nand g16 (n_217, A[2], B[2]);
  nand g17 (n_218, A[2], n_216);
  nand g18 (n_219, B[2], n_216);
  nand g19 (n_221, n_217, n_218, n_219);
  xor g20 (n_220, A[2], B[2]);
  xor g21 (Z[2], n_216, n_220);
  nand g22 (n_222, A[3], B[3]);
  nand g23 (n_223, A[3], n_221);
  nand g24 (n_224, B[3], n_221);
  nand g25 (n_226, n_222, n_223, n_224);
  xor g26 (n_225, A[3], B[3]);
  xor g27 (Z[3], n_221, n_225);
  nand g28 (n_227, A[4], B[4]);
  nand g29 (n_228, A[4], n_226);
  nand g30 (n_229, B[4], n_226);
  nand g31 (n_231, n_227, n_228, n_229);
  xor g32 (n_230, A[4], B[4]);
  xor g33 (Z[4], n_226, n_230);
  nand g34 (n_232, A[5], B[5]);
  nand g35 (n_233, A[5], n_231);
  nand g36 (n_234, B[5], n_231);
  nand g37 (n_236, n_232, n_233, n_234);
  xor g38 (n_235, A[5], B[5]);
  xor g39 (Z[5], n_231, n_235);
  nand g40 (n_237, A[6], B[6]);
  nand g41 (n_238, A[6], n_236);
  nand g42 (n_239, B[6], n_236);
  nand g43 (n_241, n_237, n_238, n_239);
  xor g44 (n_240, A[6], B[6]);
  xor g45 (Z[6], n_236, n_240);
  nand g46 (n_242, A[7], B[7]);
  nand g47 (n_243, A[7], n_241);
  nand g48 (n_244, B[7], n_241);
  nand g49 (n_246, n_242, n_243, n_244);
  xor g50 (n_245, A[7], B[7]);
  xor g51 (Z[7], n_241, n_245);
  nand g52 (n_247, A[8], B[8]);
  nand g53 (n_248, A[8], n_246);
  nand g54 (n_249, B[8], n_246);
  nand g55 (n_251, n_247, n_248, n_249);
  xor g56 (n_250, A[8], B[8]);
  xor g57 (Z[8], n_246, n_250);
  nand g58 (n_252, A[9], B[9]);
  nand g59 (n_253, A[9], n_251);
  nand g60 (n_254, B[9], n_251);
  nand g61 (n_256, n_252, n_253, n_254);
  xor g62 (n_255, A[9], B[9]);
  xor g63 (Z[9], n_251, n_255);
  nand g64 (n_257, A[10], B[10]);
  nand g65 (n_258, A[10], n_256);
  nand g66 (n_259, B[10], n_256);
  nand g67 (n_261, n_257, n_258, n_259);
  xor g68 (n_260, A[10], B[10]);
  xor g69 (Z[10], n_256, n_260);
  nand g70 (n_262, A[11], B[11]);
  nand g71 (n_263, A[11], n_261);
  nand g72 (n_264, B[11], n_261);
  nand g73 (n_266, n_262, n_263, n_264);
  xor g74 (n_265, A[11], B[11]);
  xor g75 (Z[11], n_261, n_265);
  nand g76 (n_267, A[12], B[12]);
  nand g77 (n_268, A[12], n_266);
  nand g78 (n_269, B[12], n_266);
  nand g79 (n_271, n_267, n_268, n_269);
  xor g80 (n_270, A[12], B[12]);
  xor g81 (Z[12], n_266, n_270);
  nand g82 (n_272, A[13], B[13]);
  nand g83 (n_273, A[13], n_271);
  nand g84 (n_274, B[13], n_271);
  nand g85 (n_276, n_272, n_273, n_274);
  xor g86 (n_275, A[13], B[13]);
  xor g87 (Z[13], n_271, n_275);
  nand g88 (n_277, A[14], B[14]);
  nand g89 (n_278, A[14], n_276);
  nand g90 (n_279, B[14], n_276);
  nand g91 (n_281, n_277, n_278, n_279);
  xor g92 (n_280, A[14], B[14]);
  xor g93 (Z[14], n_276, n_280);
  nand g94 (n_282, A[15], B[15]);
  nand g95 (n_283, A[15], n_281);
  nand g96 (n_284, B[15], n_281);
  nand g97 (n_286, n_282, n_283, n_284);
  xor g98 (n_285, A[15], B[15]);
  xor g99 (Z[15], n_281, n_285);
  nand g100 (n_287, A[16], B[16]);
  nand g101 (n_288, A[16], n_286);
  nand g102 (n_289, B[16], n_286);
  nand g103 (n_291, n_287, n_288, n_289);
  xor g104 (n_290, A[16], B[16]);
  xor g105 (Z[16], n_286, n_290);
  nand g106 (n_292, A[17], B[17]);
  nand g107 (n_293, A[17], n_291);
  nand g108 (n_294, B[17], n_291);
  nand g109 (n_296, n_292, n_293, n_294);
  xor g110 (n_295, A[17], B[17]);
  xor g111 (Z[17], n_291, n_295);
  nand g112 (n_297, A[18], B[18]);
  nand g113 (n_298, A[18], n_296);
  nand g114 (n_299, B[18], n_296);
  nand g115 (n_301, n_297, n_298, n_299);
  xor g116 (n_300, A[18], B[18]);
  xor g117 (Z[18], n_296, n_300);
  nand g118 (n_302, A[19], B[19]);
  nand g119 (n_303, A[19], n_301);
  nand g120 (n_304, B[19], n_301);
  nand g121 (n_306, n_302, n_303, n_304);
  xor g122 (n_305, A[19], B[19]);
  xor g123 (Z[19], n_301, n_305);
  nand g124 (n_307, A[20], B[20]);
  nand g125 (n_308, A[20], n_306);
  nand g126 (n_309, B[20], n_306);
  nand g127 (n_311, n_307, n_308, n_309);
  xor g128 (n_310, A[20], B[20]);
  xor g129 (Z[20], n_306, n_310);
  nand g130 (n_312, A[21], B[21]);
  nand g131 (n_313, A[21], n_311);
  nand g132 (n_314, B[21], n_311);
  nand g133 (n_316, n_312, n_313, n_314);
  xor g134 (n_315, A[21], B[21]);
  xor g135 (Z[21], n_311, n_315);
  nand g136 (n_317, A[22], B[22]);
  nand g137 (n_318, A[22], n_316);
  nand g138 (n_319, B[22], n_316);
  nand g139 (n_321, n_317, n_318, n_319);
  xor g140 (n_320, A[22], B[22]);
  xor g141 (Z[22], n_316, n_320);
  nand g142 (n_322, A[23], B[23]);
  nand g143 (n_323, A[23], n_321);
  nand g144 (n_324, B[23], n_321);
  nand g145 (n_326, n_322, n_323, n_324);
  xor g146 (n_325, A[23], B[23]);
  xor g147 (Z[23], n_321, n_325);
  nand g148 (n_327, A[24], B[24]);
  nand g149 (n_328, A[24], n_326);
  nand g150 (n_329, B[24], n_326);
  nand g151 (n_331, n_327, n_328, n_329);
  xor g152 (n_330, A[24], B[24]);
  xor g153 (Z[24], n_326, n_330);
  nand g154 (n_332, A[25], B[25]);
  nand g155 (n_333, A[25], n_331);
  nand g156 (n_334, B[25], n_331);
  nand g157 (n_336, n_332, n_333, n_334);
  xor g158 (n_335, A[25], B[25]);
  xor g159 (Z[25], n_331, n_335);
  nand g160 (n_337, A[26], B[26]);
  nand g161 (n_338, A[26], n_336);
  nand g162 (n_339, B[26], n_336);
  nand g163 (n_341, n_337, n_338, n_339);
  xor g164 (n_340, A[26], B[26]);
  xor g165 (Z[26], n_336, n_340);
  nand g166 (n_342, A[27], B[27]);
  nand g167 (n_343, A[27], n_341);
  nand g168 (n_344, B[27], n_341);
  nand g169 (n_346, n_342, n_343, n_344);
  xor g170 (n_345, A[27], B[27]);
  xor g171 (Z[27], n_341, n_345);
  nand g172 (n_347, A[28], B[28]);
  nand g173 (n_348, A[28], n_346);
  nand g174 (n_349, B[28], n_346);
  nand g175 (n_351, n_347, n_348, n_349);
  xor g176 (n_350, A[28], B[28]);
  xor g177 (Z[28], n_346, n_350);
  nand g178 (n_352, A[29], B[29]);
  nand g179 (n_353, A[29], n_351);
  nand g180 (n_354, B[29], n_351);
  nand g181 (n_356, n_352, n_353, n_354);
  xor g182 (n_355, A[29], B[29]);
  xor g183 (Z[29], n_351, n_355);
  nand g184 (n_357, A[30], B[30]);
  nand g185 (n_358, A[30], n_356);
  nand g186 (n_359, B[30], n_356);
  nand g187 (n_361, n_357, n_358, n_359);
  xor g188 (n_360, A[30], B[30]);
  xor g189 (Z[30], n_356, n_360);
  nand g190 (n_362, A[31], B[31]);
  nand g191 (n_363, A[31], n_361);
  nand g192 (n_364, B[31], n_361);
  nand g193 (n_366, n_362, n_363, n_364);
  xor g194 (n_365, A[31], B[31]);
  xor g195 (Z[31], n_361, n_365);
  nand g196 (n_367, A[32], B[32]);
  nand g197 (n_368, A[32], n_366);
  nand g198 (n_369, B[32], n_366);
  nand g199 (n_371, n_367, n_368, n_369);
  xor g200 (n_370, A[32], B[32]);
  xor g201 (Z[32], n_366, n_370);
  nand g202 (n_372, A[33], B[33]);
  nand g203 (n_373, A[33], n_371);
  nand g204 (n_374, B[33], n_371);
  nand g205 (n_376, n_372, n_373, n_374);
  xor g206 (n_375, A[33], B[33]);
  xor g207 (Z[33], n_371, n_375);
  nand g208 (n_377, A[34], B[34]);
  nand g209 (n_378, A[34], n_376);
  nand g210 (n_379, B[34], n_376);
  nand g211 (n_381, n_377, n_378, n_379);
  xor g212 (n_380, A[34], B[34]);
  xor g213 (Z[34], n_376, n_380);
  nand g214 (n_382, A[35], B[35]);
  nand g215 (n_383, A[35], n_381);
  nand g216 (n_384, B[35], n_381);
  nand g217 (n_386, n_382, n_383, n_384);
  xor g218 (n_385, A[35], B[35]);
  xor g219 (Z[35], n_381, n_385);
  nand g220 (n_387, A[36], B[36]);
  nand g221 (n_388, A[36], n_386);
  nand g222 (n_389, B[36], n_386);
  nand g223 (n_391, n_387, n_388, n_389);
  xor g224 (n_390, A[36], B[36]);
  xor g225 (Z[36], n_386, n_390);
  nand g226 (n_392, A[37], B[37]);
  nand g227 (n_393, A[37], n_391);
  nand g228 (n_394, B[37], n_391);
  nand g229 (n_396, n_392, n_393, n_394);
  xor g230 (n_395, A[37], B[37]);
  xor g231 (Z[37], n_391, n_395);
  nand g232 (n_397, A[38], B[38]);
  nand g233 (n_398, A[38], n_396);
  nand g234 (n_399, B[38], n_396);
  nand g235 (n_401, n_397, n_398, n_399);
  xor g236 (n_400, A[38], B[38]);
  xor g237 (Z[38], n_396, n_400);
  nand g238 (n_402, A[39], B[39]);
  nand g239 (n_403, A[39], n_401);
  nand g240 (n_404, B[39], n_401);
  nand g241 (n_406, n_402, n_403, n_404);
  xor g242 (n_405, A[39], B[39]);
  xor g243 (Z[39], n_401, n_405);
  nand g244 (n_407, A[40], B[40]);
  nand g245 (n_408, A[40], n_406);
  nand g246 (n_409, B[40], n_406);
  nand g247 (n_411, n_407, n_408, n_409);
  xor g248 (n_410, A[40], B[40]);
  xor g249 (Z[40], n_406, n_410);
  nand g250 (n_412, A[41], B[41]);
  nand g251 (n_413, A[41], n_411);
  nand g252 (n_414, B[41], n_411);
  nand g253 (n_416, n_412, n_413, n_414);
  xor g254 (n_415, A[41], B[41]);
  xor g255 (Z[41], n_411, n_415);
  nand g256 (n_417, A[42], B[42]);
  nand g257 (n_418, A[42], n_416);
  nand g258 (n_419, B[42], n_416);
  nand g259 (n_421, n_417, n_418, n_419);
  xor g260 (n_420, A[42], B[42]);
  xor g261 (Z[42], n_416, n_420);
  nand g262 (n_422, A[43], B[43]);
  nand g263 (n_423, A[43], n_421);
  nand g264 (n_424, B[43], n_421);
  nand g265 (n_426, n_422, n_423, n_424);
  xor g266 (n_425, A[43], B[43]);
  xor g267 (Z[43], n_421, n_425);
  nand g268 (n_427, A[44], B[44]);
  nand g269 (n_428, A[44], n_426);
  nand g270 (n_429, B[44], n_426);
  nand g271 (n_431, n_427, n_428, n_429);
  xor g272 (n_430, A[44], B[44]);
  xor g273 (Z[44], n_426, n_430);
  nand g274 (n_432, A[45], B[45]);
  nand g275 (n_433, A[45], n_431);
  nand g276 (n_434, B[45], n_431);
  nand g277 (n_436, n_432, n_433, n_434);
  xor g278 (n_435, A[45], B[45]);
  xor g279 (Z[45], n_431, n_435);
  nand g280 (n_437, A[46], B[46]);
  nand g281 (n_438, A[46], n_436);
  nand g282 (n_439, B[46], n_436);
  nand g283 (n_441, n_437, n_438, n_439);
  xor g284 (n_440, A[46], B[46]);
  xor g285 (Z[46], n_436, n_440);
  nand g286 (n_442, A[47], B[47]);
  nand g287 (n_443, A[47], n_441);
  nand g288 (n_444, B[47], n_441);
  nand g289 (n_446, n_442, n_443, n_444);
  xor g290 (n_445, A[47], B[47]);
  xor g291 (Z[47], n_441, n_445);
  nand g292 (n_447, A[48], B[48]);
  nand g293 (n_448, A[48], n_446);
  nand g294 (n_449, B[48], n_446);
  nand g295 (n_451, n_447, n_448, n_449);
  xor g296 (n_450, A[48], B[48]);
  xor g297 (Z[48], n_446, n_450);
  nand g298 (n_452, A[49], B[49]);
  nand g299 (n_453, A[49], n_451);
  nand g300 (n_454, B[49], n_451);
  nand g301 (n_456, n_452, n_453, n_454);
  xor g302 (n_455, A[49], B[49]);
  xor g303 (Z[49], n_451, n_455);
  nand g304 (n_457, A[50], B[50]);
  nand g305 (n_458, A[50], n_456);
  nand g306 (n_459, B[50], n_456);
  nand g307 (n_461, n_457, n_458, n_459);
  xor g308 (n_460, A[50], B[50]);
  xor g309 (Z[50], n_456, n_460);
  nand g310 (n_462, A[51], B[51]);
  nand g311 (n_463, A[51], n_461);
  nand g312 (n_464, B[51], n_461);
  nand g313 (n_466, n_462, n_463, n_464);
  xor g314 (n_465, A[51], B[51]);
  xor g315 (Z[51], n_461, n_465);
  nand g316 (n_467, A[52], B[52]);
  nand g317 (n_468, A[52], n_466);
  nand g318 (n_469, B[52], n_466);
  nand g319 (n_471, n_467, n_468, n_469);
  xor g320 (n_470, A[52], B[52]);
  xor g321 (Z[52], n_466, n_470);
  nand g322 (n_472, A[53], B[53]);
  nand g323 (n_473, A[53], n_471);
  nand g324 (n_474, B[53], n_471);
  nand g325 (n_476, n_472, n_473, n_474);
  xor g326 (n_475, A[53], B[53]);
  xor g327 (Z[53], n_471, n_475);
  nand g328 (n_477, A[54], B[54]);
  nand g329 (n_478, A[54], n_476);
  nand g330 (n_479, B[54], n_476);
  nand g331 (n_481, n_477, n_478, n_479);
  xor g332 (n_480, A[54], B[54]);
  xor g333 (Z[54], n_476, n_480);
  nand g334 (n_482, A[55], B[55]);
  nand g335 (n_483, A[55], n_481);
  nand g336 (n_484, B[55], n_481);
  nand g337 (n_486, n_482, n_483, n_484);
  xor g338 (n_485, A[55], B[55]);
  xor g339 (Z[55], n_481, n_485);
  nand g340 (n_487, A[56], B[56]);
  nand g341 (n_488, A[56], n_486);
  nand g342 (n_489, B[56], n_486);
  nand g343 (n_491, n_487, n_488, n_489);
  xor g344 (n_490, A[56], B[56]);
  xor g345 (Z[56], n_486, n_490);
  nand g346 (n_492, A[57], B[57]);
  nand g347 (n_493, A[57], n_491);
  nand g348 (n_494, B[57], n_491);
  nand g349 (n_496, n_492, n_493, n_494);
  xor g350 (n_495, A[57], B[57]);
  xor g351 (Z[57], n_491, n_495);
  nand g352 (n_497, A[58], B[58]);
  nand g353 (n_498, A[58], n_496);
  nand g354 (n_499, B[58], n_496);
  nand g355 (n_501, n_497, n_498, n_499);
  xor g356 (n_500, A[58], B[58]);
  xor g357 (Z[58], n_496, n_500);
  nand g358 (n_502, A[59], B[59]);
  nand g359 (n_503, A[59], n_501);
  nand g360 (n_504, B[59], n_501);
  nand g361 (n_506, n_502, n_503, n_504);
  xor g362 (n_505, A[59], B[59]);
  xor g363 (Z[59], n_501, n_505);
  nand g364 (n_507, A[60], B[60]);
  nand g365 (n_508, A[60], n_506);
  nand g366 (n_509, B[60], n_506);
  nand g367 (n_511, n_507, n_508, n_509);
  xor g368 (n_510, A[60], B[60]);
  xor g369 (Z[60], n_506, n_510);
  nand g370 (n_512, A[61], B[61]);
  nand g371 (n_513, A[61], n_511);
  nand g372 (n_514, B[61], n_511);
  nand g373 (n_516, n_512, n_513, n_514);
  xor g374 (n_515, A[61], B[61]);
  xor g375 (Z[61], n_511, n_515);
  nand g376 (n_517, A[62], B[62]);
  nand g377 (n_518, A[62], n_516);
  nand g378 (n_519, B[62], n_516);
  nand g379 (n_521, n_517, n_518, n_519);
  xor g380 (n_520, A[62], B[62]);
  xor g381 (Z[62], n_516, n_520);
  nand g382 (n_522, A[63], B[63]);
  nand g383 (n_523, A[63], n_521);
  nand g384 (n_524, B[63], n_521);
  nand g385 (n_526, n_522, n_523, n_524);
  xor g386 (n_525, A[63], B[63]);
  xor g387 (Z[63], n_521, n_525);
  nand g388 (n_527, A[64], B[64]);
  nand g389 (n_528, A[64], n_526);
  nand g390 (n_529, B[64], n_526);
  nand g391 (n_531, n_527, n_528, n_529);
  xor g392 (n_530, A[64], B[64]);
  xor g393 (Z[64], n_526, n_530);
  nand g394 (n_532, A[65], B[65]);
  nand g395 (n_533, A[65], n_531);
  nand g396 (n_534, B[65], n_531);
  nand g397 (n_536, n_532, n_533, n_534);
  xor g398 (n_535, A[65], B[65]);
  xor g399 (Z[65], n_531, n_535);
  nand g403 (n_206, n_537, n_538, n_539);
  xor g405 (Z[66], n_536, n_540);
  or g407 (n_537, A[66], B[66]);
  xor g408 (n_540, A[66], B[66]);
  or g409 (n_213, wc, n_207);
  not gc (wc, A[1]);
  or g410 (n_214, wc0, n_207);
  not gc0 (wc0, B[1]);
  xnor g411 (Z[1], n_207, n_215);
  or g412 (n_538, A[66], wc1);
  not gc1 (wc1, n_536);
  or g413 (n_539, B[66], wc2);
  not gc2 (wc2, n_536);
endmodule

module add_signed_1220_2_GENERIC(A, B, Z);
  input [66:0] A, B;
  output [67:0] Z;
  wire [66:0] A, B;
  wire [67:0] Z;
  add_signed_1220_2_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_1220_3_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [66:0] A, B;
  output [67:0] Z;
  wire [66:0] A, B;
  wire [67:0] Z;
  wire n_206, n_207, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540;
  not g3 (Z[67], n_206);
  nand g4 (n_207, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_212, A[1], B[1]);
  nand g13 (n_216, n_212, n_213, n_214);
  xor g14 (n_215, A[1], B[1]);
  nand g16 (n_217, A[2], B[2]);
  nand g17 (n_218, A[2], n_216);
  nand g18 (n_219, B[2], n_216);
  nand g19 (n_221, n_217, n_218, n_219);
  xor g20 (n_220, A[2], B[2]);
  xor g21 (Z[2], n_216, n_220);
  nand g22 (n_222, A[3], B[3]);
  nand g23 (n_223, A[3], n_221);
  nand g24 (n_224, B[3], n_221);
  nand g25 (n_226, n_222, n_223, n_224);
  xor g26 (n_225, A[3], B[3]);
  xor g27 (Z[3], n_221, n_225);
  nand g28 (n_227, A[4], B[4]);
  nand g29 (n_228, A[4], n_226);
  nand g30 (n_229, B[4], n_226);
  nand g31 (n_231, n_227, n_228, n_229);
  xor g32 (n_230, A[4], B[4]);
  xor g33 (Z[4], n_226, n_230);
  nand g34 (n_232, A[5], B[5]);
  nand g35 (n_233, A[5], n_231);
  nand g36 (n_234, B[5], n_231);
  nand g37 (n_236, n_232, n_233, n_234);
  xor g38 (n_235, A[5], B[5]);
  xor g39 (Z[5], n_231, n_235);
  nand g40 (n_237, A[6], B[6]);
  nand g41 (n_238, A[6], n_236);
  nand g42 (n_239, B[6], n_236);
  nand g43 (n_241, n_237, n_238, n_239);
  xor g44 (n_240, A[6], B[6]);
  xor g45 (Z[6], n_236, n_240);
  nand g46 (n_242, A[7], B[7]);
  nand g47 (n_243, A[7], n_241);
  nand g48 (n_244, B[7], n_241);
  nand g49 (n_246, n_242, n_243, n_244);
  xor g50 (n_245, A[7], B[7]);
  xor g51 (Z[7], n_241, n_245);
  nand g52 (n_247, A[8], B[8]);
  nand g53 (n_248, A[8], n_246);
  nand g54 (n_249, B[8], n_246);
  nand g55 (n_251, n_247, n_248, n_249);
  xor g56 (n_250, A[8], B[8]);
  xor g57 (Z[8], n_246, n_250);
  nand g58 (n_252, A[9], B[9]);
  nand g59 (n_253, A[9], n_251);
  nand g60 (n_254, B[9], n_251);
  nand g61 (n_256, n_252, n_253, n_254);
  xor g62 (n_255, A[9], B[9]);
  xor g63 (Z[9], n_251, n_255);
  nand g64 (n_257, A[10], B[10]);
  nand g65 (n_258, A[10], n_256);
  nand g66 (n_259, B[10], n_256);
  nand g67 (n_261, n_257, n_258, n_259);
  xor g68 (n_260, A[10], B[10]);
  xor g69 (Z[10], n_256, n_260);
  nand g70 (n_262, A[11], B[11]);
  nand g71 (n_263, A[11], n_261);
  nand g72 (n_264, B[11], n_261);
  nand g73 (n_266, n_262, n_263, n_264);
  xor g74 (n_265, A[11], B[11]);
  xor g75 (Z[11], n_261, n_265);
  nand g76 (n_267, A[12], B[12]);
  nand g77 (n_268, A[12], n_266);
  nand g78 (n_269, B[12], n_266);
  nand g79 (n_271, n_267, n_268, n_269);
  xor g80 (n_270, A[12], B[12]);
  xor g81 (Z[12], n_266, n_270);
  nand g82 (n_272, A[13], B[13]);
  nand g83 (n_273, A[13], n_271);
  nand g84 (n_274, B[13], n_271);
  nand g85 (n_276, n_272, n_273, n_274);
  xor g86 (n_275, A[13], B[13]);
  xor g87 (Z[13], n_271, n_275);
  nand g88 (n_277, A[14], B[14]);
  nand g89 (n_278, A[14], n_276);
  nand g90 (n_279, B[14], n_276);
  nand g91 (n_281, n_277, n_278, n_279);
  xor g92 (n_280, A[14], B[14]);
  xor g93 (Z[14], n_276, n_280);
  nand g94 (n_282, A[15], B[15]);
  nand g95 (n_283, A[15], n_281);
  nand g96 (n_284, B[15], n_281);
  nand g97 (n_286, n_282, n_283, n_284);
  xor g98 (n_285, A[15], B[15]);
  xor g99 (Z[15], n_281, n_285);
  nand g100 (n_287, A[16], B[16]);
  nand g101 (n_288, A[16], n_286);
  nand g102 (n_289, B[16], n_286);
  nand g103 (n_291, n_287, n_288, n_289);
  xor g104 (n_290, A[16], B[16]);
  xor g105 (Z[16], n_286, n_290);
  nand g106 (n_292, A[17], B[17]);
  nand g107 (n_293, A[17], n_291);
  nand g108 (n_294, B[17], n_291);
  nand g109 (n_296, n_292, n_293, n_294);
  xor g110 (n_295, A[17], B[17]);
  xor g111 (Z[17], n_291, n_295);
  nand g112 (n_297, A[18], B[18]);
  nand g113 (n_298, A[18], n_296);
  nand g114 (n_299, B[18], n_296);
  nand g115 (n_301, n_297, n_298, n_299);
  xor g116 (n_300, A[18], B[18]);
  xor g117 (Z[18], n_296, n_300);
  nand g118 (n_302, A[19], B[19]);
  nand g119 (n_303, A[19], n_301);
  nand g120 (n_304, B[19], n_301);
  nand g121 (n_306, n_302, n_303, n_304);
  xor g122 (n_305, A[19], B[19]);
  xor g123 (Z[19], n_301, n_305);
  nand g124 (n_307, A[20], B[20]);
  nand g125 (n_308, A[20], n_306);
  nand g126 (n_309, B[20], n_306);
  nand g127 (n_311, n_307, n_308, n_309);
  xor g128 (n_310, A[20], B[20]);
  xor g129 (Z[20], n_306, n_310);
  nand g130 (n_312, A[21], B[21]);
  nand g131 (n_313, A[21], n_311);
  nand g132 (n_314, B[21], n_311);
  nand g133 (n_316, n_312, n_313, n_314);
  xor g134 (n_315, A[21], B[21]);
  xor g135 (Z[21], n_311, n_315);
  nand g136 (n_317, A[22], B[22]);
  nand g137 (n_318, A[22], n_316);
  nand g138 (n_319, B[22], n_316);
  nand g139 (n_321, n_317, n_318, n_319);
  xor g140 (n_320, A[22], B[22]);
  xor g141 (Z[22], n_316, n_320);
  nand g142 (n_322, A[23], B[23]);
  nand g143 (n_323, A[23], n_321);
  nand g144 (n_324, B[23], n_321);
  nand g145 (n_326, n_322, n_323, n_324);
  xor g146 (n_325, A[23], B[23]);
  xor g147 (Z[23], n_321, n_325);
  nand g148 (n_327, A[24], B[24]);
  nand g149 (n_328, A[24], n_326);
  nand g150 (n_329, B[24], n_326);
  nand g151 (n_331, n_327, n_328, n_329);
  xor g152 (n_330, A[24], B[24]);
  xor g153 (Z[24], n_326, n_330);
  nand g154 (n_332, A[25], B[25]);
  nand g155 (n_333, A[25], n_331);
  nand g156 (n_334, B[25], n_331);
  nand g157 (n_336, n_332, n_333, n_334);
  xor g158 (n_335, A[25], B[25]);
  xor g159 (Z[25], n_331, n_335);
  nand g160 (n_337, A[26], B[26]);
  nand g161 (n_338, A[26], n_336);
  nand g162 (n_339, B[26], n_336);
  nand g163 (n_341, n_337, n_338, n_339);
  xor g164 (n_340, A[26], B[26]);
  xor g165 (Z[26], n_336, n_340);
  nand g166 (n_342, A[27], B[27]);
  nand g167 (n_343, A[27], n_341);
  nand g168 (n_344, B[27], n_341);
  nand g169 (n_346, n_342, n_343, n_344);
  xor g170 (n_345, A[27], B[27]);
  xor g171 (Z[27], n_341, n_345);
  nand g172 (n_347, A[28], B[28]);
  nand g173 (n_348, A[28], n_346);
  nand g174 (n_349, B[28], n_346);
  nand g175 (n_351, n_347, n_348, n_349);
  xor g176 (n_350, A[28], B[28]);
  xor g177 (Z[28], n_346, n_350);
  nand g178 (n_352, A[29], B[29]);
  nand g179 (n_353, A[29], n_351);
  nand g180 (n_354, B[29], n_351);
  nand g181 (n_356, n_352, n_353, n_354);
  xor g182 (n_355, A[29], B[29]);
  xor g183 (Z[29], n_351, n_355);
  nand g184 (n_357, A[30], B[30]);
  nand g185 (n_358, A[30], n_356);
  nand g186 (n_359, B[30], n_356);
  nand g187 (n_361, n_357, n_358, n_359);
  xor g188 (n_360, A[30], B[30]);
  xor g189 (Z[30], n_356, n_360);
  nand g190 (n_362, A[31], B[31]);
  nand g191 (n_363, A[31], n_361);
  nand g192 (n_364, B[31], n_361);
  nand g193 (n_366, n_362, n_363, n_364);
  xor g194 (n_365, A[31], B[31]);
  xor g195 (Z[31], n_361, n_365);
  nand g196 (n_367, A[32], B[32]);
  nand g197 (n_368, A[32], n_366);
  nand g198 (n_369, B[32], n_366);
  nand g199 (n_371, n_367, n_368, n_369);
  xor g200 (n_370, A[32], B[32]);
  xor g201 (Z[32], n_366, n_370);
  nand g202 (n_372, A[33], B[33]);
  nand g203 (n_373, A[33], n_371);
  nand g204 (n_374, B[33], n_371);
  nand g205 (n_376, n_372, n_373, n_374);
  xor g206 (n_375, A[33], B[33]);
  xor g207 (Z[33], n_371, n_375);
  nand g208 (n_377, A[34], B[34]);
  nand g209 (n_378, A[34], n_376);
  nand g210 (n_379, B[34], n_376);
  nand g211 (n_381, n_377, n_378, n_379);
  xor g212 (n_380, A[34], B[34]);
  xor g213 (Z[34], n_376, n_380);
  nand g214 (n_382, A[35], B[35]);
  nand g215 (n_383, A[35], n_381);
  nand g216 (n_384, B[35], n_381);
  nand g217 (n_386, n_382, n_383, n_384);
  xor g218 (n_385, A[35], B[35]);
  xor g219 (Z[35], n_381, n_385);
  nand g220 (n_387, A[36], B[36]);
  nand g221 (n_388, A[36], n_386);
  nand g222 (n_389, B[36], n_386);
  nand g223 (n_391, n_387, n_388, n_389);
  xor g224 (n_390, A[36], B[36]);
  xor g225 (Z[36], n_386, n_390);
  nand g226 (n_392, A[37], B[37]);
  nand g227 (n_393, A[37], n_391);
  nand g228 (n_394, B[37], n_391);
  nand g229 (n_396, n_392, n_393, n_394);
  xor g230 (n_395, A[37], B[37]);
  xor g231 (Z[37], n_391, n_395);
  nand g232 (n_397, A[38], B[38]);
  nand g233 (n_398, A[38], n_396);
  nand g234 (n_399, B[38], n_396);
  nand g235 (n_401, n_397, n_398, n_399);
  xor g236 (n_400, A[38], B[38]);
  xor g237 (Z[38], n_396, n_400);
  nand g238 (n_402, A[39], B[39]);
  nand g239 (n_403, A[39], n_401);
  nand g240 (n_404, B[39], n_401);
  nand g241 (n_406, n_402, n_403, n_404);
  xor g242 (n_405, A[39], B[39]);
  xor g243 (Z[39], n_401, n_405);
  nand g244 (n_407, A[40], B[40]);
  nand g245 (n_408, A[40], n_406);
  nand g246 (n_409, B[40], n_406);
  nand g247 (n_411, n_407, n_408, n_409);
  xor g248 (n_410, A[40], B[40]);
  xor g249 (Z[40], n_406, n_410);
  nand g250 (n_412, A[41], B[41]);
  nand g251 (n_413, A[41], n_411);
  nand g252 (n_414, B[41], n_411);
  nand g253 (n_416, n_412, n_413, n_414);
  xor g254 (n_415, A[41], B[41]);
  xor g255 (Z[41], n_411, n_415);
  nand g256 (n_417, A[42], B[42]);
  nand g257 (n_418, A[42], n_416);
  nand g258 (n_419, B[42], n_416);
  nand g259 (n_421, n_417, n_418, n_419);
  xor g260 (n_420, A[42], B[42]);
  xor g261 (Z[42], n_416, n_420);
  nand g262 (n_422, A[43], B[43]);
  nand g263 (n_423, A[43], n_421);
  nand g264 (n_424, B[43], n_421);
  nand g265 (n_426, n_422, n_423, n_424);
  xor g266 (n_425, A[43], B[43]);
  xor g267 (Z[43], n_421, n_425);
  nand g268 (n_427, A[44], B[44]);
  nand g269 (n_428, A[44], n_426);
  nand g270 (n_429, B[44], n_426);
  nand g271 (n_431, n_427, n_428, n_429);
  xor g272 (n_430, A[44], B[44]);
  xor g273 (Z[44], n_426, n_430);
  nand g274 (n_432, A[45], B[45]);
  nand g275 (n_433, A[45], n_431);
  nand g276 (n_434, B[45], n_431);
  nand g277 (n_436, n_432, n_433, n_434);
  xor g278 (n_435, A[45], B[45]);
  xor g279 (Z[45], n_431, n_435);
  nand g280 (n_437, A[46], B[46]);
  nand g281 (n_438, A[46], n_436);
  nand g282 (n_439, B[46], n_436);
  nand g283 (n_441, n_437, n_438, n_439);
  xor g284 (n_440, A[46], B[46]);
  xor g285 (Z[46], n_436, n_440);
  nand g286 (n_442, A[47], B[47]);
  nand g287 (n_443, A[47], n_441);
  nand g288 (n_444, B[47], n_441);
  nand g289 (n_446, n_442, n_443, n_444);
  xor g290 (n_445, A[47], B[47]);
  xor g291 (Z[47], n_441, n_445);
  nand g292 (n_447, A[48], B[48]);
  nand g293 (n_448, A[48], n_446);
  nand g294 (n_449, B[48], n_446);
  nand g295 (n_451, n_447, n_448, n_449);
  xor g296 (n_450, A[48], B[48]);
  xor g297 (Z[48], n_446, n_450);
  nand g298 (n_452, A[49], B[49]);
  nand g299 (n_453, A[49], n_451);
  nand g300 (n_454, B[49], n_451);
  nand g301 (n_456, n_452, n_453, n_454);
  xor g302 (n_455, A[49], B[49]);
  xor g303 (Z[49], n_451, n_455);
  nand g304 (n_457, A[50], B[50]);
  nand g305 (n_458, A[50], n_456);
  nand g306 (n_459, B[50], n_456);
  nand g307 (n_461, n_457, n_458, n_459);
  xor g308 (n_460, A[50], B[50]);
  xor g309 (Z[50], n_456, n_460);
  nand g310 (n_462, A[51], B[51]);
  nand g311 (n_463, A[51], n_461);
  nand g312 (n_464, B[51], n_461);
  nand g313 (n_466, n_462, n_463, n_464);
  xor g314 (n_465, A[51], B[51]);
  xor g315 (Z[51], n_461, n_465);
  nand g316 (n_467, A[52], B[52]);
  nand g317 (n_468, A[52], n_466);
  nand g318 (n_469, B[52], n_466);
  nand g319 (n_471, n_467, n_468, n_469);
  xor g320 (n_470, A[52], B[52]);
  xor g321 (Z[52], n_466, n_470);
  nand g322 (n_472, A[53], B[53]);
  nand g323 (n_473, A[53], n_471);
  nand g324 (n_474, B[53], n_471);
  nand g325 (n_476, n_472, n_473, n_474);
  xor g326 (n_475, A[53], B[53]);
  xor g327 (Z[53], n_471, n_475);
  nand g328 (n_477, A[54], B[54]);
  nand g329 (n_478, A[54], n_476);
  nand g330 (n_479, B[54], n_476);
  nand g331 (n_481, n_477, n_478, n_479);
  xor g332 (n_480, A[54], B[54]);
  xor g333 (Z[54], n_476, n_480);
  nand g334 (n_482, A[55], B[55]);
  nand g335 (n_483, A[55], n_481);
  nand g336 (n_484, B[55], n_481);
  nand g337 (n_486, n_482, n_483, n_484);
  xor g338 (n_485, A[55], B[55]);
  xor g339 (Z[55], n_481, n_485);
  nand g340 (n_487, A[56], B[56]);
  nand g341 (n_488, A[56], n_486);
  nand g342 (n_489, B[56], n_486);
  nand g343 (n_491, n_487, n_488, n_489);
  xor g344 (n_490, A[56], B[56]);
  xor g345 (Z[56], n_486, n_490);
  nand g346 (n_492, A[57], B[57]);
  nand g347 (n_493, A[57], n_491);
  nand g348 (n_494, B[57], n_491);
  nand g349 (n_496, n_492, n_493, n_494);
  xor g350 (n_495, A[57], B[57]);
  xor g351 (Z[57], n_491, n_495);
  nand g352 (n_497, A[58], B[58]);
  nand g353 (n_498, A[58], n_496);
  nand g354 (n_499, B[58], n_496);
  nand g355 (n_501, n_497, n_498, n_499);
  xor g356 (n_500, A[58], B[58]);
  xor g357 (Z[58], n_496, n_500);
  nand g358 (n_502, A[59], B[59]);
  nand g359 (n_503, A[59], n_501);
  nand g360 (n_504, B[59], n_501);
  nand g361 (n_506, n_502, n_503, n_504);
  xor g362 (n_505, A[59], B[59]);
  xor g363 (Z[59], n_501, n_505);
  nand g364 (n_507, A[60], B[60]);
  nand g365 (n_508, A[60], n_506);
  nand g366 (n_509, B[60], n_506);
  nand g367 (n_511, n_507, n_508, n_509);
  xor g368 (n_510, A[60], B[60]);
  xor g369 (Z[60], n_506, n_510);
  nand g370 (n_512, A[61], B[61]);
  nand g371 (n_513, A[61], n_511);
  nand g372 (n_514, B[61], n_511);
  nand g373 (n_516, n_512, n_513, n_514);
  xor g374 (n_515, A[61], B[61]);
  xor g375 (Z[61], n_511, n_515);
  nand g376 (n_517, A[62], B[62]);
  nand g377 (n_518, A[62], n_516);
  nand g378 (n_519, B[62], n_516);
  nand g379 (n_521, n_517, n_518, n_519);
  xor g380 (n_520, A[62], B[62]);
  xor g381 (Z[62], n_516, n_520);
  nand g382 (n_522, A[63], B[63]);
  nand g383 (n_523, A[63], n_521);
  nand g384 (n_524, B[63], n_521);
  nand g385 (n_526, n_522, n_523, n_524);
  xor g386 (n_525, A[63], B[63]);
  xor g387 (Z[63], n_521, n_525);
  nand g388 (n_527, A[64], B[64]);
  nand g389 (n_528, A[64], n_526);
  nand g390 (n_529, B[64], n_526);
  nand g391 (n_531, n_527, n_528, n_529);
  xor g392 (n_530, A[64], B[64]);
  xor g393 (Z[64], n_526, n_530);
  nand g394 (n_532, A[65], B[65]);
  nand g395 (n_533, A[65], n_531);
  nand g396 (n_534, B[65], n_531);
  nand g397 (n_536, n_532, n_533, n_534);
  xor g398 (n_535, A[65], B[65]);
  xor g399 (Z[65], n_531, n_535);
  nand g403 (n_206, n_537, n_538, n_539);
  xor g405 (Z[66], n_536, n_540);
  or g407 (n_537, A[66], B[66]);
  xor g408 (n_540, A[66], B[66]);
  or g409 (n_213, wc, n_207);
  not gc (wc, A[1]);
  or g410 (n_214, wc0, n_207);
  not gc0 (wc0, B[1]);
  xnor g411 (Z[1], n_207, n_215);
  or g412 (n_538, A[66], wc1);
  not gc1 (wc1, n_536);
  or g413 (n_539, B[66], wc2);
  not gc2 (wc2, n_536);
endmodule

module add_signed_1220_3_GENERIC(A, B, Z);
  input [66:0] A, B;
  output [67:0] Z;
  wire [66:0] A, B;
  wire [67:0] Z;
  add_signed_1220_3_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_192_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [18:0] A, B;
  output [19:0] Z;
  wire [18:0] A, B;
  wire [19:0] Z;
  wire n_62, n_63, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156;
  not g3 (Z[19], n_62);
  nand g4 (n_63, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_68, A[1], B[1]);
  nand g13 (n_72, n_68, n_69, n_70);
  xor g14 (n_71, A[1], B[1]);
  nand g16 (n_73, A[2], B[2]);
  nand g17 (n_74, A[2], n_72);
  nand g18 (n_75, B[2], n_72);
  nand g19 (n_77, n_73, n_74, n_75);
  xor g20 (n_76, A[2], B[2]);
  xor g21 (Z[2], n_72, n_76);
  nand g22 (n_78, A[3], B[3]);
  nand g23 (n_79, A[3], n_77);
  nand g24 (n_80, B[3], n_77);
  nand g25 (n_82, n_78, n_79, n_80);
  xor g26 (n_81, A[3], B[3]);
  xor g27 (Z[3], n_77, n_81);
  nand g28 (n_83, A[4], B[4]);
  nand g29 (n_84, A[4], n_82);
  nand g30 (n_85, B[4], n_82);
  nand g31 (n_87, n_83, n_84, n_85);
  xor g32 (n_86, A[4], B[4]);
  xor g33 (Z[4], n_82, n_86);
  nand g34 (n_88, A[5], B[5]);
  nand g35 (n_89, A[5], n_87);
  nand g36 (n_90, B[5], n_87);
  nand g37 (n_92, n_88, n_89, n_90);
  xor g38 (n_91, A[5], B[5]);
  xor g39 (Z[5], n_87, n_91);
  nand g40 (n_93, A[6], B[6]);
  nand g41 (n_94, A[6], n_92);
  nand g42 (n_95, B[6], n_92);
  nand g43 (n_97, n_93, n_94, n_95);
  xor g44 (n_96, A[6], B[6]);
  xor g45 (Z[6], n_92, n_96);
  nand g46 (n_98, A[7], B[7]);
  nand g47 (n_99, A[7], n_97);
  nand g48 (n_100, B[7], n_97);
  nand g49 (n_102, n_98, n_99, n_100);
  xor g50 (n_101, A[7], B[7]);
  xor g51 (Z[7], n_97, n_101);
  nand g52 (n_103, A[8], B[8]);
  nand g53 (n_104, A[8], n_102);
  nand g54 (n_105, B[8], n_102);
  nand g55 (n_107, n_103, n_104, n_105);
  xor g56 (n_106, A[8], B[8]);
  xor g57 (Z[8], n_102, n_106);
  nand g58 (n_108, A[9], B[9]);
  nand g59 (n_109, A[9], n_107);
  nand g60 (n_110, B[9], n_107);
  nand g61 (n_112, n_108, n_109, n_110);
  xor g62 (n_111, A[9], B[9]);
  xor g63 (Z[9], n_107, n_111);
  nand g64 (n_113, A[10], B[10]);
  nand g65 (n_114, A[10], n_112);
  nand g66 (n_115, B[10], n_112);
  nand g67 (n_117, n_113, n_114, n_115);
  xor g68 (n_116, A[10], B[10]);
  xor g69 (Z[10], n_112, n_116);
  nand g70 (n_118, A[11], B[11]);
  nand g71 (n_119, A[11], n_117);
  nand g72 (n_120, B[11], n_117);
  nand g73 (n_122, n_118, n_119, n_120);
  xor g74 (n_121, A[11], B[11]);
  xor g75 (Z[11], n_117, n_121);
  nand g76 (n_123, A[12], B[12]);
  nand g77 (n_124, A[12], n_122);
  nand g78 (n_125, B[12], n_122);
  nand g79 (n_127, n_123, n_124, n_125);
  xor g80 (n_126, A[12], B[12]);
  xor g81 (Z[12], n_122, n_126);
  nand g82 (n_128, A[13], B[13]);
  nand g83 (n_129, A[13], n_127);
  nand g84 (n_130, B[13], n_127);
  nand g85 (n_132, n_128, n_129, n_130);
  xor g86 (n_131, A[13], B[13]);
  xor g87 (Z[13], n_127, n_131);
  nand g88 (n_133, A[14], B[14]);
  nand g89 (n_134, A[14], n_132);
  nand g90 (n_135, B[14], n_132);
  nand g91 (n_137, n_133, n_134, n_135);
  xor g92 (n_136, A[14], B[14]);
  xor g93 (Z[14], n_132, n_136);
  nand g94 (n_138, A[15], B[15]);
  nand g95 (n_139, A[15], n_137);
  nand g96 (n_140, B[15], n_137);
  nand g97 (n_142, n_138, n_139, n_140);
  xor g98 (n_141, A[15], B[15]);
  xor g99 (Z[15], n_137, n_141);
  nand g100 (n_143, A[16], B[16]);
  nand g101 (n_144, A[16], n_142);
  nand g102 (n_145, B[16], n_142);
  nand g103 (n_147, n_143, n_144, n_145);
  xor g104 (n_146, A[16], B[16]);
  xor g105 (Z[16], n_142, n_146);
  nand g106 (n_148, A[17], B[17]);
  nand g107 (n_149, A[17], n_147);
  nand g108 (n_150, B[17], n_147);
  nand g109 (n_152, n_148, n_149, n_150);
  xor g110 (n_151, A[17], B[17]);
  xor g111 (Z[17], n_147, n_151);
  nand g115 (n_62, n_153, n_154, n_155);
  xor g117 (Z[18], n_152, n_156);
  or g119 (n_153, A[18], B[18]);
  xor g120 (n_156, A[18], B[18]);
  or g121 (n_69, wc, n_63);
  not gc (wc, A[1]);
  or g122 (n_70, wc0, n_63);
  not gc0 (wc0, B[1]);
  xnor g123 (Z[1], n_63, n_71);
  or g124 (n_154, A[18], wc1);
  not gc1 (wc1, n_152);
  or g125 (n_155, B[18], wc2);
  not gc2 (wc2, n_152);
endmodule

module add_signed_192_GENERIC(A, B, Z);
  input [18:0] A, B;
  output [19:0] Z;
  wire [18:0] A, B;
  wire [19:0] Z;
  add_signed_192_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_192_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [18:0] A, B;
  output [19:0] Z;
  wire [18:0] A, B;
  wire [19:0] Z;
  wire n_62, n_63, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156;
  not g3 (Z[19], n_62);
  nand g4 (n_63, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_68, A[1], B[1]);
  nand g13 (n_72, n_68, n_69, n_70);
  xor g14 (n_71, A[1], B[1]);
  nand g16 (n_73, A[2], B[2]);
  nand g17 (n_74, A[2], n_72);
  nand g18 (n_75, B[2], n_72);
  nand g19 (n_77, n_73, n_74, n_75);
  xor g20 (n_76, A[2], B[2]);
  xor g21 (Z[2], n_72, n_76);
  nand g22 (n_78, A[3], B[3]);
  nand g23 (n_79, A[3], n_77);
  nand g24 (n_80, B[3], n_77);
  nand g25 (n_82, n_78, n_79, n_80);
  xor g26 (n_81, A[3], B[3]);
  xor g27 (Z[3], n_77, n_81);
  nand g28 (n_83, A[4], B[4]);
  nand g29 (n_84, A[4], n_82);
  nand g30 (n_85, B[4], n_82);
  nand g31 (n_87, n_83, n_84, n_85);
  xor g32 (n_86, A[4], B[4]);
  xor g33 (Z[4], n_82, n_86);
  nand g34 (n_88, A[5], B[5]);
  nand g35 (n_89, A[5], n_87);
  nand g36 (n_90, B[5], n_87);
  nand g37 (n_92, n_88, n_89, n_90);
  xor g38 (n_91, A[5], B[5]);
  xor g39 (Z[5], n_87, n_91);
  nand g40 (n_93, A[6], B[6]);
  nand g41 (n_94, A[6], n_92);
  nand g42 (n_95, B[6], n_92);
  nand g43 (n_97, n_93, n_94, n_95);
  xor g44 (n_96, A[6], B[6]);
  xor g45 (Z[6], n_92, n_96);
  nand g46 (n_98, A[7], B[7]);
  nand g47 (n_99, A[7], n_97);
  nand g48 (n_100, B[7], n_97);
  nand g49 (n_102, n_98, n_99, n_100);
  xor g50 (n_101, A[7], B[7]);
  xor g51 (Z[7], n_97, n_101);
  nand g52 (n_103, A[8], B[8]);
  nand g53 (n_104, A[8], n_102);
  nand g54 (n_105, B[8], n_102);
  nand g55 (n_107, n_103, n_104, n_105);
  xor g56 (n_106, A[8], B[8]);
  xor g57 (Z[8], n_102, n_106);
  nand g58 (n_108, A[9], B[9]);
  nand g59 (n_109, A[9], n_107);
  nand g60 (n_110, B[9], n_107);
  nand g61 (n_112, n_108, n_109, n_110);
  xor g62 (n_111, A[9], B[9]);
  xor g63 (Z[9], n_107, n_111);
  nand g64 (n_113, A[10], B[10]);
  nand g65 (n_114, A[10], n_112);
  nand g66 (n_115, B[10], n_112);
  nand g67 (n_117, n_113, n_114, n_115);
  xor g68 (n_116, A[10], B[10]);
  xor g69 (Z[10], n_112, n_116);
  nand g70 (n_118, A[11], B[11]);
  nand g71 (n_119, A[11], n_117);
  nand g72 (n_120, B[11], n_117);
  nand g73 (n_122, n_118, n_119, n_120);
  xor g74 (n_121, A[11], B[11]);
  xor g75 (Z[11], n_117, n_121);
  nand g76 (n_123, A[12], B[12]);
  nand g77 (n_124, A[12], n_122);
  nand g78 (n_125, B[12], n_122);
  nand g79 (n_127, n_123, n_124, n_125);
  xor g80 (n_126, A[12], B[12]);
  xor g81 (Z[12], n_122, n_126);
  nand g82 (n_128, A[13], B[13]);
  nand g83 (n_129, A[13], n_127);
  nand g84 (n_130, B[13], n_127);
  nand g85 (n_132, n_128, n_129, n_130);
  xor g86 (n_131, A[13], B[13]);
  xor g87 (Z[13], n_127, n_131);
  nand g88 (n_133, A[14], B[14]);
  nand g89 (n_134, A[14], n_132);
  nand g90 (n_135, B[14], n_132);
  nand g91 (n_137, n_133, n_134, n_135);
  xor g92 (n_136, A[14], B[14]);
  xor g93 (Z[14], n_132, n_136);
  nand g94 (n_138, A[15], B[15]);
  nand g95 (n_139, A[15], n_137);
  nand g96 (n_140, B[15], n_137);
  nand g97 (n_142, n_138, n_139, n_140);
  xor g98 (n_141, A[15], B[15]);
  xor g99 (Z[15], n_137, n_141);
  nand g100 (n_143, A[16], B[16]);
  nand g101 (n_144, A[16], n_142);
  nand g102 (n_145, B[16], n_142);
  nand g103 (n_147, n_143, n_144, n_145);
  xor g104 (n_146, A[16], B[16]);
  xor g105 (Z[16], n_142, n_146);
  nand g106 (n_148, A[17], B[17]);
  nand g107 (n_149, A[17], n_147);
  nand g108 (n_150, B[17], n_147);
  nand g109 (n_152, n_148, n_149, n_150);
  xor g110 (n_151, A[17], B[17]);
  xor g111 (Z[17], n_147, n_151);
  nand g115 (n_62, n_153, n_154, n_155);
  xor g117 (Z[18], n_152, n_156);
  or g119 (n_153, A[18], B[18]);
  xor g120 (n_156, A[18], B[18]);
  or g121 (n_69, wc, n_63);
  not gc (wc, A[1]);
  or g122 (n_70, wc0, n_63);
  not gc0 (wc0, B[1]);
  xnor g123 (Z[1], n_63, n_71);
  or g124 (n_154, A[18], wc1);
  not gc1 (wc1, n_152);
  or g125 (n_155, B[18], wc2);
  not gc2 (wc2, n_152);
endmodule

module add_signed_192_2_GENERIC(A, B, Z);
  input [18:0] A, B;
  output [19:0] Z;
  wire [18:0] A, B;
  wire [19:0] Z;
  add_signed_192_2_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_2443_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [65:0] A, B;
  output [66:0] Z;
  wire [65:0] A, B;
  wire [66:0] Z;
  wire n_203, n_204, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502;
  wire n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510;
  wire n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518;
  wire n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526;
  wire n_527, n_528, n_529, n_530, n_531, n_532;
  not g3 (Z[66], n_203);
  nand g4 (n_204, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_209, A[1], B[1]);
  nand g13 (n_213, n_209, n_210, n_211);
  xor g14 (n_212, A[1], B[1]);
  nand g16 (n_214, A[2], B[2]);
  nand g17 (n_215, A[2], n_213);
  nand g18 (n_216, B[2], n_213);
  nand g19 (n_218, n_214, n_215, n_216);
  xor g20 (n_217, A[2], B[2]);
  xor g21 (Z[2], n_213, n_217);
  nand g22 (n_219, A[3], B[3]);
  nand g23 (n_220, A[3], n_218);
  nand g24 (n_221, B[3], n_218);
  nand g25 (n_223, n_219, n_220, n_221);
  xor g26 (n_222, A[3], B[3]);
  xor g27 (Z[3], n_218, n_222);
  nand g28 (n_224, A[4], B[4]);
  nand g29 (n_225, A[4], n_223);
  nand g30 (n_226, B[4], n_223);
  nand g31 (n_228, n_224, n_225, n_226);
  xor g32 (n_227, A[4], B[4]);
  xor g33 (Z[4], n_223, n_227);
  nand g34 (n_229, A[5], B[5]);
  nand g35 (n_230, A[5], n_228);
  nand g36 (n_231, B[5], n_228);
  nand g37 (n_233, n_229, n_230, n_231);
  xor g38 (n_232, A[5], B[5]);
  xor g39 (Z[5], n_228, n_232);
  nand g40 (n_234, A[6], B[6]);
  nand g41 (n_235, A[6], n_233);
  nand g42 (n_236, B[6], n_233);
  nand g43 (n_238, n_234, n_235, n_236);
  xor g44 (n_237, A[6], B[6]);
  xor g45 (Z[6], n_233, n_237);
  nand g46 (n_239, A[7], B[7]);
  nand g47 (n_240, A[7], n_238);
  nand g48 (n_241, B[7], n_238);
  nand g49 (n_243, n_239, n_240, n_241);
  xor g50 (n_242, A[7], B[7]);
  xor g51 (Z[7], n_238, n_242);
  nand g52 (n_244, A[8], B[8]);
  nand g53 (n_245, A[8], n_243);
  nand g54 (n_246, B[8], n_243);
  nand g55 (n_248, n_244, n_245, n_246);
  xor g56 (n_247, A[8], B[8]);
  xor g57 (Z[8], n_243, n_247);
  nand g58 (n_249, A[9], B[9]);
  nand g59 (n_250, A[9], n_248);
  nand g60 (n_251, B[9], n_248);
  nand g61 (n_253, n_249, n_250, n_251);
  xor g62 (n_252, A[9], B[9]);
  xor g63 (Z[9], n_248, n_252);
  nand g64 (n_254, A[10], B[10]);
  nand g65 (n_255, A[10], n_253);
  nand g66 (n_256, B[10], n_253);
  nand g67 (n_258, n_254, n_255, n_256);
  xor g68 (n_257, A[10], B[10]);
  xor g69 (Z[10], n_253, n_257);
  nand g70 (n_259, A[11], B[11]);
  nand g71 (n_260, A[11], n_258);
  nand g72 (n_261, B[11], n_258);
  nand g73 (n_263, n_259, n_260, n_261);
  xor g74 (n_262, A[11], B[11]);
  xor g75 (Z[11], n_258, n_262);
  nand g76 (n_264, A[12], B[12]);
  nand g77 (n_265, A[12], n_263);
  nand g78 (n_266, B[12], n_263);
  nand g79 (n_268, n_264, n_265, n_266);
  xor g80 (n_267, A[12], B[12]);
  xor g81 (Z[12], n_263, n_267);
  nand g82 (n_269, A[13], B[13]);
  nand g83 (n_270, A[13], n_268);
  nand g84 (n_271, B[13], n_268);
  nand g85 (n_273, n_269, n_270, n_271);
  xor g86 (n_272, A[13], B[13]);
  xor g87 (Z[13], n_268, n_272);
  nand g88 (n_274, A[14], B[14]);
  nand g89 (n_275, A[14], n_273);
  nand g90 (n_276, B[14], n_273);
  nand g91 (n_278, n_274, n_275, n_276);
  xor g92 (n_277, A[14], B[14]);
  xor g93 (Z[14], n_273, n_277);
  nand g94 (n_279, A[15], B[15]);
  nand g95 (n_280, A[15], n_278);
  nand g96 (n_281, B[15], n_278);
  nand g97 (n_283, n_279, n_280, n_281);
  xor g98 (n_282, A[15], B[15]);
  xor g99 (Z[15], n_278, n_282);
  nand g100 (n_284, A[16], B[16]);
  nand g101 (n_285, A[16], n_283);
  nand g102 (n_286, B[16], n_283);
  nand g103 (n_288, n_284, n_285, n_286);
  xor g104 (n_287, A[16], B[16]);
  xor g105 (Z[16], n_283, n_287);
  nand g106 (n_289, A[17], B[17]);
  nand g107 (n_290, A[17], n_288);
  nand g108 (n_291, B[17], n_288);
  nand g109 (n_293, n_289, n_290, n_291);
  xor g110 (n_292, A[17], B[17]);
  xor g111 (Z[17], n_288, n_292);
  nand g112 (n_294, A[18], B[18]);
  nand g113 (n_295, A[18], n_293);
  nand g114 (n_296, B[18], n_293);
  nand g115 (n_298, n_294, n_295, n_296);
  xor g116 (n_297, A[18], B[18]);
  xor g117 (Z[18], n_293, n_297);
  nand g118 (n_299, A[19], B[19]);
  nand g119 (n_300, A[19], n_298);
  nand g120 (n_301, B[19], n_298);
  nand g121 (n_303, n_299, n_300, n_301);
  xor g122 (n_302, A[19], B[19]);
  xor g123 (Z[19], n_298, n_302);
  nand g124 (n_304, A[20], B[20]);
  nand g125 (n_305, A[20], n_303);
  nand g126 (n_306, B[20], n_303);
  nand g127 (n_308, n_304, n_305, n_306);
  xor g128 (n_307, A[20], B[20]);
  xor g129 (Z[20], n_303, n_307);
  nand g130 (n_309, A[21], B[21]);
  nand g131 (n_310, A[21], n_308);
  nand g132 (n_311, B[21], n_308);
  nand g133 (n_313, n_309, n_310, n_311);
  xor g134 (n_312, A[21], B[21]);
  xor g135 (Z[21], n_308, n_312);
  nand g136 (n_314, A[22], B[22]);
  nand g137 (n_315, A[22], n_313);
  nand g138 (n_316, B[22], n_313);
  nand g139 (n_318, n_314, n_315, n_316);
  xor g140 (n_317, A[22], B[22]);
  xor g141 (Z[22], n_313, n_317);
  nand g142 (n_319, A[23], B[23]);
  nand g143 (n_320, A[23], n_318);
  nand g144 (n_321, B[23], n_318);
  nand g145 (n_323, n_319, n_320, n_321);
  xor g146 (n_322, A[23], B[23]);
  xor g147 (Z[23], n_318, n_322);
  nand g148 (n_324, A[24], B[24]);
  nand g149 (n_325, A[24], n_323);
  nand g150 (n_326, B[24], n_323);
  nand g151 (n_328, n_324, n_325, n_326);
  xor g152 (n_327, A[24], B[24]);
  xor g153 (Z[24], n_323, n_327);
  nand g154 (n_329, A[25], B[25]);
  nand g155 (n_330, A[25], n_328);
  nand g156 (n_331, B[25], n_328);
  nand g157 (n_333, n_329, n_330, n_331);
  xor g158 (n_332, A[25], B[25]);
  xor g159 (Z[25], n_328, n_332);
  nand g160 (n_334, A[26], B[26]);
  nand g161 (n_335, A[26], n_333);
  nand g162 (n_336, B[26], n_333);
  nand g163 (n_338, n_334, n_335, n_336);
  xor g164 (n_337, A[26], B[26]);
  xor g165 (Z[26], n_333, n_337);
  nand g166 (n_339, A[27], B[27]);
  nand g167 (n_340, A[27], n_338);
  nand g168 (n_341, B[27], n_338);
  nand g169 (n_343, n_339, n_340, n_341);
  xor g170 (n_342, A[27], B[27]);
  xor g171 (Z[27], n_338, n_342);
  nand g172 (n_344, A[28], B[28]);
  nand g173 (n_345, A[28], n_343);
  nand g174 (n_346, B[28], n_343);
  nand g175 (n_348, n_344, n_345, n_346);
  xor g176 (n_347, A[28], B[28]);
  xor g177 (Z[28], n_343, n_347);
  nand g178 (n_349, A[29], B[29]);
  nand g179 (n_350, A[29], n_348);
  nand g180 (n_351, B[29], n_348);
  nand g181 (n_353, n_349, n_350, n_351);
  xor g182 (n_352, A[29], B[29]);
  xor g183 (Z[29], n_348, n_352);
  nand g184 (n_354, A[30], B[30]);
  nand g185 (n_355, A[30], n_353);
  nand g186 (n_356, B[30], n_353);
  nand g187 (n_358, n_354, n_355, n_356);
  xor g188 (n_357, A[30], B[30]);
  xor g189 (Z[30], n_353, n_357);
  nand g190 (n_359, A[31], B[31]);
  nand g191 (n_360, A[31], n_358);
  nand g192 (n_361, B[31], n_358);
  nand g193 (n_363, n_359, n_360, n_361);
  xor g194 (n_362, A[31], B[31]);
  xor g195 (Z[31], n_358, n_362);
  nand g196 (n_364, A[32], B[32]);
  nand g197 (n_365, A[32], n_363);
  nand g198 (n_366, B[32], n_363);
  nand g199 (n_368, n_364, n_365, n_366);
  xor g200 (n_367, A[32], B[32]);
  xor g201 (Z[32], n_363, n_367);
  nand g202 (n_369, A[33], B[33]);
  nand g203 (n_370, A[33], n_368);
  nand g204 (n_371, B[33], n_368);
  nand g205 (n_373, n_369, n_370, n_371);
  xor g206 (n_372, A[33], B[33]);
  xor g207 (Z[33], n_368, n_372);
  nand g208 (n_374, A[34], B[34]);
  nand g209 (n_375, A[34], n_373);
  nand g210 (n_376, B[34], n_373);
  nand g211 (n_378, n_374, n_375, n_376);
  xor g212 (n_377, A[34], B[34]);
  xor g213 (Z[34], n_373, n_377);
  nand g214 (n_379, A[35], B[35]);
  nand g215 (n_380, A[35], n_378);
  nand g216 (n_381, B[35], n_378);
  nand g217 (n_383, n_379, n_380, n_381);
  xor g218 (n_382, A[35], B[35]);
  xor g219 (Z[35], n_378, n_382);
  nand g220 (n_384, A[36], B[36]);
  nand g221 (n_385, A[36], n_383);
  nand g222 (n_386, B[36], n_383);
  nand g223 (n_388, n_384, n_385, n_386);
  xor g224 (n_387, A[36], B[36]);
  xor g225 (Z[36], n_383, n_387);
  nand g226 (n_389, A[37], B[37]);
  nand g227 (n_390, A[37], n_388);
  nand g228 (n_391, B[37], n_388);
  nand g229 (n_393, n_389, n_390, n_391);
  xor g230 (n_392, A[37], B[37]);
  xor g231 (Z[37], n_388, n_392);
  nand g232 (n_394, A[38], B[38]);
  nand g233 (n_395, A[38], n_393);
  nand g234 (n_396, B[38], n_393);
  nand g235 (n_398, n_394, n_395, n_396);
  xor g236 (n_397, A[38], B[38]);
  xor g237 (Z[38], n_393, n_397);
  nand g238 (n_399, A[39], B[39]);
  nand g239 (n_400, A[39], n_398);
  nand g240 (n_401, B[39], n_398);
  nand g241 (n_403, n_399, n_400, n_401);
  xor g242 (n_402, A[39], B[39]);
  xor g243 (Z[39], n_398, n_402);
  nand g244 (n_404, A[40], B[40]);
  nand g245 (n_405, A[40], n_403);
  nand g246 (n_406, B[40], n_403);
  nand g247 (n_408, n_404, n_405, n_406);
  xor g248 (n_407, A[40], B[40]);
  xor g249 (Z[40], n_403, n_407);
  nand g250 (n_409, A[41], B[41]);
  nand g251 (n_410, A[41], n_408);
  nand g252 (n_411, B[41], n_408);
  nand g253 (n_413, n_409, n_410, n_411);
  xor g254 (n_412, A[41], B[41]);
  xor g255 (Z[41], n_408, n_412);
  nand g256 (n_414, A[42], B[42]);
  nand g257 (n_415, A[42], n_413);
  nand g258 (n_416, B[42], n_413);
  nand g259 (n_418, n_414, n_415, n_416);
  xor g260 (n_417, A[42], B[42]);
  xor g261 (Z[42], n_413, n_417);
  nand g262 (n_419, A[43], B[43]);
  nand g263 (n_420, A[43], n_418);
  nand g264 (n_421, B[43], n_418);
  nand g265 (n_423, n_419, n_420, n_421);
  xor g266 (n_422, A[43], B[43]);
  xor g267 (Z[43], n_418, n_422);
  nand g268 (n_424, A[44], B[44]);
  nand g269 (n_425, A[44], n_423);
  nand g270 (n_426, B[44], n_423);
  nand g271 (n_428, n_424, n_425, n_426);
  xor g272 (n_427, A[44], B[44]);
  xor g273 (Z[44], n_423, n_427);
  nand g274 (n_429, A[45], B[45]);
  nand g275 (n_430, A[45], n_428);
  nand g276 (n_431, B[45], n_428);
  nand g277 (n_433, n_429, n_430, n_431);
  xor g278 (n_432, A[45], B[45]);
  xor g279 (Z[45], n_428, n_432);
  nand g280 (n_434, A[46], B[46]);
  nand g281 (n_435, A[46], n_433);
  nand g282 (n_436, B[46], n_433);
  nand g283 (n_438, n_434, n_435, n_436);
  xor g284 (n_437, A[46], B[46]);
  xor g285 (Z[46], n_433, n_437);
  nand g286 (n_439, A[47], B[47]);
  nand g287 (n_440, A[47], n_438);
  nand g288 (n_441, B[47], n_438);
  nand g289 (n_443, n_439, n_440, n_441);
  xor g290 (n_442, A[47], B[47]);
  xor g291 (Z[47], n_438, n_442);
  nand g292 (n_444, A[48], B[48]);
  nand g293 (n_445, A[48], n_443);
  nand g294 (n_446, B[48], n_443);
  nand g295 (n_448, n_444, n_445, n_446);
  xor g296 (n_447, A[48], B[48]);
  xor g297 (Z[48], n_443, n_447);
  nand g298 (n_449, A[49], B[49]);
  nand g299 (n_450, A[49], n_448);
  nand g300 (n_451, B[49], n_448);
  nand g301 (n_453, n_449, n_450, n_451);
  xor g302 (n_452, A[49], B[49]);
  xor g303 (Z[49], n_448, n_452);
  nand g304 (n_454, A[50], B[50]);
  nand g305 (n_455, A[50], n_453);
  nand g306 (n_456, B[50], n_453);
  nand g307 (n_458, n_454, n_455, n_456);
  xor g308 (n_457, A[50], B[50]);
  xor g309 (Z[50], n_453, n_457);
  nand g310 (n_459, A[51], B[51]);
  nand g311 (n_460, A[51], n_458);
  nand g312 (n_461, B[51], n_458);
  nand g313 (n_463, n_459, n_460, n_461);
  xor g314 (n_462, A[51], B[51]);
  xor g315 (Z[51], n_458, n_462);
  nand g316 (n_464, A[52], B[52]);
  nand g317 (n_465, A[52], n_463);
  nand g318 (n_466, B[52], n_463);
  nand g319 (n_468, n_464, n_465, n_466);
  xor g320 (n_467, A[52], B[52]);
  xor g321 (Z[52], n_463, n_467);
  nand g322 (n_469, A[53], B[53]);
  nand g323 (n_470, A[53], n_468);
  nand g324 (n_471, B[53], n_468);
  nand g325 (n_473, n_469, n_470, n_471);
  xor g326 (n_472, A[53], B[53]);
  xor g327 (Z[53], n_468, n_472);
  nand g328 (n_474, A[54], B[54]);
  nand g329 (n_475, A[54], n_473);
  nand g330 (n_476, B[54], n_473);
  nand g331 (n_478, n_474, n_475, n_476);
  xor g332 (n_477, A[54], B[54]);
  xor g333 (Z[54], n_473, n_477);
  nand g334 (n_479, A[55], B[55]);
  nand g335 (n_480, A[55], n_478);
  nand g336 (n_481, B[55], n_478);
  nand g337 (n_483, n_479, n_480, n_481);
  xor g338 (n_482, A[55], B[55]);
  xor g339 (Z[55], n_478, n_482);
  nand g340 (n_484, A[56], B[56]);
  nand g341 (n_485, A[56], n_483);
  nand g342 (n_486, B[56], n_483);
  nand g343 (n_488, n_484, n_485, n_486);
  xor g344 (n_487, A[56], B[56]);
  xor g345 (Z[56], n_483, n_487);
  nand g346 (n_489, A[57], B[57]);
  nand g347 (n_490, A[57], n_488);
  nand g348 (n_491, B[57], n_488);
  nand g349 (n_493, n_489, n_490, n_491);
  xor g350 (n_492, A[57], B[57]);
  xor g351 (Z[57], n_488, n_492);
  nand g352 (n_494, A[58], B[58]);
  nand g353 (n_495, A[58], n_493);
  nand g354 (n_496, B[58], n_493);
  nand g355 (n_498, n_494, n_495, n_496);
  xor g356 (n_497, A[58], B[58]);
  xor g357 (Z[58], n_493, n_497);
  nand g358 (n_499, A[59], B[59]);
  nand g359 (n_500, A[59], n_498);
  nand g360 (n_501, B[59], n_498);
  nand g361 (n_503, n_499, n_500, n_501);
  xor g362 (n_502, A[59], B[59]);
  xor g363 (Z[59], n_498, n_502);
  nand g364 (n_504, A[60], B[60]);
  nand g365 (n_505, A[60], n_503);
  nand g366 (n_506, B[60], n_503);
  nand g367 (n_508, n_504, n_505, n_506);
  xor g368 (n_507, A[60], B[60]);
  xor g369 (Z[60], n_503, n_507);
  nand g370 (n_509, A[61], B[61]);
  nand g371 (n_510, A[61], n_508);
  nand g372 (n_511, B[61], n_508);
  nand g373 (n_513, n_509, n_510, n_511);
  xor g374 (n_512, A[61], B[61]);
  xor g375 (Z[61], n_508, n_512);
  nand g376 (n_514, A[62], B[62]);
  nand g377 (n_515, A[62], n_513);
  nand g378 (n_516, B[62], n_513);
  nand g379 (n_518, n_514, n_515, n_516);
  xor g380 (n_517, A[62], B[62]);
  xor g381 (Z[62], n_513, n_517);
  nand g382 (n_519, A[63], B[63]);
  nand g383 (n_520, A[63], n_518);
  nand g384 (n_521, B[63], n_518);
  nand g385 (n_523, n_519, n_520, n_521);
  xor g386 (n_522, A[63], B[63]);
  xor g387 (Z[63], n_518, n_522);
  nand g388 (n_524, A[64], B[64]);
  nand g389 (n_525, A[64], n_523);
  nand g390 (n_526, B[64], n_523);
  nand g391 (n_528, n_524, n_525, n_526);
  xor g392 (n_527, A[64], B[64]);
  xor g393 (Z[64], n_523, n_527);
  nand g397 (n_203, n_529, n_530, n_531);
  xor g399 (Z[65], n_528, n_532);
  or g401 (n_529, A[65], B[65]);
  xor g402 (n_532, A[65], B[65]);
  or g403 (n_210, wc, n_204);
  not gc (wc, A[1]);
  or g404 (n_211, wc0, n_204);
  not gc0 (wc0, B[1]);
  xnor g405 (Z[1], n_204, n_212);
  or g406 (n_530, A[65], wc1);
  not gc1 (wc1, n_528);
  or g407 (n_531, B[65], wc2);
  not gc2 (wc2, n_528);
endmodule

module add_signed_2443_GENERIC(A, B, Z);
  input [65:0] A, B;
  output [66:0] Z;
  wire [65:0] A, B;
  wire [66:0] Z;
  add_signed_2443_GENERIC_REAL g1(.A ({A[65:2], A[0], A[0]}), .B (B),
       .Z (Z));
endmodule

module add_signed_2443_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [65:0] A, B;
  output [66:0] Z;
  wire [65:0] A, B;
  wire [66:0] Z;
  wire n_203, n_204, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502;
  wire n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510;
  wire n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518;
  wire n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526;
  wire n_527, n_528, n_529, n_530, n_531, n_532;
  not g3 (Z[66], n_203);
  nand g4 (n_204, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_209, A[1], B[1]);
  nand g13 (n_213, n_209, n_210, n_211);
  xor g14 (n_212, A[1], B[1]);
  nand g16 (n_214, A[2], B[2]);
  nand g17 (n_215, A[2], n_213);
  nand g18 (n_216, B[2], n_213);
  nand g19 (n_218, n_214, n_215, n_216);
  xor g20 (n_217, A[2], B[2]);
  xor g21 (Z[2], n_213, n_217);
  nand g22 (n_219, A[3], B[3]);
  nand g23 (n_220, A[3], n_218);
  nand g24 (n_221, B[3], n_218);
  nand g25 (n_223, n_219, n_220, n_221);
  xor g26 (n_222, A[3], B[3]);
  xor g27 (Z[3], n_218, n_222);
  nand g28 (n_224, A[4], B[4]);
  nand g29 (n_225, A[4], n_223);
  nand g30 (n_226, B[4], n_223);
  nand g31 (n_228, n_224, n_225, n_226);
  xor g32 (n_227, A[4], B[4]);
  xor g33 (Z[4], n_223, n_227);
  nand g34 (n_229, A[5], B[5]);
  nand g35 (n_230, A[5], n_228);
  nand g36 (n_231, B[5], n_228);
  nand g37 (n_233, n_229, n_230, n_231);
  xor g38 (n_232, A[5], B[5]);
  xor g39 (Z[5], n_228, n_232);
  nand g40 (n_234, A[6], B[6]);
  nand g41 (n_235, A[6], n_233);
  nand g42 (n_236, B[6], n_233);
  nand g43 (n_238, n_234, n_235, n_236);
  xor g44 (n_237, A[6], B[6]);
  xor g45 (Z[6], n_233, n_237);
  nand g46 (n_239, A[7], B[7]);
  nand g47 (n_240, A[7], n_238);
  nand g48 (n_241, B[7], n_238);
  nand g49 (n_243, n_239, n_240, n_241);
  xor g50 (n_242, A[7], B[7]);
  xor g51 (Z[7], n_238, n_242);
  nand g52 (n_244, A[8], B[8]);
  nand g53 (n_245, A[8], n_243);
  nand g54 (n_246, B[8], n_243);
  nand g55 (n_248, n_244, n_245, n_246);
  xor g56 (n_247, A[8], B[8]);
  xor g57 (Z[8], n_243, n_247);
  nand g58 (n_249, A[9], B[9]);
  nand g59 (n_250, A[9], n_248);
  nand g60 (n_251, B[9], n_248);
  nand g61 (n_253, n_249, n_250, n_251);
  xor g62 (n_252, A[9], B[9]);
  xor g63 (Z[9], n_248, n_252);
  nand g64 (n_254, A[10], B[10]);
  nand g65 (n_255, A[10], n_253);
  nand g66 (n_256, B[10], n_253);
  nand g67 (n_258, n_254, n_255, n_256);
  xor g68 (n_257, A[10], B[10]);
  xor g69 (Z[10], n_253, n_257);
  nand g70 (n_259, A[11], B[11]);
  nand g71 (n_260, A[11], n_258);
  nand g72 (n_261, B[11], n_258);
  nand g73 (n_263, n_259, n_260, n_261);
  xor g74 (n_262, A[11], B[11]);
  xor g75 (Z[11], n_258, n_262);
  nand g76 (n_264, A[12], B[12]);
  nand g77 (n_265, A[12], n_263);
  nand g78 (n_266, B[12], n_263);
  nand g79 (n_268, n_264, n_265, n_266);
  xor g80 (n_267, A[12], B[12]);
  xor g81 (Z[12], n_263, n_267);
  nand g82 (n_269, A[13], B[13]);
  nand g83 (n_270, A[13], n_268);
  nand g84 (n_271, B[13], n_268);
  nand g85 (n_273, n_269, n_270, n_271);
  xor g86 (n_272, A[13], B[13]);
  xor g87 (Z[13], n_268, n_272);
  nand g88 (n_274, A[14], B[14]);
  nand g89 (n_275, A[14], n_273);
  nand g90 (n_276, B[14], n_273);
  nand g91 (n_278, n_274, n_275, n_276);
  xor g92 (n_277, A[14], B[14]);
  xor g93 (Z[14], n_273, n_277);
  nand g94 (n_279, A[15], B[15]);
  nand g95 (n_280, A[15], n_278);
  nand g96 (n_281, B[15], n_278);
  nand g97 (n_283, n_279, n_280, n_281);
  xor g98 (n_282, A[15], B[15]);
  xor g99 (Z[15], n_278, n_282);
  nand g100 (n_284, A[16], B[16]);
  nand g101 (n_285, A[16], n_283);
  nand g102 (n_286, B[16], n_283);
  nand g103 (n_288, n_284, n_285, n_286);
  xor g104 (n_287, A[16], B[16]);
  xor g105 (Z[16], n_283, n_287);
  nand g106 (n_289, A[17], B[17]);
  nand g107 (n_290, A[17], n_288);
  nand g108 (n_291, B[17], n_288);
  nand g109 (n_293, n_289, n_290, n_291);
  xor g110 (n_292, A[17], B[17]);
  xor g111 (Z[17], n_288, n_292);
  nand g112 (n_294, A[18], B[18]);
  nand g113 (n_295, A[18], n_293);
  nand g114 (n_296, B[18], n_293);
  nand g115 (n_298, n_294, n_295, n_296);
  xor g116 (n_297, A[18], B[18]);
  xor g117 (Z[18], n_293, n_297);
  nand g118 (n_299, A[19], B[19]);
  nand g119 (n_300, A[19], n_298);
  nand g120 (n_301, B[19], n_298);
  nand g121 (n_303, n_299, n_300, n_301);
  xor g122 (n_302, A[19], B[19]);
  xor g123 (Z[19], n_298, n_302);
  nand g124 (n_304, A[20], B[20]);
  nand g125 (n_305, A[20], n_303);
  nand g126 (n_306, B[20], n_303);
  nand g127 (n_308, n_304, n_305, n_306);
  xor g128 (n_307, A[20], B[20]);
  xor g129 (Z[20], n_303, n_307);
  nand g130 (n_309, A[21], B[21]);
  nand g131 (n_310, A[21], n_308);
  nand g132 (n_311, B[21], n_308);
  nand g133 (n_313, n_309, n_310, n_311);
  xor g134 (n_312, A[21], B[21]);
  xor g135 (Z[21], n_308, n_312);
  nand g136 (n_314, A[22], B[22]);
  nand g137 (n_315, A[22], n_313);
  nand g138 (n_316, B[22], n_313);
  nand g139 (n_318, n_314, n_315, n_316);
  xor g140 (n_317, A[22], B[22]);
  xor g141 (Z[22], n_313, n_317);
  nand g142 (n_319, A[23], B[23]);
  nand g143 (n_320, A[23], n_318);
  nand g144 (n_321, B[23], n_318);
  nand g145 (n_323, n_319, n_320, n_321);
  xor g146 (n_322, A[23], B[23]);
  xor g147 (Z[23], n_318, n_322);
  nand g148 (n_324, A[24], B[24]);
  nand g149 (n_325, A[24], n_323);
  nand g150 (n_326, B[24], n_323);
  nand g151 (n_328, n_324, n_325, n_326);
  xor g152 (n_327, A[24], B[24]);
  xor g153 (Z[24], n_323, n_327);
  nand g154 (n_329, A[25], B[25]);
  nand g155 (n_330, A[25], n_328);
  nand g156 (n_331, B[25], n_328);
  nand g157 (n_333, n_329, n_330, n_331);
  xor g158 (n_332, A[25], B[25]);
  xor g159 (Z[25], n_328, n_332);
  nand g160 (n_334, A[26], B[26]);
  nand g161 (n_335, A[26], n_333);
  nand g162 (n_336, B[26], n_333);
  nand g163 (n_338, n_334, n_335, n_336);
  xor g164 (n_337, A[26], B[26]);
  xor g165 (Z[26], n_333, n_337);
  nand g166 (n_339, A[27], B[27]);
  nand g167 (n_340, A[27], n_338);
  nand g168 (n_341, B[27], n_338);
  nand g169 (n_343, n_339, n_340, n_341);
  xor g170 (n_342, A[27], B[27]);
  xor g171 (Z[27], n_338, n_342);
  nand g172 (n_344, A[28], B[28]);
  nand g173 (n_345, A[28], n_343);
  nand g174 (n_346, B[28], n_343);
  nand g175 (n_348, n_344, n_345, n_346);
  xor g176 (n_347, A[28], B[28]);
  xor g177 (Z[28], n_343, n_347);
  nand g178 (n_349, A[29], B[29]);
  nand g179 (n_350, A[29], n_348);
  nand g180 (n_351, B[29], n_348);
  nand g181 (n_353, n_349, n_350, n_351);
  xor g182 (n_352, A[29], B[29]);
  xor g183 (Z[29], n_348, n_352);
  nand g184 (n_354, A[30], B[30]);
  nand g185 (n_355, A[30], n_353);
  nand g186 (n_356, B[30], n_353);
  nand g187 (n_358, n_354, n_355, n_356);
  xor g188 (n_357, A[30], B[30]);
  xor g189 (Z[30], n_353, n_357);
  nand g190 (n_359, A[31], B[31]);
  nand g191 (n_360, A[31], n_358);
  nand g192 (n_361, B[31], n_358);
  nand g193 (n_363, n_359, n_360, n_361);
  xor g194 (n_362, A[31], B[31]);
  xor g195 (Z[31], n_358, n_362);
  nand g196 (n_364, A[32], B[32]);
  nand g197 (n_365, A[32], n_363);
  nand g198 (n_366, B[32], n_363);
  nand g199 (n_368, n_364, n_365, n_366);
  xor g200 (n_367, A[32], B[32]);
  xor g201 (Z[32], n_363, n_367);
  nand g202 (n_369, A[33], B[33]);
  nand g203 (n_370, A[33], n_368);
  nand g204 (n_371, B[33], n_368);
  nand g205 (n_373, n_369, n_370, n_371);
  xor g206 (n_372, A[33], B[33]);
  xor g207 (Z[33], n_368, n_372);
  nand g208 (n_374, A[34], B[34]);
  nand g209 (n_375, A[34], n_373);
  nand g210 (n_376, B[34], n_373);
  nand g211 (n_378, n_374, n_375, n_376);
  xor g212 (n_377, A[34], B[34]);
  xor g213 (Z[34], n_373, n_377);
  nand g214 (n_379, A[35], B[35]);
  nand g215 (n_380, A[35], n_378);
  nand g216 (n_381, B[35], n_378);
  nand g217 (n_383, n_379, n_380, n_381);
  xor g218 (n_382, A[35], B[35]);
  xor g219 (Z[35], n_378, n_382);
  nand g220 (n_384, A[36], B[36]);
  nand g221 (n_385, A[36], n_383);
  nand g222 (n_386, B[36], n_383);
  nand g223 (n_388, n_384, n_385, n_386);
  xor g224 (n_387, A[36], B[36]);
  xor g225 (Z[36], n_383, n_387);
  nand g226 (n_389, A[37], B[37]);
  nand g227 (n_390, A[37], n_388);
  nand g228 (n_391, B[37], n_388);
  nand g229 (n_393, n_389, n_390, n_391);
  xor g230 (n_392, A[37], B[37]);
  xor g231 (Z[37], n_388, n_392);
  nand g232 (n_394, A[38], B[38]);
  nand g233 (n_395, A[38], n_393);
  nand g234 (n_396, B[38], n_393);
  nand g235 (n_398, n_394, n_395, n_396);
  xor g236 (n_397, A[38], B[38]);
  xor g237 (Z[38], n_393, n_397);
  nand g238 (n_399, A[39], B[39]);
  nand g239 (n_400, A[39], n_398);
  nand g240 (n_401, B[39], n_398);
  nand g241 (n_403, n_399, n_400, n_401);
  xor g242 (n_402, A[39], B[39]);
  xor g243 (Z[39], n_398, n_402);
  nand g244 (n_404, A[40], B[40]);
  nand g245 (n_405, A[40], n_403);
  nand g246 (n_406, B[40], n_403);
  nand g247 (n_408, n_404, n_405, n_406);
  xor g248 (n_407, A[40], B[40]);
  xor g249 (Z[40], n_403, n_407);
  nand g250 (n_409, A[41], B[41]);
  nand g251 (n_410, A[41], n_408);
  nand g252 (n_411, B[41], n_408);
  nand g253 (n_413, n_409, n_410, n_411);
  xor g254 (n_412, A[41], B[41]);
  xor g255 (Z[41], n_408, n_412);
  nand g256 (n_414, A[42], B[42]);
  nand g257 (n_415, A[42], n_413);
  nand g258 (n_416, B[42], n_413);
  nand g259 (n_418, n_414, n_415, n_416);
  xor g260 (n_417, A[42], B[42]);
  xor g261 (Z[42], n_413, n_417);
  nand g262 (n_419, A[43], B[43]);
  nand g263 (n_420, A[43], n_418);
  nand g264 (n_421, B[43], n_418);
  nand g265 (n_423, n_419, n_420, n_421);
  xor g266 (n_422, A[43], B[43]);
  xor g267 (Z[43], n_418, n_422);
  nand g268 (n_424, A[44], B[44]);
  nand g269 (n_425, A[44], n_423);
  nand g270 (n_426, B[44], n_423);
  nand g271 (n_428, n_424, n_425, n_426);
  xor g272 (n_427, A[44], B[44]);
  xor g273 (Z[44], n_423, n_427);
  nand g274 (n_429, A[45], B[45]);
  nand g275 (n_430, A[45], n_428);
  nand g276 (n_431, B[45], n_428);
  nand g277 (n_433, n_429, n_430, n_431);
  xor g278 (n_432, A[45], B[45]);
  xor g279 (Z[45], n_428, n_432);
  nand g280 (n_434, A[46], B[46]);
  nand g281 (n_435, A[46], n_433);
  nand g282 (n_436, B[46], n_433);
  nand g283 (n_438, n_434, n_435, n_436);
  xor g284 (n_437, A[46], B[46]);
  xor g285 (Z[46], n_433, n_437);
  nand g286 (n_439, A[47], B[47]);
  nand g287 (n_440, A[47], n_438);
  nand g288 (n_441, B[47], n_438);
  nand g289 (n_443, n_439, n_440, n_441);
  xor g290 (n_442, A[47], B[47]);
  xor g291 (Z[47], n_438, n_442);
  nand g292 (n_444, A[48], B[48]);
  nand g293 (n_445, A[48], n_443);
  nand g294 (n_446, B[48], n_443);
  nand g295 (n_448, n_444, n_445, n_446);
  xor g296 (n_447, A[48], B[48]);
  xor g297 (Z[48], n_443, n_447);
  nand g298 (n_449, A[49], B[49]);
  nand g299 (n_450, A[49], n_448);
  nand g300 (n_451, B[49], n_448);
  nand g301 (n_453, n_449, n_450, n_451);
  xor g302 (n_452, A[49], B[49]);
  xor g303 (Z[49], n_448, n_452);
  nand g304 (n_454, A[50], B[50]);
  nand g305 (n_455, A[50], n_453);
  nand g306 (n_456, B[50], n_453);
  nand g307 (n_458, n_454, n_455, n_456);
  xor g308 (n_457, A[50], B[50]);
  xor g309 (Z[50], n_453, n_457);
  nand g310 (n_459, A[51], B[51]);
  nand g311 (n_460, A[51], n_458);
  nand g312 (n_461, B[51], n_458);
  nand g313 (n_463, n_459, n_460, n_461);
  xor g314 (n_462, A[51], B[51]);
  xor g315 (Z[51], n_458, n_462);
  nand g316 (n_464, A[52], B[52]);
  nand g317 (n_465, A[52], n_463);
  nand g318 (n_466, B[52], n_463);
  nand g319 (n_468, n_464, n_465, n_466);
  xor g320 (n_467, A[52], B[52]);
  xor g321 (Z[52], n_463, n_467);
  nand g322 (n_469, A[53], B[53]);
  nand g323 (n_470, A[53], n_468);
  nand g324 (n_471, B[53], n_468);
  nand g325 (n_473, n_469, n_470, n_471);
  xor g326 (n_472, A[53], B[53]);
  xor g327 (Z[53], n_468, n_472);
  nand g328 (n_474, A[54], B[54]);
  nand g329 (n_475, A[54], n_473);
  nand g330 (n_476, B[54], n_473);
  nand g331 (n_478, n_474, n_475, n_476);
  xor g332 (n_477, A[54], B[54]);
  xor g333 (Z[54], n_473, n_477);
  nand g334 (n_479, A[55], B[55]);
  nand g335 (n_480, A[55], n_478);
  nand g336 (n_481, B[55], n_478);
  nand g337 (n_483, n_479, n_480, n_481);
  xor g338 (n_482, A[55], B[55]);
  xor g339 (Z[55], n_478, n_482);
  nand g340 (n_484, A[56], B[56]);
  nand g341 (n_485, A[56], n_483);
  nand g342 (n_486, B[56], n_483);
  nand g343 (n_488, n_484, n_485, n_486);
  xor g344 (n_487, A[56], B[56]);
  xor g345 (Z[56], n_483, n_487);
  nand g346 (n_489, A[57], B[57]);
  nand g347 (n_490, A[57], n_488);
  nand g348 (n_491, B[57], n_488);
  nand g349 (n_493, n_489, n_490, n_491);
  xor g350 (n_492, A[57], B[57]);
  xor g351 (Z[57], n_488, n_492);
  nand g352 (n_494, A[58], B[58]);
  nand g353 (n_495, A[58], n_493);
  nand g354 (n_496, B[58], n_493);
  nand g355 (n_498, n_494, n_495, n_496);
  xor g356 (n_497, A[58], B[58]);
  xor g357 (Z[58], n_493, n_497);
  nand g358 (n_499, A[59], B[59]);
  nand g359 (n_500, A[59], n_498);
  nand g360 (n_501, B[59], n_498);
  nand g361 (n_503, n_499, n_500, n_501);
  xor g362 (n_502, A[59], B[59]);
  xor g363 (Z[59], n_498, n_502);
  nand g364 (n_504, A[60], B[60]);
  nand g365 (n_505, A[60], n_503);
  nand g366 (n_506, B[60], n_503);
  nand g367 (n_508, n_504, n_505, n_506);
  xor g368 (n_507, A[60], B[60]);
  xor g369 (Z[60], n_503, n_507);
  nand g370 (n_509, A[61], B[61]);
  nand g371 (n_510, A[61], n_508);
  nand g372 (n_511, B[61], n_508);
  nand g373 (n_513, n_509, n_510, n_511);
  xor g374 (n_512, A[61], B[61]);
  xor g375 (Z[61], n_508, n_512);
  nand g376 (n_514, A[62], B[62]);
  nand g377 (n_515, A[62], n_513);
  nand g378 (n_516, B[62], n_513);
  nand g379 (n_518, n_514, n_515, n_516);
  xor g380 (n_517, A[62], B[62]);
  xor g381 (Z[62], n_513, n_517);
  nand g382 (n_519, A[63], B[63]);
  nand g383 (n_520, A[63], n_518);
  nand g384 (n_521, B[63], n_518);
  nand g385 (n_523, n_519, n_520, n_521);
  xor g386 (n_522, A[63], B[63]);
  xor g387 (Z[63], n_518, n_522);
  nand g388 (n_524, A[64], B[64]);
  nand g389 (n_525, A[64], n_523);
  nand g390 (n_526, B[64], n_523);
  nand g391 (n_528, n_524, n_525, n_526);
  xor g392 (n_527, A[64], B[64]);
  xor g393 (Z[64], n_523, n_527);
  nand g397 (n_203, n_529, n_530, n_531);
  xor g399 (Z[65], n_528, n_532);
  or g401 (n_529, A[65], B[65]);
  xor g402 (n_532, A[65], B[65]);
  or g403 (n_210, wc, n_204);
  not gc (wc, A[1]);
  or g404 (n_211, wc0, n_204);
  not gc0 (wc0, B[1]);
  xnor g405 (Z[1], n_204, n_212);
  or g406 (n_530, A[65], wc1);
  not gc1 (wc1, n_528);
  or g407 (n_531, B[65], wc2);
  not gc2 (wc2, n_528);
endmodule

module add_signed_2443_1_GENERIC(A, B, Z);
  input [65:0] A, B;
  output [66:0] Z;
  wire [65:0] A, B;
  wire [66:0] Z;
  add_signed_2443_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3032_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [63:0] A, B;
  output [64:0] Z;
  wire [63:0] A, B;
  wire [64:0] Z;
  wire n_197, n_198, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516;
  not g3 (Z[64], n_197);
  nand g4 (n_198, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_203, A[1], B[1]);
  nand g13 (n_207, n_203, n_204, n_205);
  xor g14 (n_206, A[1], B[1]);
  nand g16 (n_208, A[2], B[2]);
  nand g17 (n_209, A[2], n_207);
  nand g18 (n_210, B[2], n_207);
  nand g19 (n_212, n_208, n_209, n_210);
  xor g20 (n_211, A[2], B[2]);
  xor g21 (Z[2], n_207, n_211);
  nand g22 (n_213, A[3], B[3]);
  nand g23 (n_214, A[3], n_212);
  nand g24 (n_215, B[3], n_212);
  nand g25 (n_217, n_213, n_214, n_215);
  xor g26 (n_216, A[3], B[3]);
  xor g27 (Z[3], n_212, n_216);
  nand g28 (n_218, A[4], B[4]);
  nand g29 (n_219, A[4], n_217);
  nand g30 (n_220, B[4], n_217);
  nand g31 (n_222, n_218, n_219, n_220);
  xor g32 (n_221, A[4], B[4]);
  xor g33 (Z[4], n_217, n_221);
  nand g34 (n_223, A[5], B[5]);
  nand g35 (n_224, A[5], n_222);
  nand g36 (n_225, B[5], n_222);
  nand g37 (n_227, n_223, n_224, n_225);
  xor g38 (n_226, A[5], B[5]);
  xor g39 (Z[5], n_222, n_226);
  nand g40 (n_228, A[6], B[6]);
  nand g41 (n_229, A[6], n_227);
  nand g42 (n_230, B[6], n_227);
  nand g43 (n_232, n_228, n_229, n_230);
  xor g44 (n_231, A[6], B[6]);
  xor g45 (Z[6], n_227, n_231);
  nand g46 (n_233, A[7], B[7]);
  nand g47 (n_234, A[7], n_232);
  nand g48 (n_235, B[7], n_232);
  nand g49 (n_237, n_233, n_234, n_235);
  xor g50 (n_236, A[7], B[7]);
  xor g51 (Z[7], n_232, n_236);
  nand g52 (n_238, A[8], B[8]);
  nand g53 (n_239, A[8], n_237);
  nand g54 (n_240, B[8], n_237);
  nand g55 (n_242, n_238, n_239, n_240);
  xor g56 (n_241, A[8], B[8]);
  xor g57 (Z[8], n_237, n_241);
  nand g58 (n_243, A[9], B[9]);
  nand g59 (n_244, A[9], n_242);
  nand g60 (n_245, B[9], n_242);
  nand g61 (n_247, n_243, n_244, n_245);
  xor g62 (n_246, A[9], B[9]);
  xor g63 (Z[9], n_242, n_246);
  nand g64 (n_248, A[10], B[10]);
  nand g65 (n_249, A[10], n_247);
  nand g66 (n_250, B[10], n_247);
  nand g67 (n_252, n_248, n_249, n_250);
  xor g68 (n_251, A[10], B[10]);
  xor g69 (Z[10], n_247, n_251);
  nand g70 (n_253, A[11], B[11]);
  nand g71 (n_254, A[11], n_252);
  nand g72 (n_255, B[11], n_252);
  nand g73 (n_257, n_253, n_254, n_255);
  xor g74 (n_256, A[11], B[11]);
  xor g75 (Z[11], n_252, n_256);
  nand g76 (n_258, A[12], B[12]);
  nand g77 (n_259, A[12], n_257);
  nand g78 (n_260, B[12], n_257);
  nand g79 (n_262, n_258, n_259, n_260);
  xor g80 (n_261, A[12], B[12]);
  xor g81 (Z[12], n_257, n_261);
  nand g82 (n_263, A[13], B[13]);
  nand g83 (n_264, A[13], n_262);
  nand g84 (n_265, B[13], n_262);
  nand g85 (n_267, n_263, n_264, n_265);
  xor g86 (n_266, A[13], B[13]);
  xor g87 (Z[13], n_262, n_266);
  nand g88 (n_268, A[14], B[14]);
  nand g89 (n_269, A[14], n_267);
  nand g90 (n_270, B[14], n_267);
  nand g91 (n_272, n_268, n_269, n_270);
  xor g92 (n_271, A[14], B[14]);
  xor g93 (Z[14], n_267, n_271);
  nand g94 (n_273, A[15], B[15]);
  nand g95 (n_274, A[15], n_272);
  nand g96 (n_275, B[15], n_272);
  nand g97 (n_277, n_273, n_274, n_275);
  xor g98 (n_276, A[15], B[15]);
  xor g99 (Z[15], n_272, n_276);
  nand g100 (n_278, A[16], B[16]);
  nand g101 (n_279, A[16], n_277);
  nand g102 (n_280, B[16], n_277);
  nand g103 (n_282, n_278, n_279, n_280);
  xor g104 (n_281, A[16], B[16]);
  xor g105 (Z[16], n_277, n_281);
  nand g106 (n_283, A[17], B[17]);
  nand g107 (n_284, A[17], n_282);
  nand g108 (n_285, B[17], n_282);
  nand g109 (n_287, n_283, n_284, n_285);
  xor g110 (n_286, A[17], B[17]);
  xor g111 (Z[17], n_282, n_286);
  nand g112 (n_288, A[18], B[18]);
  nand g113 (n_289, A[18], n_287);
  nand g114 (n_290, B[18], n_287);
  nand g115 (n_292, n_288, n_289, n_290);
  xor g116 (n_291, A[18], B[18]);
  xor g117 (Z[18], n_287, n_291);
  nand g118 (n_293, A[19], B[19]);
  nand g119 (n_294, A[19], n_292);
  nand g120 (n_295, B[19], n_292);
  nand g121 (n_297, n_293, n_294, n_295);
  xor g122 (n_296, A[19], B[19]);
  xor g123 (Z[19], n_292, n_296);
  nand g124 (n_298, A[20], B[20]);
  nand g125 (n_299, A[20], n_297);
  nand g126 (n_300, B[20], n_297);
  nand g127 (n_302, n_298, n_299, n_300);
  xor g128 (n_301, A[20], B[20]);
  xor g129 (Z[20], n_297, n_301);
  nand g130 (n_303, A[21], B[21]);
  nand g131 (n_304, A[21], n_302);
  nand g132 (n_305, B[21], n_302);
  nand g133 (n_307, n_303, n_304, n_305);
  xor g134 (n_306, A[21], B[21]);
  xor g135 (Z[21], n_302, n_306);
  nand g136 (n_308, A[22], B[22]);
  nand g137 (n_309, A[22], n_307);
  nand g138 (n_310, B[22], n_307);
  nand g139 (n_312, n_308, n_309, n_310);
  xor g140 (n_311, A[22], B[22]);
  xor g141 (Z[22], n_307, n_311);
  nand g142 (n_313, A[23], B[23]);
  nand g143 (n_314, A[23], n_312);
  nand g144 (n_315, B[23], n_312);
  nand g145 (n_317, n_313, n_314, n_315);
  xor g146 (n_316, A[23], B[23]);
  xor g147 (Z[23], n_312, n_316);
  nand g148 (n_318, A[24], B[24]);
  nand g149 (n_319, A[24], n_317);
  nand g150 (n_320, B[24], n_317);
  nand g151 (n_322, n_318, n_319, n_320);
  xor g152 (n_321, A[24], B[24]);
  xor g153 (Z[24], n_317, n_321);
  nand g154 (n_323, A[25], B[25]);
  nand g155 (n_324, A[25], n_322);
  nand g156 (n_325, B[25], n_322);
  nand g157 (n_327, n_323, n_324, n_325);
  xor g158 (n_326, A[25], B[25]);
  xor g159 (Z[25], n_322, n_326);
  nand g160 (n_328, A[26], B[26]);
  nand g161 (n_329, A[26], n_327);
  nand g162 (n_330, B[26], n_327);
  nand g163 (n_332, n_328, n_329, n_330);
  xor g164 (n_331, A[26], B[26]);
  xor g165 (Z[26], n_327, n_331);
  nand g166 (n_333, A[27], B[27]);
  nand g167 (n_334, A[27], n_332);
  nand g168 (n_335, B[27], n_332);
  nand g169 (n_337, n_333, n_334, n_335);
  xor g170 (n_336, A[27], B[27]);
  xor g171 (Z[27], n_332, n_336);
  nand g172 (n_338, A[28], B[28]);
  nand g173 (n_339, A[28], n_337);
  nand g174 (n_340, B[28], n_337);
  nand g175 (n_342, n_338, n_339, n_340);
  xor g176 (n_341, A[28], B[28]);
  xor g177 (Z[28], n_337, n_341);
  nand g178 (n_343, A[29], B[29]);
  nand g179 (n_344, A[29], n_342);
  nand g180 (n_345, B[29], n_342);
  nand g181 (n_347, n_343, n_344, n_345);
  xor g182 (n_346, A[29], B[29]);
  xor g183 (Z[29], n_342, n_346);
  nand g184 (n_348, A[30], B[30]);
  nand g185 (n_349, A[30], n_347);
  nand g186 (n_350, B[30], n_347);
  nand g187 (n_352, n_348, n_349, n_350);
  xor g188 (n_351, A[30], B[30]);
  xor g189 (Z[30], n_347, n_351);
  nand g190 (n_353, A[31], B[31]);
  nand g191 (n_354, A[31], n_352);
  nand g192 (n_355, B[31], n_352);
  nand g193 (n_357, n_353, n_354, n_355);
  xor g194 (n_356, A[31], B[31]);
  xor g195 (Z[31], n_352, n_356);
  nand g196 (n_358, A[32], B[32]);
  nand g197 (n_359, A[32], n_357);
  nand g198 (n_360, B[32], n_357);
  nand g199 (n_362, n_358, n_359, n_360);
  xor g200 (n_361, A[32], B[32]);
  xor g201 (Z[32], n_357, n_361);
  nand g202 (n_363, A[33], B[33]);
  nand g203 (n_364, A[33], n_362);
  nand g204 (n_365, B[33], n_362);
  nand g205 (n_367, n_363, n_364, n_365);
  xor g206 (n_366, A[33], B[33]);
  xor g207 (Z[33], n_362, n_366);
  nand g208 (n_368, A[34], B[34]);
  nand g209 (n_369, A[34], n_367);
  nand g210 (n_370, B[34], n_367);
  nand g211 (n_372, n_368, n_369, n_370);
  xor g212 (n_371, A[34], B[34]);
  xor g213 (Z[34], n_367, n_371);
  nand g214 (n_373, A[35], B[35]);
  nand g215 (n_374, A[35], n_372);
  nand g216 (n_375, B[35], n_372);
  nand g217 (n_377, n_373, n_374, n_375);
  xor g218 (n_376, A[35], B[35]);
  xor g219 (Z[35], n_372, n_376);
  nand g220 (n_378, A[36], B[36]);
  nand g221 (n_379, A[36], n_377);
  nand g222 (n_380, B[36], n_377);
  nand g223 (n_382, n_378, n_379, n_380);
  xor g224 (n_381, A[36], B[36]);
  xor g225 (Z[36], n_377, n_381);
  nand g226 (n_383, A[37], B[37]);
  nand g227 (n_384, A[37], n_382);
  nand g228 (n_385, B[37], n_382);
  nand g229 (n_387, n_383, n_384, n_385);
  xor g230 (n_386, A[37], B[37]);
  xor g231 (Z[37], n_382, n_386);
  nand g232 (n_388, A[38], B[38]);
  nand g233 (n_389, A[38], n_387);
  nand g234 (n_390, B[38], n_387);
  nand g235 (n_392, n_388, n_389, n_390);
  xor g236 (n_391, A[38], B[38]);
  xor g237 (Z[38], n_387, n_391);
  nand g238 (n_393, A[39], B[39]);
  nand g239 (n_394, A[39], n_392);
  nand g240 (n_395, B[39], n_392);
  nand g241 (n_397, n_393, n_394, n_395);
  xor g242 (n_396, A[39], B[39]);
  xor g243 (Z[39], n_392, n_396);
  nand g244 (n_398, A[40], B[40]);
  nand g245 (n_399, A[40], n_397);
  nand g246 (n_400, B[40], n_397);
  nand g247 (n_402, n_398, n_399, n_400);
  xor g248 (n_401, A[40], B[40]);
  xor g249 (Z[40], n_397, n_401);
  nand g250 (n_403, A[41], B[41]);
  nand g251 (n_404, A[41], n_402);
  nand g252 (n_405, B[41], n_402);
  nand g253 (n_407, n_403, n_404, n_405);
  xor g254 (n_406, A[41], B[41]);
  xor g255 (Z[41], n_402, n_406);
  nand g256 (n_408, A[42], B[42]);
  nand g257 (n_409, A[42], n_407);
  nand g258 (n_410, B[42], n_407);
  nand g259 (n_412, n_408, n_409, n_410);
  xor g260 (n_411, A[42], B[42]);
  xor g261 (Z[42], n_407, n_411);
  nand g262 (n_413, A[43], B[43]);
  nand g263 (n_414, A[43], n_412);
  nand g264 (n_415, B[43], n_412);
  nand g265 (n_417, n_413, n_414, n_415);
  xor g266 (n_416, A[43], B[43]);
  xor g267 (Z[43], n_412, n_416);
  nand g268 (n_418, A[44], B[44]);
  nand g269 (n_419, A[44], n_417);
  nand g270 (n_420, B[44], n_417);
  nand g271 (n_422, n_418, n_419, n_420);
  xor g272 (n_421, A[44], B[44]);
  xor g273 (Z[44], n_417, n_421);
  nand g274 (n_423, A[45], B[45]);
  nand g275 (n_424, A[45], n_422);
  nand g276 (n_425, B[45], n_422);
  nand g277 (n_427, n_423, n_424, n_425);
  xor g278 (n_426, A[45], B[45]);
  xor g279 (Z[45], n_422, n_426);
  nand g280 (n_428, A[46], B[46]);
  nand g281 (n_429, A[46], n_427);
  nand g282 (n_430, B[46], n_427);
  nand g283 (n_432, n_428, n_429, n_430);
  xor g284 (n_431, A[46], B[46]);
  xor g285 (Z[46], n_427, n_431);
  nand g286 (n_433, A[47], B[47]);
  nand g287 (n_434, A[47], n_432);
  nand g288 (n_435, B[47], n_432);
  nand g289 (n_437, n_433, n_434, n_435);
  xor g290 (n_436, A[47], B[47]);
  xor g291 (Z[47], n_432, n_436);
  nand g292 (n_438, A[48], B[48]);
  nand g293 (n_439, A[48], n_437);
  nand g294 (n_440, B[48], n_437);
  nand g295 (n_442, n_438, n_439, n_440);
  xor g296 (n_441, A[48], B[48]);
  xor g297 (Z[48], n_437, n_441);
  nand g298 (n_443, A[49], B[49]);
  nand g299 (n_444, A[49], n_442);
  nand g300 (n_445, B[49], n_442);
  nand g301 (n_447, n_443, n_444, n_445);
  xor g302 (n_446, A[49], B[49]);
  xor g303 (Z[49], n_442, n_446);
  nand g304 (n_448, A[50], B[50]);
  nand g305 (n_449, A[50], n_447);
  nand g306 (n_450, B[50], n_447);
  nand g307 (n_452, n_448, n_449, n_450);
  xor g308 (n_451, A[50], B[50]);
  xor g309 (Z[50], n_447, n_451);
  nand g310 (n_453, A[51], B[51]);
  nand g311 (n_454, A[51], n_452);
  nand g312 (n_455, B[51], n_452);
  nand g313 (n_457, n_453, n_454, n_455);
  xor g314 (n_456, A[51], B[51]);
  xor g315 (Z[51], n_452, n_456);
  nand g316 (n_458, A[52], B[52]);
  nand g317 (n_459, A[52], n_457);
  nand g318 (n_460, B[52], n_457);
  nand g319 (n_462, n_458, n_459, n_460);
  xor g320 (n_461, A[52], B[52]);
  xor g321 (Z[52], n_457, n_461);
  nand g322 (n_463, A[53], B[53]);
  nand g323 (n_464, A[53], n_462);
  nand g324 (n_465, B[53], n_462);
  nand g325 (n_467, n_463, n_464, n_465);
  xor g326 (n_466, A[53], B[53]);
  xor g327 (Z[53], n_462, n_466);
  nand g328 (n_468, A[54], B[54]);
  nand g329 (n_469, A[54], n_467);
  nand g330 (n_470, B[54], n_467);
  nand g331 (n_472, n_468, n_469, n_470);
  xor g332 (n_471, A[54], B[54]);
  xor g333 (Z[54], n_467, n_471);
  nand g334 (n_473, A[55], B[55]);
  nand g335 (n_474, A[55], n_472);
  nand g336 (n_475, B[55], n_472);
  nand g337 (n_477, n_473, n_474, n_475);
  xor g338 (n_476, A[55], B[55]);
  xor g339 (Z[55], n_472, n_476);
  nand g340 (n_478, A[56], B[56]);
  nand g341 (n_479, A[56], n_477);
  nand g342 (n_480, B[56], n_477);
  nand g343 (n_482, n_478, n_479, n_480);
  xor g344 (n_481, A[56], B[56]);
  xor g345 (Z[56], n_477, n_481);
  nand g346 (n_483, A[57], B[57]);
  nand g347 (n_484, A[57], n_482);
  nand g348 (n_485, B[57], n_482);
  nand g349 (n_487, n_483, n_484, n_485);
  xor g350 (n_486, A[57], B[57]);
  xor g351 (Z[57], n_482, n_486);
  nand g352 (n_488, A[58], B[58]);
  nand g353 (n_489, A[58], n_487);
  nand g354 (n_490, B[58], n_487);
  nand g355 (n_492, n_488, n_489, n_490);
  xor g356 (n_491, A[58], B[58]);
  xor g357 (Z[58], n_487, n_491);
  nand g358 (n_493, A[59], B[59]);
  nand g359 (n_494, A[59], n_492);
  nand g360 (n_495, B[59], n_492);
  nand g361 (n_497, n_493, n_494, n_495);
  xor g362 (n_496, A[59], B[59]);
  xor g363 (Z[59], n_492, n_496);
  nand g364 (n_498, A[60], B[60]);
  nand g365 (n_499, A[60], n_497);
  nand g366 (n_500, B[60], n_497);
  nand g367 (n_502, n_498, n_499, n_500);
  xor g368 (n_501, A[60], B[60]);
  xor g369 (Z[60], n_497, n_501);
  nand g370 (n_503, A[61], B[61]);
  nand g371 (n_504, A[61], n_502);
  nand g372 (n_505, B[61], n_502);
  nand g373 (n_507, n_503, n_504, n_505);
  xor g374 (n_506, A[61], B[61]);
  xor g375 (Z[61], n_502, n_506);
  nand g376 (n_508, A[62], B[62]);
  nand g377 (n_509, A[62], n_507);
  nand g378 (n_510, B[62], n_507);
  nand g379 (n_512, n_508, n_509, n_510);
  xor g380 (n_511, A[62], B[62]);
  xor g381 (Z[62], n_507, n_511);
  nand g385 (n_197, n_513, n_514, n_515);
  xor g387 (Z[63], n_512, n_516);
  or g389 (n_513, A[63], B[63]);
  xor g390 (n_516, A[63], B[63]);
  or g391 (n_204, wc, n_198);
  not gc (wc, A[1]);
  or g392 (n_205, wc0, n_198);
  not gc0 (wc0, B[1]);
  xnor g393 (Z[1], n_198, n_206);
  or g394 (n_514, A[63], wc1);
  not gc1 (wc1, n_512);
  or g395 (n_515, B[63], wc2);
  not gc2 (wc2, n_512);
endmodule

module add_signed_3032_GENERIC(A, B, Z);
  input [63:0] A, B;
  output [64:0] Z;
  wire [63:0] A, B;
  wire [64:0] Z;
  add_signed_3032_GENERIC_REAL g1(.A ({A[63:2], A[0], A[0]}), .B (B),
       .Z (Z));
endmodule

module add_signed_3032_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [63:0] A, B;
  output [64:0] Z;
  wire [63:0] A, B;
  wire [64:0] Z;
  wire n_197, n_198, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516;
  not g3 (Z[64], n_197);
  nand g4 (n_198, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_203, A[1], B[1]);
  nand g13 (n_207, n_203, n_204, n_205);
  xor g14 (n_206, A[1], B[1]);
  nand g16 (n_208, A[2], B[2]);
  nand g17 (n_209, A[2], n_207);
  nand g18 (n_210, B[2], n_207);
  nand g19 (n_212, n_208, n_209, n_210);
  xor g20 (n_211, A[2], B[2]);
  xor g21 (Z[2], n_207, n_211);
  nand g22 (n_213, A[3], B[3]);
  nand g23 (n_214, A[3], n_212);
  nand g24 (n_215, B[3], n_212);
  nand g25 (n_217, n_213, n_214, n_215);
  xor g26 (n_216, A[3], B[3]);
  xor g27 (Z[3], n_212, n_216);
  nand g28 (n_218, A[4], B[4]);
  nand g29 (n_219, A[4], n_217);
  nand g30 (n_220, B[4], n_217);
  nand g31 (n_222, n_218, n_219, n_220);
  xor g32 (n_221, A[4], B[4]);
  xor g33 (Z[4], n_217, n_221);
  nand g34 (n_223, A[5], B[5]);
  nand g35 (n_224, A[5], n_222);
  nand g36 (n_225, B[5], n_222);
  nand g37 (n_227, n_223, n_224, n_225);
  xor g38 (n_226, A[5], B[5]);
  xor g39 (Z[5], n_222, n_226);
  nand g40 (n_228, A[6], B[6]);
  nand g41 (n_229, A[6], n_227);
  nand g42 (n_230, B[6], n_227);
  nand g43 (n_232, n_228, n_229, n_230);
  xor g44 (n_231, A[6], B[6]);
  xor g45 (Z[6], n_227, n_231);
  nand g46 (n_233, A[7], B[7]);
  nand g47 (n_234, A[7], n_232);
  nand g48 (n_235, B[7], n_232);
  nand g49 (n_237, n_233, n_234, n_235);
  xor g50 (n_236, A[7], B[7]);
  xor g51 (Z[7], n_232, n_236);
  nand g52 (n_238, A[8], B[8]);
  nand g53 (n_239, A[8], n_237);
  nand g54 (n_240, B[8], n_237);
  nand g55 (n_242, n_238, n_239, n_240);
  xor g56 (n_241, A[8], B[8]);
  xor g57 (Z[8], n_237, n_241);
  nand g58 (n_243, A[9], B[9]);
  nand g59 (n_244, A[9], n_242);
  nand g60 (n_245, B[9], n_242);
  nand g61 (n_247, n_243, n_244, n_245);
  xor g62 (n_246, A[9], B[9]);
  xor g63 (Z[9], n_242, n_246);
  nand g64 (n_248, A[10], B[10]);
  nand g65 (n_249, A[10], n_247);
  nand g66 (n_250, B[10], n_247);
  nand g67 (n_252, n_248, n_249, n_250);
  xor g68 (n_251, A[10], B[10]);
  xor g69 (Z[10], n_247, n_251);
  nand g70 (n_253, A[11], B[11]);
  nand g71 (n_254, A[11], n_252);
  nand g72 (n_255, B[11], n_252);
  nand g73 (n_257, n_253, n_254, n_255);
  xor g74 (n_256, A[11], B[11]);
  xor g75 (Z[11], n_252, n_256);
  nand g76 (n_258, A[12], B[12]);
  nand g77 (n_259, A[12], n_257);
  nand g78 (n_260, B[12], n_257);
  nand g79 (n_262, n_258, n_259, n_260);
  xor g80 (n_261, A[12], B[12]);
  xor g81 (Z[12], n_257, n_261);
  nand g82 (n_263, A[13], B[13]);
  nand g83 (n_264, A[13], n_262);
  nand g84 (n_265, B[13], n_262);
  nand g85 (n_267, n_263, n_264, n_265);
  xor g86 (n_266, A[13], B[13]);
  xor g87 (Z[13], n_262, n_266);
  nand g88 (n_268, A[14], B[14]);
  nand g89 (n_269, A[14], n_267);
  nand g90 (n_270, B[14], n_267);
  nand g91 (n_272, n_268, n_269, n_270);
  xor g92 (n_271, A[14], B[14]);
  xor g93 (Z[14], n_267, n_271);
  nand g94 (n_273, A[15], B[15]);
  nand g95 (n_274, A[15], n_272);
  nand g96 (n_275, B[15], n_272);
  nand g97 (n_277, n_273, n_274, n_275);
  xor g98 (n_276, A[15], B[15]);
  xor g99 (Z[15], n_272, n_276);
  nand g100 (n_278, A[16], B[16]);
  nand g101 (n_279, A[16], n_277);
  nand g102 (n_280, B[16], n_277);
  nand g103 (n_282, n_278, n_279, n_280);
  xor g104 (n_281, A[16], B[16]);
  xor g105 (Z[16], n_277, n_281);
  nand g106 (n_283, A[17], B[17]);
  nand g107 (n_284, A[17], n_282);
  nand g108 (n_285, B[17], n_282);
  nand g109 (n_287, n_283, n_284, n_285);
  xor g110 (n_286, A[17], B[17]);
  xor g111 (Z[17], n_282, n_286);
  nand g112 (n_288, A[18], B[18]);
  nand g113 (n_289, A[18], n_287);
  nand g114 (n_290, B[18], n_287);
  nand g115 (n_292, n_288, n_289, n_290);
  xor g116 (n_291, A[18], B[18]);
  xor g117 (Z[18], n_287, n_291);
  nand g118 (n_293, A[19], B[19]);
  nand g119 (n_294, A[19], n_292);
  nand g120 (n_295, B[19], n_292);
  nand g121 (n_297, n_293, n_294, n_295);
  xor g122 (n_296, A[19], B[19]);
  xor g123 (Z[19], n_292, n_296);
  nand g124 (n_298, A[20], B[20]);
  nand g125 (n_299, A[20], n_297);
  nand g126 (n_300, B[20], n_297);
  nand g127 (n_302, n_298, n_299, n_300);
  xor g128 (n_301, A[20], B[20]);
  xor g129 (Z[20], n_297, n_301);
  nand g130 (n_303, A[21], B[21]);
  nand g131 (n_304, A[21], n_302);
  nand g132 (n_305, B[21], n_302);
  nand g133 (n_307, n_303, n_304, n_305);
  xor g134 (n_306, A[21], B[21]);
  xor g135 (Z[21], n_302, n_306);
  nand g136 (n_308, A[22], B[22]);
  nand g137 (n_309, A[22], n_307);
  nand g138 (n_310, B[22], n_307);
  nand g139 (n_312, n_308, n_309, n_310);
  xor g140 (n_311, A[22], B[22]);
  xor g141 (Z[22], n_307, n_311);
  nand g142 (n_313, A[23], B[23]);
  nand g143 (n_314, A[23], n_312);
  nand g144 (n_315, B[23], n_312);
  nand g145 (n_317, n_313, n_314, n_315);
  xor g146 (n_316, A[23], B[23]);
  xor g147 (Z[23], n_312, n_316);
  nand g148 (n_318, A[24], B[24]);
  nand g149 (n_319, A[24], n_317);
  nand g150 (n_320, B[24], n_317);
  nand g151 (n_322, n_318, n_319, n_320);
  xor g152 (n_321, A[24], B[24]);
  xor g153 (Z[24], n_317, n_321);
  nand g154 (n_323, A[25], B[25]);
  nand g155 (n_324, A[25], n_322);
  nand g156 (n_325, B[25], n_322);
  nand g157 (n_327, n_323, n_324, n_325);
  xor g158 (n_326, A[25], B[25]);
  xor g159 (Z[25], n_322, n_326);
  nand g160 (n_328, A[26], B[26]);
  nand g161 (n_329, A[26], n_327);
  nand g162 (n_330, B[26], n_327);
  nand g163 (n_332, n_328, n_329, n_330);
  xor g164 (n_331, A[26], B[26]);
  xor g165 (Z[26], n_327, n_331);
  nand g166 (n_333, A[27], B[27]);
  nand g167 (n_334, A[27], n_332);
  nand g168 (n_335, B[27], n_332);
  nand g169 (n_337, n_333, n_334, n_335);
  xor g170 (n_336, A[27], B[27]);
  xor g171 (Z[27], n_332, n_336);
  nand g172 (n_338, A[28], B[28]);
  nand g173 (n_339, A[28], n_337);
  nand g174 (n_340, B[28], n_337);
  nand g175 (n_342, n_338, n_339, n_340);
  xor g176 (n_341, A[28], B[28]);
  xor g177 (Z[28], n_337, n_341);
  nand g178 (n_343, A[29], B[29]);
  nand g179 (n_344, A[29], n_342);
  nand g180 (n_345, B[29], n_342);
  nand g181 (n_347, n_343, n_344, n_345);
  xor g182 (n_346, A[29], B[29]);
  xor g183 (Z[29], n_342, n_346);
  nand g184 (n_348, A[30], B[30]);
  nand g185 (n_349, A[30], n_347);
  nand g186 (n_350, B[30], n_347);
  nand g187 (n_352, n_348, n_349, n_350);
  xor g188 (n_351, A[30], B[30]);
  xor g189 (Z[30], n_347, n_351);
  nand g190 (n_353, A[31], B[31]);
  nand g191 (n_354, A[31], n_352);
  nand g192 (n_355, B[31], n_352);
  nand g193 (n_357, n_353, n_354, n_355);
  xor g194 (n_356, A[31], B[31]);
  xor g195 (Z[31], n_352, n_356);
  nand g196 (n_358, A[32], B[32]);
  nand g197 (n_359, A[32], n_357);
  nand g198 (n_360, B[32], n_357);
  nand g199 (n_362, n_358, n_359, n_360);
  xor g200 (n_361, A[32], B[32]);
  xor g201 (Z[32], n_357, n_361);
  nand g202 (n_363, A[33], B[33]);
  nand g203 (n_364, A[33], n_362);
  nand g204 (n_365, B[33], n_362);
  nand g205 (n_367, n_363, n_364, n_365);
  xor g206 (n_366, A[33], B[33]);
  xor g207 (Z[33], n_362, n_366);
  nand g208 (n_368, A[34], B[34]);
  nand g209 (n_369, A[34], n_367);
  nand g210 (n_370, B[34], n_367);
  nand g211 (n_372, n_368, n_369, n_370);
  xor g212 (n_371, A[34], B[34]);
  xor g213 (Z[34], n_367, n_371);
  nand g214 (n_373, A[35], B[35]);
  nand g215 (n_374, A[35], n_372);
  nand g216 (n_375, B[35], n_372);
  nand g217 (n_377, n_373, n_374, n_375);
  xor g218 (n_376, A[35], B[35]);
  xor g219 (Z[35], n_372, n_376);
  nand g220 (n_378, A[36], B[36]);
  nand g221 (n_379, A[36], n_377);
  nand g222 (n_380, B[36], n_377);
  nand g223 (n_382, n_378, n_379, n_380);
  xor g224 (n_381, A[36], B[36]);
  xor g225 (Z[36], n_377, n_381);
  nand g226 (n_383, A[37], B[37]);
  nand g227 (n_384, A[37], n_382);
  nand g228 (n_385, B[37], n_382);
  nand g229 (n_387, n_383, n_384, n_385);
  xor g230 (n_386, A[37], B[37]);
  xor g231 (Z[37], n_382, n_386);
  nand g232 (n_388, A[38], B[38]);
  nand g233 (n_389, A[38], n_387);
  nand g234 (n_390, B[38], n_387);
  nand g235 (n_392, n_388, n_389, n_390);
  xor g236 (n_391, A[38], B[38]);
  xor g237 (Z[38], n_387, n_391);
  nand g238 (n_393, A[39], B[39]);
  nand g239 (n_394, A[39], n_392);
  nand g240 (n_395, B[39], n_392);
  nand g241 (n_397, n_393, n_394, n_395);
  xor g242 (n_396, A[39], B[39]);
  xor g243 (Z[39], n_392, n_396);
  nand g244 (n_398, A[40], B[40]);
  nand g245 (n_399, A[40], n_397);
  nand g246 (n_400, B[40], n_397);
  nand g247 (n_402, n_398, n_399, n_400);
  xor g248 (n_401, A[40], B[40]);
  xor g249 (Z[40], n_397, n_401);
  nand g250 (n_403, A[41], B[41]);
  nand g251 (n_404, A[41], n_402);
  nand g252 (n_405, B[41], n_402);
  nand g253 (n_407, n_403, n_404, n_405);
  xor g254 (n_406, A[41], B[41]);
  xor g255 (Z[41], n_402, n_406);
  nand g256 (n_408, A[42], B[42]);
  nand g257 (n_409, A[42], n_407);
  nand g258 (n_410, B[42], n_407);
  nand g259 (n_412, n_408, n_409, n_410);
  xor g260 (n_411, A[42], B[42]);
  xor g261 (Z[42], n_407, n_411);
  nand g262 (n_413, A[43], B[43]);
  nand g263 (n_414, A[43], n_412);
  nand g264 (n_415, B[43], n_412);
  nand g265 (n_417, n_413, n_414, n_415);
  xor g266 (n_416, A[43], B[43]);
  xor g267 (Z[43], n_412, n_416);
  nand g268 (n_418, A[44], B[44]);
  nand g269 (n_419, A[44], n_417);
  nand g270 (n_420, B[44], n_417);
  nand g271 (n_422, n_418, n_419, n_420);
  xor g272 (n_421, A[44], B[44]);
  xor g273 (Z[44], n_417, n_421);
  nand g274 (n_423, A[45], B[45]);
  nand g275 (n_424, A[45], n_422);
  nand g276 (n_425, B[45], n_422);
  nand g277 (n_427, n_423, n_424, n_425);
  xor g278 (n_426, A[45], B[45]);
  xor g279 (Z[45], n_422, n_426);
  nand g280 (n_428, A[46], B[46]);
  nand g281 (n_429, A[46], n_427);
  nand g282 (n_430, B[46], n_427);
  nand g283 (n_432, n_428, n_429, n_430);
  xor g284 (n_431, A[46], B[46]);
  xor g285 (Z[46], n_427, n_431);
  nand g286 (n_433, A[47], B[47]);
  nand g287 (n_434, A[47], n_432);
  nand g288 (n_435, B[47], n_432);
  nand g289 (n_437, n_433, n_434, n_435);
  xor g290 (n_436, A[47], B[47]);
  xor g291 (Z[47], n_432, n_436);
  nand g292 (n_438, A[48], B[48]);
  nand g293 (n_439, A[48], n_437);
  nand g294 (n_440, B[48], n_437);
  nand g295 (n_442, n_438, n_439, n_440);
  xor g296 (n_441, A[48], B[48]);
  xor g297 (Z[48], n_437, n_441);
  nand g298 (n_443, A[49], B[49]);
  nand g299 (n_444, A[49], n_442);
  nand g300 (n_445, B[49], n_442);
  nand g301 (n_447, n_443, n_444, n_445);
  xor g302 (n_446, A[49], B[49]);
  xor g303 (Z[49], n_442, n_446);
  nand g304 (n_448, A[50], B[50]);
  nand g305 (n_449, A[50], n_447);
  nand g306 (n_450, B[50], n_447);
  nand g307 (n_452, n_448, n_449, n_450);
  xor g308 (n_451, A[50], B[50]);
  xor g309 (Z[50], n_447, n_451);
  nand g310 (n_453, A[51], B[51]);
  nand g311 (n_454, A[51], n_452);
  nand g312 (n_455, B[51], n_452);
  nand g313 (n_457, n_453, n_454, n_455);
  xor g314 (n_456, A[51], B[51]);
  xor g315 (Z[51], n_452, n_456);
  nand g316 (n_458, A[52], B[52]);
  nand g317 (n_459, A[52], n_457);
  nand g318 (n_460, B[52], n_457);
  nand g319 (n_462, n_458, n_459, n_460);
  xor g320 (n_461, A[52], B[52]);
  xor g321 (Z[52], n_457, n_461);
  nand g322 (n_463, A[53], B[53]);
  nand g323 (n_464, A[53], n_462);
  nand g324 (n_465, B[53], n_462);
  nand g325 (n_467, n_463, n_464, n_465);
  xor g326 (n_466, A[53], B[53]);
  xor g327 (Z[53], n_462, n_466);
  nand g328 (n_468, A[54], B[54]);
  nand g329 (n_469, A[54], n_467);
  nand g330 (n_470, B[54], n_467);
  nand g331 (n_472, n_468, n_469, n_470);
  xor g332 (n_471, A[54], B[54]);
  xor g333 (Z[54], n_467, n_471);
  nand g334 (n_473, A[55], B[55]);
  nand g335 (n_474, A[55], n_472);
  nand g336 (n_475, B[55], n_472);
  nand g337 (n_477, n_473, n_474, n_475);
  xor g338 (n_476, A[55], B[55]);
  xor g339 (Z[55], n_472, n_476);
  nand g340 (n_478, A[56], B[56]);
  nand g341 (n_479, A[56], n_477);
  nand g342 (n_480, B[56], n_477);
  nand g343 (n_482, n_478, n_479, n_480);
  xor g344 (n_481, A[56], B[56]);
  xor g345 (Z[56], n_477, n_481);
  nand g346 (n_483, A[57], B[57]);
  nand g347 (n_484, A[57], n_482);
  nand g348 (n_485, B[57], n_482);
  nand g349 (n_487, n_483, n_484, n_485);
  xor g350 (n_486, A[57], B[57]);
  xor g351 (Z[57], n_482, n_486);
  nand g352 (n_488, A[58], B[58]);
  nand g353 (n_489, A[58], n_487);
  nand g354 (n_490, B[58], n_487);
  nand g355 (n_492, n_488, n_489, n_490);
  xor g356 (n_491, A[58], B[58]);
  xor g357 (Z[58], n_487, n_491);
  nand g358 (n_493, A[59], B[59]);
  nand g359 (n_494, A[59], n_492);
  nand g360 (n_495, B[59], n_492);
  nand g361 (n_497, n_493, n_494, n_495);
  xor g362 (n_496, A[59], B[59]);
  xor g363 (Z[59], n_492, n_496);
  nand g364 (n_498, A[60], B[60]);
  nand g365 (n_499, A[60], n_497);
  nand g366 (n_500, B[60], n_497);
  nand g367 (n_502, n_498, n_499, n_500);
  xor g368 (n_501, A[60], B[60]);
  xor g369 (Z[60], n_497, n_501);
  nand g370 (n_503, A[61], B[61]);
  nand g371 (n_504, A[61], n_502);
  nand g372 (n_505, B[61], n_502);
  nand g373 (n_507, n_503, n_504, n_505);
  xor g374 (n_506, A[61], B[61]);
  xor g375 (Z[61], n_502, n_506);
  nand g376 (n_508, A[62], B[62]);
  nand g377 (n_509, A[62], n_507);
  nand g378 (n_510, B[62], n_507);
  nand g379 (n_512, n_508, n_509, n_510);
  xor g380 (n_511, A[62], B[62]);
  xor g381 (Z[62], n_507, n_511);
  nand g385 (n_197, n_513, n_514, n_515);
  xor g387 (Z[63], n_512, n_516);
  or g389 (n_513, A[63], B[63]);
  xor g390 (n_516, A[63], B[63]);
  or g391 (n_204, wc, n_198);
  not gc (wc, A[1]);
  or g392 (n_205, wc0, n_198);
  not gc0 (wc0, B[1]);
  xnor g393 (Z[1], n_198, n_206);
  or g394 (n_514, A[63], wc1);
  not gc1 (wc1, n_512);
  or g395 (n_515, B[63], wc2);
  not gc2 (wc2, n_512);
endmodule

module add_signed_3032_1_GENERIC(A, B, Z);
  input [63:0] A, B;
  output [64:0] Z;
  wire [63:0] A, B;
  wire [64:0] Z;
  add_signed_3032_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_342_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [47:0] A, B;
  output [48:0] Z;
  wire [47:0] A, B;
  wire [48:0] Z;
  wire n_149, n_150, n_153, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_163, n_164, n_165, n_166, n_167, n_169, n_170;
  wire n_171, n_172, n_173, n_175, n_176, n_177, n_178, n_179;
  wire n_181, n_182, n_183, n_184, n_185, n_187, n_188, n_189;
  wire n_190, n_191, n_193, n_194, n_195, n_196, n_197, n_199;
  wire n_200, n_201, n_202, n_203, n_205, n_206, n_207, n_208;
  wire n_209, n_211, n_212, n_213, n_214, n_215, n_217, n_218;
  wire n_219, n_220, n_221, n_223, n_224, n_225, n_226, n_227;
  wire n_229, n_230, n_231, n_232, n_233, n_235, n_236, n_237;
  wire n_238, n_239, n_241, n_242, n_243, n_244, n_245, n_247;
  wire n_248, n_249, n_250, n_251, n_253, n_254, n_255, n_256;
  wire n_257, n_259, n_260, n_261, n_262, n_263, n_265, n_266;
  wire n_267, n_268, n_269, n_271, n_272, n_273, n_274, n_275;
  wire n_277, n_278, n_279, n_280, n_281, n_283, n_284, n_285;
  wire n_286, n_287, n_289, n_290, n_291, n_292, n_293, n_295;
  wire n_296, n_298, n_299, n_300, n_301, n_302, n_303, n_305;
  wire n_307, n_309, n_310, n_312, n_313, n_315, n_317, n_319;
  wire n_320, n_322, n_323, n_325, n_327, n_329, n_330, n_332;
  wire n_333, n_335, n_337, n_339, n_340, n_342, n_343, n_345;
  wire n_347, n_349, n_350, n_352, n_353, n_355, n_357, n_359;
  wire n_360, n_362, n_363, n_365, n_367, n_369, n_370, n_372;
  wire n_373, n_375, n_377, n_379, n_380, n_382, n_383, n_385;
  wire n_387, n_389, n_390, n_392, n_393, n_395, n_397, n_399;
  wire n_400, n_402, n_403, n_405, n_407, n_409, n_410, n_412;
  wire n_414, n_415, n_416, n_418, n_419, n_420, n_422, n_423;
  wire n_424, n_425, n_427, n_429, n_431, n_432, n_433, n_435;
  wire n_436, n_437, n_439, n_440, n_442, n_444, n_446, n_447;
  wire n_448, n_450, n_451, n_452, n_454, n_455, n_457, n_459;
  wire n_461, n_462, n_463, n_465, n_466, n_467, n_469, n_470;
  wire n_472, n_474, n_476, n_477, n_478, n_480, n_481, n_482;
  wire n_484, n_485, n_487, n_489, n_491, n_492, n_493, n_495;
  wire n_496, n_497, n_499, n_501, n_502, n_503, n_505, n_506;
  wire n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515;
  wire n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_524;
  wire n_527, n_529, n_530, n_531, n_534, n_537, n_539, n_540;
  wire n_542, n_544, n_545, n_547, n_549, n_550, n_552, n_554;
  wire n_555, n_557, n_558, n_560, n_563, n_565, n_566, n_567;
  wire n_570, n_573, n_575, n_576, n_578, n_580, n_581, n_583;
  wire n_585, n_586, n_588, n_590, n_591, n_593, n_595, n_596;
  wire n_597, n_599, n_600, n_602, n_603, n_604, n_605, n_606;
  wire n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_615;
  wire n_616, n_617, n_619, n_620, n_621, n_623, n_624, n_625;
  wire n_627, n_628, n_629, n_631, n_632, n_633, n_635, n_636;
  wire n_637, n_639, n_640, n_641, n_643, n_644, n_645, n_647;
  wire n_648, n_649, n_651, n_652, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_675, n_676;
  wire n_677, n_679, n_680, n_681, n_683, n_684, n_685, n_687;
  wire n_688, n_689, n_691, n_692, n_693, n_695, n_696, n_697;
  wire n_698, n_700, n_701, n_702, n_704, n_705, n_706, n_707;
  wire n_709, n_710, n_711, n_713, n_714, n_715, n_716, n_718;
  wire n_719, n_721, n_722, n_724, n_725, n_726, n_727, n_729;
  wire n_730, n_731, n_733, n_734, n_735, n_736, n_738, n_739;
  wire n_741, n_742, n_744, n_745, n_746, n_747, n_749, n_750;
  wire n_751, n_752, n_754, n_755, n_756, n_757, n_759, n_760;
  wire n_762, n_763, n_765, n_766, n_767, n_768, n_770, n_771;
  wire n_772, n_774, n_775, n_776, n_777, n_779, n_780, n_782;
  wire n_783, n_785, n_786, n_787, n_788, n_790, n_791, n_792;
  wire n_793, n_795, n_796, n_797, n_798, n_800, n_801, n_803;
  wire n_804, n_806, n_807, n_808, n_809, n_811, n_812;
  not g3 (Z[48], n_149);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_150, A[0], B[0]);
  nor g9 (n_153, A[1], B[1]);
  nand g10 (n_156, A[1], B[1]);
  nor g11 (n_163, A[2], B[2]);
  nand g12 (n_158, A[2], B[2]);
  nor g13 (n_159, A[3], B[3]);
  nand g14 (n_160, A[3], B[3]);
  nor g15 (n_169, A[4], B[4]);
  nand g16 (n_164, A[4], B[4]);
  nor g17 (n_165, A[5], B[5]);
  nand g18 (n_166, A[5], B[5]);
  nor g19 (n_175, A[6], B[6]);
  nand g20 (n_170, A[6], B[6]);
  nor g21 (n_171, A[7], B[7]);
  nand g22 (n_172, A[7], B[7]);
  nor g23 (n_181, A[8], B[8]);
  nand g24 (n_176, A[8], B[8]);
  nor g25 (n_177, A[9], B[9]);
  nand g26 (n_178, A[9], B[9]);
  nor g27 (n_187, A[10], B[10]);
  nand g28 (n_182, A[10], B[10]);
  nor g29 (n_183, A[11], B[11]);
  nand g30 (n_184, A[11], B[11]);
  nor g31 (n_193, A[12], B[12]);
  nand g32 (n_188, A[12], B[12]);
  nor g33 (n_189, A[13], B[13]);
  nand g34 (n_190, A[13], B[13]);
  nor g35 (n_199, A[14], B[14]);
  nand g36 (n_194, A[14], B[14]);
  nor g37 (n_195, A[15], B[15]);
  nand g38 (n_196, A[15], B[15]);
  nor g39 (n_205, A[16], B[16]);
  nand g40 (n_200, A[16], B[16]);
  nor g41 (n_201, A[17], B[17]);
  nand g42 (n_202, A[17], B[17]);
  nor g43 (n_211, A[18], B[18]);
  nand g44 (n_206, A[18], B[18]);
  nor g45 (n_207, A[19], B[19]);
  nand g46 (n_208, A[19], B[19]);
  nor g47 (n_217, A[20], B[20]);
  nand g48 (n_212, A[20], B[20]);
  nor g49 (n_213, A[21], B[21]);
  nand g50 (n_214, A[21], B[21]);
  nor g51 (n_223, A[22], B[22]);
  nand g52 (n_218, A[22], B[22]);
  nor g53 (n_219, A[23], B[23]);
  nand g54 (n_220, A[23], B[23]);
  nor g55 (n_229, A[24], B[24]);
  nand g56 (n_224, A[24], B[24]);
  nor g57 (n_225, A[25], B[25]);
  nand g58 (n_226, A[25], B[25]);
  nor g59 (n_235, A[26], B[26]);
  nand g60 (n_230, A[26], B[26]);
  nor g61 (n_231, A[27], B[27]);
  nand g62 (n_232, A[27], B[27]);
  nor g63 (n_241, A[28], B[28]);
  nand g64 (n_236, A[28], B[28]);
  nor g65 (n_237, A[29], B[29]);
  nand g66 (n_238, A[29], B[29]);
  nor g67 (n_247, A[30], B[30]);
  nand g68 (n_242, A[30], B[30]);
  nor g69 (n_243, A[31], B[31]);
  nand g70 (n_244, A[31], B[31]);
  nor g71 (n_253, A[32], B[32]);
  nand g72 (n_248, A[32], B[32]);
  nor g73 (n_249, A[33], B[33]);
  nand g74 (n_250, A[33], B[33]);
  nor g75 (n_259, A[34], B[34]);
  nand g76 (n_254, A[34], B[34]);
  nor g77 (n_255, A[35], B[35]);
  nand g78 (n_256, A[35], B[35]);
  nor g79 (n_265, A[36], B[36]);
  nand g80 (n_260, A[36], B[36]);
  nor g81 (n_261, A[37], B[37]);
  nand g82 (n_262, A[37], B[37]);
  nor g83 (n_271, A[38], B[38]);
  nand g84 (n_266, A[38], B[38]);
  nor g85 (n_267, A[39], B[39]);
  nand g86 (n_268, A[39], B[39]);
  nor g87 (n_277, A[40], B[40]);
  nand g88 (n_272, A[40], B[40]);
  nor g89 (n_273, A[41], B[41]);
  nand g90 (n_274, A[41], B[41]);
  nor g91 (n_283, A[42], B[42]);
  nand g92 (n_278, A[42], B[42]);
  nor g93 (n_279, A[43], B[43]);
  nand g94 (n_280, A[43], B[43]);
  nor g95 (n_289, A[44], B[44]);
  nand g96 (n_284, A[44], B[44]);
  nor g97 (n_285, A[45], B[45]);
  nand g98 (n_286, A[45], B[45]);
  nor g99 (n_295, A[46], B[46]);
  nand g100 (n_290, A[46], B[46]);
  nand g105 (n_296, n_156, n_157);
  nor g106 (n_161, n_158, n_159);
  nor g109 (n_299, n_163, n_159);
  nor g110 (n_167, n_164, n_165);
  nor g113 (n_305, n_169, n_165);
  nor g114 (n_173, n_170, n_171);
  nor g117 (n_307, n_175, n_171);
  nor g118 (n_179, n_176, n_177);
  nor g121 (n_315, n_181, n_177);
  nor g122 (n_185, n_182, n_183);
  nor g125 (n_317, n_187, n_183);
  nor g126 (n_191, n_188, n_189);
  nor g129 (n_325, n_193, n_189);
  nor g130 (n_197, n_194, n_195);
  nor g133 (n_327, n_199, n_195);
  nor g134 (n_203, n_200, n_201);
  nor g137 (n_335, n_205, n_201);
  nor g138 (n_209, n_206, n_207);
  nor g141 (n_337, n_211, n_207);
  nor g142 (n_215, n_212, n_213);
  nor g145 (n_345, n_217, n_213);
  nor g146 (n_221, n_218, n_219);
  nor g149 (n_347, n_223, n_219);
  nor g150 (n_227, n_224, n_225);
  nor g153 (n_355, n_229, n_225);
  nor g154 (n_233, n_230, n_231);
  nor g157 (n_357, n_235, n_231);
  nor g158 (n_239, n_236, n_237);
  nor g161 (n_365, n_241, n_237);
  nor g162 (n_245, n_242, n_243);
  nor g165 (n_367, n_247, n_243);
  nor g166 (n_251, n_248, n_249);
  nor g169 (n_375, n_253, n_249);
  nor g170 (n_257, n_254, n_255);
  nor g173 (n_377, n_259, n_255);
  nor g174 (n_263, n_260, n_261);
  nor g177 (n_385, n_265, n_261);
  nor g178 (n_269, n_266, n_267);
  nor g181 (n_387, n_271, n_267);
  nor g182 (n_275, n_272, n_273);
  nor g185 (n_395, n_277, n_273);
  nor g186 (n_281, n_278, n_279);
  nor g189 (n_397, n_283, n_279);
  nor g190 (n_287, n_284, n_285);
  nor g193 (n_405, n_289, n_285);
  nor g194 (n_293, n_290, n_291);
  nor g197 (n_407, n_295, n_291);
  nand g200 (n_700, n_158, n_298);
  nand g201 (n_301, n_299, n_296);
  nand g202 (n_412, n_300, n_301);
  nor g203 (n_303, n_175, n_302);
  nand g212 (n_420, n_305, n_307);
  nor g213 (n_313, n_187, n_312);
  nand g222 (n_427, n_315, n_317);
  nor g223 (n_323, n_199, n_322);
  nand g232 (n_435, n_325, n_327);
  nor g233 (n_333, n_211, n_332);
  nand g242 (n_442, n_335, n_337);
  nor g243 (n_343, n_223, n_342);
  nand g252 (n_450, n_345, n_347);
  nor g253 (n_353, n_235, n_352);
  nand g262 (n_457, n_355, n_357);
  nor g263 (n_363, n_247, n_362);
  nand g272 (n_465, n_365, n_367);
  nor g273 (n_373, n_259, n_372);
  nand g282 (n_472, n_375, n_377);
  nor g283 (n_383, n_271, n_382);
  nand g292 (n_480, n_385, n_387);
  nor g293 (n_393, n_283, n_392);
  nand g302 (n_487, n_395, n_397);
  nor g303 (n_403, n_295, n_402);
  nand g312 (n_495, n_405, n_407);
  nand g315 (n_704, n_164, n_414);
  nand g316 (n_415, n_305, n_412);
  nand g317 (n_706, n_302, n_415);
  nand g320 (n_709, n_418, n_419);
  nand g323 (n_499, n_422, n_423);
  nor g324 (n_425, n_193, n_424);
  nor g327 (n_509, n_193, n_427);
  nor g333 (n_433, n_431, n_424);
  nor g336 (n_515, n_427, n_431);
  nor g337 (n_437, n_435, n_424);
  nor g340 (n_518, n_427, n_435);
  nor g341 (n_440, n_217, n_439);
  nor g344 (n_603, n_217, n_442);
  nor g350 (n_448, n_446, n_439);
  nor g353 (n_609, n_442, n_446);
  nor g354 (n_452, n_450, n_439);
  nor g357 (n_524, n_442, n_450);
  nor g358 (n_455, n_241, n_454);
  nor g361 (n_537, n_241, n_457);
  nor g367 (n_463, n_461, n_454);
  nor g370 (n_547, n_457, n_461);
  nor g371 (n_467, n_465, n_454);
  nor g374 (n_552, n_457, n_465);
  nor g375 (n_470, n_265, n_469);
  nor g378 (n_655, n_265, n_472);
  nor g384 (n_478, n_476, n_469);
  nor g387 (n_661, n_472, n_476);
  nor g388 (n_482, n_480, n_469);
  nor g391 (n_560, n_472, n_480);
  nor g392 (n_485, n_289, n_484);
  nor g395 (n_573, n_289, n_487);
  nor g401 (n_493, n_491, n_484);
  nor g404 (n_583, n_487, n_491);
  nor g405 (n_497, n_495, n_484);
  nor g408 (n_588, n_487, n_495);
  nand g411 (n_713, n_176, n_501);
  nand g412 (n_502, n_315, n_499);
  nand g413 (n_715, n_312, n_502);
  nand g416 (n_718, n_505, n_506);
  nand g419 (n_721, n_424, n_508);
  nand g420 (n_511, n_509, n_499);
  nand g421 (n_724, n_510, n_511);
  nand g422 (n_514, n_512, n_499);
  nand g423 (n_726, n_513, n_514);
  nand g424 (n_517, n_515, n_499);
  nand g425 (n_729, n_516, n_517);
  nand g426 (n_520, n_518, n_499);
  nand g427 (n_593, n_519, n_520);
  nor g428 (n_522, n_229, n_521);
  nand g437 (n_617, n_355, n_524);
  nor g438 (n_531, n_529, n_521);
  nor g443 (n_534, n_457, n_521);
  nand g452 (n_629, n_524, n_537);
  nand g457 (n_633, n_524, n_542);
  nand g462 (n_637, n_524, n_547);
  nand g467 (n_641, n_524, n_552);
  nor g468 (n_558, n_277, n_557);
  nand g477 (n_669, n_395, n_560);
  nor g478 (n_567, n_565, n_557);
  nor g483 (n_570, n_487, n_557);
  nand g492 (n_681, n_560, n_573);
  nand g497 (n_685, n_560, n_578);
  nand g502 (n_689, n_560, n_583);
  nand g507 (n_693, n_560, n_588);
  nand g510 (n_733, n_200, n_595);
  nand g511 (n_596, n_335, n_593);
  nand g512 (n_735, n_332, n_596);
  nand g515 (n_738, n_599, n_600);
  nand g518 (n_741, n_439, n_602);
  nand g519 (n_605, n_603, n_593);
  nand g520 (n_744, n_604, n_605);
  nand g521 (n_608, n_606, n_593);
  nand g522 (n_746, n_607, n_608);
  nand g523 (n_611, n_609, n_593);
  nand g524 (n_749, n_610, n_611);
  nand g525 (n_612, n_524, n_593);
  nand g526 (n_751, n_521, n_612);
  nand g529 (n_754, n_615, n_616);
  nand g532 (n_756, n_619, n_620);
  nand g535 (n_759, n_623, n_624);
  nand g538 (n_762, n_627, n_628);
  nand g541 (n_765, n_631, n_632);
  nand g544 (n_767, n_635, n_636);
  nand g547 (n_770, n_639, n_640);
  nand g550 (n_645, n_643, n_644);
  nand g553 (n_774, n_248, n_647);
  nand g554 (n_648, n_375, n_645);
  nand g555 (n_776, n_372, n_648);
  nand g558 (n_779, n_651, n_652);
  nand g561 (n_782, n_469, n_654);
  nand g562 (n_657, n_655, n_645);
  nand g563 (n_785, n_656, n_657);
  nand g564 (n_660, n_658, n_645);
  nand g565 (n_787, n_659, n_660);
  nand g566 (n_663, n_661, n_645);
  nand g567 (n_790, n_662, n_663);
  nand g568 (n_664, n_560, n_645);
  nand g569 (n_792, n_557, n_664);
  nand g572 (n_795, n_667, n_668);
  nand g575 (n_797, n_671, n_672);
  nand g578 (n_800, n_675, n_676);
  nand g581 (n_803, n_679, n_680);
  nand g584 (n_806, n_683, n_684);
  nand g587 (n_808, n_687, n_688);
  nand g590 (n_811, n_691, n_692);
  nand g593 (n_149, n_695, n_696);
  xnor g597 (Z[2], n_296, n_698);
  xnor g600 (Z[3], n_700, n_701);
  xnor g602 (Z[4], n_412, n_702);
  xnor g605 (Z[5], n_704, n_705);
  xnor g607 (Z[6], n_706, n_707);
  xnor g610 (Z[7], n_709, n_710);
  xnor g612 (Z[8], n_499, n_711);
  xnor g615 (Z[9], n_713, n_714);
  xnor g617 (Z[10], n_715, n_716);
  xnor g620 (Z[11], n_718, n_719);
  xnor g623 (Z[12], n_721, n_722);
  xnor g626 (Z[13], n_724, n_725);
  xnor g628 (Z[14], n_726, n_727);
  xnor g631 (Z[15], n_729, n_730);
  xnor g633 (Z[16], n_593, n_731);
  xnor g636 (Z[17], n_733, n_734);
  xnor g638 (Z[18], n_735, n_736);
  xnor g641 (Z[19], n_738, n_739);
  xnor g644 (Z[20], n_741, n_742);
  xnor g647 (Z[21], n_744, n_745);
  xnor g649 (Z[22], n_746, n_747);
  xnor g652 (Z[23], n_749, n_750);
  xnor g654 (Z[24], n_751, n_752);
  xnor g657 (Z[25], n_754, n_755);
  xnor g659 (Z[26], n_756, n_757);
  xnor g662 (Z[27], n_759, n_760);
  xnor g665 (Z[28], n_762, n_763);
  xnor g668 (Z[29], n_765, n_766);
  xnor g670 (Z[30], n_767, n_768);
  xnor g673 (Z[31], n_770, n_771);
  xnor g675 (Z[32], n_645, n_772);
  xnor g678 (Z[33], n_774, n_775);
  xnor g680 (Z[34], n_776, n_777);
  xnor g683 (Z[35], n_779, n_780);
  xnor g686 (Z[36], n_782, n_783);
  xnor g689 (Z[37], n_785, n_786);
  xnor g691 (Z[38], n_787, n_788);
  xnor g694 (Z[39], n_790, n_791);
  xnor g696 (Z[40], n_792, n_793);
  xnor g699 (Z[41], n_795, n_796);
  xnor g701 (Z[42], n_797, n_798);
  xnor g704 (Z[43], n_800, n_801);
  xnor g707 (Z[44], n_803, n_804);
  xnor g710 (Z[45], n_806, n_807);
  xnor g712 (Z[46], n_808, n_809);
  xnor g715 (Z[47], n_811, n_812);
  and g718 (n_291, A[47], B[47]);
  or g719 (n_292, A[47], B[47]);
  and g720 (n_372, wc, n_250);
  not gc (wc, n_251);
  and g721 (n_379, wc0, n_256);
  not gc0 (wc0, n_257);
  and g722 (n_382, wc1, n_262);
  not gc1 (wc1, n_263);
  and g723 (n_389, wc2, n_268);
  not gc2 (wc2, n_269);
  and g724 (n_392, wc3, n_274);
  not gc3 (wc3, n_275);
  and g725 (n_399, wc4, n_280);
  not gc4 (wc4, n_281);
  and g726 (n_402, wc5, n_286);
  not gc5 (wc5, n_287);
  and g727 (n_332, wc6, n_202);
  not gc6 (wc6, n_203);
  and g728 (n_339, wc7, n_208);
  not gc7 (wc7, n_209);
  and g729 (n_342, wc8, n_214);
  not gc8 (wc8, n_215);
  and g730 (n_349, wc9, n_220);
  not gc9 (wc9, n_221);
  and g731 (n_352, wc10, n_226);
  not gc10 (wc10, n_227);
  and g732 (n_359, wc11, n_232);
  not gc11 (wc11, n_233);
  and g733 (n_362, wc12, n_238);
  not gc12 (wc12, n_239);
  and g734 (n_369, wc13, n_244);
  not gc13 (wc13, n_245);
  and g735 (n_312, wc14, n_178);
  not gc14 (wc14, n_179);
  and g736 (n_319, wc15, n_184);
  not gc15 (wc15, n_185);
  and g737 (n_322, wc16, n_190);
  not gc16 (wc16, n_191);
  and g738 (n_329, wc17, n_196);
  not gc17 (wc17, n_197);
  and g739 (n_302, wc18, n_166);
  not gc18 (wc18, n_167);
  and g740 (n_309, wc19, n_172);
  not gc19 (wc19, n_173);
  and g741 (n_300, wc20, n_160);
  not gc20 (wc20, n_161);
  or g742 (n_157, n_150, n_153);
  or g743 (n_416, wc21, n_175);
  not gc21 (wc21, n_305);
  or g744 (n_503, wc22, n_187);
  not gc22 (wc22, n_315);
  or g745 (n_431, wc23, n_199);
  not gc23 (wc23, n_325);
  or g746 (n_597, wc24, n_211);
  not gc24 (wc24, n_335);
  or g747 (n_446, wc25, n_223);
  not gc25 (wc25, n_345);
  or g748 (n_529, wc26, n_235);
  not gc26 (wc26, n_355);
  or g749 (n_461, wc27, n_247);
  not gc27 (wc27, n_365);
  or g750 (n_649, wc28, n_259);
  not gc28 (wc28, n_375);
  or g751 (n_476, wc29, n_271);
  not gc29 (wc29, n_385);
  or g752 (n_565, wc30, n_283);
  not gc30 (wc30, n_395);
  or g753 (n_491, wc31, n_295);
  not gc31 (wc31, n_405);
  or g754 (n_697, wc32, n_153);
  not gc32 (wc32, n_156);
  or g755 (n_698, wc33, n_163);
  not gc33 (wc33, n_158);
  or g756 (n_701, wc34, n_159);
  not gc34 (wc34, n_160);
  or g757 (n_702, wc35, n_169);
  not gc35 (wc35, n_164);
  or g758 (n_705, wc36, n_165);
  not gc36 (wc36, n_166);
  or g759 (n_707, wc37, n_175);
  not gc37 (wc37, n_170);
  or g760 (n_710, wc38, n_171);
  not gc38 (wc38, n_172);
  or g761 (n_711, wc39, n_181);
  not gc39 (wc39, n_176);
  or g762 (n_714, wc40, n_177);
  not gc40 (wc40, n_178);
  or g763 (n_716, wc41, n_187);
  not gc41 (wc41, n_182);
  or g764 (n_719, wc42, n_183);
  not gc42 (wc42, n_184);
  or g765 (n_722, wc43, n_193);
  not gc43 (wc43, n_188);
  or g766 (n_725, wc44, n_189);
  not gc44 (wc44, n_190);
  or g767 (n_727, wc45, n_199);
  not gc45 (wc45, n_194);
  or g768 (n_730, wc46, n_195);
  not gc46 (wc46, n_196);
  or g769 (n_731, wc47, n_205);
  not gc47 (wc47, n_200);
  or g770 (n_734, wc48, n_201);
  not gc48 (wc48, n_202);
  or g771 (n_736, wc49, n_211);
  not gc49 (wc49, n_206);
  or g772 (n_739, wc50, n_207);
  not gc50 (wc50, n_208);
  or g773 (n_742, wc51, n_217);
  not gc51 (wc51, n_212);
  or g774 (n_745, wc52, n_213);
  not gc52 (wc52, n_214);
  or g775 (n_747, wc53, n_223);
  not gc53 (wc53, n_218);
  or g776 (n_750, wc54, n_219);
  not gc54 (wc54, n_220);
  or g777 (n_752, wc55, n_229);
  not gc55 (wc55, n_224);
  or g778 (n_755, wc56, n_225);
  not gc56 (wc56, n_226);
  or g779 (n_757, wc57, n_235);
  not gc57 (wc57, n_230);
  or g780 (n_760, wc58, n_231);
  not gc58 (wc58, n_232);
  or g781 (n_763, wc59, n_241);
  not gc59 (wc59, n_236);
  or g782 (n_766, wc60, n_237);
  not gc60 (wc60, n_238);
  or g783 (n_768, wc61, n_247);
  not gc61 (wc61, n_242);
  or g784 (n_771, wc62, n_243);
  not gc62 (wc62, n_244);
  or g785 (n_772, wc63, n_253);
  not gc63 (wc63, n_248);
  or g786 (n_775, wc64, n_249);
  not gc64 (wc64, n_250);
  or g787 (n_777, wc65, n_259);
  not gc65 (wc65, n_254);
  or g788 (n_780, wc66, n_255);
  not gc66 (wc66, n_256);
  or g789 (n_783, wc67, n_265);
  not gc67 (wc67, n_260);
  or g790 (n_786, wc68, n_261);
  not gc68 (wc68, n_262);
  or g791 (n_788, wc69, n_271);
  not gc69 (wc69, n_266);
  or g792 (n_791, wc70, n_267);
  not gc70 (wc70, n_268);
  or g793 (n_793, wc71, n_277);
  not gc71 (wc71, n_272);
  or g794 (n_796, wc72, n_273);
  not gc72 (wc72, n_274);
  or g795 (n_798, wc73, n_283);
  not gc73 (wc73, n_278);
  or g796 (n_801, wc74, n_279);
  not gc74 (wc74, n_280);
  or g797 (n_804, wc75, n_289);
  not gc75 (wc75, n_284);
  or g798 (n_807, wc76, n_285);
  not gc76 (wc76, n_286);
  or g799 (n_809, wc77, n_295);
  not gc77 (wc77, n_290);
  and g800 (n_380, wc78, n_377);
  not gc78 (wc78, n_372);
  and g801 (n_390, wc79, n_387);
  not gc79 (wc79, n_382);
  and g802 (n_400, wc80, n_397);
  not gc80 (wc80, n_392);
  and g803 (n_409, n_292, wc81);
  not gc81 (wc81, n_293);
  and g804 (n_340, wc82, n_337);
  not gc82 (wc82, n_332);
  and g805 (n_350, wc83, n_347);
  not gc83 (wc83, n_342);
  and g806 (n_360, wc84, n_357);
  not gc84 (wc84, n_352);
  and g807 (n_370, wc85, n_367);
  not gc85 (wc85, n_362);
  and g808 (n_320, wc86, n_317);
  not gc86 (wc86, n_312);
  and g809 (n_330, wc87, n_327);
  not gc87 (wc87, n_322);
  and g810 (n_310, wc88, n_307);
  not gc88 (wc88, n_302);
  and g811 (n_512, wc89, n_325);
  not gc89 (wc89, n_427);
  and g812 (n_606, wc90, n_345);
  not gc90 (wc90, n_442);
  and g813 (n_542, wc91, n_365);
  not gc91 (wc91, n_457);
  and g814 (n_658, wc92, n_385);
  not gc92 (wc92, n_472);
  and g815 (n_578, wc93, n_405);
  not gc93 (wc93, n_487);
  xor g816 (Z[1], n_150, n_697);
  or g817 (n_812, wc94, n_291);
  not gc94 (wc94, n_292);
  and g818 (n_469, wc95, n_379);
  not gc95 (wc95, n_380);
  and g819 (n_481, wc96, n_389);
  not gc96 (wc96, n_390);
  and g820 (n_484, wc97, n_399);
  not gc97 (wc97, n_400);
  and g821 (n_410, wc98, n_407);
  not gc98 (wc98, n_402);
  and g822 (n_439, wc99, n_339);
  not gc99 (wc99, n_340);
  and g823 (n_451, wc100, n_349);
  not gc100 (wc100, n_350);
  and g824 (n_454, wc101, n_359);
  not gc101 (wc101, n_360);
  and g825 (n_466, wc102, n_369);
  not gc102 (wc102, n_370);
  and g826 (n_424, wc103, n_319);
  not gc103 (wc103, n_320);
  and g827 (n_436, wc104, n_329);
  not gc104 (wc104, n_330);
  and g828 (n_422, wc105, n_309);
  not gc105 (wc105, n_310);
  or g829 (n_298, wc106, n_163);
  not gc106 (wc106, n_296);
  and g830 (n_418, wc107, n_170);
  not gc107 (wc107, n_303);
  and g831 (n_505, wc108, n_182);
  not gc108 (wc108, n_313);
  and g832 (n_432, wc109, n_194);
  not gc109 (wc109, n_323);
  and g833 (n_599, wc110, n_206);
  not gc110 (wc110, n_333);
  and g834 (n_447, wc111, n_218);
  not gc111 (wc111, n_343);
  and g835 (n_530, wc112, n_230);
  not gc112 (wc112, n_353);
  and g836 (n_462, wc113, n_242);
  not gc113 (wc113, n_363);
  and g837 (n_651, wc114, n_254);
  not gc114 (wc114, n_373);
  and g838 (n_477, wc115, n_266);
  not gc115 (wc115, n_383);
  and g839 (n_566, wc116, n_278);
  not gc116 (wc116, n_393);
  and g840 (n_492, wc117, n_290);
  not gc117 (wc117, n_403);
  or g841 (n_613, wc118, n_229);
  not gc118 (wc118, n_524);
  or g842 (n_621, n_529, wc119);
  not gc119 (wc119, n_524);
  or g843 (n_625, wc120, n_457);
  not gc120 (wc120, n_524);
  or g844 (n_665, wc121, n_277);
  not gc121 (wc121, n_560);
  or g845 (n_673, n_565, wc122);
  not gc122 (wc122, n_560);
  or g846 (n_677, wc123, n_487);
  not gc123 (wc123, n_560);
  and g847 (n_496, wc124, n_409);
  not gc124 (wc124, n_410);
  and g848 (n_429, wc125, n_325);
  not gc125 (wc125, n_424);
  and g849 (n_444, wc126, n_345);
  not gc126 (wc126, n_439);
  and g850 (n_459, wc127, n_365);
  not gc127 (wc127, n_454);
  and g851 (n_474, wc128, n_385);
  not gc128 (wc128, n_469);
  and g852 (n_489, wc129, n_405);
  not gc129 (wc129, n_484);
  and g853 (n_557, n_481, wc130);
  not gc130 (wc130, n_482);
  and g854 (n_521, n_451, wc131);
  not gc131 (wc131, n_452);
  and g855 (n_554, n_466, wc132);
  not gc132 (wc132, n_467);
  and g856 (n_519, n_436, wc133);
  not gc133 (wc133, n_437);
  or g857 (n_423, n_420, wc134);
  not gc134 (wc134, n_412);
  or g858 (n_414, wc135, n_169);
  not gc135 (wc135, n_412);
  or g859 (n_419, n_416, wc136);
  not gc136 (wc136, n_412);
  and g860 (n_510, wc137, n_188);
  not gc137 (wc137, n_425);
  and g861 (n_513, wc138, n_322);
  not gc138 (wc138, n_429);
  and g862 (n_516, n_432, wc139);
  not gc139 (wc139, n_433);
  and g863 (n_604, wc140, n_212);
  not gc140 (wc140, n_440);
  and g864 (n_607, wc141, n_342);
  not gc141 (wc141, n_444);
  and g865 (n_610, n_447, wc142);
  not gc142 (wc142, n_448);
  and g866 (n_539, wc143, n_236);
  not gc143 (wc143, n_455);
  and g867 (n_544, wc144, n_362);
  not gc144 (wc144, n_459);
  and g868 (n_549, n_462, wc145);
  not gc145 (wc145, n_463);
  and g869 (n_656, wc146, n_260);
  not gc146 (wc146, n_470);
  and g870 (n_659, wc147, n_382);
  not gc147 (wc147, n_474);
  and g871 (n_662, n_477, wc148);
  not gc148 (wc148, n_478);
  and g872 (n_575, wc149, n_284);
  not gc149 (wc149, n_485);
  and g873 (n_580, wc150, n_402);
  not gc150 (wc150, n_489);
  and g874 (n_585, n_492, wc151);
  not gc151 (wc151, n_493);
  and g875 (n_591, wc152, n_588);
  not gc152 (wc152, n_557);
  and g876 (n_590, n_496, wc153);
  not gc153 (wc153, n_497);
  and g877 (n_555, wc154, n_552);
  not gc154 (wc154, n_521);
  and g878 (n_527, wc155, n_355);
  not gc155 (wc155, n_521);
  and g879 (n_540, wc156, n_537);
  not gc156 (wc156, n_521);
  and g880 (n_545, wc157, n_542);
  not gc157 (wc157, n_521);
  and g881 (n_550, wc158, n_547);
  not gc158 (wc158, n_521);
  and g882 (n_563, wc159, n_395);
  not gc159 (wc159, n_557);
  and g883 (n_576, wc160, n_573);
  not gc160 (wc160, n_557);
  and g884 (n_581, wc161, n_578);
  not gc161 (wc161, n_557);
  and g885 (n_586, wc162, n_583);
  not gc162 (wc162, n_557);
  and g886 (n_643, wc163, n_554);
  not gc163 (wc163, n_555);
  or g887 (n_501, wc164, n_181);
  not gc164 (wc164, n_499);
  or g888 (n_506, n_503, wc165);
  not gc165 (wc165, n_499);
  or g889 (n_508, wc166, n_427);
  not gc166 (wc166, n_499);
  and g890 (n_615, wc167, n_224);
  not gc167 (wc167, n_522);
  and g891 (n_619, wc168, n_352);
  not gc168 (wc168, n_527);
  and g892 (n_623, n_530, wc169);
  not gc169 (wc169, n_531);
  and g893 (n_627, n_454, wc170);
  not gc170 (wc170, n_534);
  and g894 (n_631, wc171, n_539);
  not gc171 (wc171, n_540);
  and g895 (n_635, wc172, n_544);
  not gc172 (wc172, n_545);
  and g896 (n_639, wc173, n_549);
  not gc173 (wc173, n_550);
  and g897 (n_667, wc174, n_272);
  not gc174 (wc174, n_558);
  and g898 (n_671, wc175, n_392);
  not gc175 (wc175, n_563);
  and g899 (n_675, n_566, wc176);
  not gc176 (wc176, n_567);
  and g900 (n_679, n_484, wc177);
  not gc177 (wc177, n_570);
  and g901 (n_683, wc178, n_575);
  not gc178 (wc178, n_576);
  and g902 (n_687, wc179, n_580);
  not gc179 (wc179, n_581);
  and g903 (n_691, wc180, n_585);
  not gc180 (wc180, n_586);
  and g904 (n_695, n_590, wc181);
  not gc181 (wc181, n_591);
  or g905 (n_644, n_641, wc182);
  not gc182 (wc182, n_593);
  or g906 (n_595, wc183, n_205);
  not gc183 (wc183, n_593);
  or g907 (n_600, n_597, wc184);
  not gc184 (wc184, n_593);
  or g908 (n_602, wc185, n_442);
  not gc185 (wc185, n_593);
  or g909 (n_616, n_613, wc186);
  not gc186 (wc186, n_593);
  or g910 (n_620, n_617, wc187);
  not gc187 (wc187, n_593);
  or g911 (n_624, n_621, wc188);
  not gc188 (wc188, n_593);
  or g912 (n_628, n_625, wc189);
  not gc189 (wc189, n_593);
  or g913 (n_632, n_629, wc190);
  not gc190 (wc190, n_593);
  or g914 (n_636, n_633, wc191);
  not gc191 (wc191, n_593);
  or g915 (n_640, n_637, wc192);
  not gc192 (wc192, n_593);
  or g916 (n_696, wc193, n_693);
  not gc193 (wc193, n_645);
  or g917 (n_647, wc194, n_253);
  not gc194 (wc194, n_645);
  or g918 (n_652, n_649, wc195);
  not gc195 (wc195, n_645);
  or g919 (n_654, wc196, n_472);
  not gc196 (wc196, n_645);
  or g920 (n_668, n_665, wc197);
  not gc197 (wc197, n_645);
  or g921 (n_672, wc198, n_669);
  not gc198 (wc198, n_645);
  or g922 (n_676, n_673, wc199);
  not gc199 (wc199, n_645);
  or g923 (n_680, n_677, wc200);
  not gc200 (wc200, n_645);
  or g924 (n_684, wc201, n_681);
  not gc201 (wc201, n_645);
  or g925 (n_688, wc202, n_685);
  not gc202 (wc202, n_645);
  or g926 (n_692, wc203, n_689);
  not gc203 (wc203, n_645);
endmodule

module add_signed_342_GENERIC(A, B, Z);
  input [47:0] A, B;
  output [48:0] Z;
  wire [47:0] A, B;
  wire [48:0] Z;
  add_signed_342_GENERIC_REAL g1(.A ({A[46], A[46:0]}), .B ({B[46],
       B[46:0]}), .Z (Z));
endmodule

module add_signed_342_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [47:0] A, B;
  output [48:0] Z;
  wire [47:0] A, B;
  wire [48:0] Z;
  wire n_149, n_150, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388;
  not g3 (Z[48], n_149);
  nand g4 (n_150, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_155, A[1], B[1]);
  nand g13 (n_159, n_155, n_156, n_157);
  xor g14 (n_158, A[1], B[1]);
  nand g16 (n_160, A[2], B[2]);
  nand g17 (n_161, A[2], n_159);
  nand g18 (n_162, B[2], n_159);
  nand g19 (n_164, n_160, n_161, n_162);
  xor g20 (n_163, A[2], B[2]);
  xor g21 (Z[2], n_159, n_163);
  nand g22 (n_165, A[3], B[3]);
  nand g23 (n_166, A[3], n_164);
  nand g24 (n_167, B[3], n_164);
  nand g25 (n_169, n_165, n_166, n_167);
  xor g26 (n_168, A[3], B[3]);
  xor g27 (Z[3], n_164, n_168);
  nand g28 (n_170, A[4], B[4]);
  nand g29 (n_171, A[4], n_169);
  nand g30 (n_172, B[4], n_169);
  nand g31 (n_174, n_170, n_171, n_172);
  xor g32 (n_173, A[4], B[4]);
  xor g33 (Z[4], n_169, n_173);
  nand g34 (n_175, A[5], B[5]);
  nand g35 (n_176, A[5], n_174);
  nand g36 (n_177, B[5], n_174);
  nand g37 (n_179, n_175, n_176, n_177);
  xor g38 (n_178, A[5], B[5]);
  xor g39 (Z[5], n_174, n_178);
  nand g40 (n_180, A[6], B[6]);
  nand g41 (n_181, A[6], n_179);
  nand g42 (n_182, B[6], n_179);
  nand g43 (n_184, n_180, n_181, n_182);
  xor g44 (n_183, A[6], B[6]);
  xor g45 (Z[6], n_179, n_183);
  nand g46 (n_185, A[7], B[7]);
  nand g47 (n_186, A[7], n_184);
  nand g48 (n_187, B[7], n_184);
  nand g49 (n_189, n_185, n_186, n_187);
  xor g50 (n_188, A[7], B[7]);
  xor g51 (Z[7], n_184, n_188);
  nand g52 (n_190, A[8], B[8]);
  nand g53 (n_191, A[8], n_189);
  nand g54 (n_192, B[8], n_189);
  nand g55 (n_194, n_190, n_191, n_192);
  xor g56 (n_193, A[8], B[8]);
  xor g57 (Z[8], n_189, n_193);
  nand g58 (n_195, A[9], B[9]);
  nand g59 (n_196, A[9], n_194);
  nand g60 (n_197, B[9], n_194);
  nand g61 (n_199, n_195, n_196, n_197);
  xor g62 (n_198, A[9], B[9]);
  xor g63 (Z[9], n_194, n_198);
  nand g64 (n_200, A[10], B[10]);
  nand g65 (n_201, A[10], n_199);
  nand g66 (n_202, B[10], n_199);
  nand g67 (n_204, n_200, n_201, n_202);
  xor g68 (n_203, A[10], B[10]);
  xor g69 (Z[10], n_199, n_203);
  nand g70 (n_205, A[11], B[11]);
  nand g71 (n_206, A[11], n_204);
  nand g72 (n_207, B[11], n_204);
  nand g73 (n_209, n_205, n_206, n_207);
  xor g74 (n_208, A[11], B[11]);
  xor g75 (Z[11], n_204, n_208);
  nand g76 (n_210, A[12], B[12]);
  nand g77 (n_211, A[12], n_209);
  nand g78 (n_212, B[12], n_209);
  nand g79 (n_214, n_210, n_211, n_212);
  xor g80 (n_213, A[12], B[12]);
  xor g81 (Z[12], n_209, n_213);
  nand g82 (n_215, A[13], B[13]);
  nand g83 (n_216, A[13], n_214);
  nand g84 (n_217, B[13], n_214);
  nand g85 (n_219, n_215, n_216, n_217);
  xor g86 (n_218, A[13], B[13]);
  xor g87 (Z[13], n_214, n_218);
  nand g88 (n_220, A[14], B[14]);
  nand g89 (n_221, A[14], n_219);
  nand g90 (n_222, B[14], n_219);
  nand g91 (n_224, n_220, n_221, n_222);
  xor g92 (n_223, A[14], B[14]);
  xor g93 (Z[14], n_219, n_223);
  nand g94 (n_225, A[15], B[15]);
  nand g95 (n_226, A[15], n_224);
  nand g96 (n_227, B[15], n_224);
  nand g97 (n_229, n_225, n_226, n_227);
  xor g98 (n_228, A[15], B[15]);
  xor g99 (Z[15], n_224, n_228);
  nand g100 (n_230, A[16], B[16]);
  nand g101 (n_231, A[16], n_229);
  nand g102 (n_232, B[16], n_229);
  nand g103 (n_234, n_230, n_231, n_232);
  xor g104 (n_233, A[16], B[16]);
  xor g105 (Z[16], n_229, n_233);
  nand g106 (n_235, A[17], B[17]);
  nand g107 (n_236, A[17], n_234);
  nand g108 (n_237, B[17], n_234);
  nand g109 (n_239, n_235, n_236, n_237);
  xor g110 (n_238, A[17], B[17]);
  xor g111 (Z[17], n_234, n_238);
  nand g112 (n_240, A[18], B[18]);
  nand g113 (n_241, A[18], n_239);
  nand g114 (n_242, B[18], n_239);
  nand g115 (n_244, n_240, n_241, n_242);
  xor g116 (n_243, A[18], B[18]);
  xor g117 (Z[18], n_239, n_243);
  nand g118 (n_245, A[19], B[19]);
  nand g119 (n_246, A[19], n_244);
  nand g120 (n_247, B[19], n_244);
  nand g121 (n_249, n_245, n_246, n_247);
  xor g122 (n_248, A[19], B[19]);
  xor g123 (Z[19], n_244, n_248);
  nand g124 (n_250, A[20], B[20]);
  nand g125 (n_251, A[20], n_249);
  nand g126 (n_252, B[20], n_249);
  nand g127 (n_254, n_250, n_251, n_252);
  xor g128 (n_253, A[20], B[20]);
  xor g129 (Z[20], n_249, n_253);
  nand g130 (n_255, A[21], B[21]);
  nand g131 (n_256, A[21], n_254);
  nand g132 (n_257, B[21], n_254);
  nand g133 (n_259, n_255, n_256, n_257);
  xor g134 (n_258, A[21], B[21]);
  xor g135 (Z[21], n_254, n_258);
  nand g136 (n_260, A[22], B[22]);
  nand g137 (n_261, A[22], n_259);
  nand g138 (n_262, B[22], n_259);
  nand g139 (n_264, n_260, n_261, n_262);
  xor g140 (n_263, A[22], B[22]);
  xor g141 (Z[22], n_259, n_263);
  nand g142 (n_265, A[23], B[23]);
  nand g143 (n_266, A[23], n_264);
  nand g144 (n_267, B[23], n_264);
  nand g145 (n_269, n_265, n_266, n_267);
  xor g146 (n_268, A[23], B[23]);
  xor g147 (Z[23], n_264, n_268);
  nand g148 (n_270, A[24], B[24]);
  nand g149 (n_271, A[24], n_269);
  nand g150 (n_272, B[24], n_269);
  nand g151 (n_274, n_270, n_271, n_272);
  xor g152 (n_273, A[24], B[24]);
  xor g153 (Z[24], n_269, n_273);
  nand g154 (n_275, A[25], B[25]);
  nand g155 (n_276, A[25], n_274);
  nand g156 (n_277, B[25], n_274);
  nand g157 (n_279, n_275, n_276, n_277);
  xor g158 (n_278, A[25], B[25]);
  xor g159 (Z[25], n_274, n_278);
  nand g160 (n_280, A[26], B[26]);
  nand g161 (n_281, A[26], n_279);
  nand g162 (n_282, B[26], n_279);
  nand g163 (n_284, n_280, n_281, n_282);
  xor g164 (n_283, A[26], B[26]);
  xor g165 (Z[26], n_279, n_283);
  nand g166 (n_285, A[27], B[27]);
  nand g167 (n_286, A[27], n_284);
  nand g168 (n_287, B[27], n_284);
  nand g169 (n_289, n_285, n_286, n_287);
  xor g170 (n_288, A[27], B[27]);
  xor g171 (Z[27], n_284, n_288);
  nand g172 (n_290, A[28], B[28]);
  nand g173 (n_291, A[28], n_289);
  nand g174 (n_292, B[28], n_289);
  nand g175 (n_294, n_290, n_291, n_292);
  xor g176 (n_293, A[28], B[28]);
  xor g177 (Z[28], n_289, n_293);
  nand g178 (n_295, A[29], B[29]);
  nand g179 (n_296, A[29], n_294);
  nand g180 (n_297, B[29], n_294);
  nand g181 (n_299, n_295, n_296, n_297);
  xor g182 (n_298, A[29], B[29]);
  xor g183 (Z[29], n_294, n_298);
  nand g184 (n_300, A[30], B[30]);
  nand g185 (n_301, A[30], n_299);
  nand g186 (n_302, B[30], n_299);
  nand g187 (n_304, n_300, n_301, n_302);
  xor g188 (n_303, A[30], B[30]);
  xor g189 (Z[30], n_299, n_303);
  nand g190 (n_305, A[31], B[31]);
  nand g191 (n_306, A[31], n_304);
  nand g192 (n_307, B[31], n_304);
  nand g193 (n_309, n_305, n_306, n_307);
  xor g194 (n_308, A[31], B[31]);
  xor g195 (Z[31], n_304, n_308);
  nand g196 (n_310, A[32], B[32]);
  nand g197 (n_311, A[32], n_309);
  nand g198 (n_312, B[32], n_309);
  nand g199 (n_314, n_310, n_311, n_312);
  xor g200 (n_313, A[32], B[32]);
  xor g201 (Z[32], n_309, n_313);
  nand g202 (n_315, A[33], B[33]);
  nand g203 (n_316, A[33], n_314);
  nand g204 (n_317, B[33], n_314);
  nand g205 (n_319, n_315, n_316, n_317);
  xor g206 (n_318, A[33], B[33]);
  xor g207 (Z[33], n_314, n_318);
  nand g208 (n_320, A[34], B[34]);
  nand g209 (n_321, A[34], n_319);
  nand g210 (n_322, B[34], n_319);
  nand g211 (n_324, n_320, n_321, n_322);
  xor g212 (n_323, A[34], B[34]);
  xor g213 (Z[34], n_319, n_323);
  nand g214 (n_325, A[35], B[35]);
  nand g215 (n_326, A[35], n_324);
  nand g216 (n_327, B[35], n_324);
  nand g217 (n_329, n_325, n_326, n_327);
  xor g218 (n_328, A[35], B[35]);
  xor g219 (Z[35], n_324, n_328);
  nand g220 (n_330, A[36], B[36]);
  nand g221 (n_331, A[36], n_329);
  nand g222 (n_332, B[36], n_329);
  nand g223 (n_334, n_330, n_331, n_332);
  xor g224 (n_333, A[36], B[36]);
  xor g225 (Z[36], n_329, n_333);
  nand g226 (n_335, A[37], B[37]);
  nand g227 (n_336, A[37], n_334);
  nand g228 (n_337, B[37], n_334);
  nand g229 (n_339, n_335, n_336, n_337);
  xor g230 (n_338, A[37], B[37]);
  xor g231 (Z[37], n_334, n_338);
  nand g232 (n_340, A[38], B[38]);
  nand g233 (n_341, A[38], n_339);
  nand g234 (n_342, B[38], n_339);
  nand g235 (n_344, n_340, n_341, n_342);
  xor g236 (n_343, A[38], B[38]);
  xor g237 (Z[38], n_339, n_343);
  nand g238 (n_345, A[39], B[39]);
  nand g239 (n_346, A[39], n_344);
  nand g240 (n_347, B[39], n_344);
  nand g241 (n_349, n_345, n_346, n_347);
  xor g242 (n_348, A[39], B[39]);
  xor g243 (Z[39], n_344, n_348);
  nand g244 (n_350, A[40], B[40]);
  nand g245 (n_351, A[40], n_349);
  nand g246 (n_352, B[40], n_349);
  nand g247 (n_354, n_350, n_351, n_352);
  xor g248 (n_353, A[40], B[40]);
  xor g249 (Z[40], n_349, n_353);
  nand g250 (n_355, A[41], B[41]);
  nand g251 (n_356, A[41], n_354);
  nand g252 (n_357, B[41], n_354);
  nand g253 (n_359, n_355, n_356, n_357);
  xor g254 (n_358, A[41], B[41]);
  xor g255 (Z[41], n_354, n_358);
  nand g256 (n_360, A[42], B[42]);
  nand g257 (n_361, A[42], n_359);
  nand g258 (n_362, B[42], n_359);
  nand g259 (n_364, n_360, n_361, n_362);
  xor g260 (n_363, A[42], B[42]);
  xor g261 (Z[42], n_359, n_363);
  nand g262 (n_365, A[43], B[43]);
  nand g263 (n_366, A[43], n_364);
  nand g264 (n_367, B[43], n_364);
  nand g265 (n_369, n_365, n_366, n_367);
  xor g266 (n_368, A[43], B[43]);
  xor g267 (Z[43], n_364, n_368);
  nand g268 (n_370, A[44], B[44]);
  nand g269 (n_371, A[44], n_369);
  nand g270 (n_372, B[44], n_369);
  nand g271 (n_374, n_370, n_371, n_372);
  xor g272 (n_373, A[44], B[44]);
  xor g273 (Z[44], n_369, n_373);
  nand g274 (n_375, A[45], B[45]);
  nand g275 (n_376, A[45], n_374);
  nand g276 (n_377, B[45], n_374);
  nand g277 (n_379, n_375, n_376, n_377);
  xor g278 (n_378, A[45], B[45]);
  xor g279 (Z[45], n_374, n_378);
  nand g280 (n_380, A[46], B[46]);
  nand g281 (n_381, A[46], n_379);
  nand g282 (n_382, B[46], n_379);
  nand g283 (n_384, n_380, n_381, n_382);
  xor g284 (n_383, A[46], B[46]);
  xor g285 (Z[46], n_379, n_383);
  nand g289 (n_149, n_385, n_386, n_387);
  xor g291 (Z[47], n_384, n_388);
  or g293 (n_385, A[47], B[47]);
  xor g294 (n_388, A[47], B[47]);
  or g295 (n_156, wc, n_150);
  not gc (wc, A[1]);
  or g296 (n_157, wc0, n_150);
  not gc0 (wc0, B[1]);
  xnor g297 (Z[1], n_150, n_158);
  or g298 (n_386, A[47], wc1);
  not gc1 (wc1, n_384);
  or g299 (n_387, B[47], wc2);
  not gc2 (wc2, n_384);
endmodule

module add_signed_342_1_GENERIC(A, B, Z);
  input [47:0] A, B;
  output [48:0] Z;
  wire [47:0] A, B;
  wire [48:0] Z;
  add_signed_342_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_342_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [47:0] A, B;
  output [48:0] Z;
  wire [47:0] A, B;
  wire [48:0] Z;
  wire n_149, n_150, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388;
  not g3 (Z[48], n_149);
  nand g4 (n_150, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_155, A[1], B[1]);
  nand g13 (n_159, n_155, n_156, n_157);
  xor g14 (n_158, A[1], B[1]);
  nand g16 (n_160, A[2], B[2]);
  nand g17 (n_161, A[2], n_159);
  nand g18 (n_162, B[2], n_159);
  nand g19 (n_164, n_160, n_161, n_162);
  xor g20 (n_163, A[2], B[2]);
  xor g21 (Z[2], n_159, n_163);
  nand g22 (n_165, A[3], B[3]);
  nand g23 (n_166, A[3], n_164);
  nand g24 (n_167, B[3], n_164);
  nand g25 (n_169, n_165, n_166, n_167);
  xor g26 (n_168, A[3], B[3]);
  xor g27 (Z[3], n_164, n_168);
  nand g28 (n_170, A[4], B[4]);
  nand g29 (n_171, A[4], n_169);
  nand g30 (n_172, B[4], n_169);
  nand g31 (n_174, n_170, n_171, n_172);
  xor g32 (n_173, A[4], B[4]);
  xor g33 (Z[4], n_169, n_173);
  nand g34 (n_175, A[5], B[5]);
  nand g35 (n_176, A[5], n_174);
  nand g36 (n_177, B[5], n_174);
  nand g37 (n_179, n_175, n_176, n_177);
  xor g38 (n_178, A[5], B[5]);
  xor g39 (Z[5], n_174, n_178);
  nand g40 (n_180, A[6], B[6]);
  nand g41 (n_181, A[6], n_179);
  nand g42 (n_182, B[6], n_179);
  nand g43 (n_184, n_180, n_181, n_182);
  xor g44 (n_183, A[6], B[6]);
  xor g45 (Z[6], n_179, n_183);
  nand g46 (n_185, A[7], B[7]);
  nand g47 (n_186, A[7], n_184);
  nand g48 (n_187, B[7], n_184);
  nand g49 (n_189, n_185, n_186, n_187);
  xor g50 (n_188, A[7], B[7]);
  xor g51 (Z[7], n_184, n_188);
  nand g52 (n_190, A[8], B[8]);
  nand g53 (n_191, A[8], n_189);
  nand g54 (n_192, B[8], n_189);
  nand g55 (n_194, n_190, n_191, n_192);
  xor g56 (n_193, A[8], B[8]);
  xor g57 (Z[8], n_189, n_193);
  nand g58 (n_195, A[9], B[9]);
  nand g59 (n_196, A[9], n_194);
  nand g60 (n_197, B[9], n_194);
  nand g61 (n_199, n_195, n_196, n_197);
  xor g62 (n_198, A[9], B[9]);
  xor g63 (Z[9], n_194, n_198);
  nand g64 (n_200, A[10], B[10]);
  nand g65 (n_201, A[10], n_199);
  nand g66 (n_202, B[10], n_199);
  nand g67 (n_204, n_200, n_201, n_202);
  xor g68 (n_203, A[10], B[10]);
  xor g69 (Z[10], n_199, n_203);
  nand g70 (n_205, A[11], B[11]);
  nand g71 (n_206, A[11], n_204);
  nand g72 (n_207, B[11], n_204);
  nand g73 (n_209, n_205, n_206, n_207);
  xor g74 (n_208, A[11], B[11]);
  xor g75 (Z[11], n_204, n_208);
  nand g76 (n_210, A[12], B[12]);
  nand g77 (n_211, A[12], n_209);
  nand g78 (n_212, B[12], n_209);
  nand g79 (n_214, n_210, n_211, n_212);
  xor g80 (n_213, A[12], B[12]);
  xor g81 (Z[12], n_209, n_213);
  nand g82 (n_215, A[13], B[13]);
  nand g83 (n_216, A[13], n_214);
  nand g84 (n_217, B[13], n_214);
  nand g85 (n_219, n_215, n_216, n_217);
  xor g86 (n_218, A[13], B[13]);
  xor g87 (Z[13], n_214, n_218);
  nand g88 (n_220, A[14], B[14]);
  nand g89 (n_221, A[14], n_219);
  nand g90 (n_222, B[14], n_219);
  nand g91 (n_224, n_220, n_221, n_222);
  xor g92 (n_223, A[14], B[14]);
  xor g93 (Z[14], n_219, n_223);
  nand g94 (n_225, A[15], B[15]);
  nand g95 (n_226, A[15], n_224);
  nand g96 (n_227, B[15], n_224);
  nand g97 (n_229, n_225, n_226, n_227);
  xor g98 (n_228, A[15], B[15]);
  xor g99 (Z[15], n_224, n_228);
  nand g100 (n_230, A[16], B[16]);
  nand g101 (n_231, A[16], n_229);
  nand g102 (n_232, B[16], n_229);
  nand g103 (n_234, n_230, n_231, n_232);
  xor g104 (n_233, A[16], B[16]);
  xor g105 (Z[16], n_229, n_233);
  nand g106 (n_235, A[17], B[17]);
  nand g107 (n_236, A[17], n_234);
  nand g108 (n_237, B[17], n_234);
  nand g109 (n_239, n_235, n_236, n_237);
  xor g110 (n_238, A[17], B[17]);
  xor g111 (Z[17], n_234, n_238);
  nand g112 (n_240, A[18], B[18]);
  nand g113 (n_241, A[18], n_239);
  nand g114 (n_242, B[18], n_239);
  nand g115 (n_244, n_240, n_241, n_242);
  xor g116 (n_243, A[18], B[18]);
  xor g117 (Z[18], n_239, n_243);
  nand g118 (n_245, A[19], B[19]);
  nand g119 (n_246, A[19], n_244);
  nand g120 (n_247, B[19], n_244);
  nand g121 (n_249, n_245, n_246, n_247);
  xor g122 (n_248, A[19], B[19]);
  xor g123 (Z[19], n_244, n_248);
  nand g124 (n_250, A[20], B[20]);
  nand g125 (n_251, A[20], n_249);
  nand g126 (n_252, B[20], n_249);
  nand g127 (n_254, n_250, n_251, n_252);
  xor g128 (n_253, A[20], B[20]);
  xor g129 (Z[20], n_249, n_253);
  nand g130 (n_255, A[21], B[21]);
  nand g131 (n_256, A[21], n_254);
  nand g132 (n_257, B[21], n_254);
  nand g133 (n_259, n_255, n_256, n_257);
  xor g134 (n_258, A[21], B[21]);
  xor g135 (Z[21], n_254, n_258);
  nand g136 (n_260, A[22], B[22]);
  nand g137 (n_261, A[22], n_259);
  nand g138 (n_262, B[22], n_259);
  nand g139 (n_264, n_260, n_261, n_262);
  xor g140 (n_263, A[22], B[22]);
  xor g141 (Z[22], n_259, n_263);
  nand g142 (n_265, A[23], B[23]);
  nand g143 (n_266, A[23], n_264);
  nand g144 (n_267, B[23], n_264);
  nand g145 (n_269, n_265, n_266, n_267);
  xor g146 (n_268, A[23], B[23]);
  xor g147 (Z[23], n_264, n_268);
  nand g148 (n_270, A[24], B[24]);
  nand g149 (n_271, A[24], n_269);
  nand g150 (n_272, B[24], n_269);
  nand g151 (n_274, n_270, n_271, n_272);
  xor g152 (n_273, A[24], B[24]);
  xor g153 (Z[24], n_269, n_273);
  nand g154 (n_275, A[25], B[25]);
  nand g155 (n_276, A[25], n_274);
  nand g156 (n_277, B[25], n_274);
  nand g157 (n_279, n_275, n_276, n_277);
  xor g158 (n_278, A[25], B[25]);
  xor g159 (Z[25], n_274, n_278);
  nand g160 (n_280, A[26], B[26]);
  nand g161 (n_281, A[26], n_279);
  nand g162 (n_282, B[26], n_279);
  nand g163 (n_284, n_280, n_281, n_282);
  xor g164 (n_283, A[26], B[26]);
  xor g165 (Z[26], n_279, n_283);
  nand g166 (n_285, A[27], B[27]);
  nand g167 (n_286, A[27], n_284);
  nand g168 (n_287, B[27], n_284);
  nand g169 (n_289, n_285, n_286, n_287);
  xor g170 (n_288, A[27], B[27]);
  xor g171 (Z[27], n_284, n_288);
  nand g172 (n_290, A[28], B[28]);
  nand g173 (n_291, A[28], n_289);
  nand g174 (n_292, B[28], n_289);
  nand g175 (n_294, n_290, n_291, n_292);
  xor g176 (n_293, A[28], B[28]);
  xor g177 (Z[28], n_289, n_293);
  nand g178 (n_295, A[29], B[29]);
  nand g179 (n_296, A[29], n_294);
  nand g180 (n_297, B[29], n_294);
  nand g181 (n_299, n_295, n_296, n_297);
  xor g182 (n_298, A[29], B[29]);
  xor g183 (Z[29], n_294, n_298);
  nand g184 (n_300, A[30], B[30]);
  nand g185 (n_301, A[30], n_299);
  nand g186 (n_302, B[30], n_299);
  nand g187 (n_304, n_300, n_301, n_302);
  xor g188 (n_303, A[30], B[30]);
  xor g189 (Z[30], n_299, n_303);
  nand g190 (n_305, A[31], B[31]);
  nand g191 (n_306, A[31], n_304);
  nand g192 (n_307, B[31], n_304);
  nand g193 (n_309, n_305, n_306, n_307);
  xor g194 (n_308, A[31], B[31]);
  xor g195 (Z[31], n_304, n_308);
  nand g196 (n_310, A[32], B[32]);
  nand g197 (n_311, A[32], n_309);
  nand g198 (n_312, B[32], n_309);
  nand g199 (n_314, n_310, n_311, n_312);
  xor g200 (n_313, A[32], B[32]);
  xor g201 (Z[32], n_309, n_313);
  nand g202 (n_315, A[33], B[33]);
  nand g203 (n_316, A[33], n_314);
  nand g204 (n_317, B[33], n_314);
  nand g205 (n_319, n_315, n_316, n_317);
  xor g206 (n_318, A[33], B[33]);
  xor g207 (Z[33], n_314, n_318);
  nand g208 (n_320, A[34], B[34]);
  nand g209 (n_321, A[34], n_319);
  nand g210 (n_322, B[34], n_319);
  nand g211 (n_324, n_320, n_321, n_322);
  xor g212 (n_323, A[34], B[34]);
  xor g213 (Z[34], n_319, n_323);
  nand g214 (n_325, A[35], B[35]);
  nand g215 (n_326, A[35], n_324);
  nand g216 (n_327, B[35], n_324);
  nand g217 (n_329, n_325, n_326, n_327);
  xor g218 (n_328, A[35], B[35]);
  xor g219 (Z[35], n_324, n_328);
  nand g220 (n_330, A[36], B[36]);
  nand g221 (n_331, A[36], n_329);
  nand g222 (n_332, B[36], n_329);
  nand g223 (n_334, n_330, n_331, n_332);
  xor g224 (n_333, A[36], B[36]);
  xor g225 (Z[36], n_329, n_333);
  nand g226 (n_335, A[37], B[37]);
  nand g227 (n_336, A[37], n_334);
  nand g228 (n_337, B[37], n_334);
  nand g229 (n_339, n_335, n_336, n_337);
  xor g230 (n_338, A[37], B[37]);
  xor g231 (Z[37], n_334, n_338);
  nand g232 (n_340, A[38], B[38]);
  nand g233 (n_341, A[38], n_339);
  nand g234 (n_342, B[38], n_339);
  nand g235 (n_344, n_340, n_341, n_342);
  xor g236 (n_343, A[38], B[38]);
  xor g237 (Z[38], n_339, n_343);
  nand g238 (n_345, A[39], B[39]);
  nand g239 (n_346, A[39], n_344);
  nand g240 (n_347, B[39], n_344);
  nand g241 (n_349, n_345, n_346, n_347);
  xor g242 (n_348, A[39], B[39]);
  xor g243 (Z[39], n_344, n_348);
  nand g244 (n_350, A[40], B[40]);
  nand g245 (n_351, A[40], n_349);
  nand g246 (n_352, B[40], n_349);
  nand g247 (n_354, n_350, n_351, n_352);
  xor g248 (n_353, A[40], B[40]);
  xor g249 (Z[40], n_349, n_353);
  nand g250 (n_355, A[41], B[41]);
  nand g251 (n_356, A[41], n_354);
  nand g252 (n_357, B[41], n_354);
  nand g253 (n_359, n_355, n_356, n_357);
  xor g254 (n_358, A[41], B[41]);
  xor g255 (Z[41], n_354, n_358);
  nand g256 (n_360, A[42], B[42]);
  nand g257 (n_361, A[42], n_359);
  nand g258 (n_362, B[42], n_359);
  nand g259 (n_364, n_360, n_361, n_362);
  xor g260 (n_363, A[42], B[42]);
  xor g261 (Z[42], n_359, n_363);
  nand g262 (n_365, A[43], B[43]);
  nand g263 (n_366, A[43], n_364);
  nand g264 (n_367, B[43], n_364);
  nand g265 (n_369, n_365, n_366, n_367);
  xor g266 (n_368, A[43], B[43]);
  xor g267 (Z[43], n_364, n_368);
  nand g268 (n_370, A[44], B[44]);
  nand g269 (n_371, A[44], n_369);
  nand g270 (n_372, B[44], n_369);
  nand g271 (n_374, n_370, n_371, n_372);
  xor g272 (n_373, A[44], B[44]);
  xor g273 (Z[44], n_369, n_373);
  nand g274 (n_375, A[45], B[45]);
  nand g275 (n_376, A[45], n_374);
  nand g276 (n_377, B[45], n_374);
  nand g277 (n_379, n_375, n_376, n_377);
  xor g278 (n_378, A[45], B[45]);
  xor g279 (Z[45], n_374, n_378);
  nand g280 (n_380, A[46], B[46]);
  nand g281 (n_381, A[46], n_379);
  nand g282 (n_382, B[46], n_379);
  nand g283 (n_384, n_380, n_381, n_382);
  xor g284 (n_383, A[46], B[46]);
  xor g285 (Z[46], n_379, n_383);
  nand g289 (n_149, n_385, n_386, n_387);
  xor g291 (Z[47], n_384, n_388);
  or g293 (n_385, A[47], B[47]);
  xor g294 (n_388, A[47], B[47]);
  or g295 (n_156, wc, n_150);
  not gc (wc, A[1]);
  or g296 (n_157, wc0, n_150);
  not gc0 (wc0, B[1]);
  xnor g297 (Z[1], n_150, n_158);
  or g298 (n_386, A[47], wc1);
  not gc1 (wc1, n_384);
  or g299 (n_387, B[47], wc2);
  not gc2 (wc2, n_384);
endmodule

module add_signed_342_2_GENERIC(A, B, Z);
  input [47:0] A, B;
  output [48:0] Z;
  wire [47:0] A, B;
  wire [48:0] Z;
  add_signed_342_2_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_356_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [46:0] A, B;
  output [47:0] Z;
  wire [46:0] A, B;
  wire [47:0] Z;
  wire n_146, n_147, n_150, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_160, n_161, n_162, n_163, n_164, n_166, n_167;
  wire n_168, n_169, n_170, n_172, n_173, n_174, n_175, n_176;
  wire n_178, n_179, n_180, n_181, n_182, n_184, n_185, n_186;
  wire n_187, n_188, n_190, n_191, n_192, n_193, n_194, n_196;
  wire n_197, n_198, n_199, n_200, n_202, n_203, n_204, n_205;
  wire n_206, n_208, n_209, n_210, n_211, n_212, n_214, n_215;
  wire n_216, n_217, n_218, n_220, n_221, n_222, n_223, n_224;
  wire n_226, n_227, n_228, n_229, n_230, n_232, n_233, n_234;
  wire n_235, n_236, n_238, n_239, n_240, n_241, n_242, n_244;
  wire n_245, n_246, n_247, n_248, n_250, n_251, n_252, n_253;
  wire n_254, n_256, n_257, n_258, n_259, n_260, n_262, n_263;
  wire n_264, n_265, n_266, n_268, n_269, n_270, n_271, n_272;
  wire n_274, n_275, n_276, n_277, n_278, n_280, n_281, n_282;
  wire n_283, n_284, n_286, n_287, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_296, n_298, n_300, n_301, n_303, n_304;
  wire n_306, n_308, n_310, n_311, n_313, n_314, n_316, n_318;
  wire n_320, n_321, n_323, n_324, n_326, n_328, n_330, n_331;
  wire n_333, n_334, n_336, n_338, n_340, n_341, n_343, n_344;
  wire n_346, n_348, n_350, n_351, n_353, n_354, n_356, n_358;
  wire n_360, n_361, n_363, n_364, n_366, n_368, n_370, n_371;
  wire n_373, n_374, n_376, n_378, n_380, n_381, n_383, n_384;
  wire n_386, n_388, n_390, n_391, n_393, n_394, n_395, n_396;
  wire n_398, n_400, n_402, n_403, n_404, n_406, n_407, n_408;
  wire n_410, n_411, n_412, n_413, n_415, n_417, n_419, n_420;
  wire n_421, n_423, n_424, n_425, n_427, n_428, n_430, n_432;
  wire n_434, n_435, n_436, n_438, n_439, n_440, n_442, n_443;
  wire n_445, n_447, n_449, n_450, n_451, n_453, n_454, n_455;
  wire n_457, n_458, n_460, n_462, n_464, n_465, n_466, n_468;
  wire n_469, n_470, n_472, n_473, n_475, n_477, n_479, n_480;
  wire n_481, n_483, n_485, n_486, n_487, n_489, n_490, n_492;
  wire n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500;
  wire n_501, n_502, n_503, n_504, n_505, n_506, n_508, n_511;
  wire n_513, n_514, n_515, n_518, n_521, n_523, n_524, n_526;
  wire n_528, n_529, n_531, n_533, n_534, n_536, n_538, n_539;
  wire n_541, n_542, n_544, n_547, n_549, n_550, n_551, n_554;
  wire n_557, n_559, n_560, n_562, n_564, n_565, n_567, n_569;
  wire n_570, n_572, n_574, n_575, n_576, n_578, n_579, n_581;
  wire n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589;
  wire n_590, n_591, n_592, n_594, n_595, n_596, n_598, n_599;
  wire n_600, n_602, n_603, n_604, n_606, n_607, n_608, n_610;
  wire n_611, n_612, n_614, n_615, n_616, n_618, n_619, n_620;
  wire n_622, n_623, n_624, n_626, n_627, n_628, n_630, n_631;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_643, n_644, n_646, n_647, n_648, n_650;
  wire n_651, n_652, n_654, n_655, n_656, n_658, n_659, n_660;
  wire n_662, n_663, n_664, n_666, n_667, n_668, n_670, n_671;
  wire n_672, n_673, n_675, n_676, n_677, n_679, n_680, n_681;
  wire n_682, n_684, n_685, n_686, n_688, n_689, n_690, n_691;
  wire n_693, n_694, n_696, n_697, n_699, n_700, n_701, n_702;
  wire n_704, n_705, n_706, n_708, n_709, n_710, n_711, n_713;
  wire n_714, n_716, n_717, n_719, n_720, n_721, n_722, n_724;
  wire n_725, n_726, n_727, n_729, n_730, n_731, n_732, n_734;
  wire n_735, n_737, n_738, n_740, n_741, n_742, n_743, n_745;
  wire n_746, n_747, n_749, n_750, n_751, n_752, n_754, n_755;
  wire n_757, n_758, n_760, n_761, n_762, n_763, n_765, n_766;
  wire n_767, n_768, n_770, n_771, n_772, n_773, n_775, n_776;
  wire n_778, n_779, n_781, n_782, n_783, n_784;
  not g3 (Z[47], n_146);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_147, A[0], B[0]);
  nor g9 (n_150, A[1], B[1]);
  nand g10 (n_153, A[1], B[1]);
  nor g11 (n_160, A[2], B[2]);
  nand g12 (n_155, A[2], B[2]);
  nor g13 (n_156, A[3], B[3]);
  nand g14 (n_157, A[3], B[3]);
  nor g15 (n_166, A[4], B[4]);
  nand g16 (n_161, A[4], B[4]);
  nor g17 (n_162, A[5], B[5]);
  nand g18 (n_163, A[5], B[5]);
  nor g19 (n_172, A[6], B[6]);
  nand g20 (n_167, A[6], B[6]);
  nor g21 (n_168, A[7], B[7]);
  nand g22 (n_169, A[7], B[7]);
  nor g23 (n_178, A[8], B[8]);
  nand g24 (n_173, A[8], B[8]);
  nor g25 (n_174, A[9], B[9]);
  nand g26 (n_175, A[9], B[9]);
  nor g27 (n_184, A[10], B[10]);
  nand g28 (n_179, A[10], B[10]);
  nor g29 (n_180, A[11], B[11]);
  nand g30 (n_181, A[11], B[11]);
  nor g31 (n_190, A[12], B[12]);
  nand g32 (n_185, A[12], B[12]);
  nor g33 (n_186, A[13], B[13]);
  nand g34 (n_187, A[13], B[13]);
  nor g35 (n_196, A[14], B[14]);
  nand g36 (n_191, A[14], B[14]);
  nor g37 (n_192, A[15], B[15]);
  nand g38 (n_193, A[15], B[15]);
  nor g39 (n_202, A[16], B[16]);
  nand g40 (n_197, A[16], B[16]);
  nor g41 (n_198, A[17], B[17]);
  nand g42 (n_199, A[17], B[17]);
  nor g43 (n_208, A[18], B[18]);
  nand g44 (n_203, A[18], B[18]);
  nor g45 (n_204, A[19], B[19]);
  nand g46 (n_205, A[19], B[19]);
  nor g47 (n_214, A[20], B[20]);
  nand g48 (n_209, A[20], B[20]);
  nor g49 (n_210, A[21], B[21]);
  nand g50 (n_211, A[21], B[21]);
  nor g51 (n_220, A[22], B[22]);
  nand g52 (n_215, A[22], B[22]);
  nor g53 (n_216, A[23], B[23]);
  nand g54 (n_217, A[23], B[23]);
  nor g55 (n_226, A[24], B[24]);
  nand g56 (n_221, A[24], B[24]);
  nor g57 (n_222, A[25], B[25]);
  nand g58 (n_223, A[25], B[25]);
  nor g59 (n_232, A[26], B[26]);
  nand g60 (n_227, A[26], B[26]);
  nor g61 (n_228, A[27], B[27]);
  nand g62 (n_229, A[27], B[27]);
  nor g63 (n_238, A[28], B[28]);
  nand g64 (n_233, A[28], B[28]);
  nor g65 (n_234, A[29], B[29]);
  nand g66 (n_235, A[29], B[29]);
  nor g67 (n_244, A[30], B[30]);
  nand g68 (n_239, A[30], B[30]);
  nor g69 (n_240, A[31], B[31]);
  nand g70 (n_241, A[31], B[31]);
  nor g71 (n_250, A[32], B[32]);
  nand g72 (n_245, A[32], B[32]);
  nor g73 (n_246, A[33], B[33]);
  nand g74 (n_247, A[33], B[33]);
  nor g75 (n_256, A[34], B[34]);
  nand g76 (n_251, A[34], B[34]);
  nor g77 (n_252, A[35], B[35]);
  nand g78 (n_253, A[35], B[35]);
  nor g79 (n_262, A[36], B[36]);
  nand g80 (n_257, A[36], B[36]);
  nor g81 (n_258, A[37], B[37]);
  nand g82 (n_259, A[37], B[37]);
  nor g83 (n_268, A[38], B[38]);
  nand g84 (n_263, A[38], B[38]);
  nor g85 (n_264, A[39], B[39]);
  nand g86 (n_265, A[39], B[39]);
  nor g87 (n_274, A[40], B[40]);
  nand g88 (n_269, A[40], B[40]);
  nor g89 (n_270, A[41], B[41]);
  nand g90 (n_271, A[41], B[41]);
  nor g91 (n_280, A[42], B[42]);
  nand g92 (n_275, A[42], B[42]);
  nor g93 (n_276, A[43], B[43]);
  nand g94 (n_277, A[43], B[43]);
  nor g95 (n_286, A[44], B[44]);
  nand g96 (n_281, A[44], B[44]);
  nor g97 (n_282, A[45], B[45]);
  nand g98 (n_283, A[45], B[45]);
  nand g103 (n_287, n_153, n_154);
  nor g104 (n_158, n_155, n_156);
  nor g107 (n_290, n_160, n_156);
  nor g108 (n_164, n_161, n_162);
  nor g111 (n_296, n_166, n_162);
  nor g112 (n_170, n_167, n_168);
  nor g115 (n_298, n_172, n_168);
  nor g116 (n_176, n_173, n_174);
  nor g119 (n_306, n_178, n_174);
  nor g120 (n_182, n_179, n_180);
  nor g123 (n_308, n_184, n_180);
  nor g124 (n_188, n_185, n_186);
  nor g127 (n_316, n_190, n_186);
  nor g128 (n_194, n_191, n_192);
  nor g131 (n_318, n_196, n_192);
  nor g132 (n_200, n_197, n_198);
  nor g135 (n_326, n_202, n_198);
  nor g136 (n_206, n_203, n_204);
  nor g139 (n_328, n_208, n_204);
  nor g140 (n_212, n_209, n_210);
  nor g143 (n_336, n_214, n_210);
  nor g144 (n_218, n_215, n_216);
  nor g147 (n_338, n_220, n_216);
  nor g148 (n_224, n_221, n_222);
  nor g151 (n_346, n_226, n_222);
  nor g152 (n_230, n_227, n_228);
  nor g155 (n_348, n_232, n_228);
  nor g156 (n_236, n_233, n_234);
  nor g159 (n_356, n_238, n_234);
  nor g160 (n_242, n_239, n_240);
  nor g163 (n_358, n_244, n_240);
  nor g164 (n_248, n_245, n_246);
  nor g167 (n_366, n_250, n_246);
  nor g168 (n_254, n_251, n_252);
  nor g171 (n_368, n_256, n_252);
  nor g172 (n_260, n_257, n_258);
  nor g175 (n_376, n_262, n_258);
  nor g176 (n_266, n_263, n_264);
  nor g179 (n_378, n_268, n_264);
  nor g180 (n_272, n_269, n_270);
  nor g183 (n_386, n_274, n_270);
  nor g184 (n_278, n_275, n_276);
  nor g187 (n_388, n_280, n_276);
  nor g188 (n_284, n_281, n_282);
  nor g191 (n_398, n_286, n_282);
  nand g194 (n_675, n_155, n_289);
  nand g195 (n_292, n_290, n_287);
  nand g196 (n_400, n_291, n_292);
  nor g197 (n_294, n_172, n_293);
  nand g206 (n_408, n_296, n_298);
  nor g207 (n_304, n_184, n_303);
  nand g216 (n_415, n_306, n_308);
  nor g217 (n_314, n_196, n_313);
  nand g226 (n_423, n_316, n_318);
  nor g227 (n_324, n_208, n_323);
  nand g236 (n_430, n_326, n_328);
  nor g237 (n_334, n_220, n_333);
  nand g246 (n_438, n_336, n_338);
  nor g247 (n_344, n_232, n_343);
  nand g256 (n_445, n_346, n_348);
  nor g257 (n_354, n_244, n_353);
  nand g266 (n_453, n_356, n_358);
  nor g267 (n_364, n_256, n_363);
  nand g276 (n_460, n_366, n_368);
  nor g277 (n_374, n_268, n_373);
  nand g286 (n_468, n_376, n_378);
  nor g287 (n_384, n_280, n_383);
  nand g296 (n_475, n_386, n_388);
  nor g297 (n_396, n_393, n_394);
  nand g304 (n_679, n_161, n_402);
  nand g305 (n_403, n_296, n_400);
  nand g306 (n_681, n_293, n_403);
  nand g309 (n_684, n_406, n_407);
  nand g312 (n_483, n_410, n_411);
  nor g313 (n_413, n_190, n_412);
  nor g316 (n_493, n_190, n_415);
  nor g322 (n_421, n_419, n_412);
  nor g325 (n_499, n_415, n_419);
  nor g326 (n_425, n_423, n_412);
  nor g329 (n_502, n_415, n_423);
  nor g330 (n_428, n_214, n_427);
  nor g333 (n_582, n_214, n_430);
  nor g339 (n_436, n_434, n_427);
  nor g342 (n_588, n_430, n_434);
  nor g343 (n_440, n_438, n_427);
  nor g346 (n_508, n_430, n_438);
  nor g347 (n_443, n_238, n_442);
  nor g350 (n_521, n_238, n_445);
  nor g356 (n_451, n_449, n_442);
  nor g359 (n_531, n_445, n_449);
  nor g360 (n_455, n_453, n_442);
  nor g363 (n_536, n_445, n_453);
  nor g364 (n_458, n_262, n_457);
  nor g367 (n_634, n_262, n_460);
  nor g373 (n_466, n_464, n_457);
  nor g376 (n_640, n_460, n_464);
  nor g377 (n_470, n_468, n_457);
  nor g380 (n_544, n_460, n_468);
  nor g381 (n_473, n_286, n_472);
  nor g384 (n_557, n_286, n_475);
  nor g390 (n_481, n_479, n_472);
  nor g393 (n_567, n_475, n_479);
  nand g396 (n_688, n_173, n_485);
  nand g397 (n_486, n_306, n_483);
  nand g398 (n_690, n_303, n_486);
  nand g401 (n_693, n_489, n_490);
  nand g404 (n_696, n_412, n_492);
  nand g405 (n_495, n_493, n_483);
  nand g406 (n_699, n_494, n_495);
  nand g407 (n_498, n_496, n_483);
  nand g408 (n_701, n_497, n_498);
  nand g409 (n_501, n_499, n_483);
  nand g410 (n_704, n_500, n_501);
  nand g411 (n_504, n_502, n_483);
  nand g412 (n_572, n_503, n_504);
  nor g413 (n_506, n_226, n_505);
  nand g422 (n_596, n_346, n_508);
  nor g423 (n_515, n_513, n_505);
  nor g428 (n_518, n_445, n_505);
  nand g437 (n_608, n_508, n_521);
  nand g442 (n_612, n_508, n_526);
  nand g447 (n_616, n_508, n_531);
  nand g452 (n_620, n_508, n_536);
  nor g453 (n_542, n_274, n_541);
  nand g462 (n_648, n_386, n_544);
  nor g463 (n_551, n_549, n_541);
  nor g468 (n_554, n_475, n_541);
  nand g477 (n_660, n_544, n_557);
  nand g482 (n_664, n_544, n_562);
  nand g487 (n_668, n_544, n_567);
  nand g490 (n_708, n_197, n_574);
  nand g491 (n_575, n_326, n_572);
  nand g492 (n_710, n_323, n_575);
  nand g495 (n_713, n_578, n_579);
  nand g498 (n_716, n_427, n_581);
  nand g499 (n_584, n_582, n_572);
  nand g500 (n_719, n_583, n_584);
  nand g501 (n_587, n_585, n_572);
  nand g502 (n_721, n_586, n_587);
  nand g503 (n_590, n_588, n_572);
  nand g504 (n_724, n_589, n_590);
  nand g505 (n_591, n_508, n_572);
  nand g506 (n_726, n_505, n_591);
  nand g509 (n_729, n_594, n_595);
  nand g512 (n_731, n_598, n_599);
  nand g515 (n_734, n_602, n_603);
  nand g518 (n_737, n_606, n_607);
  nand g521 (n_740, n_610, n_611);
  nand g524 (n_742, n_614, n_615);
  nand g527 (n_745, n_618, n_619);
  nand g530 (n_624, n_622, n_623);
  nand g533 (n_749, n_245, n_626);
  nand g534 (n_627, n_366, n_624);
  nand g535 (n_751, n_363, n_627);
  nand g538 (n_754, n_630, n_631);
  nand g541 (n_757, n_457, n_633);
  nand g542 (n_636, n_634, n_624);
  nand g543 (n_760, n_635, n_636);
  nand g544 (n_639, n_637, n_624);
  nand g545 (n_762, n_638, n_639);
  nand g546 (n_642, n_640, n_624);
  nand g547 (n_765, n_641, n_642);
  nand g548 (n_643, n_544, n_624);
  nand g549 (n_767, n_541, n_643);
  nand g552 (n_770, n_646, n_647);
  nand g555 (n_772, n_650, n_651);
  nand g558 (n_775, n_654, n_655);
  nand g561 (n_778, n_658, n_659);
  nand g564 (n_781, n_662, n_663);
  nand g567 (n_783, n_666, n_667);
  nand g570 (n_146, n_670, n_671);
  xnor g574 (Z[2], n_287, n_673);
  xnor g577 (Z[3], n_675, n_676);
  xnor g579 (Z[4], n_400, n_677);
  xnor g582 (Z[5], n_679, n_680);
  xnor g584 (Z[6], n_681, n_682);
  xnor g587 (Z[7], n_684, n_685);
  xnor g589 (Z[8], n_483, n_686);
  xnor g592 (Z[9], n_688, n_689);
  xnor g594 (Z[10], n_690, n_691);
  xnor g597 (Z[11], n_693, n_694);
  xnor g600 (Z[12], n_696, n_697);
  xnor g603 (Z[13], n_699, n_700);
  xnor g605 (Z[14], n_701, n_702);
  xnor g608 (Z[15], n_704, n_705);
  xnor g610 (Z[16], n_572, n_706);
  xnor g613 (Z[17], n_708, n_709);
  xnor g615 (Z[18], n_710, n_711);
  xnor g618 (Z[19], n_713, n_714);
  xnor g621 (Z[20], n_716, n_717);
  xnor g624 (Z[21], n_719, n_720);
  xnor g626 (Z[22], n_721, n_722);
  xnor g629 (Z[23], n_724, n_725);
  xnor g631 (Z[24], n_726, n_727);
  xnor g634 (Z[25], n_729, n_730);
  xnor g636 (Z[26], n_731, n_732);
  xnor g639 (Z[27], n_734, n_735);
  xnor g642 (Z[28], n_737, n_738);
  xnor g645 (Z[29], n_740, n_741);
  xnor g647 (Z[30], n_742, n_743);
  xnor g650 (Z[31], n_745, n_746);
  xnor g652 (Z[32], n_624, n_747);
  xnor g655 (Z[33], n_749, n_750);
  xnor g657 (Z[34], n_751, n_752);
  xnor g660 (Z[35], n_754, n_755);
  xnor g663 (Z[36], n_757, n_758);
  xnor g666 (Z[37], n_760, n_761);
  xnor g668 (Z[38], n_762, n_763);
  xnor g671 (Z[39], n_765, n_766);
  xnor g673 (Z[40], n_767, n_768);
  xnor g676 (Z[41], n_770, n_771);
  xnor g678 (Z[42], n_772, n_773);
  xnor g681 (Z[43], n_775, n_776);
  xnor g684 (Z[44], n_778, n_779);
  xnor g687 (Z[45], n_781, n_782);
  xnor g689 (Z[46], n_783, n_784);
  and g692 (n_393, A[46], B[46]);
  or g693 (n_395, A[46], B[46]);
  and g694 (n_363, wc, n_247);
  not gc (wc, n_248);
  and g695 (n_370, wc0, n_253);
  not gc0 (wc0, n_254);
  and g696 (n_373, wc1, n_259);
  not gc1 (wc1, n_260);
  and g697 (n_380, wc2, n_265);
  not gc2 (wc2, n_266);
  and g698 (n_383, wc3, n_271);
  not gc3 (wc3, n_272);
  and g699 (n_390, wc4, n_277);
  not gc4 (wc4, n_278);
  and g700 (n_394, wc5, n_283);
  not gc5 (wc5, n_284);
  and g701 (n_323, wc6, n_199);
  not gc6 (wc6, n_200);
  and g702 (n_330, wc7, n_205);
  not gc7 (wc7, n_206);
  and g703 (n_333, wc8, n_211);
  not gc8 (wc8, n_212);
  and g704 (n_340, wc9, n_217);
  not gc9 (wc9, n_218);
  and g705 (n_343, wc10, n_223);
  not gc10 (wc10, n_224);
  and g706 (n_350, wc11, n_229);
  not gc11 (wc11, n_230);
  and g707 (n_353, wc12, n_235);
  not gc12 (wc12, n_236);
  and g708 (n_360, wc13, n_241);
  not gc13 (wc13, n_242);
  and g709 (n_303, wc14, n_175);
  not gc14 (wc14, n_176);
  and g710 (n_310, wc15, n_181);
  not gc15 (wc15, n_182);
  and g711 (n_313, wc16, n_187);
  not gc16 (wc16, n_188);
  and g712 (n_320, wc17, n_193);
  not gc17 (wc17, n_194);
  and g713 (n_293, wc18, n_163);
  not gc18 (wc18, n_164);
  and g714 (n_300, wc19, n_169);
  not gc19 (wc19, n_170);
  and g715 (n_291, wc20, n_157);
  not gc20 (wc20, n_158);
  or g716 (n_154, n_147, n_150);
  or g717 (n_404, wc21, n_172);
  not gc21 (wc21, n_296);
  or g718 (n_487, wc22, n_184);
  not gc22 (wc22, n_306);
  or g719 (n_419, wc23, n_196);
  not gc23 (wc23, n_316);
  or g720 (n_576, wc24, n_208);
  not gc24 (wc24, n_326);
  or g721 (n_434, wc25, n_220);
  not gc25 (wc25, n_336);
  or g722 (n_513, wc26, n_232);
  not gc26 (wc26, n_346);
  or g723 (n_449, wc27, n_244);
  not gc27 (wc27, n_356);
  or g724 (n_628, wc28, n_256);
  not gc28 (wc28, n_366);
  or g725 (n_464, wc29, n_268);
  not gc29 (wc29, n_376);
  or g726 (n_549, wc30, n_280);
  not gc30 (wc30, n_386);
  or g727 (n_672, wc31, n_150);
  not gc31 (wc31, n_153);
  or g728 (n_673, wc32, n_160);
  not gc32 (wc32, n_155);
  or g729 (n_676, wc33, n_156);
  not gc33 (wc33, n_157);
  or g730 (n_677, wc34, n_166);
  not gc34 (wc34, n_161);
  or g731 (n_680, wc35, n_162);
  not gc35 (wc35, n_163);
  or g732 (n_682, wc36, n_172);
  not gc36 (wc36, n_167);
  or g733 (n_685, wc37, n_168);
  not gc37 (wc37, n_169);
  or g734 (n_686, wc38, n_178);
  not gc38 (wc38, n_173);
  or g735 (n_689, wc39, n_174);
  not gc39 (wc39, n_175);
  or g736 (n_691, wc40, n_184);
  not gc40 (wc40, n_179);
  or g737 (n_694, wc41, n_180);
  not gc41 (wc41, n_181);
  or g738 (n_697, wc42, n_190);
  not gc42 (wc42, n_185);
  or g739 (n_700, wc43, n_186);
  not gc43 (wc43, n_187);
  or g740 (n_702, wc44, n_196);
  not gc44 (wc44, n_191);
  or g741 (n_705, wc45, n_192);
  not gc45 (wc45, n_193);
  or g742 (n_706, wc46, n_202);
  not gc46 (wc46, n_197);
  or g743 (n_709, wc47, n_198);
  not gc47 (wc47, n_199);
  or g744 (n_711, wc48, n_208);
  not gc48 (wc48, n_203);
  or g745 (n_714, wc49, n_204);
  not gc49 (wc49, n_205);
  or g746 (n_717, wc50, n_214);
  not gc50 (wc50, n_209);
  or g747 (n_720, wc51, n_210);
  not gc51 (wc51, n_211);
  or g748 (n_722, wc52, n_220);
  not gc52 (wc52, n_215);
  or g749 (n_725, wc53, n_216);
  not gc53 (wc53, n_217);
  or g750 (n_727, wc54, n_226);
  not gc54 (wc54, n_221);
  or g751 (n_730, wc55, n_222);
  not gc55 (wc55, n_223);
  or g752 (n_732, wc56, n_232);
  not gc56 (wc56, n_227);
  or g753 (n_735, wc57, n_228);
  not gc57 (wc57, n_229);
  or g754 (n_738, wc58, n_238);
  not gc58 (wc58, n_233);
  or g755 (n_741, wc59, n_234);
  not gc59 (wc59, n_235);
  or g756 (n_743, wc60, n_244);
  not gc60 (wc60, n_239);
  or g757 (n_746, wc61, n_240);
  not gc61 (wc61, n_241);
  or g758 (n_747, wc62, n_250);
  not gc62 (wc62, n_245);
  or g759 (n_750, wc63, n_246);
  not gc63 (wc63, n_247);
  or g760 (n_752, wc64, n_256);
  not gc64 (wc64, n_251);
  or g761 (n_755, wc65, n_252);
  not gc65 (wc65, n_253);
  or g762 (n_758, wc66, n_262);
  not gc66 (wc66, n_257);
  or g763 (n_761, wc67, n_258);
  not gc67 (wc67, n_259);
  or g764 (n_763, wc68, n_268);
  not gc68 (wc68, n_263);
  or g765 (n_766, wc69, n_264);
  not gc69 (wc69, n_265);
  or g766 (n_768, wc70, n_274);
  not gc70 (wc70, n_269);
  or g767 (n_771, wc71, n_270);
  not gc71 (wc71, n_271);
  or g768 (n_773, wc72, n_280);
  not gc72 (wc72, n_275);
  or g769 (n_776, wc73, n_276);
  not gc73 (wc73, n_277);
  or g770 (n_779, wc74, n_286);
  not gc74 (wc74, n_281);
  or g771 (n_782, wc75, n_282);
  not gc75 (wc75, n_283);
  and g772 (n_371, wc76, n_368);
  not gc76 (wc76, n_363);
  and g773 (n_381, wc77, n_378);
  not gc77 (wc77, n_373);
  or g774 (n_479, n_393, wc78);
  not gc78 (wc78, n_398);
  and g775 (n_391, wc79, n_388);
  not gc79 (wc79, n_383);
  and g776 (n_331, wc80, n_328);
  not gc80 (wc80, n_323);
  and g777 (n_341, wc81, n_338);
  not gc81 (wc81, n_333);
  and g778 (n_351, wc82, n_348);
  not gc82 (wc82, n_343);
  and g779 (n_361, wc83, n_358);
  not gc83 (wc83, n_353);
  and g780 (n_311, wc84, n_308);
  not gc84 (wc84, n_303);
  and g781 (n_321, wc85, n_318);
  not gc85 (wc85, n_313);
  and g782 (n_301, wc86, n_298);
  not gc86 (wc86, n_293);
  and g783 (n_496, wc87, n_316);
  not gc87 (wc87, n_415);
  and g784 (n_585, wc88, n_336);
  not gc88 (wc88, n_430);
  and g785 (n_526, wc89, n_356);
  not gc89 (wc89, n_445);
  and g786 (n_637, wc90, n_376);
  not gc90 (wc90, n_460);
  and g787 (n_562, wc91, n_398);
  not gc91 (wc91, n_475);
  xor g788 (Z[1], n_147, n_672);
  or g789 (n_784, wc92, n_393);
  not gc92 (wc92, n_395);
  and g790 (n_457, wc93, n_370);
  not gc93 (wc93, n_371);
  and g791 (n_469, wc94, n_380);
  not gc94 (wc94, n_381);
  and g792 (n_472, wc95, n_390);
  not gc95 (wc95, n_391);
  and g793 (n_480, n_395, wc96);
  not gc96 (wc96, n_396);
  and g794 (n_427, wc97, n_330);
  not gc97 (wc97, n_331);
  and g795 (n_439, wc98, n_340);
  not gc98 (wc98, n_341);
  and g796 (n_442, wc99, n_350);
  not gc99 (wc99, n_351);
  and g797 (n_454, wc100, n_360);
  not gc100 (wc100, n_361);
  and g798 (n_412, wc101, n_310);
  not gc101 (wc101, n_311);
  and g799 (n_424, wc102, n_320);
  not gc102 (wc102, n_321);
  and g800 (n_410, wc103, n_300);
  not gc103 (wc103, n_301);
  or g801 (n_289, wc104, n_160);
  not gc104 (wc104, n_287);
  and g802 (n_406, wc105, n_167);
  not gc105 (wc105, n_294);
  and g803 (n_489, wc106, n_179);
  not gc106 (wc106, n_304);
  and g804 (n_420, wc107, n_191);
  not gc107 (wc107, n_314);
  and g805 (n_578, wc108, n_203);
  not gc108 (wc108, n_324);
  and g806 (n_435, wc109, n_215);
  not gc109 (wc109, n_334);
  and g807 (n_514, wc110, n_227);
  not gc110 (wc110, n_344);
  and g808 (n_450, wc111, n_239);
  not gc111 (wc111, n_354);
  and g809 (n_630, wc112, n_251);
  not gc112 (wc112, n_364);
  and g810 (n_465, wc113, n_263);
  not gc113 (wc113, n_374);
  and g811 (n_550, wc114, n_275);
  not gc114 (wc114, n_384);
  or g812 (n_592, wc115, n_226);
  not gc115 (wc115, n_508);
  or g813 (n_600, n_513, wc116);
  not gc116 (wc116, n_508);
  or g814 (n_604, wc117, n_445);
  not gc117 (wc117, n_508);
  or g815 (n_644, wc118, n_274);
  not gc118 (wc118, n_544);
  or g816 (n_652, n_549, wc119);
  not gc119 (wc119, n_544);
  or g817 (n_656, wc120, n_475);
  not gc120 (wc120, n_544);
  and g818 (n_417, wc121, n_316);
  not gc121 (wc121, n_412);
  and g819 (n_432, wc122, n_336);
  not gc122 (wc122, n_427);
  and g820 (n_447, wc123, n_356);
  not gc123 (wc123, n_442);
  and g821 (n_462, wc124, n_376);
  not gc124 (wc124, n_457);
  and g822 (n_477, wc125, n_398);
  not gc125 (wc125, n_472);
  and g823 (n_541, n_469, wc126);
  not gc126 (wc126, n_470);
  and g824 (n_569, n_480, wc127);
  not gc127 (wc127, n_481);
  and g825 (n_505, n_439, wc128);
  not gc128 (wc128, n_440);
  and g826 (n_538, n_454, wc129);
  not gc129 (wc129, n_455);
  and g827 (n_503, n_424, wc130);
  not gc130 (wc130, n_425);
  or g828 (n_411, n_408, wc131);
  not gc131 (wc131, n_400);
  or g829 (n_402, wc132, n_166);
  not gc132 (wc132, n_400);
  or g830 (n_407, n_404, wc133);
  not gc133 (wc133, n_400);
  and g831 (n_494, wc134, n_185);
  not gc134 (wc134, n_413);
  and g832 (n_497, wc135, n_313);
  not gc135 (wc135, n_417);
  and g833 (n_500, n_420, wc136);
  not gc136 (wc136, n_421);
  and g834 (n_583, wc137, n_209);
  not gc137 (wc137, n_428);
  and g835 (n_586, wc138, n_333);
  not gc138 (wc138, n_432);
  and g836 (n_589, n_435, wc139);
  not gc139 (wc139, n_436);
  and g837 (n_523, wc140, n_233);
  not gc140 (wc140, n_443);
  and g838 (n_528, wc141, n_353);
  not gc141 (wc141, n_447);
  and g839 (n_533, n_450, wc142);
  not gc142 (wc142, n_451);
  and g840 (n_635, wc143, n_257);
  not gc143 (wc143, n_458);
  and g841 (n_638, wc144, n_373);
  not gc144 (wc144, n_462);
  and g842 (n_641, n_465, wc145);
  not gc145 (wc145, n_466);
  and g843 (n_559, wc146, n_281);
  not gc146 (wc146, n_473);
  and g844 (n_564, wc147, n_394);
  not gc147 (wc147, n_477);
  and g845 (n_570, wc148, n_567);
  not gc148 (wc148, n_541);
  and g846 (n_539, wc149, n_536);
  not gc149 (wc149, n_505);
  and g847 (n_511, wc150, n_346);
  not gc150 (wc150, n_505);
  and g848 (n_524, wc151, n_521);
  not gc151 (wc151, n_505);
  and g849 (n_529, wc152, n_526);
  not gc152 (wc152, n_505);
  and g850 (n_534, wc153, n_531);
  not gc153 (wc153, n_505);
  and g851 (n_547, wc154, n_386);
  not gc154 (wc154, n_541);
  and g852 (n_560, wc155, n_557);
  not gc155 (wc155, n_541);
  and g853 (n_565, wc156, n_562);
  not gc156 (wc156, n_541);
  and g854 (n_670, wc157, n_569);
  not gc157 (wc157, n_570);
  and g855 (n_622, wc158, n_538);
  not gc158 (wc158, n_539);
  or g856 (n_485, wc159, n_178);
  not gc159 (wc159, n_483);
  or g857 (n_490, n_487, wc160);
  not gc160 (wc160, n_483);
  or g858 (n_492, wc161, n_415);
  not gc161 (wc161, n_483);
  and g859 (n_594, wc162, n_221);
  not gc162 (wc162, n_506);
  and g860 (n_598, wc163, n_343);
  not gc163 (wc163, n_511);
  and g861 (n_602, n_514, wc164);
  not gc164 (wc164, n_515);
  and g862 (n_606, n_442, wc165);
  not gc165 (wc165, n_518);
  and g863 (n_610, wc166, n_523);
  not gc166 (wc166, n_524);
  and g864 (n_614, wc167, n_528);
  not gc167 (wc167, n_529);
  and g865 (n_618, wc168, n_533);
  not gc168 (wc168, n_534);
  and g866 (n_646, wc169, n_269);
  not gc169 (wc169, n_542);
  and g867 (n_650, wc170, n_383);
  not gc170 (wc170, n_547);
  and g868 (n_654, n_550, wc171);
  not gc171 (wc171, n_551);
  and g869 (n_658, n_472, wc172);
  not gc172 (wc172, n_554);
  and g870 (n_662, wc173, n_559);
  not gc173 (wc173, n_560);
  and g871 (n_666, wc174, n_564);
  not gc174 (wc174, n_565);
  or g872 (n_623, n_620, wc175);
  not gc175 (wc175, n_572);
  or g873 (n_574, wc176, n_202);
  not gc176 (wc176, n_572);
  or g874 (n_579, n_576, wc177);
  not gc177 (wc177, n_572);
  or g875 (n_581, wc178, n_430);
  not gc178 (wc178, n_572);
  or g876 (n_595, n_592, wc179);
  not gc179 (wc179, n_572);
  or g877 (n_599, n_596, wc180);
  not gc180 (wc180, n_572);
  or g878 (n_603, n_600, wc181);
  not gc181 (wc181, n_572);
  or g879 (n_607, n_604, wc182);
  not gc182 (wc182, n_572);
  or g880 (n_611, n_608, wc183);
  not gc183 (wc183, n_572);
  or g881 (n_615, n_612, wc184);
  not gc184 (wc184, n_572);
  or g882 (n_619, n_616, wc185);
  not gc185 (wc185, n_572);
  or g883 (n_671, wc186, n_668);
  not gc186 (wc186, n_624);
  or g884 (n_626, wc187, n_250);
  not gc187 (wc187, n_624);
  or g885 (n_631, n_628, wc188);
  not gc188 (wc188, n_624);
  or g886 (n_633, wc189, n_460);
  not gc189 (wc189, n_624);
  or g887 (n_647, n_644, wc190);
  not gc190 (wc190, n_624);
  or g888 (n_651, wc191, n_648);
  not gc191 (wc191, n_624);
  or g889 (n_655, n_652, wc192);
  not gc192 (wc192, n_624);
  or g890 (n_659, n_656, wc193);
  not gc193 (wc193, n_624);
  or g891 (n_663, wc194, n_660);
  not gc194 (wc194, n_624);
  or g892 (n_667, wc195, n_664);
  not gc195 (wc195, n_624);
endmodule

module add_signed_356_GENERIC(A, B, Z);
  input [46:0] A, B;
  output [47:0] Z;
  wire [46:0] A, B;
  wire [47:0] Z;
  add_signed_356_GENERIC_REAL g1(.A ({A[45], A[45:0]}), .B ({B[45],
       B[45:0]}), .Z (Z));
endmodule

module add_signed_356_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [46:0] A, B;
  output [47:0] Z;
  wire [46:0] A, B;
  wire [47:0] Z;
  wire n_146, n_147, n_152, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213;
  wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253;
  wire n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261;
  wire n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269;
  wire n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285;
  wire n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_380;
  not g3 (Z[47], n_146);
  nand g4 (n_147, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_152, A[1], B[1]);
  nand g13 (n_156, n_152, n_153, n_154);
  xor g14 (n_155, A[1], B[1]);
  nand g16 (n_157, A[2], B[2]);
  nand g17 (n_158, A[2], n_156);
  nand g18 (n_159, B[2], n_156);
  nand g19 (n_161, n_157, n_158, n_159);
  xor g20 (n_160, A[2], B[2]);
  xor g21 (Z[2], n_156, n_160);
  nand g22 (n_162, A[3], B[3]);
  nand g23 (n_163, A[3], n_161);
  nand g24 (n_164, B[3], n_161);
  nand g25 (n_166, n_162, n_163, n_164);
  xor g26 (n_165, A[3], B[3]);
  xor g27 (Z[3], n_161, n_165);
  nand g28 (n_167, A[4], B[4]);
  nand g29 (n_168, A[4], n_166);
  nand g30 (n_169, B[4], n_166);
  nand g31 (n_171, n_167, n_168, n_169);
  xor g32 (n_170, A[4], B[4]);
  xor g33 (Z[4], n_166, n_170);
  nand g34 (n_172, A[5], B[5]);
  nand g35 (n_173, A[5], n_171);
  nand g36 (n_174, B[5], n_171);
  nand g37 (n_176, n_172, n_173, n_174);
  xor g38 (n_175, A[5], B[5]);
  xor g39 (Z[5], n_171, n_175);
  nand g40 (n_177, A[6], B[6]);
  nand g41 (n_178, A[6], n_176);
  nand g42 (n_179, B[6], n_176);
  nand g43 (n_181, n_177, n_178, n_179);
  xor g44 (n_180, A[6], B[6]);
  xor g45 (Z[6], n_176, n_180);
  nand g46 (n_182, A[7], B[7]);
  nand g47 (n_183, A[7], n_181);
  nand g48 (n_184, B[7], n_181);
  nand g49 (n_186, n_182, n_183, n_184);
  xor g50 (n_185, A[7], B[7]);
  xor g51 (Z[7], n_181, n_185);
  nand g52 (n_187, A[8], B[8]);
  nand g53 (n_188, A[8], n_186);
  nand g54 (n_189, B[8], n_186);
  nand g55 (n_191, n_187, n_188, n_189);
  xor g56 (n_190, A[8], B[8]);
  xor g57 (Z[8], n_186, n_190);
  nand g58 (n_192, A[9], B[9]);
  nand g59 (n_193, A[9], n_191);
  nand g60 (n_194, B[9], n_191);
  nand g61 (n_196, n_192, n_193, n_194);
  xor g62 (n_195, A[9], B[9]);
  xor g63 (Z[9], n_191, n_195);
  nand g64 (n_197, A[10], B[10]);
  nand g65 (n_198, A[10], n_196);
  nand g66 (n_199, B[10], n_196);
  nand g67 (n_201, n_197, n_198, n_199);
  xor g68 (n_200, A[10], B[10]);
  xor g69 (Z[10], n_196, n_200);
  nand g70 (n_202, A[11], B[11]);
  nand g71 (n_203, A[11], n_201);
  nand g72 (n_204, B[11], n_201);
  nand g73 (n_206, n_202, n_203, n_204);
  xor g74 (n_205, A[11], B[11]);
  xor g75 (Z[11], n_201, n_205);
  nand g76 (n_207, A[12], B[12]);
  nand g77 (n_208, A[12], n_206);
  nand g78 (n_209, B[12], n_206);
  nand g79 (n_211, n_207, n_208, n_209);
  xor g80 (n_210, A[12], B[12]);
  xor g81 (Z[12], n_206, n_210);
  nand g82 (n_212, A[13], B[13]);
  nand g83 (n_213, A[13], n_211);
  nand g84 (n_214, B[13], n_211);
  nand g85 (n_216, n_212, n_213, n_214);
  xor g86 (n_215, A[13], B[13]);
  xor g87 (Z[13], n_211, n_215);
  nand g88 (n_217, A[14], B[14]);
  nand g89 (n_218, A[14], n_216);
  nand g90 (n_219, B[14], n_216);
  nand g91 (n_221, n_217, n_218, n_219);
  xor g92 (n_220, A[14], B[14]);
  xor g93 (Z[14], n_216, n_220);
  nand g94 (n_222, A[15], B[15]);
  nand g95 (n_223, A[15], n_221);
  nand g96 (n_224, B[15], n_221);
  nand g97 (n_226, n_222, n_223, n_224);
  xor g98 (n_225, A[15], B[15]);
  xor g99 (Z[15], n_221, n_225);
  nand g100 (n_227, A[16], B[16]);
  nand g101 (n_228, A[16], n_226);
  nand g102 (n_229, B[16], n_226);
  nand g103 (n_231, n_227, n_228, n_229);
  xor g104 (n_230, A[16], B[16]);
  xor g105 (Z[16], n_226, n_230);
  nand g106 (n_232, A[17], B[17]);
  nand g107 (n_233, A[17], n_231);
  nand g108 (n_234, B[17], n_231);
  nand g109 (n_236, n_232, n_233, n_234);
  xor g110 (n_235, A[17], B[17]);
  xor g111 (Z[17], n_231, n_235);
  nand g112 (n_237, A[18], B[18]);
  nand g113 (n_238, A[18], n_236);
  nand g114 (n_239, B[18], n_236);
  nand g115 (n_241, n_237, n_238, n_239);
  xor g116 (n_240, A[18], B[18]);
  xor g117 (Z[18], n_236, n_240);
  nand g118 (n_242, A[19], B[19]);
  nand g119 (n_243, A[19], n_241);
  nand g120 (n_244, B[19], n_241);
  nand g121 (n_246, n_242, n_243, n_244);
  xor g122 (n_245, A[19], B[19]);
  xor g123 (Z[19], n_241, n_245);
  nand g124 (n_247, A[20], B[20]);
  nand g125 (n_248, A[20], n_246);
  nand g126 (n_249, B[20], n_246);
  nand g127 (n_251, n_247, n_248, n_249);
  xor g128 (n_250, A[20], B[20]);
  xor g129 (Z[20], n_246, n_250);
  nand g130 (n_252, A[21], B[21]);
  nand g131 (n_253, A[21], n_251);
  nand g132 (n_254, B[21], n_251);
  nand g133 (n_256, n_252, n_253, n_254);
  xor g134 (n_255, A[21], B[21]);
  xor g135 (Z[21], n_251, n_255);
  nand g136 (n_257, A[22], B[22]);
  nand g137 (n_258, A[22], n_256);
  nand g138 (n_259, B[22], n_256);
  nand g139 (n_261, n_257, n_258, n_259);
  xor g140 (n_260, A[22], B[22]);
  xor g141 (Z[22], n_256, n_260);
  nand g142 (n_262, A[23], B[23]);
  nand g143 (n_263, A[23], n_261);
  nand g144 (n_264, B[23], n_261);
  nand g145 (n_266, n_262, n_263, n_264);
  xor g146 (n_265, A[23], B[23]);
  xor g147 (Z[23], n_261, n_265);
  nand g148 (n_267, A[24], B[24]);
  nand g149 (n_268, A[24], n_266);
  nand g150 (n_269, B[24], n_266);
  nand g151 (n_271, n_267, n_268, n_269);
  xor g152 (n_270, A[24], B[24]);
  xor g153 (Z[24], n_266, n_270);
  nand g154 (n_272, A[25], B[25]);
  nand g155 (n_273, A[25], n_271);
  nand g156 (n_274, B[25], n_271);
  nand g157 (n_276, n_272, n_273, n_274);
  xor g158 (n_275, A[25], B[25]);
  xor g159 (Z[25], n_271, n_275);
  nand g160 (n_277, A[26], B[26]);
  nand g161 (n_278, A[26], n_276);
  nand g162 (n_279, B[26], n_276);
  nand g163 (n_281, n_277, n_278, n_279);
  xor g164 (n_280, A[26], B[26]);
  xor g165 (Z[26], n_276, n_280);
  nand g166 (n_282, A[27], B[27]);
  nand g167 (n_283, A[27], n_281);
  nand g168 (n_284, B[27], n_281);
  nand g169 (n_286, n_282, n_283, n_284);
  xor g170 (n_285, A[27], B[27]);
  xor g171 (Z[27], n_281, n_285);
  nand g172 (n_287, A[28], B[28]);
  nand g173 (n_288, A[28], n_286);
  nand g174 (n_289, B[28], n_286);
  nand g175 (n_291, n_287, n_288, n_289);
  xor g176 (n_290, A[28], B[28]);
  xor g177 (Z[28], n_286, n_290);
  nand g178 (n_292, A[29], B[29]);
  nand g179 (n_293, A[29], n_291);
  nand g180 (n_294, B[29], n_291);
  nand g181 (n_296, n_292, n_293, n_294);
  xor g182 (n_295, A[29], B[29]);
  xor g183 (Z[29], n_291, n_295);
  nand g184 (n_297, A[30], B[30]);
  nand g185 (n_298, A[30], n_296);
  nand g186 (n_299, B[30], n_296);
  nand g187 (n_301, n_297, n_298, n_299);
  xor g188 (n_300, A[30], B[30]);
  xor g189 (Z[30], n_296, n_300);
  nand g190 (n_302, A[31], B[31]);
  nand g191 (n_303, A[31], n_301);
  nand g192 (n_304, B[31], n_301);
  nand g193 (n_306, n_302, n_303, n_304);
  xor g194 (n_305, A[31], B[31]);
  xor g195 (Z[31], n_301, n_305);
  nand g196 (n_307, A[32], B[32]);
  nand g197 (n_308, A[32], n_306);
  nand g198 (n_309, B[32], n_306);
  nand g199 (n_311, n_307, n_308, n_309);
  xor g200 (n_310, A[32], B[32]);
  xor g201 (Z[32], n_306, n_310);
  nand g202 (n_312, A[33], B[33]);
  nand g203 (n_313, A[33], n_311);
  nand g204 (n_314, B[33], n_311);
  nand g205 (n_316, n_312, n_313, n_314);
  xor g206 (n_315, A[33], B[33]);
  xor g207 (Z[33], n_311, n_315);
  nand g208 (n_317, A[34], B[34]);
  nand g209 (n_318, A[34], n_316);
  nand g210 (n_319, B[34], n_316);
  nand g211 (n_321, n_317, n_318, n_319);
  xor g212 (n_320, A[34], B[34]);
  xor g213 (Z[34], n_316, n_320);
  nand g214 (n_322, A[35], B[35]);
  nand g215 (n_323, A[35], n_321);
  nand g216 (n_324, B[35], n_321);
  nand g217 (n_326, n_322, n_323, n_324);
  xor g218 (n_325, A[35], B[35]);
  xor g219 (Z[35], n_321, n_325);
  nand g220 (n_327, A[36], B[36]);
  nand g221 (n_328, A[36], n_326);
  nand g222 (n_329, B[36], n_326);
  nand g223 (n_331, n_327, n_328, n_329);
  xor g224 (n_330, A[36], B[36]);
  xor g225 (Z[36], n_326, n_330);
  nand g226 (n_332, A[37], B[37]);
  nand g227 (n_333, A[37], n_331);
  nand g228 (n_334, B[37], n_331);
  nand g229 (n_336, n_332, n_333, n_334);
  xor g230 (n_335, A[37], B[37]);
  xor g231 (Z[37], n_331, n_335);
  nand g232 (n_337, A[38], B[38]);
  nand g233 (n_338, A[38], n_336);
  nand g234 (n_339, B[38], n_336);
  nand g235 (n_341, n_337, n_338, n_339);
  xor g236 (n_340, A[38], B[38]);
  xor g237 (Z[38], n_336, n_340);
  nand g238 (n_342, A[39], B[39]);
  nand g239 (n_343, A[39], n_341);
  nand g240 (n_344, B[39], n_341);
  nand g241 (n_346, n_342, n_343, n_344);
  xor g242 (n_345, A[39], B[39]);
  xor g243 (Z[39], n_341, n_345);
  nand g244 (n_347, A[40], B[40]);
  nand g245 (n_348, A[40], n_346);
  nand g246 (n_349, B[40], n_346);
  nand g247 (n_351, n_347, n_348, n_349);
  xor g248 (n_350, A[40], B[40]);
  xor g249 (Z[40], n_346, n_350);
  nand g250 (n_352, A[41], B[41]);
  nand g251 (n_353, A[41], n_351);
  nand g252 (n_354, B[41], n_351);
  nand g253 (n_356, n_352, n_353, n_354);
  xor g254 (n_355, A[41], B[41]);
  xor g255 (Z[41], n_351, n_355);
  nand g256 (n_357, A[42], B[42]);
  nand g257 (n_358, A[42], n_356);
  nand g258 (n_359, B[42], n_356);
  nand g259 (n_361, n_357, n_358, n_359);
  xor g260 (n_360, A[42], B[42]);
  xor g261 (Z[42], n_356, n_360);
  nand g262 (n_362, A[43], B[43]);
  nand g263 (n_363, A[43], n_361);
  nand g264 (n_364, B[43], n_361);
  nand g265 (n_366, n_362, n_363, n_364);
  xor g266 (n_365, A[43], B[43]);
  xor g267 (Z[43], n_361, n_365);
  nand g268 (n_367, A[44], B[44]);
  nand g269 (n_368, A[44], n_366);
  nand g270 (n_369, B[44], n_366);
  nand g271 (n_371, n_367, n_368, n_369);
  xor g272 (n_370, A[44], B[44]);
  xor g273 (Z[44], n_366, n_370);
  nand g274 (n_372, A[45], B[45]);
  nand g275 (n_373, A[45], n_371);
  nand g276 (n_374, B[45], n_371);
  nand g277 (n_376, n_372, n_373, n_374);
  xor g278 (n_375, A[45], B[45]);
  xor g279 (Z[45], n_371, n_375);
  nand g283 (n_146, n_377, n_378, n_379);
  xor g285 (Z[46], n_376, n_380);
  or g287 (n_377, A[46], B[46]);
  xor g288 (n_380, A[46], B[46]);
  or g289 (n_153, wc, n_147);
  not gc (wc, A[1]);
  or g290 (n_154, wc0, n_147);
  not gc0 (wc0, B[1]);
  xnor g291 (Z[1], n_147, n_155);
  or g292 (n_378, A[46], wc1);
  not gc1 (wc1, n_376);
  or g293 (n_379, B[46], wc2);
  not gc2 (wc2, n_376);
endmodule

module add_signed_356_1_GENERIC(A, B, Z);
  input [46:0] A, B;
  output [47:0] Z;
  wire [46:0] A, B;
  wire [47:0] Z;
  add_signed_356_1_GENERIC_REAL g1(.A ({A[46:2], A[0], A[0]}), .B (B),
       .Z (Z));
endmodule

module add_signed_356_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [46:0] A, B;
  output [47:0] Z;
  wire [46:0] A, B;
  wire [47:0] Z;
  wire n_146, n_147, n_152, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213;
  wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253;
  wire n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261;
  wire n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269;
  wire n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285;
  wire n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_380;
  not g3 (Z[47], n_146);
  nand g4 (n_147, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_152, A[1], B[1]);
  nand g13 (n_156, n_152, n_153, n_154);
  xor g14 (n_155, A[1], B[1]);
  nand g16 (n_157, A[2], B[2]);
  nand g17 (n_158, A[2], n_156);
  nand g18 (n_159, B[2], n_156);
  nand g19 (n_161, n_157, n_158, n_159);
  xor g20 (n_160, A[2], B[2]);
  xor g21 (Z[2], n_156, n_160);
  nand g22 (n_162, A[3], B[3]);
  nand g23 (n_163, A[3], n_161);
  nand g24 (n_164, B[3], n_161);
  nand g25 (n_166, n_162, n_163, n_164);
  xor g26 (n_165, A[3], B[3]);
  xor g27 (Z[3], n_161, n_165);
  nand g28 (n_167, A[4], B[4]);
  nand g29 (n_168, A[4], n_166);
  nand g30 (n_169, B[4], n_166);
  nand g31 (n_171, n_167, n_168, n_169);
  xor g32 (n_170, A[4], B[4]);
  xor g33 (Z[4], n_166, n_170);
  nand g34 (n_172, A[5], B[5]);
  nand g35 (n_173, A[5], n_171);
  nand g36 (n_174, B[5], n_171);
  nand g37 (n_176, n_172, n_173, n_174);
  xor g38 (n_175, A[5], B[5]);
  xor g39 (Z[5], n_171, n_175);
  nand g40 (n_177, A[6], B[6]);
  nand g41 (n_178, A[6], n_176);
  nand g42 (n_179, B[6], n_176);
  nand g43 (n_181, n_177, n_178, n_179);
  xor g44 (n_180, A[6], B[6]);
  xor g45 (Z[6], n_176, n_180);
  nand g46 (n_182, A[7], B[7]);
  nand g47 (n_183, A[7], n_181);
  nand g48 (n_184, B[7], n_181);
  nand g49 (n_186, n_182, n_183, n_184);
  xor g50 (n_185, A[7], B[7]);
  xor g51 (Z[7], n_181, n_185);
  nand g52 (n_187, A[8], B[8]);
  nand g53 (n_188, A[8], n_186);
  nand g54 (n_189, B[8], n_186);
  nand g55 (n_191, n_187, n_188, n_189);
  xor g56 (n_190, A[8], B[8]);
  xor g57 (Z[8], n_186, n_190);
  nand g58 (n_192, A[9], B[9]);
  nand g59 (n_193, A[9], n_191);
  nand g60 (n_194, B[9], n_191);
  nand g61 (n_196, n_192, n_193, n_194);
  xor g62 (n_195, A[9], B[9]);
  xor g63 (Z[9], n_191, n_195);
  nand g64 (n_197, A[10], B[10]);
  nand g65 (n_198, A[10], n_196);
  nand g66 (n_199, B[10], n_196);
  nand g67 (n_201, n_197, n_198, n_199);
  xor g68 (n_200, A[10], B[10]);
  xor g69 (Z[10], n_196, n_200);
  nand g70 (n_202, A[11], B[11]);
  nand g71 (n_203, A[11], n_201);
  nand g72 (n_204, B[11], n_201);
  nand g73 (n_206, n_202, n_203, n_204);
  xor g74 (n_205, A[11], B[11]);
  xor g75 (Z[11], n_201, n_205);
  nand g76 (n_207, A[12], B[12]);
  nand g77 (n_208, A[12], n_206);
  nand g78 (n_209, B[12], n_206);
  nand g79 (n_211, n_207, n_208, n_209);
  xor g80 (n_210, A[12], B[12]);
  xor g81 (Z[12], n_206, n_210);
  nand g82 (n_212, A[13], B[13]);
  nand g83 (n_213, A[13], n_211);
  nand g84 (n_214, B[13], n_211);
  nand g85 (n_216, n_212, n_213, n_214);
  xor g86 (n_215, A[13], B[13]);
  xor g87 (Z[13], n_211, n_215);
  nand g88 (n_217, A[14], B[14]);
  nand g89 (n_218, A[14], n_216);
  nand g90 (n_219, B[14], n_216);
  nand g91 (n_221, n_217, n_218, n_219);
  xor g92 (n_220, A[14], B[14]);
  xor g93 (Z[14], n_216, n_220);
  nand g94 (n_222, A[15], B[15]);
  nand g95 (n_223, A[15], n_221);
  nand g96 (n_224, B[15], n_221);
  nand g97 (n_226, n_222, n_223, n_224);
  xor g98 (n_225, A[15], B[15]);
  xor g99 (Z[15], n_221, n_225);
  nand g100 (n_227, A[16], B[16]);
  nand g101 (n_228, A[16], n_226);
  nand g102 (n_229, B[16], n_226);
  nand g103 (n_231, n_227, n_228, n_229);
  xor g104 (n_230, A[16], B[16]);
  xor g105 (Z[16], n_226, n_230);
  nand g106 (n_232, A[17], B[17]);
  nand g107 (n_233, A[17], n_231);
  nand g108 (n_234, B[17], n_231);
  nand g109 (n_236, n_232, n_233, n_234);
  xor g110 (n_235, A[17], B[17]);
  xor g111 (Z[17], n_231, n_235);
  nand g112 (n_237, A[18], B[18]);
  nand g113 (n_238, A[18], n_236);
  nand g114 (n_239, B[18], n_236);
  nand g115 (n_241, n_237, n_238, n_239);
  xor g116 (n_240, A[18], B[18]);
  xor g117 (Z[18], n_236, n_240);
  nand g118 (n_242, A[19], B[19]);
  nand g119 (n_243, A[19], n_241);
  nand g120 (n_244, B[19], n_241);
  nand g121 (n_246, n_242, n_243, n_244);
  xor g122 (n_245, A[19], B[19]);
  xor g123 (Z[19], n_241, n_245);
  nand g124 (n_247, A[20], B[20]);
  nand g125 (n_248, A[20], n_246);
  nand g126 (n_249, B[20], n_246);
  nand g127 (n_251, n_247, n_248, n_249);
  xor g128 (n_250, A[20], B[20]);
  xor g129 (Z[20], n_246, n_250);
  nand g130 (n_252, A[21], B[21]);
  nand g131 (n_253, A[21], n_251);
  nand g132 (n_254, B[21], n_251);
  nand g133 (n_256, n_252, n_253, n_254);
  xor g134 (n_255, A[21], B[21]);
  xor g135 (Z[21], n_251, n_255);
  nand g136 (n_257, A[22], B[22]);
  nand g137 (n_258, A[22], n_256);
  nand g138 (n_259, B[22], n_256);
  nand g139 (n_261, n_257, n_258, n_259);
  xor g140 (n_260, A[22], B[22]);
  xor g141 (Z[22], n_256, n_260);
  nand g142 (n_262, A[23], B[23]);
  nand g143 (n_263, A[23], n_261);
  nand g144 (n_264, B[23], n_261);
  nand g145 (n_266, n_262, n_263, n_264);
  xor g146 (n_265, A[23], B[23]);
  xor g147 (Z[23], n_261, n_265);
  nand g148 (n_267, A[24], B[24]);
  nand g149 (n_268, A[24], n_266);
  nand g150 (n_269, B[24], n_266);
  nand g151 (n_271, n_267, n_268, n_269);
  xor g152 (n_270, A[24], B[24]);
  xor g153 (Z[24], n_266, n_270);
  nand g154 (n_272, A[25], B[25]);
  nand g155 (n_273, A[25], n_271);
  nand g156 (n_274, B[25], n_271);
  nand g157 (n_276, n_272, n_273, n_274);
  xor g158 (n_275, A[25], B[25]);
  xor g159 (Z[25], n_271, n_275);
  nand g160 (n_277, A[26], B[26]);
  nand g161 (n_278, A[26], n_276);
  nand g162 (n_279, B[26], n_276);
  nand g163 (n_281, n_277, n_278, n_279);
  xor g164 (n_280, A[26], B[26]);
  xor g165 (Z[26], n_276, n_280);
  nand g166 (n_282, A[27], B[27]);
  nand g167 (n_283, A[27], n_281);
  nand g168 (n_284, B[27], n_281);
  nand g169 (n_286, n_282, n_283, n_284);
  xor g170 (n_285, A[27], B[27]);
  xor g171 (Z[27], n_281, n_285);
  nand g172 (n_287, A[28], B[28]);
  nand g173 (n_288, A[28], n_286);
  nand g174 (n_289, B[28], n_286);
  nand g175 (n_291, n_287, n_288, n_289);
  xor g176 (n_290, A[28], B[28]);
  xor g177 (Z[28], n_286, n_290);
  nand g178 (n_292, A[29], B[29]);
  nand g179 (n_293, A[29], n_291);
  nand g180 (n_294, B[29], n_291);
  nand g181 (n_296, n_292, n_293, n_294);
  xor g182 (n_295, A[29], B[29]);
  xor g183 (Z[29], n_291, n_295);
  nand g184 (n_297, A[30], B[30]);
  nand g185 (n_298, A[30], n_296);
  nand g186 (n_299, B[30], n_296);
  nand g187 (n_301, n_297, n_298, n_299);
  xor g188 (n_300, A[30], B[30]);
  xor g189 (Z[30], n_296, n_300);
  nand g190 (n_302, A[31], B[31]);
  nand g191 (n_303, A[31], n_301);
  nand g192 (n_304, B[31], n_301);
  nand g193 (n_306, n_302, n_303, n_304);
  xor g194 (n_305, A[31], B[31]);
  xor g195 (Z[31], n_301, n_305);
  nand g196 (n_307, A[32], B[32]);
  nand g197 (n_308, A[32], n_306);
  nand g198 (n_309, B[32], n_306);
  nand g199 (n_311, n_307, n_308, n_309);
  xor g200 (n_310, A[32], B[32]);
  xor g201 (Z[32], n_306, n_310);
  nand g202 (n_312, A[33], B[33]);
  nand g203 (n_313, A[33], n_311);
  nand g204 (n_314, B[33], n_311);
  nand g205 (n_316, n_312, n_313, n_314);
  xor g206 (n_315, A[33], B[33]);
  xor g207 (Z[33], n_311, n_315);
  nand g208 (n_317, A[34], B[34]);
  nand g209 (n_318, A[34], n_316);
  nand g210 (n_319, B[34], n_316);
  nand g211 (n_321, n_317, n_318, n_319);
  xor g212 (n_320, A[34], B[34]);
  xor g213 (Z[34], n_316, n_320);
  nand g214 (n_322, A[35], B[35]);
  nand g215 (n_323, A[35], n_321);
  nand g216 (n_324, B[35], n_321);
  nand g217 (n_326, n_322, n_323, n_324);
  xor g218 (n_325, A[35], B[35]);
  xor g219 (Z[35], n_321, n_325);
  nand g220 (n_327, A[36], B[36]);
  nand g221 (n_328, A[36], n_326);
  nand g222 (n_329, B[36], n_326);
  nand g223 (n_331, n_327, n_328, n_329);
  xor g224 (n_330, A[36], B[36]);
  xor g225 (Z[36], n_326, n_330);
  nand g226 (n_332, A[37], B[37]);
  nand g227 (n_333, A[37], n_331);
  nand g228 (n_334, B[37], n_331);
  nand g229 (n_336, n_332, n_333, n_334);
  xor g230 (n_335, A[37], B[37]);
  xor g231 (Z[37], n_331, n_335);
  nand g232 (n_337, A[38], B[38]);
  nand g233 (n_338, A[38], n_336);
  nand g234 (n_339, B[38], n_336);
  nand g235 (n_341, n_337, n_338, n_339);
  xor g236 (n_340, A[38], B[38]);
  xor g237 (Z[38], n_336, n_340);
  nand g238 (n_342, A[39], B[39]);
  nand g239 (n_343, A[39], n_341);
  nand g240 (n_344, B[39], n_341);
  nand g241 (n_346, n_342, n_343, n_344);
  xor g242 (n_345, A[39], B[39]);
  xor g243 (Z[39], n_341, n_345);
  nand g244 (n_347, A[40], B[40]);
  nand g245 (n_348, A[40], n_346);
  nand g246 (n_349, B[40], n_346);
  nand g247 (n_351, n_347, n_348, n_349);
  xor g248 (n_350, A[40], B[40]);
  xor g249 (Z[40], n_346, n_350);
  nand g250 (n_352, A[41], B[41]);
  nand g251 (n_353, A[41], n_351);
  nand g252 (n_354, B[41], n_351);
  nand g253 (n_356, n_352, n_353, n_354);
  xor g254 (n_355, A[41], B[41]);
  xor g255 (Z[41], n_351, n_355);
  nand g256 (n_357, A[42], B[42]);
  nand g257 (n_358, A[42], n_356);
  nand g258 (n_359, B[42], n_356);
  nand g259 (n_361, n_357, n_358, n_359);
  xor g260 (n_360, A[42], B[42]);
  xor g261 (Z[42], n_356, n_360);
  nand g262 (n_362, A[43], B[43]);
  nand g263 (n_363, A[43], n_361);
  nand g264 (n_364, B[43], n_361);
  nand g265 (n_366, n_362, n_363, n_364);
  xor g266 (n_365, A[43], B[43]);
  xor g267 (Z[43], n_361, n_365);
  nand g268 (n_367, A[44], B[44]);
  nand g269 (n_368, A[44], n_366);
  nand g270 (n_369, B[44], n_366);
  nand g271 (n_371, n_367, n_368, n_369);
  xor g272 (n_370, A[44], B[44]);
  xor g273 (Z[44], n_366, n_370);
  nand g274 (n_372, A[45], B[45]);
  nand g275 (n_373, A[45], n_371);
  nand g276 (n_374, B[45], n_371);
  nand g277 (n_376, n_372, n_373, n_374);
  xor g278 (n_375, A[45], B[45]);
  xor g279 (Z[45], n_371, n_375);
  nand g283 (n_146, n_377, n_378, n_379);
  xor g285 (Z[46], n_376, n_380);
  or g287 (n_377, A[46], B[46]);
  xor g288 (n_380, A[46], B[46]);
  or g289 (n_153, wc, n_147);
  not gc (wc, A[1]);
  or g290 (n_154, wc0, n_147);
  not gc0 (wc0, B[1]);
  xnor g291 (Z[1], n_147, n_155);
  or g292 (n_378, A[46], wc1);
  not gc1 (wc1, n_376);
  or g293 (n_379, B[46], wc2);
  not gc2 (wc2, n_376);
endmodule

module add_signed_356_2_GENERIC(A, B, Z);
  input [46:0] A, B;
  output [47:0] Z;
  wire [46:0] A, B;
  wire [47:0] Z;
  add_signed_356_2_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3603_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [61:0] A, B;
  output [62:0] Z;
  wire [61:0] A, B;
  wire [62:0] Z;
  wire n_191, n_192, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500;
  not g3 (Z[62], n_191);
  nand g4 (n_192, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_197, A[1], B[1]);
  nand g13 (n_201, n_197, n_198, n_199);
  xor g14 (n_200, A[1], B[1]);
  nand g16 (n_202, A[2], B[2]);
  nand g17 (n_203, A[2], n_201);
  nand g18 (n_204, B[2], n_201);
  nand g19 (n_206, n_202, n_203, n_204);
  xor g20 (n_205, A[2], B[2]);
  xor g21 (Z[2], n_201, n_205);
  nand g22 (n_207, A[3], B[3]);
  nand g23 (n_208, A[3], n_206);
  nand g24 (n_209, B[3], n_206);
  nand g25 (n_211, n_207, n_208, n_209);
  xor g26 (n_210, A[3], B[3]);
  xor g27 (Z[3], n_206, n_210);
  nand g28 (n_212, A[4], B[4]);
  nand g29 (n_213, A[4], n_211);
  nand g30 (n_214, B[4], n_211);
  nand g31 (n_216, n_212, n_213, n_214);
  xor g32 (n_215, A[4], B[4]);
  xor g33 (Z[4], n_211, n_215);
  nand g34 (n_217, A[5], B[5]);
  nand g35 (n_218, A[5], n_216);
  nand g36 (n_219, B[5], n_216);
  nand g37 (n_221, n_217, n_218, n_219);
  xor g38 (n_220, A[5], B[5]);
  xor g39 (Z[5], n_216, n_220);
  nand g40 (n_222, A[6], B[6]);
  nand g41 (n_223, A[6], n_221);
  nand g42 (n_224, B[6], n_221);
  nand g43 (n_226, n_222, n_223, n_224);
  xor g44 (n_225, A[6], B[6]);
  xor g45 (Z[6], n_221, n_225);
  nand g46 (n_227, A[7], B[7]);
  nand g47 (n_228, A[7], n_226);
  nand g48 (n_229, B[7], n_226);
  nand g49 (n_231, n_227, n_228, n_229);
  xor g50 (n_230, A[7], B[7]);
  xor g51 (Z[7], n_226, n_230);
  nand g52 (n_232, A[8], B[8]);
  nand g53 (n_233, A[8], n_231);
  nand g54 (n_234, B[8], n_231);
  nand g55 (n_236, n_232, n_233, n_234);
  xor g56 (n_235, A[8], B[8]);
  xor g57 (Z[8], n_231, n_235);
  nand g58 (n_237, A[9], B[9]);
  nand g59 (n_238, A[9], n_236);
  nand g60 (n_239, B[9], n_236);
  nand g61 (n_241, n_237, n_238, n_239);
  xor g62 (n_240, A[9], B[9]);
  xor g63 (Z[9], n_236, n_240);
  nand g64 (n_242, A[10], B[10]);
  nand g65 (n_243, A[10], n_241);
  nand g66 (n_244, B[10], n_241);
  nand g67 (n_246, n_242, n_243, n_244);
  xor g68 (n_245, A[10], B[10]);
  xor g69 (Z[10], n_241, n_245);
  nand g70 (n_247, A[11], B[11]);
  nand g71 (n_248, A[11], n_246);
  nand g72 (n_249, B[11], n_246);
  nand g73 (n_251, n_247, n_248, n_249);
  xor g74 (n_250, A[11], B[11]);
  xor g75 (Z[11], n_246, n_250);
  nand g76 (n_252, A[12], B[12]);
  nand g77 (n_253, A[12], n_251);
  nand g78 (n_254, B[12], n_251);
  nand g79 (n_256, n_252, n_253, n_254);
  xor g80 (n_255, A[12], B[12]);
  xor g81 (Z[12], n_251, n_255);
  nand g82 (n_257, A[13], B[13]);
  nand g83 (n_258, A[13], n_256);
  nand g84 (n_259, B[13], n_256);
  nand g85 (n_261, n_257, n_258, n_259);
  xor g86 (n_260, A[13], B[13]);
  xor g87 (Z[13], n_256, n_260);
  nand g88 (n_262, A[14], B[14]);
  nand g89 (n_263, A[14], n_261);
  nand g90 (n_264, B[14], n_261);
  nand g91 (n_266, n_262, n_263, n_264);
  xor g92 (n_265, A[14], B[14]);
  xor g93 (Z[14], n_261, n_265);
  nand g94 (n_267, A[15], B[15]);
  nand g95 (n_268, A[15], n_266);
  nand g96 (n_269, B[15], n_266);
  nand g97 (n_271, n_267, n_268, n_269);
  xor g98 (n_270, A[15], B[15]);
  xor g99 (Z[15], n_266, n_270);
  nand g100 (n_272, A[16], B[16]);
  nand g101 (n_273, A[16], n_271);
  nand g102 (n_274, B[16], n_271);
  nand g103 (n_276, n_272, n_273, n_274);
  xor g104 (n_275, A[16], B[16]);
  xor g105 (Z[16], n_271, n_275);
  nand g106 (n_277, A[17], B[17]);
  nand g107 (n_278, A[17], n_276);
  nand g108 (n_279, B[17], n_276);
  nand g109 (n_281, n_277, n_278, n_279);
  xor g110 (n_280, A[17], B[17]);
  xor g111 (Z[17], n_276, n_280);
  nand g112 (n_282, A[18], B[18]);
  nand g113 (n_283, A[18], n_281);
  nand g114 (n_284, B[18], n_281);
  nand g115 (n_286, n_282, n_283, n_284);
  xor g116 (n_285, A[18], B[18]);
  xor g117 (Z[18], n_281, n_285);
  nand g118 (n_287, A[19], B[19]);
  nand g119 (n_288, A[19], n_286);
  nand g120 (n_289, B[19], n_286);
  nand g121 (n_291, n_287, n_288, n_289);
  xor g122 (n_290, A[19], B[19]);
  xor g123 (Z[19], n_286, n_290);
  nand g124 (n_292, A[20], B[20]);
  nand g125 (n_293, A[20], n_291);
  nand g126 (n_294, B[20], n_291);
  nand g127 (n_296, n_292, n_293, n_294);
  xor g128 (n_295, A[20], B[20]);
  xor g129 (Z[20], n_291, n_295);
  nand g130 (n_297, A[21], B[21]);
  nand g131 (n_298, A[21], n_296);
  nand g132 (n_299, B[21], n_296);
  nand g133 (n_301, n_297, n_298, n_299);
  xor g134 (n_300, A[21], B[21]);
  xor g135 (Z[21], n_296, n_300);
  nand g136 (n_302, A[22], B[22]);
  nand g137 (n_303, A[22], n_301);
  nand g138 (n_304, B[22], n_301);
  nand g139 (n_306, n_302, n_303, n_304);
  xor g140 (n_305, A[22], B[22]);
  xor g141 (Z[22], n_301, n_305);
  nand g142 (n_307, A[23], B[23]);
  nand g143 (n_308, A[23], n_306);
  nand g144 (n_309, B[23], n_306);
  nand g145 (n_311, n_307, n_308, n_309);
  xor g146 (n_310, A[23], B[23]);
  xor g147 (Z[23], n_306, n_310);
  nand g148 (n_312, A[24], B[24]);
  nand g149 (n_313, A[24], n_311);
  nand g150 (n_314, B[24], n_311);
  nand g151 (n_316, n_312, n_313, n_314);
  xor g152 (n_315, A[24], B[24]);
  xor g153 (Z[24], n_311, n_315);
  nand g154 (n_317, A[25], B[25]);
  nand g155 (n_318, A[25], n_316);
  nand g156 (n_319, B[25], n_316);
  nand g157 (n_321, n_317, n_318, n_319);
  xor g158 (n_320, A[25], B[25]);
  xor g159 (Z[25], n_316, n_320);
  nand g160 (n_322, A[26], B[26]);
  nand g161 (n_323, A[26], n_321);
  nand g162 (n_324, B[26], n_321);
  nand g163 (n_326, n_322, n_323, n_324);
  xor g164 (n_325, A[26], B[26]);
  xor g165 (Z[26], n_321, n_325);
  nand g166 (n_327, A[27], B[27]);
  nand g167 (n_328, A[27], n_326);
  nand g168 (n_329, B[27], n_326);
  nand g169 (n_331, n_327, n_328, n_329);
  xor g170 (n_330, A[27], B[27]);
  xor g171 (Z[27], n_326, n_330);
  nand g172 (n_332, A[28], B[28]);
  nand g173 (n_333, A[28], n_331);
  nand g174 (n_334, B[28], n_331);
  nand g175 (n_336, n_332, n_333, n_334);
  xor g176 (n_335, A[28], B[28]);
  xor g177 (Z[28], n_331, n_335);
  nand g178 (n_337, A[29], B[29]);
  nand g179 (n_338, A[29], n_336);
  nand g180 (n_339, B[29], n_336);
  nand g181 (n_341, n_337, n_338, n_339);
  xor g182 (n_340, A[29], B[29]);
  xor g183 (Z[29], n_336, n_340);
  nand g184 (n_342, A[30], B[30]);
  nand g185 (n_343, A[30], n_341);
  nand g186 (n_344, B[30], n_341);
  nand g187 (n_346, n_342, n_343, n_344);
  xor g188 (n_345, A[30], B[30]);
  xor g189 (Z[30], n_341, n_345);
  nand g190 (n_347, A[31], B[31]);
  nand g191 (n_348, A[31], n_346);
  nand g192 (n_349, B[31], n_346);
  nand g193 (n_351, n_347, n_348, n_349);
  xor g194 (n_350, A[31], B[31]);
  xor g195 (Z[31], n_346, n_350);
  nand g196 (n_352, A[32], B[32]);
  nand g197 (n_353, A[32], n_351);
  nand g198 (n_354, B[32], n_351);
  nand g199 (n_356, n_352, n_353, n_354);
  xor g200 (n_355, A[32], B[32]);
  xor g201 (Z[32], n_351, n_355);
  nand g202 (n_357, A[33], B[33]);
  nand g203 (n_358, A[33], n_356);
  nand g204 (n_359, B[33], n_356);
  nand g205 (n_361, n_357, n_358, n_359);
  xor g206 (n_360, A[33], B[33]);
  xor g207 (Z[33], n_356, n_360);
  nand g208 (n_362, A[34], B[34]);
  nand g209 (n_363, A[34], n_361);
  nand g210 (n_364, B[34], n_361);
  nand g211 (n_366, n_362, n_363, n_364);
  xor g212 (n_365, A[34], B[34]);
  xor g213 (Z[34], n_361, n_365);
  nand g214 (n_367, A[35], B[35]);
  nand g215 (n_368, A[35], n_366);
  nand g216 (n_369, B[35], n_366);
  nand g217 (n_371, n_367, n_368, n_369);
  xor g218 (n_370, A[35], B[35]);
  xor g219 (Z[35], n_366, n_370);
  nand g220 (n_372, A[36], B[36]);
  nand g221 (n_373, A[36], n_371);
  nand g222 (n_374, B[36], n_371);
  nand g223 (n_376, n_372, n_373, n_374);
  xor g224 (n_375, A[36], B[36]);
  xor g225 (Z[36], n_371, n_375);
  nand g226 (n_377, A[37], B[37]);
  nand g227 (n_378, A[37], n_376);
  nand g228 (n_379, B[37], n_376);
  nand g229 (n_381, n_377, n_378, n_379);
  xor g230 (n_380, A[37], B[37]);
  xor g231 (Z[37], n_376, n_380);
  nand g232 (n_382, A[38], B[38]);
  nand g233 (n_383, A[38], n_381);
  nand g234 (n_384, B[38], n_381);
  nand g235 (n_386, n_382, n_383, n_384);
  xor g236 (n_385, A[38], B[38]);
  xor g237 (Z[38], n_381, n_385);
  nand g238 (n_387, A[39], B[39]);
  nand g239 (n_388, A[39], n_386);
  nand g240 (n_389, B[39], n_386);
  nand g241 (n_391, n_387, n_388, n_389);
  xor g242 (n_390, A[39], B[39]);
  xor g243 (Z[39], n_386, n_390);
  nand g244 (n_392, A[40], B[40]);
  nand g245 (n_393, A[40], n_391);
  nand g246 (n_394, B[40], n_391);
  nand g247 (n_396, n_392, n_393, n_394);
  xor g248 (n_395, A[40], B[40]);
  xor g249 (Z[40], n_391, n_395);
  nand g250 (n_397, A[41], B[41]);
  nand g251 (n_398, A[41], n_396);
  nand g252 (n_399, B[41], n_396);
  nand g253 (n_401, n_397, n_398, n_399);
  xor g254 (n_400, A[41], B[41]);
  xor g255 (Z[41], n_396, n_400);
  nand g256 (n_402, A[42], B[42]);
  nand g257 (n_403, A[42], n_401);
  nand g258 (n_404, B[42], n_401);
  nand g259 (n_406, n_402, n_403, n_404);
  xor g260 (n_405, A[42], B[42]);
  xor g261 (Z[42], n_401, n_405);
  nand g262 (n_407, A[43], B[43]);
  nand g263 (n_408, A[43], n_406);
  nand g264 (n_409, B[43], n_406);
  nand g265 (n_411, n_407, n_408, n_409);
  xor g266 (n_410, A[43], B[43]);
  xor g267 (Z[43], n_406, n_410);
  nand g268 (n_412, A[44], B[44]);
  nand g269 (n_413, A[44], n_411);
  nand g270 (n_414, B[44], n_411);
  nand g271 (n_416, n_412, n_413, n_414);
  xor g272 (n_415, A[44], B[44]);
  xor g273 (Z[44], n_411, n_415);
  nand g274 (n_417, A[45], B[45]);
  nand g275 (n_418, A[45], n_416);
  nand g276 (n_419, B[45], n_416);
  nand g277 (n_421, n_417, n_418, n_419);
  xor g278 (n_420, A[45], B[45]);
  xor g279 (Z[45], n_416, n_420);
  nand g280 (n_422, A[46], B[46]);
  nand g281 (n_423, A[46], n_421);
  nand g282 (n_424, B[46], n_421);
  nand g283 (n_426, n_422, n_423, n_424);
  xor g284 (n_425, A[46], B[46]);
  xor g285 (Z[46], n_421, n_425);
  nand g286 (n_427, A[47], B[47]);
  nand g287 (n_428, A[47], n_426);
  nand g288 (n_429, B[47], n_426);
  nand g289 (n_431, n_427, n_428, n_429);
  xor g290 (n_430, A[47], B[47]);
  xor g291 (Z[47], n_426, n_430);
  nand g292 (n_432, A[48], B[48]);
  nand g293 (n_433, A[48], n_431);
  nand g294 (n_434, B[48], n_431);
  nand g295 (n_436, n_432, n_433, n_434);
  xor g296 (n_435, A[48], B[48]);
  xor g297 (Z[48], n_431, n_435);
  nand g298 (n_437, A[49], B[49]);
  nand g299 (n_438, A[49], n_436);
  nand g300 (n_439, B[49], n_436);
  nand g301 (n_441, n_437, n_438, n_439);
  xor g302 (n_440, A[49], B[49]);
  xor g303 (Z[49], n_436, n_440);
  nand g304 (n_442, A[50], B[50]);
  nand g305 (n_443, A[50], n_441);
  nand g306 (n_444, B[50], n_441);
  nand g307 (n_446, n_442, n_443, n_444);
  xor g308 (n_445, A[50], B[50]);
  xor g309 (Z[50], n_441, n_445);
  nand g310 (n_447, A[51], B[51]);
  nand g311 (n_448, A[51], n_446);
  nand g312 (n_449, B[51], n_446);
  nand g313 (n_451, n_447, n_448, n_449);
  xor g314 (n_450, A[51], B[51]);
  xor g315 (Z[51], n_446, n_450);
  nand g316 (n_452, A[52], B[52]);
  nand g317 (n_453, A[52], n_451);
  nand g318 (n_454, B[52], n_451);
  nand g319 (n_456, n_452, n_453, n_454);
  xor g320 (n_455, A[52], B[52]);
  xor g321 (Z[52], n_451, n_455);
  nand g322 (n_457, A[53], B[53]);
  nand g323 (n_458, A[53], n_456);
  nand g324 (n_459, B[53], n_456);
  nand g325 (n_461, n_457, n_458, n_459);
  xor g326 (n_460, A[53], B[53]);
  xor g327 (Z[53], n_456, n_460);
  nand g328 (n_462, A[54], B[54]);
  nand g329 (n_463, A[54], n_461);
  nand g330 (n_464, B[54], n_461);
  nand g331 (n_466, n_462, n_463, n_464);
  xor g332 (n_465, A[54], B[54]);
  xor g333 (Z[54], n_461, n_465);
  nand g334 (n_467, A[55], B[55]);
  nand g335 (n_468, A[55], n_466);
  nand g336 (n_469, B[55], n_466);
  nand g337 (n_471, n_467, n_468, n_469);
  xor g338 (n_470, A[55], B[55]);
  xor g339 (Z[55], n_466, n_470);
  nand g340 (n_472, A[56], B[56]);
  nand g341 (n_473, A[56], n_471);
  nand g342 (n_474, B[56], n_471);
  nand g343 (n_476, n_472, n_473, n_474);
  xor g344 (n_475, A[56], B[56]);
  xor g345 (Z[56], n_471, n_475);
  nand g346 (n_477, A[57], B[57]);
  nand g347 (n_478, A[57], n_476);
  nand g348 (n_479, B[57], n_476);
  nand g349 (n_481, n_477, n_478, n_479);
  xor g350 (n_480, A[57], B[57]);
  xor g351 (Z[57], n_476, n_480);
  nand g352 (n_482, A[58], B[58]);
  nand g353 (n_483, A[58], n_481);
  nand g354 (n_484, B[58], n_481);
  nand g355 (n_486, n_482, n_483, n_484);
  xor g356 (n_485, A[58], B[58]);
  xor g357 (Z[58], n_481, n_485);
  nand g358 (n_487, A[59], B[59]);
  nand g359 (n_488, A[59], n_486);
  nand g360 (n_489, B[59], n_486);
  nand g361 (n_491, n_487, n_488, n_489);
  xor g362 (n_490, A[59], B[59]);
  xor g363 (Z[59], n_486, n_490);
  nand g364 (n_492, A[60], B[60]);
  nand g365 (n_493, A[60], n_491);
  nand g366 (n_494, B[60], n_491);
  nand g367 (n_496, n_492, n_493, n_494);
  xor g368 (n_495, A[60], B[60]);
  xor g369 (Z[60], n_491, n_495);
  nand g373 (n_191, n_497, n_498, n_499);
  xor g375 (Z[61], n_496, n_500);
  or g377 (n_497, A[61], B[61]);
  xor g378 (n_500, A[61], B[61]);
  or g379 (n_198, wc, n_192);
  not gc (wc, A[1]);
  or g380 (n_199, wc0, n_192);
  not gc0 (wc0, B[1]);
  xnor g381 (Z[1], n_192, n_200);
  or g382 (n_498, A[61], wc1);
  not gc1 (wc1, n_496);
  or g383 (n_499, B[61], wc2);
  not gc2 (wc2, n_496);
endmodule

module add_signed_3603_GENERIC(A, B, Z);
  input [61:0] A, B;
  output [62:0] Z;
  wire [61:0] A, B;
  wire [62:0] Z;
  add_signed_3603_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3603_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [61:0] A, B;
  output [62:0] Z;
  wire [61:0] A, B;
  wire [62:0] Z;
  wire n_191, n_192, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500;
  not g3 (Z[62], n_191);
  nand g4 (n_192, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_197, A[1], B[1]);
  nand g13 (n_201, n_197, n_198, n_199);
  xor g14 (n_200, A[1], B[1]);
  nand g16 (n_202, A[2], B[2]);
  nand g17 (n_203, A[2], n_201);
  nand g18 (n_204, B[2], n_201);
  nand g19 (n_206, n_202, n_203, n_204);
  xor g20 (n_205, A[2], B[2]);
  xor g21 (Z[2], n_201, n_205);
  nand g22 (n_207, A[3], B[3]);
  nand g23 (n_208, A[3], n_206);
  nand g24 (n_209, B[3], n_206);
  nand g25 (n_211, n_207, n_208, n_209);
  xor g26 (n_210, A[3], B[3]);
  xor g27 (Z[3], n_206, n_210);
  nand g28 (n_212, A[4], B[4]);
  nand g29 (n_213, A[4], n_211);
  nand g30 (n_214, B[4], n_211);
  nand g31 (n_216, n_212, n_213, n_214);
  xor g32 (n_215, A[4], B[4]);
  xor g33 (Z[4], n_211, n_215);
  nand g34 (n_217, A[5], B[5]);
  nand g35 (n_218, A[5], n_216);
  nand g36 (n_219, B[5], n_216);
  nand g37 (n_221, n_217, n_218, n_219);
  xor g38 (n_220, A[5], B[5]);
  xor g39 (Z[5], n_216, n_220);
  nand g40 (n_222, A[6], B[6]);
  nand g41 (n_223, A[6], n_221);
  nand g42 (n_224, B[6], n_221);
  nand g43 (n_226, n_222, n_223, n_224);
  xor g44 (n_225, A[6], B[6]);
  xor g45 (Z[6], n_221, n_225);
  nand g46 (n_227, A[7], B[7]);
  nand g47 (n_228, A[7], n_226);
  nand g48 (n_229, B[7], n_226);
  nand g49 (n_231, n_227, n_228, n_229);
  xor g50 (n_230, A[7], B[7]);
  xor g51 (Z[7], n_226, n_230);
  nand g52 (n_232, A[8], B[8]);
  nand g53 (n_233, A[8], n_231);
  nand g54 (n_234, B[8], n_231);
  nand g55 (n_236, n_232, n_233, n_234);
  xor g56 (n_235, A[8], B[8]);
  xor g57 (Z[8], n_231, n_235);
  nand g58 (n_237, A[9], B[9]);
  nand g59 (n_238, A[9], n_236);
  nand g60 (n_239, B[9], n_236);
  nand g61 (n_241, n_237, n_238, n_239);
  xor g62 (n_240, A[9], B[9]);
  xor g63 (Z[9], n_236, n_240);
  nand g64 (n_242, A[10], B[10]);
  nand g65 (n_243, A[10], n_241);
  nand g66 (n_244, B[10], n_241);
  nand g67 (n_246, n_242, n_243, n_244);
  xor g68 (n_245, A[10], B[10]);
  xor g69 (Z[10], n_241, n_245);
  nand g70 (n_247, A[11], B[11]);
  nand g71 (n_248, A[11], n_246);
  nand g72 (n_249, B[11], n_246);
  nand g73 (n_251, n_247, n_248, n_249);
  xor g74 (n_250, A[11], B[11]);
  xor g75 (Z[11], n_246, n_250);
  nand g76 (n_252, A[12], B[12]);
  nand g77 (n_253, A[12], n_251);
  nand g78 (n_254, B[12], n_251);
  nand g79 (n_256, n_252, n_253, n_254);
  xor g80 (n_255, A[12], B[12]);
  xor g81 (Z[12], n_251, n_255);
  nand g82 (n_257, A[13], B[13]);
  nand g83 (n_258, A[13], n_256);
  nand g84 (n_259, B[13], n_256);
  nand g85 (n_261, n_257, n_258, n_259);
  xor g86 (n_260, A[13], B[13]);
  xor g87 (Z[13], n_256, n_260);
  nand g88 (n_262, A[14], B[14]);
  nand g89 (n_263, A[14], n_261);
  nand g90 (n_264, B[14], n_261);
  nand g91 (n_266, n_262, n_263, n_264);
  xor g92 (n_265, A[14], B[14]);
  xor g93 (Z[14], n_261, n_265);
  nand g94 (n_267, A[15], B[15]);
  nand g95 (n_268, A[15], n_266);
  nand g96 (n_269, B[15], n_266);
  nand g97 (n_271, n_267, n_268, n_269);
  xor g98 (n_270, A[15], B[15]);
  xor g99 (Z[15], n_266, n_270);
  nand g100 (n_272, A[16], B[16]);
  nand g101 (n_273, A[16], n_271);
  nand g102 (n_274, B[16], n_271);
  nand g103 (n_276, n_272, n_273, n_274);
  xor g104 (n_275, A[16], B[16]);
  xor g105 (Z[16], n_271, n_275);
  nand g106 (n_277, A[17], B[17]);
  nand g107 (n_278, A[17], n_276);
  nand g108 (n_279, B[17], n_276);
  nand g109 (n_281, n_277, n_278, n_279);
  xor g110 (n_280, A[17], B[17]);
  xor g111 (Z[17], n_276, n_280);
  nand g112 (n_282, A[18], B[18]);
  nand g113 (n_283, A[18], n_281);
  nand g114 (n_284, B[18], n_281);
  nand g115 (n_286, n_282, n_283, n_284);
  xor g116 (n_285, A[18], B[18]);
  xor g117 (Z[18], n_281, n_285);
  nand g118 (n_287, A[19], B[19]);
  nand g119 (n_288, A[19], n_286);
  nand g120 (n_289, B[19], n_286);
  nand g121 (n_291, n_287, n_288, n_289);
  xor g122 (n_290, A[19], B[19]);
  xor g123 (Z[19], n_286, n_290);
  nand g124 (n_292, A[20], B[20]);
  nand g125 (n_293, A[20], n_291);
  nand g126 (n_294, B[20], n_291);
  nand g127 (n_296, n_292, n_293, n_294);
  xor g128 (n_295, A[20], B[20]);
  xor g129 (Z[20], n_291, n_295);
  nand g130 (n_297, A[21], B[21]);
  nand g131 (n_298, A[21], n_296);
  nand g132 (n_299, B[21], n_296);
  nand g133 (n_301, n_297, n_298, n_299);
  xor g134 (n_300, A[21], B[21]);
  xor g135 (Z[21], n_296, n_300);
  nand g136 (n_302, A[22], B[22]);
  nand g137 (n_303, A[22], n_301);
  nand g138 (n_304, B[22], n_301);
  nand g139 (n_306, n_302, n_303, n_304);
  xor g140 (n_305, A[22], B[22]);
  xor g141 (Z[22], n_301, n_305);
  nand g142 (n_307, A[23], B[23]);
  nand g143 (n_308, A[23], n_306);
  nand g144 (n_309, B[23], n_306);
  nand g145 (n_311, n_307, n_308, n_309);
  xor g146 (n_310, A[23], B[23]);
  xor g147 (Z[23], n_306, n_310);
  nand g148 (n_312, A[24], B[24]);
  nand g149 (n_313, A[24], n_311);
  nand g150 (n_314, B[24], n_311);
  nand g151 (n_316, n_312, n_313, n_314);
  xor g152 (n_315, A[24], B[24]);
  xor g153 (Z[24], n_311, n_315);
  nand g154 (n_317, A[25], B[25]);
  nand g155 (n_318, A[25], n_316);
  nand g156 (n_319, B[25], n_316);
  nand g157 (n_321, n_317, n_318, n_319);
  xor g158 (n_320, A[25], B[25]);
  xor g159 (Z[25], n_316, n_320);
  nand g160 (n_322, A[26], B[26]);
  nand g161 (n_323, A[26], n_321);
  nand g162 (n_324, B[26], n_321);
  nand g163 (n_326, n_322, n_323, n_324);
  xor g164 (n_325, A[26], B[26]);
  xor g165 (Z[26], n_321, n_325);
  nand g166 (n_327, A[27], B[27]);
  nand g167 (n_328, A[27], n_326);
  nand g168 (n_329, B[27], n_326);
  nand g169 (n_331, n_327, n_328, n_329);
  xor g170 (n_330, A[27], B[27]);
  xor g171 (Z[27], n_326, n_330);
  nand g172 (n_332, A[28], B[28]);
  nand g173 (n_333, A[28], n_331);
  nand g174 (n_334, B[28], n_331);
  nand g175 (n_336, n_332, n_333, n_334);
  xor g176 (n_335, A[28], B[28]);
  xor g177 (Z[28], n_331, n_335);
  nand g178 (n_337, A[29], B[29]);
  nand g179 (n_338, A[29], n_336);
  nand g180 (n_339, B[29], n_336);
  nand g181 (n_341, n_337, n_338, n_339);
  xor g182 (n_340, A[29], B[29]);
  xor g183 (Z[29], n_336, n_340);
  nand g184 (n_342, A[30], B[30]);
  nand g185 (n_343, A[30], n_341);
  nand g186 (n_344, B[30], n_341);
  nand g187 (n_346, n_342, n_343, n_344);
  xor g188 (n_345, A[30], B[30]);
  xor g189 (Z[30], n_341, n_345);
  nand g190 (n_347, A[31], B[31]);
  nand g191 (n_348, A[31], n_346);
  nand g192 (n_349, B[31], n_346);
  nand g193 (n_351, n_347, n_348, n_349);
  xor g194 (n_350, A[31], B[31]);
  xor g195 (Z[31], n_346, n_350);
  nand g196 (n_352, A[32], B[32]);
  nand g197 (n_353, A[32], n_351);
  nand g198 (n_354, B[32], n_351);
  nand g199 (n_356, n_352, n_353, n_354);
  xor g200 (n_355, A[32], B[32]);
  xor g201 (Z[32], n_351, n_355);
  nand g202 (n_357, A[33], B[33]);
  nand g203 (n_358, A[33], n_356);
  nand g204 (n_359, B[33], n_356);
  nand g205 (n_361, n_357, n_358, n_359);
  xor g206 (n_360, A[33], B[33]);
  xor g207 (Z[33], n_356, n_360);
  nand g208 (n_362, A[34], B[34]);
  nand g209 (n_363, A[34], n_361);
  nand g210 (n_364, B[34], n_361);
  nand g211 (n_366, n_362, n_363, n_364);
  xor g212 (n_365, A[34], B[34]);
  xor g213 (Z[34], n_361, n_365);
  nand g214 (n_367, A[35], B[35]);
  nand g215 (n_368, A[35], n_366);
  nand g216 (n_369, B[35], n_366);
  nand g217 (n_371, n_367, n_368, n_369);
  xor g218 (n_370, A[35], B[35]);
  xor g219 (Z[35], n_366, n_370);
  nand g220 (n_372, A[36], B[36]);
  nand g221 (n_373, A[36], n_371);
  nand g222 (n_374, B[36], n_371);
  nand g223 (n_376, n_372, n_373, n_374);
  xor g224 (n_375, A[36], B[36]);
  xor g225 (Z[36], n_371, n_375);
  nand g226 (n_377, A[37], B[37]);
  nand g227 (n_378, A[37], n_376);
  nand g228 (n_379, B[37], n_376);
  nand g229 (n_381, n_377, n_378, n_379);
  xor g230 (n_380, A[37], B[37]);
  xor g231 (Z[37], n_376, n_380);
  nand g232 (n_382, A[38], B[38]);
  nand g233 (n_383, A[38], n_381);
  nand g234 (n_384, B[38], n_381);
  nand g235 (n_386, n_382, n_383, n_384);
  xor g236 (n_385, A[38], B[38]);
  xor g237 (Z[38], n_381, n_385);
  nand g238 (n_387, A[39], B[39]);
  nand g239 (n_388, A[39], n_386);
  nand g240 (n_389, B[39], n_386);
  nand g241 (n_391, n_387, n_388, n_389);
  xor g242 (n_390, A[39], B[39]);
  xor g243 (Z[39], n_386, n_390);
  nand g244 (n_392, A[40], B[40]);
  nand g245 (n_393, A[40], n_391);
  nand g246 (n_394, B[40], n_391);
  nand g247 (n_396, n_392, n_393, n_394);
  xor g248 (n_395, A[40], B[40]);
  xor g249 (Z[40], n_391, n_395);
  nand g250 (n_397, A[41], B[41]);
  nand g251 (n_398, A[41], n_396);
  nand g252 (n_399, B[41], n_396);
  nand g253 (n_401, n_397, n_398, n_399);
  xor g254 (n_400, A[41], B[41]);
  xor g255 (Z[41], n_396, n_400);
  nand g256 (n_402, A[42], B[42]);
  nand g257 (n_403, A[42], n_401);
  nand g258 (n_404, B[42], n_401);
  nand g259 (n_406, n_402, n_403, n_404);
  xor g260 (n_405, A[42], B[42]);
  xor g261 (Z[42], n_401, n_405);
  nand g262 (n_407, A[43], B[43]);
  nand g263 (n_408, A[43], n_406);
  nand g264 (n_409, B[43], n_406);
  nand g265 (n_411, n_407, n_408, n_409);
  xor g266 (n_410, A[43], B[43]);
  xor g267 (Z[43], n_406, n_410);
  nand g268 (n_412, A[44], B[44]);
  nand g269 (n_413, A[44], n_411);
  nand g270 (n_414, B[44], n_411);
  nand g271 (n_416, n_412, n_413, n_414);
  xor g272 (n_415, A[44], B[44]);
  xor g273 (Z[44], n_411, n_415);
  nand g274 (n_417, A[45], B[45]);
  nand g275 (n_418, A[45], n_416);
  nand g276 (n_419, B[45], n_416);
  nand g277 (n_421, n_417, n_418, n_419);
  xor g278 (n_420, A[45], B[45]);
  xor g279 (Z[45], n_416, n_420);
  nand g280 (n_422, A[46], B[46]);
  nand g281 (n_423, A[46], n_421);
  nand g282 (n_424, B[46], n_421);
  nand g283 (n_426, n_422, n_423, n_424);
  xor g284 (n_425, A[46], B[46]);
  xor g285 (Z[46], n_421, n_425);
  nand g286 (n_427, A[47], B[47]);
  nand g287 (n_428, A[47], n_426);
  nand g288 (n_429, B[47], n_426);
  nand g289 (n_431, n_427, n_428, n_429);
  xor g290 (n_430, A[47], B[47]);
  xor g291 (Z[47], n_426, n_430);
  nand g292 (n_432, A[48], B[48]);
  nand g293 (n_433, A[48], n_431);
  nand g294 (n_434, B[48], n_431);
  nand g295 (n_436, n_432, n_433, n_434);
  xor g296 (n_435, A[48], B[48]);
  xor g297 (Z[48], n_431, n_435);
  nand g298 (n_437, A[49], B[49]);
  nand g299 (n_438, A[49], n_436);
  nand g300 (n_439, B[49], n_436);
  nand g301 (n_441, n_437, n_438, n_439);
  xor g302 (n_440, A[49], B[49]);
  xor g303 (Z[49], n_436, n_440);
  nand g304 (n_442, A[50], B[50]);
  nand g305 (n_443, A[50], n_441);
  nand g306 (n_444, B[50], n_441);
  nand g307 (n_446, n_442, n_443, n_444);
  xor g308 (n_445, A[50], B[50]);
  xor g309 (Z[50], n_441, n_445);
  nand g310 (n_447, A[51], B[51]);
  nand g311 (n_448, A[51], n_446);
  nand g312 (n_449, B[51], n_446);
  nand g313 (n_451, n_447, n_448, n_449);
  xor g314 (n_450, A[51], B[51]);
  xor g315 (Z[51], n_446, n_450);
  nand g316 (n_452, A[52], B[52]);
  nand g317 (n_453, A[52], n_451);
  nand g318 (n_454, B[52], n_451);
  nand g319 (n_456, n_452, n_453, n_454);
  xor g320 (n_455, A[52], B[52]);
  xor g321 (Z[52], n_451, n_455);
  nand g322 (n_457, A[53], B[53]);
  nand g323 (n_458, A[53], n_456);
  nand g324 (n_459, B[53], n_456);
  nand g325 (n_461, n_457, n_458, n_459);
  xor g326 (n_460, A[53], B[53]);
  xor g327 (Z[53], n_456, n_460);
  nand g328 (n_462, A[54], B[54]);
  nand g329 (n_463, A[54], n_461);
  nand g330 (n_464, B[54], n_461);
  nand g331 (n_466, n_462, n_463, n_464);
  xor g332 (n_465, A[54], B[54]);
  xor g333 (Z[54], n_461, n_465);
  nand g334 (n_467, A[55], B[55]);
  nand g335 (n_468, A[55], n_466);
  nand g336 (n_469, B[55], n_466);
  nand g337 (n_471, n_467, n_468, n_469);
  xor g338 (n_470, A[55], B[55]);
  xor g339 (Z[55], n_466, n_470);
  nand g340 (n_472, A[56], B[56]);
  nand g341 (n_473, A[56], n_471);
  nand g342 (n_474, B[56], n_471);
  nand g343 (n_476, n_472, n_473, n_474);
  xor g344 (n_475, A[56], B[56]);
  xor g345 (Z[56], n_471, n_475);
  nand g346 (n_477, A[57], B[57]);
  nand g347 (n_478, A[57], n_476);
  nand g348 (n_479, B[57], n_476);
  nand g349 (n_481, n_477, n_478, n_479);
  xor g350 (n_480, A[57], B[57]);
  xor g351 (Z[57], n_476, n_480);
  nand g352 (n_482, A[58], B[58]);
  nand g353 (n_483, A[58], n_481);
  nand g354 (n_484, B[58], n_481);
  nand g355 (n_486, n_482, n_483, n_484);
  xor g356 (n_485, A[58], B[58]);
  xor g357 (Z[58], n_481, n_485);
  nand g358 (n_487, A[59], B[59]);
  nand g359 (n_488, A[59], n_486);
  nand g360 (n_489, B[59], n_486);
  nand g361 (n_491, n_487, n_488, n_489);
  xor g362 (n_490, A[59], B[59]);
  xor g363 (Z[59], n_486, n_490);
  nand g364 (n_492, A[60], B[60]);
  nand g365 (n_493, A[60], n_491);
  nand g366 (n_494, B[60], n_491);
  nand g367 (n_496, n_492, n_493, n_494);
  xor g368 (n_495, A[60], B[60]);
  xor g369 (Z[60], n_491, n_495);
  nand g373 (n_191, n_497, n_498, n_499);
  xor g375 (Z[61], n_496, n_500);
  or g377 (n_497, A[61], B[61]);
  xor g378 (n_500, A[61], B[61]);
  or g379 (n_198, wc, n_192);
  not gc (wc, A[1]);
  or g380 (n_199, wc0, n_192);
  not gc0 (wc0, B[1]);
  xnor g381 (Z[1], n_192, n_200);
  or g382 (n_498, A[61], wc1);
  not gc1 (wc1, n_496);
  or g383 (n_499, B[61], wc2);
  not gc2 (wc2, n_496);
endmodule

module add_signed_3603_1_GENERIC(A, B, Z);
  input [61:0] A, B;
  output [62:0] Z;
  wire [61:0] A, B;
  wire [62:0] Z;
  add_signed_3603_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_370_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [45:0] A, B;
  output [46:0] Z;
  wire [45:0] A, B;
  wire [46:0] Z;
  wire n_143, n_144, n_147, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_157, n_158, n_159, n_160, n_161, n_163, n_164;
  wire n_165, n_166, n_167, n_169, n_170, n_171, n_172, n_173;
  wire n_175, n_176, n_177, n_178, n_179, n_181, n_182, n_183;
  wire n_184, n_185, n_187, n_188, n_189, n_190, n_191, n_193;
  wire n_194, n_195, n_196, n_197, n_199, n_200, n_201, n_202;
  wire n_203, n_205, n_206, n_207, n_208, n_209, n_211, n_212;
  wire n_213, n_214, n_215, n_217, n_218, n_219, n_220, n_221;
  wire n_223, n_224, n_225, n_226, n_227, n_229, n_230, n_231;
  wire n_232, n_233, n_235, n_236, n_237, n_238, n_239, n_241;
  wire n_242, n_243, n_244, n_245, n_247, n_248, n_249, n_250;
  wire n_251, n_253, n_254, n_255, n_256, n_257, n_259, n_260;
  wire n_261, n_262, n_263, n_265, n_266, n_267, n_268, n_269;
  wire n_271, n_272, n_273, n_274, n_275, n_277, n_278, n_279;
  wire n_280, n_281, n_283, n_284, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_293, n_295, n_297, n_298, n_300, n_301;
  wire n_303, n_305, n_307, n_308, n_310, n_311, n_313, n_315;
  wire n_317, n_318, n_320, n_321, n_323, n_325, n_327, n_328;
  wire n_330, n_331, n_333, n_335, n_337, n_338, n_340, n_341;
  wire n_343, n_345, n_347, n_348, n_350, n_351, n_353, n_355;
  wire n_357, n_358, n_360, n_361, n_363, n_365, n_367, n_368;
  wire n_370, n_371, n_373, n_375, n_377, n_378, n_380, n_381;
  wire n_383, n_385, n_387, n_388, n_390, n_392, n_393, n_394;
  wire n_396, n_397, n_398, n_400, n_401, n_402, n_403, n_405;
  wire n_407, n_409, n_410, n_411, n_413, n_414, n_415, n_417;
  wire n_418, n_420, n_422, n_424, n_425, n_426, n_428, n_429;
  wire n_430, n_432, n_433, n_435, n_437, n_439, n_440, n_441;
  wire n_443, n_444, n_445, n_447, n_448, n_450, n_452, n_454;
  wire n_455, n_456, n_458, n_459, n_460, n_462, n_463, n_465;
  wire n_466, n_468, n_469, n_471, n_473, n_474, n_475, n_477;
  wire n_478, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_496, n_499, n_501, n_502, n_503, n_506, n_509, n_511;
  wire n_512, n_514, n_516, n_517, n_519, n_521, n_522, n_524;
  wire n_526, n_527, n_529, n_530, n_532, n_535, n_537, n_538;
  wire n_539, n_542, n_545, n_547, n_548, n_550, n_552, n_553;
  wire n_555, n_557, n_558, n_559, n_561, n_562, n_564, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_585, n_586, n_587, n_589, n_590, n_591, n_593, n_594;
  wire n_595, n_597, n_598, n_599, n_601, n_602, n_603, n_605;
  wire n_606, n_607, n_609, n_610, n_611, n_613, n_614, n_616;
  wire n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_629, n_630, n_631, n_633, n_634;
  wire n_635, n_637, n_638, n_639, n_641, n_642, n_643, n_645;
  wire n_646, n_647, n_649, n_650, n_651, n_652, n_654, n_655;
  wire n_656, n_658, n_659, n_660, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_670, n_672, n_673, n_675, n_676;
  wire n_678, n_679, n_680, n_681, n_683, n_684, n_685, n_687;
  wire n_688, n_689, n_690, n_692, n_693, n_695, n_696, n_698;
  wire n_699, n_700, n_701, n_703, n_704, n_705, n_706, n_708;
  wire n_709, n_710, n_711, n_713, n_714, n_716, n_717, n_719;
  wire n_720, n_721, n_722, n_724, n_725, n_726, n_728, n_729;
  wire n_730, n_731, n_733, n_734, n_736, n_737, n_739, n_740;
  wire n_741, n_742, n_744, n_745, n_746, n_747, n_749, n_750;
  wire n_751, n_752, n_754, n_755, n_757, n_758, n_760, n_761;
  not g3 (Z[46], n_143);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_144, A[0], B[0]);
  nor g9 (n_147, A[1], B[1]);
  nand g10 (n_150, A[1], B[1]);
  nor g11 (n_157, A[2], B[2]);
  nand g12 (n_152, A[2], B[2]);
  nor g13 (n_153, A[3], B[3]);
  nand g14 (n_154, A[3], B[3]);
  nor g15 (n_163, A[4], B[4]);
  nand g16 (n_158, A[4], B[4]);
  nor g17 (n_159, A[5], B[5]);
  nand g18 (n_160, A[5], B[5]);
  nor g19 (n_169, A[6], B[6]);
  nand g20 (n_164, A[6], B[6]);
  nor g21 (n_165, A[7], B[7]);
  nand g22 (n_166, A[7], B[7]);
  nor g23 (n_175, A[8], B[8]);
  nand g24 (n_170, A[8], B[8]);
  nor g25 (n_171, A[9], B[9]);
  nand g26 (n_172, A[9], B[9]);
  nor g27 (n_181, A[10], B[10]);
  nand g28 (n_176, A[10], B[10]);
  nor g29 (n_177, A[11], B[11]);
  nand g30 (n_178, A[11], B[11]);
  nor g31 (n_187, A[12], B[12]);
  nand g32 (n_182, A[12], B[12]);
  nor g33 (n_183, A[13], B[13]);
  nand g34 (n_184, A[13], B[13]);
  nor g35 (n_193, A[14], B[14]);
  nand g36 (n_188, A[14], B[14]);
  nor g37 (n_189, A[15], B[15]);
  nand g38 (n_190, A[15], B[15]);
  nor g39 (n_199, A[16], B[16]);
  nand g40 (n_194, A[16], B[16]);
  nor g41 (n_195, A[17], B[17]);
  nand g42 (n_196, A[17], B[17]);
  nor g43 (n_205, A[18], B[18]);
  nand g44 (n_200, A[18], B[18]);
  nor g45 (n_201, A[19], B[19]);
  nand g46 (n_202, A[19], B[19]);
  nor g47 (n_211, A[20], B[20]);
  nand g48 (n_206, A[20], B[20]);
  nor g49 (n_207, A[21], B[21]);
  nand g50 (n_208, A[21], B[21]);
  nor g51 (n_217, A[22], B[22]);
  nand g52 (n_212, A[22], B[22]);
  nor g53 (n_213, A[23], B[23]);
  nand g54 (n_214, A[23], B[23]);
  nor g55 (n_223, A[24], B[24]);
  nand g56 (n_218, A[24], B[24]);
  nor g57 (n_219, A[25], B[25]);
  nand g58 (n_220, A[25], B[25]);
  nor g59 (n_229, A[26], B[26]);
  nand g60 (n_224, A[26], B[26]);
  nor g61 (n_225, A[27], B[27]);
  nand g62 (n_226, A[27], B[27]);
  nor g63 (n_235, A[28], B[28]);
  nand g64 (n_230, A[28], B[28]);
  nor g65 (n_231, A[29], B[29]);
  nand g66 (n_232, A[29], B[29]);
  nor g67 (n_241, A[30], B[30]);
  nand g68 (n_236, A[30], B[30]);
  nor g69 (n_237, A[31], B[31]);
  nand g70 (n_238, A[31], B[31]);
  nor g71 (n_247, A[32], B[32]);
  nand g72 (n_242, A[32], B[32]);
  nor g73 (n_243, A[33], B[33]);
  nand g74 (n_244, A[33], B[33]);
  nor g75 (n_253, A[34], B[34]);
  nand g76 (n_248, A[34], B[34]);
  nor g77 (n_249, A[35], B[35]);
  nand g78 (n_250, A[35], B[35]);
  nor g79 (n_259, A[36], B[36]);
  nand g80 (n_254, A[36], B[36]);
  nor g81 (n_255, A[37], B[37]);
  nand g82 (n_256, A[37], B[37]);
  nor g83 (n_265, A[38], B[38]);
  nand g84 (n_260, A[38], B[38]);
  nor g85 (n_261, A[39], B[39]);
  nand g86 (n_262, A[39], B[39]);
  nor g87 (n_271, A[40], B[40]);
  nand g88 (n_266, A[40], B[40]);
  nor g89 (n_267, A[41], B[41]);
  nand g90 (n_268, A[41], B[41]);
  nor g91 (n_277, A[42], B[42]);
  nand g92 (n_272, A[42], B[42]);
  nor g93 (n_273, A[43], B[43]);
  nand g94 (n_274, A[43], B[43]);
  nor g95 (n_283, A[44], B[44]);
  nand g96 (n_278, A[44], B[44]);
  nand g101 (n_284, n_150, n_151);
  nor g102 (n_155, n_152, n_153);
  nor g105 (n_287, n_157, n_153);
  nor g106 (n_161, n_158, n_159);
  nor g109 (n_293, n_163, n_159);
  nor g110 (n_167, n_164, n_165);
  nor g113 (n_295, n_169, n_165);
  nor g114 (n_173, n_170, n_171);
  nor g117 (n_303, n_175, n_171);
  nor g118 (n_179, n_176, n_177);
  nor g121 (n_305, n_181, n_177);
  nor g122 (n_185, n_182, n_183);
  nor g125 (n_313, n_187, n_183);
  nor g126 (n_191, n_188, n_189);
  nor g129 (n_315, n_193, n_189);
  nor g130 (n_197, n_194, n_195);
  nor g133 (n_323, n_199, n_195);
  nor g134 (n_203, n_200, n_201);
  nor g137 (n_325, n_205, n_201);
  nor g138 (n_209, n_206, n_207);
  nor g141 (n_333, n_211, n_207);
  nor g142 (n_215, n_212, n_213);
  nor g145 (n_335, n_217, n_213);
  nor g146 (n_221, n_218, n_219);
  nor g149 (n_343, n_223, n_219);
  nor g150 (n_227, n_224, n_225);
  nor g153 (n_345, n_229, n_225);
  nor g154 (n_233, n_230, n_231);
  nor g157 (n_353, n_235, n_231);
  nor g158 (n_239, n_236, n_237);
  nor g161 (n_355, n_241, n_237);
  nor g162 (n_245, n_242, n_243);
  nor g165 (n_363, n_247, n_243);
  nor g166 (n_251, n_248, n_249);
  nor g169 (n_365, n_253, n_249);
  nor g170 (n_257, n_254, n_255);
  nor g173 (n_373, n_259, n_255);
  nor g174 (n_263, n_260, n_261);
  nor g177 (n_375, n_265, n_261);
  nor g178 (n_269, n_266, n_267);
  nor g181 (n_383, n_271, n_267);
  nor g182 (n_275, n_272, n_273);
  nor g185 (n_385, n_277, n_273);
  nor g186 (n_281, n_278, n_279);
  nor g189 (n_466, n_283, n_279);
  nand g192 (n_654, n_152, n_286);
  nand g193 (n_289, n_287, n_284);
  nand g194 (n_390, n_288, n_289);
  nor g195 (n_291, n_169, n_290);
  nand g204 (n_398, n_293, n_295);
  nor g205 (n_301, n_181, n_300);
  nand g214 (n_405, n_303, n_305);
  nor g215 (n_311, n_193, n_310);
  nand g224 (n_413, n_313, n_315);
  nor g225 (n_321, n_205, n_320);
  nand g234 (n_420, n_323, n_325);
  nor g235 (n_331, n_217, n_330);
  nand g244 (n_428, n_333, n_335);
  nor g245 (n_341, n_229, n_340);
  nand g254 (n_435, n_343, n_345);
  nor g255 (n_351, n_241, n_350);
  nand g264 (n_443, n_353, n_355);
  nor g265 (n_361, n_253, n_360);
  nand g274 (n_450, n_363, n_365);
  nor g275 (n_371, n_265, n_370);
  nand g284 (n_458, n_373, n_375);
  nor g285 (n_381, n_277, n_380);
  nand g294 (n_465, n_383, n_385);
  nand g297 (n_658, n_158, n_392);
  nand g298 (n_393, n_293, n_390);
  nand g299 (n_660, n_290, n_393);
  nand g302 (n_663, n_396, n_397);
  nand g305 (n_471, n_400, n_401);
  nor g306 (n_403, n_187, n_402);
  nor g309 (n_481, n_187, n_405);
  nor g315 (n_411, n_409, n_402);
  nor g318 (n_487, n_405, n_409);
  nor g319 (n_415, n_413, n_402);
  nor g322 (n_490, n_405, n_413);
  nor g323 (n_418, n_211, n_417);
  nor g326 (n_565, n_211, n_420);
  nor g332 (n_426, n_424, n_417);
  nor g335 (n_571, n_420, n_424);
  nor g336 (n_430, n_428, n_417);
  nor g339 (n_496, n_420, n_428);
  nor g340 (n_433, n_235, n_432);
  nor g343 (n_509, n_235, n_435);
  nor g349 (n_441, n_439, n_432);
  nor g352 (n_519, n_435, n_439);
  nor g353 (n_445, n_443, n_432);
  nor g356 (n_524, n_435, n_443);
  nor g357 (n_448, n_259, n_447);
  nor g360 (n_617, n_259, n_450);
  nor g366 (n_456, n_454, n_447);
  nor g369 (n_623, n_450, n_454);
  nor g370 (n_460, n_458, n_447);
  nor g373 (n_532, n_450, n_458);
  nor g374 (n_463, n_283, n_462);
  nor g377 (n_545, n_283, n_465);
  nand g385 (n_667, n_170, n_473);
  nand g386 (n_474, n_303, n_471);
  nand g387 (n_669, n_300, n_474);
  nand g390 (n_672, n_477, n_478);
  nand g393 (n_675, n_402, n_480);
  nand g394 (n_483, n_481, n_471);
  nand g395 (n_678, n_482, n_483);
  nand g396 (n_486, n_484, n_471);
  nand g397 (n_680, n_485, n_486);
  nand g398 (n_489, n_487, n_471);
  nand g399 (n_683, n_488, n_489);
  nand g400 (n_492, n_490, n_471);
  nand g401 (n_555, n_491, n_492);
  nor g402 (n_494, n_223, n_493);
  nand g411 (n_579, n_343, n_496);
  nor g412 (n_503, n_501, n_493);
  nor g417 (n_506, n_435, n_493);
  nand g426 (n_591, n_496, n_509);
  nand g431 (n_595, n_496, n_514);
  nand g436 (n_599, n_496, n_519);
  nand g441 (n_603, n_496, n_524);
  nor g442 (n_530, n_271, n_529);
  nand g451 (n_631, n_383, n_532);
  nor g452 (n_539, n_537, n_529);
  nor g457 (n_542, n_465, n_529);
  nand g466 (n_643, n_532, n_545);
  nand g471 (n_647, n_532, n_550);
  nand g474 (n_687, n_194, n_557);
  nand g475 (n_558, n_323, n_555);
  nand g476 (n_689, n_320, n_558);
  nand g479 (n_692, n_561, n_562);
  nand g482 (n_695, n_417, n_564);
  nand g483 (n_567, n_565, n_555);
  nand g484 (n_698, n_566, n_567);
  nand g485 (n_570, n_568, n_555);
  nand g486 (n_700, n_569, n_570);
  nand g487 (n_573, n_571, n_555);
  nand g488 (n_703, n_572, n_573);
  nand g489 (n_574, n_496, n_555);
  nand g490 (n_705, n_493, n_574);
  nand g493 (n_708, n_577, n_578);
  nand g496 (n_710, n_581, n_582);
  nand g499 (n_713, n_585, n_586);
  nand g502 (n_716, n_589, n_590);
  nand g505 (n_719, n_593, n_594);
  nand g508 (n_721, n_597, n_598);
  nand g511 (n_724, n_601, n_602);
  nand g514 (n_607, n_605, n_606);
  nand g517 (n_728, n_242, n_609);
  nand g518 (n_610, n_363, n_607);
  nand g519 (n_730, n_360, n_610);
  nand g522 (n_733, n_613, n_614);
  nand g525 (n_736, n_447, n_616);
  nand g526 (n_619, n_617, n_607);
  nand g527 (n_739, n_618, n_619);
  nand g528 (n_622, n_620, n_607);
  nand g529 (n_741, n_621, n_622);
  nand g530 (n_625, n_623, n_607);
  nand g531 (n_744, n_624, n_625);
  nand g532 (n_626, n_532, n_607);
  nand g533 (n_746, n_529, n_626);
  nand g536 (n_749, n_629, n_630);
  nand g539 (n_751, n_633, n_634);
  nand g542 (n_754, n_637, n_638);
  nand g545 (n_757, n_641, n_642);
  nand g548 (n_760, n_645, n_646);
  nand g551 (n_143, n_649, n_650);
  xnor g555 (Z[2], n_284, n_652);
  xnor g558 (Z[3], n_654, n_655);
  xnor g560 (Z[4], n_390, n_656);
  xnor g563 (Z[5], n_658, n_659);
  xnor g565 (Z[6], n_660, n_661);
  xnor g568 (Z[7], n_663, n_664);
  xnor g570 (Z[8], n_471, n_665);
  xnor g573 (Z[9], n_667, n_668);
  xnor g575 (Z[10], n_669, n_670);
  xnor g578 (Z[11], n_672, n_673);
  xnor g581 (Z[12], n_675, n_676);
  xnor g584 (Z[13], n_678, n_679);
  xnor g586 (Z[14], n_680, n_681);
  xnor g589 (Z[15], n_683, n_684);
  xnor g591 (Z[16], n_555, n_685);
  xnor g594 (Z[17], n_687, n_688);
  xnor g596 (Z[18], n_689, n_690);
  xnor g599 (Z[19], n_692, n_693);
  xnor g602 (Z[20], n_695, n_696);
  xnor g605 (Z[21], n_698, n_699);
  xnor g607 (Z[22], n_700, n_701);
  xnor g610 (Z[23], n_703, n_704);
  xnor g612 (Z[24], n_705, n_706);
  xnor g615 (Z[25], n_708, n_709);
  xnor g617 (Z[26], n_710, n_711);
  xnor g620 (Z[27], n_713, n_714);
  xnor g623 (Z[28], n_716, n_717);
  xnor g626 (Z[29], n_719, n_720);
  xnor g628 (Z[30], n_721, n_722);
  xnor g631 (Z[31], n_724, n_725);
  xnor g633 (Z[32], n_607, n_726);
  xnor g636 (Z[33], n_728, n_729);
  xnor g638 (Z[34], n_730, n_731);
  xnor g641 (Z[35], n_733, n_734);
  xnor g644 (Z[36], n_736, n_737);
  xnor g647 (Z[37], n_739, n_740);
  xnor g649 (Z[38], n_741, n_742);
  xnor g652 (Z[39], n_744, n_745);
  xnor g654 (Z[40], n_746, n_747);
  xnor g657 (Z[41], n_749, n_750);
  xnor g659 (Z[42], n_751, n_752);
  xnor g662 (Z[43], n_754, n_755);
  xnor g665 (Z[44], n_757, n_758);
  xnor g668 (Z[45], n_760, n_761);
  and g671 (n_279, A[45], B[45]);
  or g672 (n_280, A[45], B[45]);
  and g673 (n_360, wc, n_244);
  not gc (wc, n_245);
  and g674 (n_367, wc0, n_250);
  not gc0 (wc0, n_251);
  and g675 (n_370, wc1, n_256);
  not gc1 (wc1, n_257);
  and g676 (n_377, wc2, n_262);
  not gc2 (wc2, n_263);
  and g677 (n_380, wc3, n_268);
  not gc3 (wc3, n_269);
  and g678 (n_387, wc4, n_274);
  not gc4 (wc4, n_275);
  and g679 (n_320, wc5, n_196);
  not gc5 (wc5, n_197);
  and g680 (n_327, wc6, n_202);
  not gc6 (wc6, n_203);
  and g681 (n_330, wc7, n_208);
  not gc7 (wc7, n_209);
  and g682 (n_337, wc8, n_214);
  not gc8 (wc8, n_215);
  and g683 (n_340, wc9, n_220);
  not gc9 (wc9, n_221);
  and g684 (n_347, wc10, n_226);
  not gc10 (wc10, n_227);
  and g685 (n_350, wc11, n_232);
  not gc11 (wc11, n_233);
  and g686 (n_357, wc12, n_238);
  not gc12 (wc12, n_239);
  and g687 (n_300, wc13, n_172);
  not gc13 (wc13, n_173);
  and g688 (n_307, wc14, n_178);
  not gc14 (wc14, n_179);
  and g689 (n_310, wc15, n_184);
  not gc15 (wc15, n_185);
  and g690 (n_317, wc16, n_190);
  not gc16 (wc16, n_191);
  and g691 (n_290, wc17, n_160);
  not gc17 (wc17, n_161);
  and g692 (n_297, wc18, n_166);
  not gc18 (wc18, n_167);
  and g693 (n_288, wc19, n_154);
  not gc19 (wc19, n_155);
  or g694 (n_151, n_144, n_147);
  or g695 (n_394, wc20, n_169);
  not gc20 (wc20, n_293);
  or g696 (n_475, wc21, n_181);
  not gc21 (wc21, n_303);
  or g697 (n_409, wc22, n_193);
  not gc22 (wc22, n_313);
  or g698 (n_559, wc23, n_205);
  not gc23 (wc23, n_323);
  or g699 (n_424, wc24, n_217);
  not gc24 (wc24, n_333);
  or g700 (n_501, wc25, n_229);
  not gc25 (wc25, n_343);
  or g701 (n_439, wc26, n_241);
  not gc26 (wc26, n_353);
  or g702 (n_611, wc27, n_253);
  not gc27 (wc27, n_363);
  or g703 (n_454, wc28, n_265);
  not gc28 (wc28, n_373);
  or g704 (n_537, wc29, n_277);
  not gc29 (wc29, n_383);
  or g705 (n_651, wc30, n_147);
  not gc30 (wc30, n_150);
  or g706 (n_652, wc31, n_157);
  not gc31 (wc31, n_152);
  or g707 (n_655, wc32, n_153);
  not gc32 (wc32, n_154);
  or g708 (n_656, wc33, n_163);
  not gc33 (wc33, n_158);
  or g709 (n_659, wc34, n_159);
  not gc34 (wc34, n_160);
  or g710 (n_661, wc35, n_169);
  not gc35 (wc35, n_164);
  or g711 (n_664, wc36, n_165);
  not gc36 (wc36, n_166);
  or g712 (n_665, wc37, n_175);
  not gc37 (wc37, n_170);
  or g713 (n_668, wc38, n_171);
  not gc38 (wc38, n_172);
  or g714 (n_670, wc39, n_181);
  not gc39 (wc39, n_176);
  or g715 (n_673, wc40, n_177);
  not gc40 (wc40, n_178);
  or g716 (n_676, wc41, n_187);
  not gc41 (wc41, n_182);
  or g717 (n_679, wc42, n_183);
  not gc42 (wc42, n_184);
  or g718 (n_681, wc43, n_193);
  not gc43 (wc43, n_188);
  or g719 (n_684, wc44, n_189);
  not gc44 (wc44, n_190);
  or g720 (n_685, wc45, n_199);
  not gc45 (wc45, n_194);
  or g721 (n_688, wc46, n_195);
  not gc46 (wc46, n_196);
  or g722 (n_690, wc47, n_205);
  not gc47 (wc47, n_200);
  or g723 (n_693, wc48, n_201);
  not gc48 (wc48, n_202);
  or g724 (n_696, wc49, n_211);
  not gc49 (wc49, n_206);
  or g725 (n_699, wc50, n_207);
  not gc50 (wc50, n_208);
  or g726 (n_701, wc51, n_217);
  not gc51 (wc51, n_212);
  or g727 (n_704, wc52, n_213);
  not gc52 (wc52, n_214);
  or g728 (n_706, wc53, n_223);
  not gc53 (wc53, n_218);
  or g729 (n_709, wc54, n_219);
  not gc54 (wc54, n_220);
  or g730 (n_711, wc55, n_229);
  not gc55 (wc55, n_224);
  or g731 (n_714, wc56, n_225);
  not gc56 (wc56, n_226);
  or g732 (n_717, wc57, n_235);
  not gc57 (wc57, n_230);
  or g733 (n_720, wc58, n_231);
  not gc58 (wc58, n_232);
  or g734 (n_722, wc59, n_241);
  not gc59 (wc59, n_236);
  or g735 (n_725, wc60, n_237);
  not gc60 (wc60, n_238);
  or g736 (n_726, wc61, n_247);
  not gc61 (wc61, n_242);
  or g737 (n_729, wc62, n_243);
  not gc62 (wc62, n_244);
  or g738 (n_731, wc63, n_253);
  not gc63 (wc63, n_248);
  or g739 (n_734, wc64, n_249);
  not gc64 (wc64, n_250);
  or g740 (n_737, wc65, n_259);
  not gc65 (wc65, n_254);
  or g741 (n_740, wc66, n_255);
  not gc66 (wc66, n_256);
  or g742 (n_742, wc67, n_265);
  not gc67 (wc67, n_260);
  or g743 (n_745, wc68, n_261);
  not gc68 (wc68, n_262);
  or g744 (n_747, wc69, n_271);
  not gc69 (wc69, n_266);
  or g745 (n_750, wc70, n_267);
  not gc70 (wc70, n_268);
  or g746 (n_752, wc71, n_277);
  not gc71 (wc71, n_272);
  or g747 (n_755, wc72, n_273);
  not gc72 (wc72, n_274);
  or g748 (n_758, wc73, n_283);
  not gc73 (wc73, n_278);
  and g749 (n_368, wc74, n_365);
  not gc74 (wc74, n_360);
  and g750 (n_378, wc75, n_375);
  not gc75 (wc75, n_370);
  and g751 (n_388, wc76, n_385);
  not gc76 (wc76, n_380);
  and g752 (n_468, n_280, wc77);
  not gc77 (wc77, n_281);
  and g753 (n_328, wc78, n_325);
  not gc78 (wc78, n_320);
  and g754 (n_338, wc79, n_335);
  not gc79 (wc79, n_330);
  and g755 (n_348, wc80, n_345);
  not gc80 (wc80, n_340);
  and g756 (n_358, wc81, n_355);
  not gc81 (wc81, n_350);
  and g757 (n_308, wc82, n_305);
  not gc82 (wc82, n_300);
  and g758 (n_318, wc83, n_315);
  not gc83 (wc83, n_310);
  and g759 (n_298, wc84, n_295);
  not gc84 (wc84, n_290);
  and g760 (n_484, wc85, n_313);
  not gc85 (wc85, n_405);
  and g761 (n_568, wc86, n_333);
  not gc86 (wc86, n_420);
  and g762 (n_514, wc87, n_353);
  not gc87 (wc87, n_435);
  and g763 (n_620, wc88, n_373);
  not gc88 (wc88, n_450);
  xor g764 (Z[1], n_144, n_651);
  or g765 (n_761, wc89, n_279);
  not gc89 (wc89, n_280);
  and g766 (n_447, wc90, n_367);
  not gc90 (wc90, n_368);
  and g767 (n_459, wc91, n_377);
  not gc91 (wc91, n_378);
  and g768 (n_550, wc92, n_466);
  not gc92 (wc92, n_465);
  and g769 (n_462, wc93, n_387);
  not gc93 (wc93, n_388);
  and g770 (n_417, wc94, n_327);
  not gc94 (wc94, n_328);
  and g771 (n_429, wc95, n_337);
  not gc95 (wc95, n_338);
  and g772 (n_432, wc96, n_347);
  not gc96 (wc96, n_348);
  and g773 (n_444, wc97, n_357);
  not gc97 (wc97, n_358);
  and g774 (n_402, wc98, n_307);
  not gc98 (wc98, n_308);
  and g775 (n_414, wc99, n_317);
  not gc99 (wc99, n_318);
  and g776 (n_400, wc100, n_297);
  not gc100 (wc100, n_298);
  or g777 (n_286, wc101, n_157);
  not gc101 (wc101, n_284);
  and g778 (n_396, wc102, n_164);
  not gc102 (wc102, n_291);
  and g779 (n_477, wc103, n_176);
  not gc103 (wc103, n_301);
  and g780 (n_410, wc104, n_188);
  not gc104 (wc104, n_311);
  and g781 (n_561, wc105, n_200);
  not gc105 (wc105, n_321);
  and g782 (n_425, wc106, n_212);
  not gc106 (wc106, n_331);
  and g783 (n_502, wc107, n_224);
  not gc107 (wc107, n_341);
  and g784 (n_440, wc108, n_236);
  not gc108 (wc108, n_351);
  and g785 (n_613, wc109, n_248);
  not gc109 (wc109, n_361);
  and g786 (n_455, wc110, n_260);
  not gc110 (wc110, n_371);
  and g787 (n_538, wc111, n_272);
  not gc111 (wc111, n_381);
  or g788 (n_575, wc112, n_223);
  not gc112 (wc112, n_496);
  or g789 (n_583, n_501, wc113);
  not gc113 (wc113, n_496);
  or g790 (n_587, wc114, n_435);
  not gc114 (wc114, n_496);
  or g791 (n_627, wc115, n_271);
  not gc115 (wc115, n_532);
  or g792 (n_635, n_537, wc116);
  not gc116 (wc116, n_532);
  or g793 (n_639, wc117, n_465);
  not gc117 (wc117, n_532);
  and g794 (n_469, wc118, n_466);
  not gc118 (wc118, n_462);
  and g795 (n_407, wc119, n_313);
  not gc119 (wc119, n_402);
  and g796 (n_422, wc120, n_333);
  not gc120 (wc120, n_417);
  and g797 (n_437, wc121, n_353);
  not gc121 (wc121, n_432);
  and g798 (n_452, wc122, n_373);
  not gc122 (wc122, n_447);
  and g799 (n_529, n_459, wc123);
  not gc123 (wc123, n_460);
  and g800 (n_552, wc124, n_468);
  not gc124 (wc124, n_469);
  and g801 (n_493, n_429, wc125);
  not gc125 (wc125, n_430);
  and g802 (n_526, n_444, wc126);
  not gc126 (wc126, n_445);
  and g803 (n_491, n_414, wc127);
  not gc127 (wc127, n_415);
  or g804 (n_401, n_398, wc128);
  not gc128 (wc128, n_390);
  or g805 (n_392, wc129, n_163);
  not gc129 (wc129, n_390);
  or g806 (n_397, n_394, wc130);
  not gc130 (wc130, n_390);
  and g807 (n_482, wc131, n_182);
  not gc131 (wc131, n_403);
  and g808 (n_485, wc132, n_310);
  not gc132 (wc132, n_407);
  and g809 (n_488, n_410, wc133);
  not gc133 (wc133, n_411);
  and g810 (n_566, wc134, n_206);
  not gc134 (wc134, n_418);
  and g811 (n_569, wc135, n_330);
  not gc135 (wc135, n_422);
  and g812 (n_572, n_425, wc136);
  not gc136 (wc136, n_426);
  and g813 (n_511, wc137, n_230);
  not gc137 (wc137, n_433);
  and g814 (n_516, wc138, n_350);
  not gc138 (wc138, n_437);
  and g815 (n_521, n_440, wc139);
  not gc139 (wc139, n_441);
  and g816 (n_618, wc140, n_254);
  not gc140 (wc140, n_448);
  and g817 (n_621, wc141, n_370);
  not gc141 (wc141, n_452);
  and g818 (n_624, n_455, wc142);
  not gc142 (wc142, n_456);
  and g819 (n_547, wc143, n_278);
  not gc143 (wc143, n_463);
  and g820 (n_553, wc144, n_550);
  not gc144 (wc144, n_529);
  and g821 (n_527, wc145, n_524);
  not gc145 (wc145, n_493);
  and g822 (n_499, wc146, n_343);
  not gc146 (wc146, n_493);
  and g823 (n_512, wc147, n_509);
  not gc147 (wc147, n_493);
  and g824 (n_517, wc148, n_514);
  not gc148 (wc148, n_493);
  and g825 (n_522, wc149, n_519);
  not gc149 (wc149, n_493);
  and g826 (n_535, wc150, n_383);
  not gc150 (wc150, n_529);
  and g827 (n_548, wc151, n_545);
  not gc151 (wc151, n_529);
  and g828 (n_649, wc152, n_552);
  not gc152 (wc152, n_553);
  and g829 (n_605, wc153, n_526);
  not gc153 (wc153, n_527);
  or g830 (n_473, wc154, n_175);
  not gc154 (wc154, n_471);
  or g831 (n_478, n_475, wc155);
  not gc155 (wc155, n_471);
  or g832 (n_480, wc156, n_405);
  not gc156 (wc156, n_471);
  and g833 (n_577, wc157, n_218);
  not gc157 (wc157, n_494);
  and g834 (n_581, wc158, n_340);
  not gc158 (wc158, n_499);
  and g835 (n_585, n_502, wc159);
  not gc159 (wc159, n_503);
  and g836 (n_589, n_432, wc160);
  not gc160 (wc160, n_506);
  and g837 (n_593, wc161, n_511);
  not gc161 (wc161, n_512);
  and g838 (n_597, wc162, n_516);
  not gc162 (wc162, n_517);
  and g839 (n_601, wc163, n_521);
  not gc163 (wc163, n_522);
  and g840 (n_629, wc164, n_266);
  not gc164 (wc164, n_530);
  and g841 (n_633, wc165, n_380);
  not gc165 (wc165, n_535);
  and g842 (n_637, n_538, wc166);
  not gc166 (wc166, n_539);
  and g843 (n_641, n_462, wc167);
  not gc167 (wc167, n_542);
  and g844 (n_645, wc168, n_547);
  not gc168 (wc168, n_548);
  or g845 (n_606, n_603, wc169);
  not gc169 (wc169, n_555);
  or g846 (n_557, wc170, n_199);
  not gc170 (wc170, n_555);
  or g847 (n_562, n_559, wc171);
  not gc171 (wc171, n_555);
  or g848 (n_564, wc172, n_420);
  not gc172 (wc172, n_555);
  or g849 (n_578, n_575, wc173);
  not gc173 (wc173, n_555);
  or g850 (n_582, n_579, wc174);
  not gc174 (wc174, n_555);
  or g851 (n_586, n_583, wc175);
  not gc175 (wc175, n_555);
  or g852 (n_590, n_587, wc176);
  not gc176 (wc176, n_555);
  or g853 (n_594, n_591, wc177);
  not gc177 (wc177, n_555);
  or g854 (n_598, n_595, wc178);
  not gc178 (wc178, n_555);
  or g855 (n_602, n_599, wc179);
  not gc179 (wc179, n_555);
  or g856 (n_650, wc180, n_647);
  not gc180 (wc180, n_607);
  or g857 (n_609, wc181, n_247);
  not gc181 (wc181, n_607);
  or g858 (n_614, n_611, wc182);
  not gc182 (wc182, n_607);
  or g859 (n_616, wc183, n_450);
  not gc183 (wc183, n_607);
  or g860 (n_630, n_627, wc184);
  not gc184 (wc184, n_607);
  or g861 (n_634, wc185, n_631);
  not gc185 (wc185, n_607);
  or g862 (n_638, n_635, wc186);
  not gc186 (wc186, n_607);
  or g863 (n_642, n_639, wc187);
  not gc187 (wc187, n_607);
  or g864 (n_646, wc188, n_643);
  not gc188 (wc188, n_607);
endmodule

module add_signed_370_GENERIC(A, B, Z);
  input [45:0] A, B;
  output [46:0] Z;
  wire [45:0] A, B;
  wire [46:0] Z;
  add_signed_370_GENERIC_REAL g1(.A ({A[44], A[44:0]}), .B ({B[44],
       B[44:0]}), .Z (Z));
endmodule

module add_signed_384_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [44:0] A, B;
  output [45:0] Z;
  wire [44:0] A, B;
  wire [45:0] Z;
  wire n_140, n_141, n_144, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_154, n_155, n_156, n_157, n_158, n_160, n_161;
  wire n_162, n_163, n_164, n_166, n_167, n_168, n_169, n_170;
  wire n_172, n_173, n_174, n_175, n_176, n_178, n_179, n_180;
  wire n_181, n_182, n_184, n_185, n_186, n_187, n_188, n_190;
  wire n_191, n_192, n_193, n_194, n_196, n_197, n_198, n_199;
  wire n_200, n_202, n_203, n_204, n_205, n_206, n_208, n_209;
  wire n_210, n_211, n_212, n_214, n_215, n_216, n_217, n_218;
  wire n_220, n_221, n_222, n_223, n_224, n_226, n_227, n_228;
  wire n_229, n_230, n_232, n_233, n_234, n_235, n_236, n_238;
  wire n_239, n_240, n_241, n_242, n_244, n_245, n_246, n_247;
  wire n_248, n_250, n_251, n_252, n_253, n_254, n_256, n_257;
  wire n_258, n_259, n_260, n_262, n_263, n_264, n_265, n_266;
  wire n_268, n_269, n_270, n_271, n_272, n_274, n_275, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_284, n_286, n_288;
  wire n_289, n_291, n_292, n_294, n_296, n_298, n_299, n_301;
  wire n_302, n_304, n_306, n_308, n_309, n_311, n_312, n_314;
  wire n_316, n_318, n_319, n_321, n_322, n_324, n_326, n_328;
  wire n_329, n_331, n_332, n_334, n_336, n_338, n_339, n_341;
  wire n_342, n_344, n_346, n_348, n_349, n_351, n_352, n_354;
  wire n_356, n_358, n_359, n_361, n_362, n_364, n_366, n_368;
  wire n_369, n_371, n_372, n_374, n_376, n_378, n_379, n_381;
  wire n_383, n_384, n_385, n_387, n_388, n_389, n_391, n_392;
  wire n_393, n_394, n_396, n_398, n_400, n_401, n_402, n_404;
  wire n_405, n_406, n_408, n_409, n_411, n_413, n_415, n_416;
  wire n_417, n_419, n_420, n_421, n_423, n_424, n_426, n_428;
  wire n_430, n_431, n_432, n_434, n_435, n_436, n_438, n_439;
  wire n_441, n_443, n_445, n_446, n_447, n_449, n_450, n_451;
  wire n_453, n_454, n_455, n_456, n_458, n_459, n_461, n_462;
  wire n_463, n_465, n_466, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_484, n_487, n_489, n_490, n_491, n_494;
  wire n_497, n_499, n_500, n_502, n_504, n_505, n_507, n_509;
  wire n_510, n_512, n_514, n_515, n_517, n_518, n_520, n_523;
  wire n_525, n_526, n_527, n_530, n_533, n_535, n_536, n_538;
  wire n_540, n_541, n_542, n_544, n_545, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_560, n_561, n_562, n_564, n_565, n_566, n_568;
  wire n_569, n_570, n_572, n_573, n_574, n_576, n_577, n_578;
  wire n_580, n_581, n_582, n_584, n_585, n_586, n_588, n_589;
  wire n_590, n_592, n_593, n_594, n_596, n_597, n_599, n_600;
  wire n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608;
  wire n_609, n_610, n_612, n_613, n_614, n_616, n_617, n_618;
  wire n_620, n_621, n_622, n_624, n_625, n_626, n_628, n_629;
  wire n_630, n_631, n_633, n_634, n_635, n_637, n_638, n_639;
  wire n_640, n_642, n_643, n_644, n_646, n_647, n_648, n_649;
  wire n_651, n_652, n_654, n_655, n_657, n_658, n_659, n_660;
  wire n_662, n_663, n_664, n_666, n_667, n_668, n_669, n_671;
  wire n_672, n_674, n_675, n_677, n_678, n_679, n_680, n_682;
  wire n_683, n_684, n_685, n_687, n_688, n_689, n_690, n_692;
  wire n_693, n_695, n_696, n_698, n_699, n_700, n_701, n_703;
  wire n_704, n_705, n_707, n_708, n_709, n_710, n_712, n_713;
  wire n_715, n_716, n_718, n_719, n_720, n_721, n_723, n_724;
  wire n_725, n_726, n_728, n_729, n_730, n_731, n_733, n_734;
  wire n_736, n_737;
  not g3 (Z[45], n_140);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_141, A[0], B[0]);
  nor g9 (n_144, A[1], B[1]);
  nand g10 (n_147, A[1], B[1]);
  nor g11 (n_154, A[2], B[2]);
  nand g12 (n_149, A[2], B[2]);
  nor g13 (n_150, A[3], B[3]);
  nand g14 (n_151, A[3], B[3]);
  nor g15 (n_160, A[4], B[4]);
  nand g16 (n_155, A[4], B[4]);
  nor g17 (n_156, A[5], B[5]);
  nand g18 (n_157, A[5], B[5]);
  nor g19 (n_166, A[6], B[6]);
  nand g20 (n_161, A[6], B[6]);
  nor g21 (n_162, A[7], B[7]);
  nand g22 (n_163, A[7], B[7]);
  nor g23 (n_172, A[8], B[8]);
  nand g24 (n_167, A[8], B[8]);
  nor g25 (n_168, A[9], B[9]);
  nand g26 (n_169, A[9], B[9]);
  nor g27 (n_178, A[10], B[10]);
  nand g28 (n_173, A[10], B[10]);
  nor g29 (n_174, A[11], B[11]);
  nand g30 (n_175, A[11], B[11]);
  nor g31 (n_184, A[12], B[12]);
  nand g32 (n_179, A[12], B[12]);
  nor g33 (n_180, A[13], B[13]);
  nand g34 (n_181, A[13], B[13]);
  nor g35 (n_190, A[14], B[14]);
  nand g36 (n_185, A[14], B[14]);
  nor g37 (n_186, A[15], B[15]);
  nand g38 (n_187, A[15], B[15]);
  nor g39 (n_196, A[16], B[16]);
  nand g40 (n_191, A[16], B[16]);
  nor g41 (n_192, A[17], B[17]);
  nand g42 (n_193, A[17], B[17]);
  nor g43 (n_202, A[18], B[18]);
  nand g44 (n_197, A[18], B[18]);
  nor g45 (n_198, A[19], B[19]);
  nand g46 (n_199, A[19], B[19]);
  nor g47 (n_208, A[20], B[20]);
  nand g48 (n_203, A[20], B[20]);
  nor g49 (n_204, A[21], B[21]);
  nand g50 (n_205, A[21], B[21]);
  nor g51 (n_214, A[22], B[22]);
  nand g52 (n_209, A[22], B[22]);
  nor g53 (n_210, A[23], B[23]);
  nand g54 (n_211, A[23], B[23]);
  nor g55 (n_220, A[24], B[24]);
  nand g56 (n_215, A[24], B[24]);
  nor g57 (n_216, A[25], B[25]);
  nand g58 (n_217, A[25], B[25]);
  nor g59 (n_226, A[26], B[26]);
  nand g60 (n_221, A[26], B[26]);
  nor g61 (n_222, A[27], B[27]);
  nand g62 (n_223, A[27], B[27]);
  nor g63 (n_232, A[28], B[28]);
  nand g64 (n_227, A[28], B[28]);
  nor g65 (n_228, A[29], B[29]);
  nand g66 (n_229, A[29], B[29]);
  nor g67 (n_238, A[30], B[30]);
  nand g68 (n_233, A[30], B[30]);
  nor g69 (n_234, A[31], B[31]);
  nand g70 (n_235, A[31], B[31]);
  nor g71 (n_244, A[32], B[32]);
  nand g72 (n_239, A[32], B[32]);
  nor g73 (n_240, A[33], B[33]);
  nand g74 (n_241, A[33], B[33]);
  nor g75 (n_250, A[34], B[34]);
  nand g76 (n_245, A[34], B[34]);
  nor g77 (n_246, A[35], B[35]);
  nand g78 (n_247, A[35], B[35]);
  nor g79 (n_256, A[36], B[36]);
  nand g80 (n_251, A[36], B[36]);
  nor g81 (n_252, A[37], B[37]);
  nand g82 (n_253, A[37], B[37]);
  nor g83 (n_262, A[38], B[38]);
  nand g84 (n_257, A[38], B[38]);
  nor g85 (n_258, A[39], B[39]);
  nand g86 (n_259, A[39], B[39]);
  nor g87 (n_268, A[40], B[40]);
  nand g88 (n_263, A[40], B[40]);
  nor g89 (n_264, A[41], B[41]);
  nand g90 (n_265, A[41], B[41]);
  nor g91 (n_274, A[42], B[42]);
  nand g92 (n_269, A[42], B[42]);
  nor g93 (n_270, A[43], B[43]);
  nand g94 (n_271, A[43], B[43]);
  nand g99 (n_275, n_147, n_148);
  nor g100 (n_152, n_149, n_150);
  nor g103 (n_278, n_154, n_150);
  nor g104 (n_158, n_155, n_156);
  nor g107 (n_284, n_160, n_156);
  nor g108 (n_164, n_161, n_162);
  nor g111 (n_286, n_166, n_162);
  nor g112 (n_170, n_167, n_168);
  nor g115 (n_294, n_172, n_168);
  nor g116 (n_176, n_173, n_174);
  nor g119 (n_296, n_178, n_174);
  nor g120 (n_182, n_179, n_180);
  nor g123 (n_304, n_184, n_180);
  nor g124 (n_188, n_185, n_186);
  nor g127 (n_306, n_190, n_186);
  nor g128 (n_194, n_191, n_192);
  nor g131 (n_314, n_196, n_192);
  nor g132 (n_200, n_197, n_198);
  nor g135 (n_316, n_202, n_198);
  nor g136 (n_206, n_203, n_204);
  nor g139 (n_324, n_208, n_204);
  nor g140 (n_212, n_209, n_210);
  nor g143 (n_326, n_214, n_210);
  nor g144 (n_218, n_215, n_216);
  nor g147 (n_334, n_220, n_216);
  nor g148 (n_224, n_221, n_222);
  nor g151 (n_336, n_226, n_222);
  nor g152 (n_230, n_227, n_228);
  nor g155 (n_344, n_232, n_228);
  nor g156 (n_236, n_233, n_234);
  nor g159 (n_346, n_238, n_234);
  nor g160 (n_242, n_239, n_240);
  nor g163 (n_354, n_244, n_240);
  nor g164 (n_248, n_245, n_246);
  nor g167 (n_356, n_250, n_246);
  nor g168 (n_254, n_251, n_252);
  nor g171 (n_364, n_256, n_252);
  nor g172 (n_260, n_257, n_258);
  nor g175 (n_366, n_262, n_258);
  nor g176 (n_266, n_263, n_264);
  nor g179 (n_374, n_268, n_264);
  nor g180 (n_272, n_269, n_270);
  nor g183 (n_376, n_274, n_270);
  nand g186 (n_633, n_149, n_277);
  nand g187 (n_280, n_278, n_275);
  nand g188 (n_381, n_279, n_280);
  nor g189 (n_282, n_166, n_281);
  nand g198 (n_389, n_284, n_286);
  nor g199 (n_292, n_178, n_291);
  nand g208 (n_396, n_294, n_296);
  nor g209 (n_302, n_190, n_301);
  nand g218 (n_404, n_304, n_306);
  nor g219 (n_312, n_202, n_311);
  nand g228 (n_411, n_314, n_316);
  nor g229 (n_322, n_214, n_321);
  nand g238 (n_419, n_324, n_326);
  nor g239 (n_332, n_226, n_331);
  nand g248 (n_426, n_334, n_336);
  nor g249 (n_342, n_238, n_341);
  nand g258 (n_434, n_344, n_346);
  nor g259 (n_352, n_250, n_351);
  nand g268 (n_441, n_354, n_356);
  nor g269 (n_362, n_262, n_361);
  nand g278 (n_449, n_364, n_366);
  nor g279 (n_372, n_274, n_371);
  nand g288 (n_458, n_374, n_376);
  nand g291 (n_637, n_155, n_383);
  nand g292 (n_384, n_284, n_381);
  nand g293 (n_639, n_281, n_384);
  nand g296 (n_642, n_387, n_388);
  nand g299 (n_459, n_391, n_392);
  nor g300 (n_394, n_184, n_393);
  nor g303 (n_469, n_184, n_396);
  nor g309 (n_402, n_400, n_393);
  nor g312 (n_475, n_396, n_400);
  nor g313 (n_406, n_404, n_393);
  nor g316 (n_478, n_396, n_404);
  nor g317 (n_409, n_208, n_408);
  nor g320 (n_548, n_208, n_411);
  nor g326 (n_417, n_415, n_408);
  nor g329 (n_554, n_411, n_415);
  nor g330 (n_421, n_419, n_408);
  nor g333 (n_484, n_411, n_419);
  nor g334 (n_424, n_232, n_423);
  nor g337 (n_497, n_232, n_426);
  nor g343 (n_432, n_430, n_423);
  nor g346 (n_507, n_426, n_430);
  nor g347 (n_436, n_434, n_423);
  nor g350 (n_512, n_426, n_434);
  nor g351 (n_439, n_256, n_438);
  nor g354 (n_600, n_256, n_441);
  nor g360 (n_447, n_445, n_438);
  nor g363 (n_606, n_441, n_445);
  nor g364 (n_451, n_449, n_438);
  nor g367 (n_520, n_441, n_449);
  nor g368 (n_456, n_453, n_454);
  nor g371 (n_533, n_453, n_458);
  nand g374 (n_646, n_167, n_461);
  nand g375 (n_462, n_294, n_459);
  nand g376 (n_648, n_291, n_462);
  nand g379 (n_651, n_465, n_466);
  nand g382 (n_654, n_393, n_468);
  nand g383 (n_471, n_469, n_459);
  nand g384 (n_657, n_470, n_471);
  nand g385 (n_474, n_472, n_459);
  nand g386 (n_659, n_473, n_474);
  nand g387 (n_477, n_475, n_459);
  nand g388 (n_662, n_476, n_477);
  nand g389 (n_480, n_478, n_459);
  nand g390 (n_538, n_479, n_480);
  nor g391 (n_482, n_220, n_481);
  nand g400 (n_562, n_334, n_484);
  nor g401 (n_491, n_489, n_481);
  nor g406 (n_494, n_426, n_481);
  nand g415 (n_574, n_484, n_497);
  nand g420 (n_578, n_484, n_502);
  nand g425 (n_582, n_484, n_507);
  nand g430 (n_586, n_484, n_512);
  nor g431 (n_518, n_268, n_517);
  nand g440 (n_614, n_374, n_520);
  nor g441 (n_527, n_525, n_517);
  nor g446 (n_530, n_458, n_517);
  nand g455 (n_626, n_520, n_533);
  nand g458 (n_666, n_191, n_540);
  nand g459 (n_541, n_314, n_538);
  nand g460 (n_668, n_311, n_541);
  nand g463 (n_671, n_544, n_545);
  nand g466 (n_674, n_408, n_547);
  nand g467 (n_550, n_548, n_538);
  nand g468 (n_677, n_549, n_550);
  nand g469 (n_553, n_551, n_538);
  nand g470 (n_679, n_552, n_553);
  nand g471 (n_556, n_554, n_538);
  nand g472 (n_682, n_555, n_556);
  nand g473 (n_557, n_484, n_538);
  nand g474 (n_684, n_481, n_557);
  nand g477 (n_687, n_560, n_561);
  nand g480 (n_689, n_564, n_565);
  nand g483 (n_692, n_568, n_569);
  nand g486 (n_695, n_572, n_573);
  nand g489 (n_698, n_576, n_577);
  nand g492 (n_700, n_580, n_581);
  nand g495 (n_703, n_584, n_585);
  nand g498 (n_590, n_588, n_589);
  nand g501 (n_707, n_239, n_592);
  nand g502 (n_593, n_354, n_590);
  nand g503 (n_709, n_351, n_593);
  nand g506 (n_712, n_596, n_597);
  nand g509 (n_715, n_438, n_599);
  nand g510 (n_602, n_600, n_590);
  nand g511 (n_718, n_601, n_602);
  nand g512 (n_605, n_603, n_590);
  nand g513 (n_720, n_604, n_605);
  nand g514 (n_608, n_606, n_590);
  nand g515 (n_723, n_607, n_608);
  nand g516 (n_609, n_520, n_590);
  nand g517 (n_725, n_517, n_609);
  nand g520 (n_728, n_612, n_613);
  nand g523 (n_730, n_616, n_617);
  nand g526 (n_733, n_620, n_621);
  nand g529 (n_736, n_624, n_625);
  nand g532 (n_140, n_628, n_629);
  xnor g536 (Z[2], n_275, n_631);
  xnor g539 (Z[3], n_633, n_634);
  xnor g541 (Z[4], n_381, n_635);
  xnor g544 (Z[5], n_637, n_638);
  xnor g546 (Z[6], n_639, n_640);
  xnor g549 (Z[7], n_642, n_643);
  xnor g551 (Z[8], n_459, n_644);
  xnor g554 (Z[9], n_646, n_647);
  xnor g556 (Z[10], n_648, n_649);
  xnor g559 (Z[11], n_651, n_652);
  xnor g562 (Z[12], n_654, n_655);
  xnor g565 (Z[13], n_657, n_658);
  xnor g567 (Z[14], n_659, n_660);
  xnor g570 (Z[15], n_662, n_663);
  xnor g572 (Z[16], n_538, n_664);
  xnor g575 (Z[17], n_666, n_667);
  xnor g577 (Z[18], n_668, n_669);
  xnor g580 (Z[19], n_671, n_672);
  xnor g583 (Z[20], n_674, n_675);
  xnor g586 (Z[21], n_677, n_678);
  xnor g588 (Z[22], n_679, n_680);
  xnor g591 (Z[23], n_682, n_683);
  xnor g593 (Z[24], n_684, n_685);
  xnor g596 (Z[25], n_687, n_688);
  xnor g598 (Z[26], n_689, n_690);
  xnor g601 (Z[27], n_692, n_693);
  xnor g604 (Z[28], n_695, n_696);
  xnor g607 (Z[29], n_698, n_699);
  xnor g609 (Z[30], n_700, n_701);
  xnor g612 (Z[31], n_703, n_704);
  xnor g614 (Z[32], n_590, n_705);
  xnor g617 (Z[33], n_707, n_708);
  xnor g619 (Z[34], n_709, n_710);
  xnor g622 (Z[35], n_712, n_713);
  xnor g625 (Z[36], n_715, n_716);
  xnor g628 (Z[37], n_718, n_719);
  xnor g630 (Z[38], n_720, n_721);
  xnor g633 (Z[39], n_723, n_724);
  xnor g635 (Z[40], n_725, n_726);
  xnor g638 (Z[41], n_728, n_729);
  xnor g640 (Z[42], n_730, n_731);
  xnor g643 (Z[43], n_733, n_734);
  xnor g646 (Z[44], n_736, n_737);
  and g649 (n_453, A[44], B[44]);
  or g650 (n_455, A[44], B[44]);
  and g651 (n_351, wc, n_241);
  not gc (wc, n_242);
  and g652 (n_358, wc0, n_247);
  not gc0 (wc0, n_248);
  and g653 (n_361, wc1, n_253);
  not gc1 (wc1, n_254);
  and g654 (n_368, wc2, n_259);
  not gc2 (wc2, n_260);
  and g655 (n_371, wc3, n_265);
  not gc3 (wc3, n_266);
  and g656 (n_378, wc4, n_271);
  not gc4 (wc4, n_272);
  and g657 (n_311, wc5, n_193);
  not gc5 (wc5, n_194);
  and g658 (n_318, wc6, n_199);
  not gc6 (wc6, n_200);
  and g659 (n_321, wc7, n_205);
  not gc7 (wc7, n_206);
  and g660 (n_328, wc8, n_211);
  not gc8 (wc8, n_212);
  and g661 (n_331, wc9, n_217);
  not gc9 (wc9, n_218);
  and g662 (n_338, wc10, n_223);
  not gc10 (wc10, n_224);
  and g663 (n_341, wc11, n_229);
  not gc11 (wc11, n_230);
  and g664 (n_348, wc12, n_235);
  not gc12 (wc12, n_236);
  and g665 (n_291, wc13, n_169);
  not gc13 (wc13, n_170);
  and g666 (n_298, wc14, n_175);
  not gc14 (wc14, n_176);
  and g667 (n_301, wc15, n_181);
  not gc15 (wc15, n_182);
  and g668 (n_308, wc16, n_187);
  not gc16 (wc16, n_188);
  and g669 (n_281, wc17, n_157);
  not gc17 (wc17, n_158);
  and g670 (n_288, wc18, n_163);
  not gc18 (wc18, n_164);
  and g671 (n_279, wc19, n_151);
  not gc19 (wc19, n_152);
  or g672 (n_148, n_141, n_144);
  or g673 (n_385, wc20, n_166);
  not gc20 (wc20, n_284);
  or g674 (n_463, wc21, n_178);
  not gc21 (wc21, n_294);
  or g675 (n_400, wc22, n_190);
  not gc22 (wc22, n_304);
  or g676 (n_542, wc23, n_202);
  not gc23 (wc23, n_314);
  or g677 (n_415, wc24, n_214);
  not gc24 (wc24, n_324);
  or g678 (n_489, wc25, n_226);
  not gc25 (wc25, n_334);
  or g679 (n_430, wc26, n_238);
  not gc26 (wc26, n_344);
  or g680 (n_594, wc27, n_250);
  not gc27 (wc27, n_354);
  or g681 (n_445, wc28, n_262);
  not gc28 (wc28, n_364);
  or g682 (n_525, wc29, n_274);
  not gc29 (wc29, n_374);
  or g683 (n_630, wc30, n_144);
  not gc30 (wc30, n_147);
  or g684 (n_631, wc31, n_154);
  not gc31 (wc31, n_149);
  or g685 (n_634, wc32, n_150);
  not gc32 (wc32, n_151);
  or g686 (n_635, wc33, n_160);
  not gc33 (wc33, n_155);
  or g687 (n_638, wc34, n_156);
  not gc34 (wc34, n_157);
  or g688 (n_640, wc35, n_166);
  not gc35 (wc35, n_161);
  or g689 (n_643, wc36, n_162);
  not gc36 (wc36, n_163);
  or g690 (n_644, wc37, n_172);
  not gc37 (wc37, n_167);
  or g691 (n_647, wc38, n_168);
  not gc38 (wc38, n_169);
  or g692 (n_649, wc39, n_178);
  not gc39 (wc39, n_173);
  or g693 (n_652, wc40, n_174);
  not gc40 (wc40, n_175);
  or g694 (n_655, wc41, n_184);
  not gc41 (wc41, n_179);
  or g695 (n_658, wc42, n_180);
  not gc42 (wc42, n_181);
  or g696 (n_660, wc43, n_190);
  not gc43 (wc43, n_185);
  or g697 (n_663, wc44, n_186);
  not gc44 (wc44, n_187);
  or g698 (n_664, wc45, n_196);
  not gc45 (wc45, n_191);
  or g699 (n_667, wc46, n_192);
  not gc46 (wc46, n_193);
  or g700 (n_669, wc47, n_202);
  not gc47 (wc47, n_197);
  or g701 (n_672, wc48, n_198);
  not gc48 (wc48, n_199);
  or g702 (n_675, wc49, n_208);
  not gc49 (wc49, n_203);
  or g703 (n_678, wc50, n_204);
  not gc50 (wc50, n_205);
  or g704 (n_680, wc51, n_214);
  not gc51 (wc51, n_209);
  or g705 (n_683, wc52, n_210);
  not gc52 (wc52, n_211);
  or g706 (n_685, wc53, n_220);
  not gc53 (wc53, n_215);
  or g707 (n_688, wc54, n_216);
  not gc54 (wc54, n_217);
  or g708 (n_690, wc55, n_226);
  not gc55 (wc55, n_221);
  or g709 (n_693, wc56, n_222);
  not gc56 (wc56, n_223);
  or g710 (n_696, wc57, n_232);
  not gc57 (wc57, n_227);
  or g711 (n_699, wc58, n_228);
  not gc58 (wc58, n_229);
  or g712 (n_701, wc59, n_238);
  not gc59 (wc59, n_233);
  or g713 (n_704, wc60, n_234);
  not gc60 (wc60, n_235);
  or g714 (n_705, wc61, n_244);
  not gc61 (wc61, n_239);
  or g715 (n_708, wc62, n_240);
  not gc62 (wc62, n_241);
  or g716 (n_710, wc63, n_250);
  not gc63 (wc63, n_245);
  or g717 (n_713, wc64, n_246);
  not gc64 (wc64, n_247);
  or g718 (n_716, wc65, n_256);
  not gc65 (wc65, n_251);
  or g719 (n_719, wc66, n_252);
  not gc66 (wc66, n_253);
  or g720 (n_721, wc67, n_262);
  not gc67 (wc67, n_257);
  or g721 (n_724, wc68, n_258);
  not gc68 (wc68, n_259);
  or g722 (n_726, wc69, n_268);
  not gc69 (wc69, n_263);
  or g723 (n_729, wc70, n_264);
  not gc70 (wc70, n_265);
  or g724 (n_731, wc71, n_274);
  not gc71 (wc71, n_269);
  or g725 (n_734, wc72, n_270);
  not gc72 (wc72, n_271);
  and g726 (n_359, wc73, n_356);
  not gc73 (wc73, n_351);
  and g727 (n_369, wc74, n_366);
  not gc74 (wc74, n_361);
  and g728 (n_379, wc75, n_376);
  not gc75 (wc75, n_371);
  and g729 (n_319, wc76, n_316);
  not gc76 (wc76, n_311);
  and g730 (n_329, wc77, n_326);
  not gc77 (wc77, n_321);
  and g731 (n_339, wc78, n_336);
  not gc78 (wc78, n_331);
  and g732 (n_349, wc79, n_346);
  not gc79 (wc79, n_341);
  and g733 (n_299, wc80, n_296);
  not gc80 (wc80, n_291);
  and g734 (n_309, wc81, n_306);
  not gc81 (wc81, n_301);
  and g735 (n_289, wc82, n_286);
  not gc82 (wc82, n_281);
  and g736 (n_472, wc83, n_304);
  not gc83 (wc83, n_396);
  and g737 (n_551, wc84, n_324);
  not gc84 (wc84, n_411);
  and g738 (n_502, wc85, n_344);
  not gc85 (wc85, n_426);
  and g739 (n_603, wc86, n_364);
  not gc86 (wc86, n_441);
  xor g740 (Z[1], n_141, n_630);
  or g741 (n_737, wc87, n_453);
  not gc87 (wc87, n_455);
  and g742 (n_438, wc88, n_358);
  not gc88 (wc88, n_359);
  and g743 (n_450, wc89, n_368);
  not gc89 (wc89, n_369);
  and g744 (n_454, wc90, n_378);
  not gc90 (wc90, n_379);
  and g745 (n_408, wc91, n_318);
  not gc91 (wc91, n_319);
  and g746 (n_420, wc92, n_328);
  not gc92 (wc92, n_329);
  and g747 (n_423, wc93, n_338);
  not gc93 (wc93, n_339);
  and g748 (n_435, wc94, n_348);
  not gc94 (wc94, n_349);
  and g749 (n_393, wc95, n_298);
  not gc95 (wc95, n_299);
  and g750 (n_405, wc96, n_308);
  not gc96 (wc96, n_309);
  and g751 (n_391, wc97, n_288);
  not gc97 (wc97, n_289);
  or g752 (n_277, wc98, n_154);
  not gc98 (wc98, n_275);
  and g753 (n_387, wc99, n_161);
  not gc99 (wc99, n_282);
  and g754 (n_465, wc100, n_173);
  not gc100 (wc100, n_292);
  and g755 (n_401, wc101, n_185);
  not gc101 (wc101, n_302);
  and g756 (n_544, wc102, n_197);
  not gc102 (wc102, n_312);
  and g757 (n_416, wc103, n_209);
  not gc103 (wc103, n_322);
  and g758 (n_490, wc104, n_221);
  not gc104 (wc104, n_332);
  and g759 (n_431, wc105, n_233);
  not gc105 (wc105, n_342);
  and g760 (n_596, wc106, n_245);
  not gc106 (wc106, n_352);
  and g761 (n_446, wc107, n_257);
  not gc107 (wc107, n_362);
  and g762 (n_526, wc108, n_269);
  not gc108 (wc108, n_372);
  or g763 (n_558, wc109, n_220);
  not gc109 (wc109, n_484);
  or g764 (n_566, n_489, wc110);
  not gc110 (wc110, n_484);
  or g765 (n_570, wc111, n_426);
  not gc111 (wc111, n_484);
  or g766 (n_610, wc112, n_268);
  not gc112 (wc112, n_520);
  or g767 (n_618, n_525, wc113);
  not gc113 (wc113, n_520);
  or g768 (n_622, wc114, n_458);
  not gc114 (wc114, n_520);
  and g769 (n_398, wc115, n_304);
  not gc115 (wc115, n_393);
  and g770 (n_413, wc116, n_324);
  not gc116 (wc116, n_408);
  and g771 (n_428, wc117, n_344);
  not gc117 (wc117, n_423);
  and g772 (n_443, wc118, n_364);
  not gc118 (wc118, n_438);
  and g773 (n_517, n_450, wc119);
  not gc119 (wc119, n_451);
  and g774 (n_535, n_455, wc120);
  not gc120 (wc120, n_456);
  and g775 (n_481, n_420, wc121);
  not gc121 (wc121, n_421);
  and g776 (n_514, n_435, wc122);
  not gc122 (wc122, n_436);
  and g777 (n_479, n_405, wc123);
  not gc123 (wc123, n_406);
  or g778 (n_392, n_389, wc124);
  not gc124 (wc124, n_381);
  or g779 (n_383, wc125, n_160);
  not gc125 (wc125, n_381);
  or g780 (n_388, n_385, wc126);
  not gc126 (wc126, n_381);
  and g781 (n_470, wc127, n_179);
  not gc127 (wc127, n_394);
  and g782 (n_473, wc128, n_301);
  not gc128 (wc128, n_398);
  and g783 (n_476, n_401, wc129);
  not gc129 (wc129, n_402);
  and g784 (n_549, wc130, n_203);
  not gc130 (wc130, n_409);
  and g785 (n_552, wc131, n_321);
  not gc131 (wc131, n_413);
  and g786 (n_555, n_416, wc132);
  not gc132 (wc132, n_417);
  and g787 (n_499, wc133, n_227);
  not gc133 (wc133, n_424);
  and g788 (n_504, wc134, n_341);
  not gc134 (wc134, n_428);
  and g789 (n_509, n_431, wc135);
  not gc135 (wc135, n_432);
  and g790 (n_601, wc136, n_251);
  not gc136 (wc136, n_439);
  and g791 (n_604, wc137, n_361);
  not gc137 (wc137, n_443);
  and g792 (n_607, n_446, wc138);
  not gc138 (wc138, n_447);
  and g793 (n_536, wc139, n_533);
  not gc139 (wc139, n_517);
  and g794 (n_515, wc140, n_512);
  not gc140 (wc140, n_481);
  and g795 (n_487, wc141, n_334);
  not gc141 (wc141, n_481);
  and g796 (n_500, wc142, n_497);
  not gc142 (wc142, n_481);
  and g797 (n_505, wc143, n_502);
  not gc143 (wc143, n_481);
  and g798 (n_510, wc144, n_507);
  not gc144 (wc144, n_481);
  and g799 (n_523, wc145, n_374);
  not gc145 (wc145, n_517);
  and g800 (n_628, wc146, n_535);
  not gc146 (wc146, n_536);
  and g801 (n_588, wc147, n_514);
  not gc147 (wc147, n_515);
  or g802 (n_461, wc148, n_172);
  not gc148 (wc148, n_459);
  or g803 (n_466, n_463, wc149);
  not gc149 (wc149, n_459);
  or g804 (n_468, wc150, n_396);
  not gc150 (wc150, n_459);
  and g805 (n_560, wc151, n_215);
  not gc151 (wc151, n_482);
  and g806 (n_564, wc152, n_331);
  not gc152 (wc152, n_487);
  and g807 (n_568, n_490, wc153);
  not gc153 (wc153, n_491);
  and g808 (n_572, n_423, wc154);
  not gc154 (wc154, n_494);
  and g809 (n_576, wc155, n_499);
  not gc155 (wc155, n_500);
  and g810 (n_580, wc156, n_504);
  not gc156 (wc156, n_505);
  and g811 (n_584, wc157, n_509);
  not gc157 (wc157, n_510);
  and g812 (n_612, wc158, n_263);
  not gc158 (wc158, n_518);
  and g813 (n_616, wc159, n_371);
  not gc159 (wc159, n_523);
  and g814 (n_620, n_526, wc160);
  not gc160 (wc160, n_527);
  and g815 (n_624, n_454, wc161);
  not gc161 (wc161, n_530);
  or g816 (n_589, n_586, wc162);
  not gc162 (wc162, n_538);
  or g817 (n_540, wc163, n_196);
  not gc163 (wc163, n_538);
  or g818 (n_545, n_542, wc164);
  not gc164 (wc164, n_538);
  or g819 (n_547, wc165, n_411);
  not gc165 (wc165, n_538);
  or g820 (n_561, n_558, wc166);
  not gc166 (wc166, n_538);
  or g821 (n_565, n_562, wc167);
  not gc167 (wc167, n_538);
  or g822 (n_569, n_566, wc168);
  not gc168 (wc168, n_538);
  or g823 (n_573, n_570, wc169);
  not gc169 (wc169, n_538);
  or g824 (n_577, n_574, wc170);
  not gc170 (wc170, n_538);
  or g825 (n_581, n_578, wc171);
  not gc171 (wc171, n_538);
  or g826 (n_585, n_582, wc172);
  not gc172 (wc172, n_538);
  or g827 (n_629, wc173, n_626);
  not gc173 (wc173, n_590);
  or g828 (n_592, wc174, n_244);
  not gc174 (wc174, n_590);
  or g829 (n_597, n_594, wc175);
  not gc175 (wc175, n_590);
  or g830 (n_599, wc176, n_441);
  not gc176 (wc176, n_590);
  or g831 (n_613, n_610, wc177);
  not gc177 (wc177, n_590);
  or g832 (n_617, wc178, n_614);
  not gc178 (wc178, n_590);
  or g833 (n_621, n_618, wc179);
  not gc179 (wc179, n_590);
  or g834 (n_625, n_622, wc180);
  not gc180 (wc180, n_590);
endmodule

module add_signed_384_GENERIC(A, B, Z);
  input [44:0] A, B;
  output [45:0] Z;
  wire [44:0] A, B;
  wire [45:0] Z;
  add_signed_384_GENERIC_REAL g1(.A ({A[43], A[43:0]}), .B ({B[43],
       B[43:0]}), .Z (Z));
endmodule

module add_signed_384_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [44:0] A, B;
  output [45:0] Z;
  wire [44:0] A, B;
  wire [45:0] Z;
  wire n_140, n_141, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361, n_362, n_363, n_364;
  not g3 (Z[45], n_140);
  nand g4 (n_141, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_146, A[1], B[1]);
  nand g13 (n_150, n_146, n_147, n_148);
  xor g14 (n_149, A[1], B[1]);
  nand g16 (n_151, A[2], B[2]);
  nand g17 (n_152, A[2], n_150);
  nand g18 (n_153, B[2], n_150);
  nand g19 (n_155, n_151, n_152, n_153);
  xor g20 (n_154, A[2], B[2]);
  xor g21 (Z[2], n_150, n_154);
  nand g22 (n_156, A[3], B[3]);
  nand g23 (n_157, A[3], n_155);
  nand g24 (n_158, B[3], n_155);
  nand g25 (n_160, n_156, n_157, n_158);
  xor g26 (n_159, A[3], B[3]);
  xor g27 (Z[3], n_155, n_159);
  nand g28 (n_161, A[4], B[4]);
  nand g29 (n_162, A[4], n_160);
  nand g30 (n_163, B[4], n_160);
  nand g31 (n_165, n_161, n_162, n_163);
  xor g32 (n_164, A[4], B[4]);
  xor g33 (Z[4], n_160, n_164);
  nand g34 (n_166, A[5], B[5]);
  nand g35 (n_167, A[5], n_165);
  nand g36 (n_168, B[5], n_165);
  nand g37 (n_170, n_166, n_167, n_168);
  xor g38 (n_169, A[5], B[5]);
  xor g39 (Z[5], n_165, n_169);
  nand g40 (n_171, A[6], B[6]);
  nand g41 (n_172, A[6], n_170);
  nand g42 (n_173, B[6], n_170);
  nand g43 (n_175, n_171, n_172, n_173);
  xor g44 (n_174, A[6], B[6]);
  xor g45 (Z[6], n_170, n_174);
  nand g46 (n_176, A[7], B[7]);
  nand g47 (n_177, A[7], n_175);
  nand g48 (n_178, B[7], n_175);
  nand g49 (n_180, n_176, n_177, n_178);
  xor g50 (n_179, A[7], B[7]);
  xor g51 (Z[7], n_175, n_179);
  nand g52 (n_181, A[8], B[8]);
  nand g53 (n_182, A[8], n_180);
  nand g54 (n_183, B[8], n_180);
  nand g55 (n_185, n_181, n_182, n_183);
  xor g56 (n_184, A[8], B[8]);
  xor g57 (Z[8], n_180, n_184);
  nand g58 (n_186, A[9], B[9]);
  nand g59 (n_187, A[9], n_185);
  nand g60 (n_188, B[9], n_185);
  nand g61 (n_190, n_186, n_187, n_188);
  xor g62 (n_189, A[9], B[9]);
  xor g63 (Z[9], n_185, n_189);
  nand g64 (n_191, A[10], B[10]);
  nand g65 (n_192, A[10], n_190);
  nand g66 (n_193, B[10], n_190);
  nand g67 (n_195, n_191, n_192, n_193);
  xor g68 (n_194, A[10], B[10]);
  xor g69 (Z[10], n_190, n_194);
  nand g70 (n_196, A[11], B[11]);
  nand g71 (n_197, A[11], n_195);
  nand g72 (n_198, B[11], n_195);
  nand g73 (n_200, n_196, n_197, n_198);
  xor g74 (n_199, A[11], B[11]);
  xor g75 (Z[11], n_195, n_199);
  nand g76 (n_201, A[12], B[12]);
  nand g77 (n_202, A[12], n_200);
  nand g78 (n_203, B[12], n_200);
  nand g79 (n_205, n_201, n_202, n_203);
  xor g80 (n_204, A[12], B[12]);
  xor g81 (Z[12], n_200, n_204);
  nand g82 (n_206, A[13], B[13]);
  nand g83 (n_207, A[13], n_205);
  nand g84 (n_208, B[13], n_205);
  nand g85 (n_210, n_206, n_207, n_208);
  xor g86 (n_209, A[13], B[13]);
  xor g87 (Z[13], n_205, n_209);
  nand g88 (n_211, A[14], B[14]);
  nand g89 (n_212, A[14], n_210);
  nand g90 (n_213, B[14], n_210);
  nand g91 (n_215, n_211, n_212, n_213);
  xor g92 (n_214, A[14], B[14]);
  xor g93 (Z[14], n_210, n_214);
  nand g94 (n_216, A[15], B[15]);
  nand g95 (n_217, A[15], n_215);
  nand g96 (n_218, B[15], n_215);
  nand g97 (n_220, n_216, n_217, n_218);
  xor g98 (n_219, A[15], B[15]);
  xor g99 (Z[15], n_215, n_219);
  nand g100 (n_221, A[16], B[16]);
  nand g101 (n_222, A[16], n_220);
  nand g102 (n_223, B[16], n_220);
  nand g103 (n_225, n_221, n_222, n_223);
  xor g104 (n_224, A[16], B[16]);
  xor g105 (Z[16], n_220, n_224);
  nand g106 (n_226, A[17], B[17]);
  nand g107 (n_227, A[17], n_225);
  nand g108 (n_228, B[17], n_225);
  nand g109 (n_230, n_226, n_227, n_228);
  xor g110 (n_229, A[17], B[17]);
  xor g111 (Z[17], n_225, n_229);
  nand g112 (n_231, A[18], B[18]);
  nand g113 (n_232, A[18], n_230);
  nand g114 (n_233, B[18], n_230);
  nand g115 (n_235, n_231, n_232, n_233);
  xor g116 (n_234, A[18], B[18]);
  xor g117 (Z[18], n_230, n_234);
  nand g118 (n_236, A[19], B[19]);
  nand g119 (n_237, A[19], n_235);
  nand g120 (n_238, B[19], n_235);
  nand g121 (n_240, n_236, n_237, n_238);
  xor g122 (n_239, A[19], B[19]);
  xor g123 (Z[19], n_235, n_239);
  nand g124 (n_241, A[20], B[20]);
  nand g125 (n_242, A[20], n_240);
  nand g126 (n_243, B[20], n_240);
  nand g127 (n_245, n_241, n_242, n_243);
  xor g128 (n_244, A[20], B[20]);
  xor g129 (Z[20], n_240, n_244);
  nand g130 (n_246, A[21], B[21]);
  nand g131 (n_247, A[21], n_245);
  nand g132 (n_248, B[21], n_245);
  nand g133 (n_250, n_246, n_247, n_248);
  xor g134 (n_249, A[21], B[21]);
  xor g135 (Z[21], n_245, n_249);
  nand g136 (n_251, A[22], B[22]);
  nand g137 (n_252, A[22], n_250);
  nand g138 (n_253, B[22], n_250);
  nand g139 (n_255, n_251, n_252, n_253);
  xor g140 (n_254, A[22], B[22]);
  xor g141 (Z[22], n_250, n_254);
  nand g142 (n_256, A[23], B[23]);
  nand g143 (n_257, A[23], n_255);
  nand g144 (n_258, B[23], n_255);
  nand g145 (n_260, n_256, n_257, n_258);
  xor g146 (n_259, A[23], B[23]);
  xor g147 (Z[23], n_255, n_259);
  nand g148 (n_261, A[24], B[24]);
  nand g149 (n_262, A[24], n_260);
  nand g150 (n_263, B[24], n_260);
  nand g151 (n_265, n_261, n_262, n_263);
  xor g152 (n_264, A[24], B[24]);
  xor g153 (Z[24], n_260, n_264);
  nand g154 (n_266, A[25], B[25]);
  nand g155 (n_267, A[25], n_265);
  nand g156 (n_268, B[25], n_265);
  nand g157 (n_270, n_266, n_267, n_268);
  xor g158 (n_269, A[25], B[25]);
  xor g159 (Z[25], n_265, n_269);
  nand g160 (n_271, A[26], B[26]);
  nand g161 (n_272, A[26], n_270);
  nand g162 (n_273, B[26], n_270);
  nand g163 (n_275, n_271, n_272, n_273);
  xor g164 (n_274, A[26], B[26]);
  xor g165 (Z[26], n_270, n_274);
  nand g166 (n_276, A[27], B[27]);
  nand g167 (n_277, A[27], n_275);
  nand g168 (n_278, B[27], n_275);
  nand g169 (n_280, n_276, n_277, n_278);
  xor g170 (n_279, A[27], B[27]);
  xor g171 (Z[27], n_275, n_279);
  nand g172 (n_281, A[28], B[28]);
  nand g173 (n_282, A[28], n_280);
  nand g174 (n_283, B[28], n_280);
  nand g175 (n_285, n_281, n_282, n_283);
  xor g176 (n_284, A[28], B[28]);
  xor g177 (Z[28], n_280, n_284);
  nand g178 (n_286, A[29], B[29]);
  nand g179 (n_287, A[29], n_285);
  nand g180 (n_288, B[29], n_285);
  nand g181 (n_290, n_286, n_287, n_288);
  xor g182 (n_289, A[29], B[29]);
  xor g183 (Z[29], n_285, n_289);
  nand g184 (n_291, A[30], B[30]);
  nand g185 (n_292, A[30], n_290);
  nand g186 (n_293, B[30], n_290);
  nand g187 (n_295, n_291, n_292, n_293);
  xor g188 (n_294, A[30], B[30]);
  xor g189 (Z[30], n_290, n_294);
  nand g190 (n_296, A[31], B[31]);
  nand g191 (n_297, A[31], n_295);
  nand g192 (n_298, B[31], n_295);
  nand g193 (n_300, n_296, n_297, n_298);
  xor g194 (n_299, A[31], B[31]);
  xor g195 (Z[31], n_295, n_299);
  nand g196 (n_301, A[32], B[32]);
  nand g197 (n_302, A[32], n_300);
  nand g198 (n_303, B[32], n_300);
  nand g199 (n_305, n_301, n_302, n_303);
  xor g200 (n_304, A[32], B[32]);
  xor g201 (Z[32], n_300, n_304);
  nand g202 (n_306, A[33], B[33]);
  nand g203 (n_307, A[33], n_305);
  nand g204 (n_308, B[33], n_305);
  nand g205 (n_310, n_306, n_307, n_308);
  xor g206 (n_309, A[33], B[33]);
  xor g207 (Z[33], n_305, n_309);
  nand g208 (n_311, A[34], B[34]);
  nand g209 (n_312, A[34], n_310);
  nand g210 (n_313, B[34], n_310);
  nand g211 (n_315, n_311, n_312, n_313);
  xor g212 (n_314, A[34], B[34]);
  xor g213 (Z[34], n_310, n_314);
  nand g214 (n_316, A[35], B[35]);
  nand g215 (n_317, A[35], n_315);
  nand g216 (n_318, B[35], n_315);
  nand g217 (n_320, n_316, n_317, n_318);
  xor g218 (n_319, A[35], B[35]);
  xor g219 (Z[35], n_315, n_319);
  nand g220 (n_321, A[36], B[36]);
  nand g221 (n_322, A[36], n_320);
  nand g222 (n_323, B[36], n_320);
  nand g223 (n_325, n_321, n_322, n_323);
  xor g224 (n_324, A[36], B[36]);
  xor g225 (Z[36], n_320, n_324);
  nand g226 (n_326, A[37], B[37]);
  nand g227 (n_327, A[37], n_325);
  nand g228 (n_328, B[37], n_325);
  nand g229 (n_330, n_326, n_327, n_328);
  xor g230 (n_329, A[37], B[37]);
  xor g231 (Z[37], n_325, n_329);
  nand g232 (n_331, A[38], B[38]);
  nand g233 (n_332, A[38], n_330);
  nand g234 (n_333, B[38], n_330);
  nand g235 (n_335, n_331, n_332, n_333);
  xor g236 (n_334, A[38], B[38]);
  xor g237 (Z[38], n_330, n_334);
  nand g238 (n_336, A[39], B[39]);
  nand g239 (n_337, A[39], n_335);
  nand g240 (n_338, B[39], n_335);
  nand g241 (n_340, n_336, n_337, n_338);
  xor g242 (n_339, A[39], B[39]);
  xor g243 (Z[39], n_335, n_339);
  nand g244 (n_341, A[40], B[40]);
  nand g245 (n_342, A[40], n_340);
  nand g246 (n_343, B[40], n_340);
  nand g247 (n_345, n_341, n_342, n_343);
  xor g248 (n_344, A[40], B[40]);
  xor g249 (Z[40], n_340, n_344);
  nand g250 (n_346, A[41], B[41]);
  nand g251 (n_347, A[41], n_345);
  nand g252 (n_348, B[41], n_345);
  nand g253 (n_350, n_346, n_347, n_348);
  xor g254 (n_349, A[41], B[41]);
  xor g255 (Z[41], n_345, n_349);
  nand g256 (n_351, A[42], B[42]);
  nand g257 (n_352, A[42], n_350);
  nand g258 (n_353, B[42], n_350);
  nand g259 (n_355, n_351, n_352, n_353);
  xor g260 (n_354, A[42], B[42]);
  xor g261 (Z[42], n_350, n_354);
  nand g262 (n_356, A[43], B[43]);
  nand g263 (n_357, A[43], n_355);
  nand g264 (n_358, B[43], n_355);
  nand g265 (n_360, n_356, n_357, n_358);
  xor g266 (n_359, A[43], B[43]);
  xor g267 (Z[43], n_355, n_359);
  nand g271 (n_140, n_361, n_362, n_363);
  xor g273 (Z[44], n_360, n_364);
  or g275 (n_361, A[44], B[44]);
  xor g276 (n_364, A[44], B[44]);
  or g277 (n_147, wc, n_141);
  not gc (wc, A[1]);
  or g278 (n_148, wc0, n_141);
  not gc0 (wc0, B[1]);
  xnor g279 (Z[1], n_141, n_149);
  or g280 (n_362, A[44], wc1);
  not gc1 (wc1, n_360);
  or g281 (n_363, B[44], wc2);
  not gc2 (wc2, n_360);
endmodule

module add_signed_384_1_GENERIC(A, B, Z);
  input [44:0] A, B;
  output [45:0] Z;
  wire [44:0] A, B;
  wire [45:0] Z;
  add_signed_384_1_GENERIC_REAL g1(.A ({A[44:2], A[0], A[0]}), .B (B),
       .Z (Z));
endmodule

module add_signed_384_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [44:0] A, B;
  output [45:0] Z;
  wire [44:0] A, B;
  wire [45:0] Z;
  wire n_140, n_141, n_144, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_154, n_155, n_156, n_157, n_158, n_160, n_161;
  wire n_162, n_163, n_164, n_166, n_167, n_168, n_169, n_170;
  wire n_172, n_173, n_174, n_175, n_176, n_178, n_179, n_180;
  wire n_181, n_182, n_184, n_185, n_186, n_187, n_188, n_190;
  wire n_191, n_192, n_193, n_194, n_196, n_197, n_198, n_199;
  wire n_200, n_202, n_203, n_204, n_205, n_206, n_208, n_209;
  wire n_210, n_211, n_212, n_214, n_215, n_216, n_217, n_218;
  wire n_220, n_221, n_222, n_223, n_224, n_226, n_227, n_228;
  wire n_229, n_230, n_232, n_233, n_234, n_235, n_236, n_238;
  wire n_239, n_240, n_241, n_242, n_244, n_245, n_246, n_247;
  wire n_248, n_250, n_251, n_252, n_253, n_254, n_256, n_257;
  wire n_258, n_259, n_260, n_262, n_263, n_264, n_265, n_266;
  wire n_268, n_269, n_270, n_271, n_272, n_274, n_275, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_284, n_286, n_288;
  wire n_289, n_291, n_292, n_294, n_296, n_298, n_299, n_301;
  wire n_302, n_304, n_306, n_308, n_309, n_311, n_312, n_314;
  wire n_316, n_318, n_319, n_321, n_322, n_324, n_326, n_328;
  wire n_329, n_331, n_332, n_334, n_336, n_338, n_339, n_341;
  wire n_342, n_344, n_346, n_348, n_349, n_351, n_352, n_354;
  wire n_356, n_358, n_359, n_361, n_362, n_364, n_366, n_368;
  wire n_369, n_371, n_372, n_374, n_376, n_378, n_379, n_381;
  wire n_383, n_384, n_385, n_387, n_388, n_389, n_391, n_392;
  wire n_393, n_394, n_396, n_398, n_400, n_401, n_402, n_404;
  wire n_405, n_406, n_408, n_409, n_411, n_413, n_415, n_416;
  wire n_417, n_419, n_420, n_421, n_423, n_424, n_426, n_428;
  wire n_430, n_431, n_432, n_434, n_435, n_436, n_438, n_439;
  wire n_441, n_443, n_445, n_446, n_447, n_449, n_450, n_451;
  wire n_453, n_454, n_455, n_456, n_458, n_459, n_461, n_462;
  wire n_463, n_465, n_466, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_484, n_487, n_489, n_490, n_491, n_494;
  wire n_497, n_499, n_500, n_502, n_504, n_505, n_507, n_509;
  wire n_510, n_512, n_514, n_515, n_517, n_518, n_520, n_523;
  wire n_525, n_526, n_527, n_530, n_533, n_535, n_536, n_538;
  wire n_540, n_541, n_542, n_544, n_545, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_560, n_561, n_562, n_564, n_565, n_566, n_568;
  wire n_569, n_570, n_572, n_573, n_574, n_576, n_577, n_578;
  wire n_580, n_581, n_582, n_584, n_585, n_586, n_588, n_589;
  wire n_590, n_592, n_593, n_594, n_596, n_597, n_599, n_600;
  wire n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608;
  wire n_609, n_610, n_612, n_613, n_614, n_616, n_617, n_618;
  wire n_620, n_621, n_622, n_624, n_625, n_626, n_628, n_629;
  wire n_630, n_631, n_633, n_634, n_635, n_637, n_638, n_639;
  wire n_640, n_642, n_643, n_644, n_646, n_647, n_648, n_649;
  wire n_651, n_652, n_654, n_655, n_657, n_658, n_659, n_660;
  wire n_662, n_663, n_664, n_666, n_667, n_668, n_669, n_671;
  wire n_672, n_674, n_675, n_677, n_678, n_679, n_680, n_682;
  wire n_683, n_684, n_685, n_687, n_688, n_689, n_690, n_692;
  wire n_693, n_695, n_696, n_698, n_699, n_700, n_701, n_703;
  wire n_704, n_705, n_707, n_708, n_709, n_710, n_712, n_713;
  wire n_715, n_716, n_718, n_719, n_720, n_721, n_723, n_724;
  wire n_725, n_726, n_728, n_729, n_730, n_731, n_733, n_734;
  wire n_736, n_737;
  not g3 (Z[45], n_140);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_141, A[0], B[0]);
  nor g9 (n_144, A[1], B[1]);
  nand g10 (n_147, A[1], B[1]);
  nor g11 (n_154, A[2], B[2]);
  nand g12 (n_149, A[2], B[2]);
  nor g13 (n_150, A[3], B[3]);
  nand g14 (n_151, A[3], B[3]);
  nor g15 (n_160, A[4], B[4]);
  nand g16 (n_155, A[4], B[4]);
  nor g17 (n_156, A[5], B[5]);
  nand g18 (n_157, A[5], B[5]);
  nor g19 (n_166, A[6], B[6]);
  nand g20 (n_161, A[6], B[6]);
  nor g21 (n_162, A[7], B[7]);
  nand g22 (n_163, A[7], B[7]);
  nor g23 (n_172, A[8], B[8]);
  nand g24 (n_167, A[8], B[8]);
  nor g25 (n_168, A[9], B[9]);
  nand g26 (n_169, A[9], B[9]);
  nor g27 (n_178, A[10], B[10]);
  nand g28 (n_173, A[10], B[10]);
  nor g29 (n_174, A[11], B[11]);
  nand g30 (n_175, A[11], B[11]);
  nor g31 (n_184, A[12], B[12]);
  nand g32 (n_179, A[12], B[12]);
  nor g33 (n_180, A[13], B[13]);
  nand g34 (n_181, A[13], B[13]);
  nor g35 (n_190, A[14], B[14]);
  nand g36 (n_185, A[14], B[14]);
  nor g37 (n_186, A[15], B[15]);
  nand g38 (n_187, A[15], B[15]);
  nor g39 (n_196, A[16], B[16]);
  nand g40 (n_191, A[16], B[16]);
  nor g41 (n_192, A[17], B[17]);
  nand g42 (n_193, A[17], B[17]);
  nor g43 (n_202, A[18], B[18]);
  nand g44 (n_197, A[18], B[18]);
  nor g45 (n_198, A[19], B[19]);
  nand g46 (n_199, A[19], B[19]);
  nor g47 (n_208, A[20], B[20]);
  nand g48 (n_203, A[20], B[20]);
  nor g49 (n_204, A[21], B[21]);
  nand g50 (n_205, A[21], B[21]);
  nor g51 (n_214, A[22], B[22]);
  nand g52 (n_209, A[22], B[22]);
  nor g53 (n_210, A[23], B[23]);
  nand g54 (n_211, A[23], B[23]);
  nor g55 (n_220, A[24], B[24]);
  nand g56 (n_215, A[24], B[24]);
  nor g57 (n_216, A[25], B[25]);
  nand g58 (n_217, A[25], B[25]);
  nor g59 (n_226, A[26], B[26]);
  nand g60 (n_221, A[26], B[26]);
  nor g61 (n_222, A[27], B[27]);
  nand g62 (n_223, A[27], B[27]);
  nor g63 (n_232, A[28], B[28]);
  nand g64 (n_227, A[28], B[28]);
  nor g65 (n_228, A[29], B[29]);
  nand g66 (n_229, A[29], B[29]);
  nor g67 (n_238, A[30], B[30]);
  nand g68 (n_233, A[30], B[30]);
  nor g69 (n_234, A[31], B[31]);
  nand g70 (n_235, A[31], B[31]);
  nor g71 (n_244, A[32], B[32]);
  nand g72 (n_239, A[32], B[32]);
  nor g73 (n_240, A[33], B[33]);
  nand g74 (n_241, A[33], B[33]);
  nor g75 (n_250, A[34], B[34]);
  nand g76 (n_245, A[34], B[34]);
  nor g77 (n_246, A[35], B[35]);
  nand g78 (n_247, A[35], B[35]);
  nor g79 (n_256, A[36], B[36]);
  nand g80 (n_251, A[36], B[36]);
  nor g81 (n_252, A[37], B[37]);
  nand g82 (n_253, A[37], B[37]);
  nor g83 (n_262, A[38], B[38]);
  nand g84 (n_257, A[38], B[38]);
  nor g85 (n_258, A[39], B[39]);
  nand g86 (n_259, A[39], B[39]);
  nor g87 (n_268, A[40], B[40]);
  nand g88 (n_263, A[40], B[40]);
  nor g89 (n_264, A[41], B[41]);
  nand g90 (n_265, A[41], B[41]);
  nor g91 (n_274, A[42], B[42]);
  nand g92 (n_269, A[42], B[42]);
  nor g93 (n_270, A[43], B[43]);
  nand g94 (n_271, A[43], B[43]);
  nand g99 (n_275, n_147, n_148);
  nor g100 (n_152, n_149, n_150);
  nor g103 (n_278, n_154, n_150);
  nor g104 (n_158, n_155, n_156);
  nor g107 (n_284, n_160, n_156);
  nor g108 (n_164, n_161, n_162);
  nor g111 (n_286, n_166, n_162);
  nor g112 (n_170, n_167, n_168);
  nor g115 (n_294, n_172, n_168);
  nor g116 (n_176, n_173, n_174);
  nor g119 (n_296, n_178, n_174);
  nor g120 (n_182, n_179, n_180);
  nor g123 (n_304, n_184, n_180);
  nor g124 (n_188, n_185, n_186);
  nor g127 (n_306, n_190, n_186);
  nor g128 (n_194, n_191, n_192);
  nor g131 (n_314, n_196, n_192);
  nor g132 (n_200, n_197, n_198);
  nor g135 (n_316, n_202, n_198);
  nor g136 (n_206, n_203, n_204);
  nor g139 (n_324, n_208, n_204);
  nor g140 (n_212, n_209, n_210);
  nor g143 (n_326, n_214, n_210);
  nor g144 (n_218, n_215, n_216);
  nor g147 (n_334, n_220, n_216);
  nor g148 (n_224, n_221, n_222);
  nor g151 (n_336, n_226, n_222);
  nor g152 (n_230, n_227, n_228);
  nor g155 (n_344, n_232, n_228);
  nor g156 (n_236, n_233, n_234);
  nor g159 (n_346, n_238, n_234);
  nor g160 (n_242, n_239, n_240);
  nor g163 (n_354, n_244, n_240);
  nor g164 (n_248, n_245, n_246);
  nor g167 (n_356, n_250, n_246);
  nor g168 (n_254, n_251, n_252);
  nor g171 (n_364, n_256, n_252);
  nor g172 (n_260, n_257, n_258);
  nor g175 (n_366, n_262, n_258);
  nor g176 (n_266, n_263, n_264);
  nor g179 (n_374, n_268, n_264);
  nor g180 (n_272, n_269, n_270);
  nor g183 (n_376, n_274, n_270);
  nand g186 (n_633, n_149, n_277);
  nand g187 (n_280, n_278, n_275);
  nand g188 (n_381, n_279, n_280);
  nor g189 (n_282, n_166, n_281);
  nand g198 (n_389, n_284, n_286);
  nor g199 (n_292, n_178, n_291);
  nand g208 (n_396, n_294, n_296);
  nor g209 (n_302, n_190, n_301);
  nand g218 (n_404, n_304, n_306);
  nor g219 (n_312, n_202, n_311);
  nand g228 (n_411, n_314, n_316);
  nor g229 (n_322, n_214, n_321);
  nand g238 (n_419, n_324, n_326);
  nor g239 (n_332, n_226, n_331);
  nand g248 (n_426, n_334, n_336);
  nor g249 (n_342, n_238, n_341);
  nand g258 (n_434, n_344, n_346);
  nor g259 (n_352, n_250, n_351);
  nand g268 (n_441, n_354, n_356);
  nor g269 (n_362, n_262, n_361);
  nand g278 (n_449, n_364, n_366);
  nor g279 (n_372, n_274, n_371);
  nand g288 (n_458, n_374, n_376);
  nand g291 (n_637, n_155, n_383);
  nand g292 (n_384, n_284, n_381);
  nand g293 (n_639, n_281, n_384);
  nand g296 (n_642, n_387, n_388);
  nand g299 (n_459, n_391, n_392);
  nor g300 (n_394, n_184, n_393);
  nor g303 (n_469, n_184, n_396);
  nor g309 (n_402, n_400, n_393);
  nor g312 (n_475, n_396, n_400);
  nor g313 (n_406, n_404, n_393);
  nor g316 (n_478, n_396, n_404);
  nor g317 (n_409, n_208, n_408);
  nor g320 (n_548, n_208, n_411);
  nor g326 (n_417, n_415, n_408);
  nor g329 (n_554, n_411, n_415);
  nor g330 (n_421, n_419, n_408);
  nor g333 (n_484, n_411, n_419);
  nor g334 (n_424, n_232, n_423);
  nor g337 (n_497, n_232, n_426);
  nor g343 (n_432, n_430, n_423);
  nor g346 (n_507, n_426, n_430);
  nor g347 (n_436, n_434, n_423);
  nor g350 (n_512, n_426, n_434);
  nor g351 (n_439, n_256, n_438);
  nor g354 (n_600, n_256, n_441);
  nor g360 (n_447, n_445, n_438);
  nor g363 (n_606, n_441, n_445);
  nor g364 (n_451, n_449, n_438);
  nor g367 (n_520, n_441, n_449);
  nor g368 (n_456, n_453, n_454);
  nor g371 (n_533, n_453, n_458);
  nand g374 (n_646, n_167, n_461);
  nand g375 (n_462, n_294, n_459);
  nand g376 (n_648, n_291, n_462);
  nand g379 (n_651, n_465, n_466);
  nand g382 (n_654, n_393, n_468);
  nand g383 (n_471, n_469, n_459);
  nand g384 (n_657, n_470, n_471);
  nand g385 (n_474, n_472, n_459);
  nand g386 (n_659, n_473, n_474);
  nand g387 (n_477, n_475, n_459);
  nand g388 (n_662, n_476, n_477);
  nand g389 (n_480, n_478, n_459);
  nand g390 (n_538, n_479, n_480);
  nor g391 (n_482, n_220, n_481);
  nand g400 (n_562, n_334, n_484);
  nor g401 (n_491, n_489, n_481);
  nor g406 (n_494, n_426, n_481);
  nand g415 (n_574, n_484, n_497);
  nand g420 (n_578, n_484, n_502);
  nand g425 (n_582, n_484, n_507);
  nand g430 (n_586, n_484, n_512);
  nor g431 (n_518, n_268, n_517);
  nand g440 (n_614, n_374, n_520);
  nor g441 (n_527, n_525, n_517);
  nor g446 (n_530, n_458, n_517);
  nand g455 (n_626, n_520, n_533);
  nand g458 (n_666, n_191, n_540);
  nand g459 (n_541, n_314, n_538);
  nand g460 (n_668, n_311, n_541);
  nand g463 (n_671, n_544, n_545);
  nand g466 (n_674, n_408, n_547);
  nand g467 (n_550, n_548, n_538);
  nand g468 (n_677, n_549, n_550);
  nand g469 (n_553, n_551, n_538);
  nand g470 (n_679, n_552, n_553);
  nand g471 (n_556, n_554, n_538);
  nand g472 (n_682, n_555, n_556);
  nand g473 (n_557, n_484, n_538);
  nand g474 (n_684, n_481, n_557);
  nand g477 (n_687, n_560, n_561);
  nand g480 (n_689, n_564, n_565);
  nand g483 (n_692, n_568, n_569);
  nand g486 (n_695, n_572, n_573);
  nand g489 (n_698, n_576, n_577);
  nand g492 (n_700, n_580, n_581);
  nand g495 (n_703, n_584, n_585);
  nand g498 (n_590, n_588, n_589);
  nand g501 (n_707, n_239, n_592);
  nand g502 (n_593, n_354, n_590);
  nand g503 (n_709, n_351, n_593);
  nand g506 (n_712, n_596, n_597);
  nand g509 (n_715, n_438, n_599);
  nand g510 (n_602, n_600, n_590);
  nand g511 (n_718, n_601, n_602);
  nand g512 (n_605, n_603, n_590);
  nand g513 (n_720, n_604, n_605);
  nand g514 (n_608, n_606, n_590);
  nand g515 (n_723, n_607, n_608);
  nand g516 (n_609, n_520, n_590);
  nand g517 (n_725, n_517, n_609);
  nand g520 (n_728, n_612, n_613);
  nand g523 (n_730, n_616, n_617);
  nand g526 (n_733, n_620, n_621);
  nand g529 (n_736, n_624, n_625);
  nand g532 (n_140, n_628, n_629);
  xnor g536 (Z[2], n_275, n_631);
  xnor g539 (Z[3], n_633, n_634);
  xnor g541 (Z[4], n_381, n_635);
  xnor g544 (Z[5], n_637, n_638);
  xnor g546 (Z[6], n_639, n_640);
  xnor g549 (Z[7], n_642, n_643);
  xnor g551 (Z[8], n_459, n_644);
  xnor g554 (Z[9], n_646, n_647);
  xnor g556 (Z[10], n_648, n_649);
  xnor g559 (Z[11], n_651, n_652);
  xnor g562 (Z[12], n_654, n_655);
  xnor g565 (Z[13], n_657, n_658);
  xnor g567 (Z[14], n_659, n_660);
  xnor g570 (Z[15], n_662, n_663);
  xnor g572 (Z[16], n_538, n_664);
  xnor g575 (Z[17], n_666, n_667);
  xnor g577 (Z[18], n_668, n_669);
  xnor g580 (Z[19], n_671, n_672);
  xnor g583 (Z[20], n_674, n_675);
  xnor g586 (Z[21], n_677, n_678);
  xnor g588 (Z[22], n_679, n_680);
  xnor g591 (Z[23], n_682, n_683);
  xnor g593 (Z[24], n_684, n_685);
  xnor g596 (Z[25], n_687, n_688);
  xnor g598 (Z[26], n_689, n_690);
  xnor g601 (Z[27], n_692, n_693);
  xnor g604 (Z[28], n_695, n_696);
  xnor g607 (Z[29], n_698, n_699);
  xnor g609 (Z[30], n_700, n_701);
  xnor g612 (Z[31], n_703, n_704);
  xnor g614 (Z[32], n_590, n_705);
  xnor g617 (Z[33], n_707, n_708);
  xnor g619 (Z[34], n_709, n_710);
  xnor g622 (Z[35], n_712, n_713);
  xnor g625 (Z[36], n_715, n_716);
  xnor g628 (Z[37], n_718, n_719);
  xnor g630 (Z[38], n_720, n_721);
  xnor g633 (Z[39], n_723, n_724);
  xnor g635 (Z[40], n_725, n_726);
  xnor g638 (Z[41], n_728, n_729);
  xnor g640 (Z[42], n_730, n_731);
  xnor g643 (Z[43], n_733, n_734);
  xnor g646 (Z[44], n_736, n_737);
  and g649 (n_453, A[44], B[44]);
  or g650 (n_455, A[44], B[44]);
  and g651 (n_351, wc, n_241);
  not gc (wc, n_242);
  and g652 (n_358, wc0, n_247);
  not gc0 (wc0, n_248);
  and g653 (n_361, wc1, n_253);
  not gc1 (wc1, n_254);
  and g654 (n_368, wc2, n_259);
  not gc2 (wc2, n_260);
  and g655 (n_371, wc3, n_265);
  not gc3 (wc3, n_266);
  and g656 (n_378, wc4, n_271);
  not gc4 (wc4, n_272);
  and g657 (n_311, wc5, n_193);
  not gc5 (wc5, n_194);
  and g658 (n_318, wc6, n_199);
  not gc6 (wc6, n_200);
  and g659 (n_321, wc7, n_205);
  not gc7 (wc7, n_206);
  and g660 (n_328, wc8, n_211);
  not gc8 (wc8, n_212);
  and g661 (n_331, wc9, n_217);
  not gc9 (wc9, n_218);
  and g662 (n_338, wc10, n_223);
  not gc10 (wc10, n_224);
  and g663 (n_341, wc11, n_229);
  not gc11 (wc11, n_230);
  and g664 (n_348, wc12, n_235);
  not gc12 (wc12, n_236);
  and g665 (n_291, wc13, n_169);
  not gc13 (wc13, n_170);
  and g666 (n_298, wc14, n_175);
  not gc14 (wc14, n_176);
  and g667 (n_301, wc15, n_181);
  not gc15 (wc15, n_182);
  and g668 (n_308, wc16, n_187);
  not gc16 (wc16, n_188);
  and g669 (n_281, wc17, n_157);
  not gc17 (wc17, n_158);
  and g670 (n_288, wc18, n_163);
  not gc18 (wc18, n_164);
  and g671 (n_279, wc19, n_151);
  not gc19 (wc19, n_152);
  or g672 (n_148, n_141, n_144);
  or g673 (n_385, wc20, n_166);
  not gc20 (wc20, n_284);
  or g674 (n_463, wc21, n_178);
  not gc21 (wc21, n_294);
  or g675 (n_400, wc22, n_190);
  not gc22 (wc22, n_304);
  or g676 (n_542, wc23, n_202);
  not gc23 (wc23, n_314);
  or g677 (n_415, wc24, n_214);
  not gc24 (wc24, n_324);
  or g678 (n_489, wc25, n_226);
  not gc25 (wc25, n_334);
  or g679 (n_430, wc26, n_238);
  not gc26 (wc26, n_344);
  or g680 (n_594, wc27, n_250);
  not gc27 (wc27, n_354);
  or g681 (n_445, wc28, n_262);
  not gc28 (wc28, n_364);
  or g682 (n_525, wc29, n_274);
  not gc29 (wc29, n_374);
  or g683 (n_630, wc30, n_144);
  not gc30 (wc30, n_147);
  or g684 (n_631, wc31, n_154);
  not gc31 (wc31, n_149);
  or g685 (n_634, wc32, n_150);
  not gc32 (wc32, n_151);
  or g686 (n_635, wc33, n_160);
  not gc33 (wc33, n_155);
  or g687 (n_638, wc34, n_156);
  not gc34 (wc34, n_157);
  or g688 (n_640, wc35, n_166);
  not gc35 (wc35, n_161);
  or g689 (n_643, wc36, n_162);
  not gc36 (wc36, n_163);
  or g690 (n_644, wc37, n_172);
  not gc37 (wc37, n_167);
  or g691 (n_647, wc38, n_168);
  not gc38 (wc38, n_169);
  or g692 (n_649, wc39, n_178);
  not gc39 (wc39, n_173);
  or g693 (n_652, wc40, n_174);
  not gc40 (wc40, n_175);
  or g694 (n_655, wc41, n_184);
  not gc41 (wc41, n_179);
  or g695 (n_658, wc42, n_180);
  not gc42 (wc42, n_181);
  or g696 (n_660, wc43, n_190);
  not gc43 (wc43, n_185);
  or g697 (n_663, wc44, n_186);
  not gc44 (wc44, n_187);
  or g698 (n_664, wc45, n_196);
  not gc45 (wc45, n_191);
  or g699 (n_667, wc46, n_192);
  not gc46 (wc46, n_193);
  or g700 (n_669, wc47, n_202);
  not gc47 (wc47, n_197);
  or g701 (n_672, wc48, n_198);
  not gc48 (wc48, n_199);
  or g702 (n_675, wc49, n_208);
  not gc49 (wc49, n_203);
  or g703 (n_678, wc50, n_204);
  not gc50 (wc50, n_205);
  or g704 (n_680, wc51, n_214);
  not gc51 (wc51, n_209);
  or g705 (n_683, wc52, n_210);
  not gc52 (wc52, n_211);
  or g706 (n_685, wc53, n_220);
  not gc53 (wc53, n_215);
  or g707 (n_688, wc54, n_216);
  not gc54 (wc54, n_217);
  or g708 (n_690, wc55, n_226);
  not gc55 (wc55, n_221);
  or g709 (n_693, wc56, n_222);
  not gc56 (wc56, n_223);
  or g710 (n_696, wc57, n_232);
  not gc57 (wc57, n_227);
  or g711 (n_699, wc58, n_228);
  not gc58 (wc58, n_229);
  or g712 (n_701, wc59, n_238);
  not gc59 (wc59, n_233);
  or g713 (n_704, wc60, n_234);
  not gc60 (wc60, n_235);
  or g714 (n_705, wc61, n_244);
  not gc61 (wc61, n_239);
  or g715 (n_708, wc62, n_240);
  not gc62 (wc62, n_241);
  or g716 (n_710, wc63, n_250);
  not gc63 (wc63, n_245);
  or g717 (n_713, wc64, n_246);
  not gc64 (wc64, n_247);
  or g718 (n_716, wc65, n_256);
  not gc65 (wc65, n_251);
  or g719 (n_719, wc66, n_252);
  not gc66 (wc66, n_253);
  or g720 (n_721, wc67, n_262);
  not gc67 (wc67, n_257);
  or g721 (n_724, wc68, n_258);
  not gc68 (wc68, n_259);
  or g722 (n_726, wc69, n_268);
  not gc69 (wc69, n_263);
  or g723 (n_729, wc70, n_264);
  not gc70 (wc70, n_265);
  or g724 (n_731, wc71, n_274);
  not gc71 (wc71, n_269);
  or g725 (n_734, wc72, n_270);
  not gc72 (wc72, n_271);
  and g726 (n_359, wc73, n_356);
  not gc73 (wc73, n_351);
  and g727 (n_369, wc74, n_366);
  not gc74 (wc74, n_361);
  and g728 (n_379, wc75, n_376);
  not gc75 (wc75, n_371);
  and g729 (n_319, wc76, n_316);
  not gc76 (wc76, n_311);
  and g730 (n_329, wc77, n_326);
  not gc77 (wc77, n_321);
  and g731 (n_339, wc78, n_336);
  not gc78 (wc78, n_331);
  and g732 (n_349, wc79, n_346);
  not gc79 (wc79, n_341);
  and g733 (n_299, wc80, n_296);
  not gc80 (wc80, n_291);
  and g734 (n_309, wc81, n_306);
  not gc81 (wc81, n_301);
  and g735 (n_289, wc82, n_286);
  not gc82 (wc82, n_281);
  and g736 (n_472, wc83, n_304);
  not gc83 (wc83, n_396);
  and g737 (n_551, wc84, n_324);
  not gc84 (wc84, n_411);
  and g738 (n_502, wc85, n_344);
  not gc85 (wc85, n_426);
  and g739 (n_603, wc86, n_364);
  not gc86 (wc86, n_441);
  xor g740 (Z[1], n_141, n_630);
  or g741 (n_737, wc87, n_453);
  not gc87 (wc87, n_455);
  and g742 (n_438, wc88, n_358);
  not gc88 (wc88, n_359);
  and g743 (n_450, wc89, n_368);
  not gc89 (wc89, n_369);
  and g744 (n_454, wc90, n_378);
  not gc90 (wc90, n_379);
  and g745 (n_408, wc91, n_318);
  not gc91 (wc91, n_319);
  and g746 (n_420, wc92, n_328);
  not gc92 (wc92, n_329);
  and g747 (n_423, wc93, n_338);
  not gc93 (wc93, n_339);
  and g748 (n_435, wc94, n_348);
  not gc94 (wc94, n_349);
  and g749 (n_393, wc95, n_298);
  not gc95 (wc95, n_299);
  and g750 (n_405, wc96, n_308);
  not gc96 (wc96, n_309);
  and g751 (n_391, wc97, n_288);
  not gc97 (wc97, n_289);
  or g752 (n_277, wc98, n_154);
  not gc98 (wc98, n_275);
  and g753 (n_387, wc99, n_161);
  not gc99 (wc99, n_282);
  and g754 (n_465, wc100, n_173);
  not gc100 (wc100, n_292);
  and g755 (n_401, wc101, n_185);
  not gc101 (wc101, n_302);
  and g756 (n_544, wc102, n_197);
  not gc102 (wc102, n_312);
  and g757 (n_416, wc103, n_209);
  not gc103 (wc103, n_322);
  and g758 (n_490, wc104, n_221);
  not gc104 (wc104, n_332);
  and g759 (n_431, wc105, n_233);
  not gc105 (wc105, n_342);
  and g760 (n_596, wc106, n_245);
  not gc106 (wc106, n_352);
  and g761 (n_446, wc107, n_257);
  not gc107 (wc107, n_362);
  and g762 (n_526, wc108, n_269);
  not gc108 (wc108, n_372);
  or g763 (n_558, wc109, n_220);
  not gc109 (wc109, n_484);
  or g764 (n_566, n_489, wc110);
  not gc110 (wc110, n_484);
  or g765 (n_570, wc111, n_426);
  not gc111 (wc111, n_484);
  or g766 (n_610, wc112, n_268);
  not gc112 (wc112, n_520);
  or g767 (n_618, n_525, wc113);
  not gc113 (wc113, n_520);
  or g768 (n_622, wc114, n_458);
  not gc114 (wc114, n_520);
  and g769 (n_398, wc115, n_304);
  not gc115 (wc115, n_393);
  and g770 (n_413, wc116, n_324);
  not gc116 (wc116, n_408);
  and g771 (n_428, wc117, n_344);
  not gc117 (wc117, n_423);
  and g772 (n_443, wc118, n_364);
  not gc118 (wc118, n_438);
  and g773 (n_517, n_450, wc119);
  not gc119 (wc119, n_451);
  and g774 (n_535, n_455, wc120);
  not gc120 (wc120, n_456);
  and g775 (n_481, n_420, wc121);
  not gc121 (wc121, n_421);
  and g776 (n_514, n_435, wc122);
  not gc122 (wc122, n_436);
  and g777 (n_479, n_405, wc123);
  not gc123 (wc123, n_406);
  or g778 (n_392, n_389, wc124);
  not gc124 (wc124, n_381);
  or g779 (n_383, wc125, n_160);
  not gc125 (wc125, n_381);
  or g780 (n_388, n_385, wc126);
  not gc126 (wc126, n_381);
  and g781 (n_470, wc127, n_179);
  not gc127 (wc127, n_394);
  and g782 (n_473, wc128, n_301);
  not gc128 (wc128, n_398);
  and g783 (n_476, n_401, wc129);
  not gc129 (wc129, n_402);
  and g784 (n_549, wc130, n_203);
  not gc130 (wc130, n_409);
  and g785 (n_552, wc131, n_321);
  not gc131 (wc131, n_413);
  and g786 (n_555, n_416, wc132);
  not gc132 (wc132, n_417);
  and g787 (n_499, wc133, n_227);
  not gc133 (wc133, n_424);
  and g788 (n_504, wc134, n_341);
  not gc134 (wc134, n_428);
  and g789 (n_509, n_431, wc135);
  not gc135 (wc135, n_432);
  and g790 (n_601, wc136, n_251);
  not gc136 (wc136, n_439);
  and g791 (n_604, wc137, n_361);
  not gc137 (wc137, n_443);
  and g792 (n_607, n_446, wc138);
  not gc138 (wc138, n_447);
  and g793 (n_536, wc139, n_533);
  not gc139 (wc139, n_517);
  and g794 (n_515, wc140, n_512);
  not gc140 (wc140, n_481);
  and g795 (n_487, wc141, n_334);
  not gc141 (wc141, n_481);
  and g796 (n_500, wc142, n_497);
  not gc142 (wc142, n_481);
  and g797 (n_505, wc143, n_502);
  not gc143 (wc143, n_481);
  and g798 (n_510, wc144, n_507);
  not gc144 (wc144, n_481);
  and g799 (n_523, wc145, n_374);
  not gc145 (wc145, n_517);
  and g800 (n_628, wc146, n_535);
  not gc146 (wc146, n_536);
  and g801 (n_588, wc147, n_514);
  not gc147 (wc147, n_515);
  or g802 (n_461, wc148, n_172);
  not gc148 (wc148, n_459);
  or g803 (n_466, n_463, wc149);
  not gc149 (wc149, n_459);
  or g804 (n_468, wc150, n_396);
  not gc150 (wc150, n_459);
  and g805 (n_560, wc151, n_215);
  not gc151 (wc151, n_482);
  and g806 (n_564, wc152, n_331);
  not gc152 (wc152, n_487);
  and g807 (n_568, n_490, wc153);
  not gc153 (wc153, n_491);
  and g808 (n_572, n_423, wc154);
  not gc154 (wc154, n_494);
  and g809 (n_576, wc155, n_499);
  not gc155 (wc155, n_500);
  and g810 (n_580, wc156, n_504);
  not gc156 (wc156, n_505);
  and g811 (n_584, wc157, n_509);
  not gc157 (wc157, n_510);
  and g812 (n_612, wc158, n_263);
  not gc158 (wc158, n_518);
  and g813 (n_616, wc159, n_371);
  not gc159 (wc159, n_523);
  and g814 (n_620, n_526, wc160);
  not gc160 (wc160, n_527);
  and g815 (n_624, n_454, wc161);
  not gc161 (wc161, n_530);
  or g816 (n_589, n_586, wc162);
  not gc162 (wc162, n_538);
  or g817 (n_540, wc163, n_196);
  not gc163 (wc163, n_538);
  or g818 (n_545, n_542, wc164);
  not gc164 (wc164, n_538);
  or g819 (n_547, wc165, n_411);
  not gc165 (wc165, n_538);
  or g820 (n_561, n_558, wc166);
  not gc166 (wc166, n_538);
  or g821 (n_565, n_562, wc167);
  not gc167 (wc167, n_538);
  or g822 (n_569, n_566, wc168);
  not gc168 (wc168, n_538);
  or g823 (n_573, n_570, wc169);
  not gc169 (wc169, n_538);
  or g824 (n_577, n_574, wc170);
  not gc170 (wc170, n_538);
  or g825 (n_581, n_578, wc171);
  not gc171 (wc171, n_538);
  or g826 (n_585, n_582, wc172);
  not gc172 (wc172, n_538);
  or g827 (n_629, wc173, n_626);
  not gc173 (wc173, n_590);
  or g828 (n_592, wc174, n_244);
  not gc174 (wc174, n_590);
  or g829 (n_597, n_594, wc175);
  not gc175 (wc175, n_590);
  or g830 (n_599, wc176, n_441);
  not gc176 (wc176, n_590);
  or g831 (n_613, n_610, wc177);
  not gc177 (wc177, n_590);
  or g832 (n_617, wc178, n_614);
  not gc178 (wc178, n_590);
  or g833 (n_621, n_618, wc179);
  not gc179 (wc179, n_590);
  or g834 (n_625, n_622, wc180);
  not gc180 (wc180, n_590);
endmodule

module add_signed_384_2_GENERIC(A, B, Z);
  input [44:0] A, B;
  output [45:0] Z;
  wire [44:0] A, B;
  wire [45:0] Z;
  add_signed_384_2_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_398_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [43:0] A, B;
  output [44:0] Z;
  wire [43:0] A, B;
  wire [44:0] Z;
  wire n_137, n_138, n_141, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_151, n_152, n_153, n_154, n_155, n_157, n_158;
  wire n_159, n_160, n_161, n_163, n_164, n_165, n_166, n_167;
  wire n_169, n_170, n_171, n_172, n_173, n_175, n_176, n_177;
  wire n_178, n_179, n_181, n_182, n_183, n_184, n_185, n_187;
  wire n_188, n_189, n_190, n_191, n_193, n_194, n_195, n_196;
  wire n_197, n_199, n_200, n_201, n_202, n_203, n_205, n_206;
  wire n_207, n_208, n_209, n_211, n_212, n_213, n_214, n_215;
  wire n_217, n_218, n_219, n_220, n_221, n_223, n_224, n_225;
  wire n_226, n_227, n_229, n_230, n_231, n_232, n_233, n_235;
  wire n_236, n_237, n_238, n_239, n_241, n_242, n_243, n_244;
  wire n_245, n_247, n_248, n_249, n_250, n_251, n_253, n_254;
  wire n_255, n_256, n_257, n_259, n_260, n_261, n_262, n_263;
  wire n_265, n_266, n_267, n_268, n_269, n_271, n_272, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_281, n_283, n_285;
  wire n_286, n_288, n_289, n_291, n_293, n_295, n_296, n_298;
  wire n_299, n_301, n_303, n_305, n_306, n_308, n_309, n_311;
  wire n_313, n_315, n_316, n_318, n_319, n_321, n_323, n_325;
  wire n_326, n_328, n_329, n_331, n_333, n_335, n_336, n_338;
  wire n_339, n_341, n_343, n_345, n_346, n_348, n_349, n_351;
  wire n_353, n_355, n_356, n_358, n_359, n_361, n_363, n_365;
  wire n_366, n_368, n_369, n_371, n_373, n_375, n_376, n_378;
  wire n_380, n_381, n_382, n_384, n_385, n_386, n_388, n_389;
  wire n_390, n_391, n_393, n_395, n_397, n_398, n_399, n_401;
  wire n_402, n_403, n_405, n_406, n_408, n_410, n_412, n_413;
  wire n_414, n_416, n_417, n_418, n_420, n_421, n_423, n_425;
  wire n_427, n_428, n_429, n_431, n_432, n_433, n_435, n_436;
  wire n_438, n_440, n_442, n_443, n_444, n_446, n_447, n_448;
  wire n_450, n_452, n_453, n_454, n_456, n_457, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_469, n_470, n_471, n_472, n_473, n_475, n_478, n_480;
  wire n_481, n_482, n_485, n_488, n_490, n_491, n_493, n_495;
  wire n_496, n_498, n_500, n_501, n_503, n_505, n_506, n_508;
  wire n_509, n_511, n_514, n_516, n_517, n_518, n_521, n_522;
  wire n_523, n_526, n_528, n_529, n_530, n_532, n_533, n_535;
  wire n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543;
  wire n_544, n_545, n_546, n_548, n_549, n_550, n_552, n_553;
  wire n_554, n_556, n_557, n_558, n_560, n_561, n_562, n_564;
  wire n_565, n_566, n_568, n_569, n_570, n_572, n_573, n_574;
  wire n_576, n_577, n_578, n_580, n_581, n_582, n_584, n_585;
  wire n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594;
  wire n_595, n_596, n_597, n_598, n_600, n_601, n_602, n_604;
  wire n_605, n_606, n_608, n_609, n_610, n_612, n_613, n_614;
  wire n_615, n_617, n_618, n_619, n_621, n_622, n_623, n_624;
  wire n_626, n_627, n_628, n_630, n_631, n_632, n_633, n_635;
  wire n_636, n_638, n_639, n_641, n_642, n_643, n_644, n_646;
  wire n_647, n_648, n_650, n_651, n_652, n_653, n_655, n_656;
  wire n_658, n_659, n_661, n_662, n_663, n_664, n_666, n_667;
  wire n_668, n_669, n_671, n_672, n_673, n_674, n_676, n_677;
  wire n_679, n_680, n_682, n_683, n_684, n_685, n_687, n_688;
  wire n_689, n_691, n_692, n_693, n_694, n_696, n_697, n_699;
  wire n_700, n_702, n_703, n_704, n_705, n_707, n_708, n_709;
  wire n_710, n_712, n_713, n_714, n_715, n_717, n_718;
  not g3 (Z[44], n_137);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_138, A[0], B[0]);
  nor g9 (n_141, A[1], B[1]);
  nand g10 (n_144, A[1], B[1]);
  nor g11 (n_151, A[2], B[2]);
  nand g12 (n_146, A[2], B[2]);
  nor g13 (n_147, A[3], B[3]);
  nand g14 (n_148, A[3], B[3]);
  nor g15 (n_157, A[4], B[4]);
  nand g16 (n_152, A[4], B[4]);
  nor g17 (n_153, A[5], B[5]);
  nand g18 (n_154, A[5], B[5]);
  nor g19 (n_163, A[6], B[6]);
  nand g20 (n_158, A[6], B[6]);
  nor g21 (n_159, A[7], B[7]);
  nand g22 (n_160, A[7], B[7]);
  nor g23 (n_169, A[8], B[8]);
  nand g24 (n_164, A[8], B[8]);
  nor g25 (n_165, A[9], B[9]);
  nand g26 (n_166, A[9], B[9]);
  nor g27 (n_175, A[10], B[10]);
  nand g28 (n_170, A[10], B[10]);
  nor g29 (n_171, A[11], B[11]);
  nand g30 (n_172, A[11], B[11]);
  nor g31 (n_181, A[12], B[12]);
  nand g32 (n_176, A[12], B[12]);
  nor g33 (n_177, A[13], B[13]);
  nand g34 (n_178, A[13], B[13]);
  nor g35 (n_187, A[14], B[14]);
  nand g36 (n_182, A[14], B[14]);
  nor g37 (n_183, A[15], B[15]);
  nand g38 (n_184, A[15], B[15]);
  nor g39 (n_193, A[16], B[16]);
  nand g40 (n_188, A[16], B[16]);
  nor g41 (n_189, A[17], B[17]);
  nand g42 (n_190, A[17], B[17]);
  nor g43 (n_199, A[18], B[18]);
  nand g44 (n_194, A[18], B[18]);
  nor g45 (n_195, A[19], B[19]);
  nand g46 (n_196, A[19], B[19]);
  nor g47 (n_205, A[20], B[20]);
  nand g48 (n_200, A[20], B[20]);
  nor g49 (n_201, A[21], B[21]);
  nand g50 (n_202, A[21], B[21]);
  nor g51 (n_211, A[22], B[22]);
  nand g52 (n_206, A[22], B[22]);
  nor g53 (n_207, A[23], B[23]);
  nand g54 (n_208, A[23], B[23]);
  nor g55 (n_217, A[24], B[24]);
  nand g56 (n_212, A[24], B[24]);
  nor g57 (n_213, A[25], B[25]);
  nand g58 (n_214, A[25], B[25]);
  nor g59 (n_223, A[26], B[26]);
  nand g60 (n_218, A[26], B[26]);
  nor g61 (n_219, A[27], B[27]);
  nand g62 (n_220, A[27], B[27]);
  nor g63 (n_229, A[28], B[28]);
  nand g64 (n_224, A[28], B[28]);
  nor g65 (n_225, A[29], B[29]);
  nand g66 (n_226, A[29], B[29]);
  nor g67 (n_235, A[30], B[30]);
  nand g68 (n_230, A[30], B[30]);
  nor g69 (n_231, A[31], B[31]);
  nand g70 (n_232, A[31], B[31]);
  nor g71 (n_241, A[32], B[32]);
  nand g72 (n_236, A[32], B[32]);
  nor g73 (n_237, A[33], B[33]);
  nand g74 (n_238, A[33], B[33]);
  nor g75 (n_247, A[34], B[34]);
  nand g76 (n_242, A[34], B[34]);
  nor g77 (n_243, A[35], B[35]);
  nand g78 (n_244, A[35], B[35]);
  nor g79 (n_253, A[36], B[36]);
  nand g80 (n_248, A[36], B[36]);
  nor g81 (n_249, A[37], B[37]);
  nand g82 (n_250, A[37], B[37]);
  nor g83 (n_259, A[38], B[38]);
  nand g84 (n_254, A[38], B[38]);
  nor g85 (n_255, A[39], B[39]);
  nand g86 (n_256, A[39], B[39]);
  nor g87 (n_265, A[40], B[40]);
  nand g88 (n_260, A[40], B[40]);
  nor g89 (n_261, A[41], B[41]);
  nand g90 (n_262, A[41], B[41]);
  nor g91 (n_271, A[42], B[42]);
  nand g92 (n_266, A[42], B[42]);
  nand g97 (n_272, n_144, n_145);
  nor g98 (n_149, n_146, n_147);
  nor g101 (n_275, n_151, n_147);
  nor g102 (n_155, n_152, n_153);
  nor g105 (n_281, n_157, n_153);
  nor g106 (n_161, n_158, n_159);
  nor g109 (n_283, n_163, n_159);
  nor g110 (n_167, n_164, n_165);
  nor g113 (n_291, n_169, n_165);
  nor g114 (n_173, n_170, n_171);
  nor g117 (n_293, n_175, n_171);
  nor g118 (n_179, n_176, n_177);
  nor g121 (n_301, n_181, n_177);
  nor g122 (n_185, n_182, n_183);
  nor g125 (n_303, n_187, n_183);
  nor g126 (n_191, n_188, n_189);
  nor g129 (n_311, n_193, n_189);
  nor g130 (n_197, n_194, n_195);
  nor g133 (n_313, n_199, n_195);
  nor g134 (n_203, n_200, n_201);
  nor g137 (n_321, n_205, n_201);
  nor g138 (n_209, n_206, n_207);
  nor g141 (n_323, n_211, n_207);
  nor g142 (n_215, n_212, n_213);
  nor g145 (n_331, n_217, n_213);
  nor g146 (n_221, n_218, n_219);
  nor g149 (n_333, n_223, n_219);
  nor g150 (n_227, n_224, n_225);
  nor g153 (n_341, n_229, n_225);
  nor g154 (n_233, n_230, n_231);
  nor g157 (n_343, n_235, n_231);
  nor g158 (n_239, n_236, n_237);
  nor g161 (n_351, n_241, n_237);
  nor g162 (n_245, n_242, n_243);
  nor g165 (n_353, n_247, n_243);
  nor g166 (n_251, n_248, n_249);
  nor g169 (n_361, n_253, n_249);
  nor g170 (n_257, n_254, n_255);
  nor g173 (n_363, n_259, n_255);
  nor g174 (n_263, n_260, n_261);
  nor g177 (n_371, n_265, n_261);
  nor g178 (n_269, n_266, n_267);
  nor g181 (n_373, n_271, n_267);
  nand g184 (n_617, n_146, n_274);
  nand g185 (n_277, n_275, n_272);
  nand g186 (n_378, n_276, n_277);
  nor g187 (n_279, n_163, n_278);
  nand g196 (n_386, n_281, n_283);
  nor g197 (n_289, n_175, n_288);
  nand g206 (n_393, n_291, n_293);
  nor g207 (n_299, n_187, n_298);
  nand g216 (n_401, n_301, n_303);
  nor g217 (n_309, n_199, n_308);
  nand g226 (n_408, n_311, n_313);
  nor g227 (n_319, n_211, n_318);
  nand g236 (n_416, n_321, n_323);
  nor g237 (n_329, n_223, n_328);
  nand g246 (n_423, n_331, n_333);
  nor g247 (n_339, n_235, n_338);
  nand g256 (n_431, n_341, n_343);
  nor g257 (n_349, n_247, n_348);
  nand g266 (n_438, n_351, n_353);
  nor g267 (n_359, n_259, n_358);
  nand g276 (n_446, n_361, n_363);
  nor g277 (n_369, n_271, n_368);
  nand g286 (n_521, n_371, n_373);
  nand g289 (n_621, n_152, n_380);
  nand g290 (n_381, n_281, n_378);
  nand g291 (n_623, n_278, n_381);
  nand g294 (n_626, n_384, n_385);
  nand g297 (n_450, n_388, n_389);
  nor g298 (n_391, n_181, n_390);
  nor g301 (n_460, n_181, n_393);
  nor g307 (n_399, n_397, n_390);
  nor g310 (n_466, n_393, n_397);
  nor g311 (n_403, n_401, n_390);
  nor g314 (n_469, n_393, n_401);
  nor g315 (n_406, n_205, n_405);
  nor g318 (n_536, n_205, n_408);
  nor g324 (n_414, n_412, n_405);
  nor g327 (n_542, n_408, n_412);
  nor g328 (n_418, n_416, n_405);
  nor g331 (n_475, n_408, n_416);
  nor g332 (n_421, n_229, n_420);
  nor g335 (n_488, n_229, n_423);
  nor g341 (n_429, n_427, n_420);
  nor g344 (n_498, n_423, n_427);
  nor g345 (n_433, n_431, n_420);
  nor g348 (n_503, n_423, n_431);
  nor g349 (n_436, n_253, n_435);
  nor g352 (n_588, n_253, n_438);
  nor g358 (n_444, n_442, n_435);
  nor g361 (n_594, n_438, n_442);
  nor g362 (n_448, n_446, n_435);
  nor g365 (n_511, n_438, n_446);
  nand g368 (n_630, n_164, n_452);
  nand g369 (n_453, n_291, n_450);
  nand g370 (n_632, n_288, n_453);
  nand g373 (n_635, n_456, n_457);
  nand g376 (n_638, n_390, n_459);
  nand g377 (n_462, n_460, n_450);
  nand g378 (n_641, n_461, n_462);
  nand g379 (n_465, n_463, n_450);
  nand g380 (n_643, n_464, n_465);
  nand g381 (n_468, n_466, n_450);
  nand g382 (n_646, n_467, n_468);
  nand g383 (n_471, n_469, n_450);
  nand g384 (n_526, n_470, n_471);
  nor g385 (n_473, n_217, n_472);
  nand g394 (n_550, n_331, n_475);
  nor g395 (n_482, n_480, n_472);
  nor g400 (n_485, n_423, n_472);
  nand g409 (n_562, n_475, n_488);
  nand g414 (n_566, n_475, n_493);
  nand g419 (n_570, n_475, n_498);
  nand g424 (n_574, n_475, n_503);
  nor g425 (n_509, n_265, n_508);
  nand g434 (n_602, n_371, n_511);
  nor g435 (n_518, n_516, n_508);
  nor g440 (n_523, n_521, n_508);
  nand g447 (n_650, n_188, n_528);
  nand g448 (n_529, n_311, n_526);
  nand g449 (n_652, n_308, n_529);
  nand g452 (n_655, n_532, n_533);
  nand g455 (n_658, n_405, n_535);
  nand g456 (n_538, n_536, n_526);
  nand g457 (n_661, n_537, n_538);
  nand g458 (n_541, n_539, n_526);
  nand g459 (n_663, n_540, n_541);
  nand g460 (n_544, n_542, n_526);
  nand g461 (n_666, n_543, n_544);
  nand g462 (n_545, n_475, n_526);
  nand g463 (n_668, n_472, n_545);
  nand g466 (n_671, n_548, n_549);
  nand g469 (n_673, n_552, n_553);
  nand g472 (n_676, n_556, n_557);
  nand g475 (n_679, n_560, n_561);
  nand g478 (n_682, n_564, n_565);
  nand g481 (n_684, n_568, n_569);
  nand g484 (n_687, n_572, n_573);
  nand g487 (n_578, n_576, n_577);
  nand g490 (n_691, n_236, n_580);
  nand g491 (n_581, n_351, n_578);
  nand g492 (n_693, n_348, n_581);
  nand g495 (n_696, n_584, n_585);
  nand g498 (n_699, n_435, n_587);
  nand g499 (n_590, n_588, n_578);
  nand g500 (n_702, n_589, n_590);
  nand g501 (n_593, n_591, n_578);
  nand g502 (n_704, n_592, n_593);
  nand g503 (n_596, n_594, n_578);
  nand g504 (n_707, n_595, n_596);
  nand g505 (n_597, n_511, n_578);
  nand g506 (n_709, n_508, n_597);
  nand g509 (n_712, n_600, n_601);
  nand g512 (n_714, n_604, n_605);
  nand g515 (n_717, n_608, n_609);
  nand g518 (n_137, n_612, n_613);
  xnor g522 (Z[2], n_272, n_615);
  xnor g525 (Z[3], n_617, n_618);
  xnor g527 (Z[4], n_378, n_619);
  xnor g530 (Z[5], n_621, n_622);
  xnor g532 (Z[6], n_623, n_624);
  xnor g535 (Z[7], n_626, n_627);
  xnor g537 (Z[8], n_450, n_628);
  xnor g540 (Z[9], n_630, n_631);
  xnor g542 (Z[10], n_632, n_633);
  xnor g545 (Z[11], n_635, n_636);
  xnor g548 (Z[12], n_638, n_639);
  xnor g551 (Z[13], n_641, n_642);
  xnor g553 (Z[14], n_643, n_644);
  xnor g556 (Z[15], n_646, n_647);
  xnor g558 (Z[16], n_526, n_648);
  xnor g561 (Z[17], n_650, n_651);
  xnor g563 (Z[18], n_652, n_653);
  xnor g566 (Z[19], n_655, n_656);
  xnor g569 (Z[20], n_658, n_659);
  xnor g572 (Z[21], n_661, n_662);
  xnor g574 (Z[22], n_663, n_664);
  xnor g577 (Z[23], n_666, n_667);
  xnor g579 (Z[24], n_668, n_669);
  xnor g582 (Z[25], n_671, n_672);
  xnor g584 (Z[26], n_673, n_674);
  xnor g587 (Z[27], n_676, n_677);
  xnor g590 (Z[28], n_679, n_680);
  xnor g593 (Z[29], n_682, n_683);
  xnor g595 (Z[30], n_684, n_685);
  xnor g598 (Z[31], n_687, n_688);
  xnor g600 (Z[32], n_578, n_689);
  xnor g603 (Z[33], n_691, n_692);
  xnor g605 (Z[34], n_693, n_694);
  xnor g608 (Z[35], n_696, n_697);
  xnor g611 (Z[36], n_699, n_700);
  xnor g614 (Z[37], n_702, n_703);
  xnor g616 (Z[38], n_704, n_705);
  xnor g619 (Z[39], n_707, n_708);
  xnor g621 (Z[40], n_709, n_710);
  xnor g624 (Z[41], n_712, n_713);
  xnor g626 (Z[42], n_714, n_715);
  xnor g629 (Z[43], n_717, n_718);
  and g632 (n_267, A[43], B[43]);
  or g633 (n_268, A[43], B[43]);
  and g634 (n_348, wc, n_238);
  not gc (wc, n_239);
  and g635 (n_355, wc0, n_244);
  not gc0 (wc0, n_245);
  and g636 (n_358, wc1, n_250);
  not gc1 (wc1, n_251);
  and g637 (n_365, wc2, n_256);
  not gc2 (wc2, n_257);
  and g638 (n_368, wc3, n_262);
  not gc3 (wc3, n_263);
  and g639 (n_308, wc4, n_190);
  not gc4 (wc4, n_191);
  and g640 (n_315, wc5, n_196);
  not gc5 (wc5, n_197);
  and g641 (n_318, wc6, n_202);
  not gc6 (wc6, n_203);
  and g642 (n_325, wc7, n_208);
  not gc7 (wc7, n_209);
  and g643 (n_328, wc8, n_214);
  not gc8 (wc8, n_215);
  and g644 (n_335, wc9, n_220);
  not gc9 (wc9, n_221);
  and g645 (n_338, wc10, n_226);
  not gc10 (wc10, n_227);
  and g646 (n_345, wc11, n_232);
  not gc11 (wc11, n_233);
  and g647 (n_288, wc12, n_166);
  not gc12 (wc12, n_167);
  and g648 (n_295, wc13, n_172);
  not gc13 (wc13, n_173);
  and g649 (n_298, wc14, n_178);
  not gc14 (wc14, n_179);
  and g650 (n_305, wc15, n_184);
  not gc15 (wc15, n_185);
  and g651 (n_278, wc16, n_154);
  not gc16 (wc16, n_155);
  and g652 (n_285, wc17, n_160);
  not gc17 (wc17, n_161);
  and g653 (n_276, wc18, n_148);
  not gc18 (wc18, n_149);
  or g654 (n_145, n_138, n_141);
  or g655 (n_382, wc19, n_163);
  not gc19 (wc19, n_281);
  or g656 (n_454, wc20, n_175);
  not gc20 (wc20, n_291);
  or g657 (n_397, wc21, n_187);
  not gc21 (wc21, n_301);
  or g658 (n_530, wc22, n_199);
  not gc22 (wc22, n_311);
  or g659 (n_412, wc23, n_211);
  not gc23 (wc23, n_321);
  or g660 (n_480, wc24, n_223);
  not gc24 (wc24, n_331);
  or g661 (n_427, wc25, n_235);
  not gc25 (wc25, n_341);
  or g662 (n_582, wc26, n_247);
  not gc26 (wc26, n_351);
  or g663 (n_442, wc27, n_259);
  not gc27 (wc27, n_361);
  or g664 (n_516, wc28, n_271);
  not gc28 (wc28, n_371);
  or g665 (n_614, wc29, n_141);
  not gc29 (wc29, n_144);
  or g666 (n_615, wc30, n_151);
  not gc30 (wc30, n_146);
  or g667 (n_618, wc31, n_147);
  not gc31 (wc31, n_148);
  or g668 (n_619, wc32, n_157);
  not gc32 (wc32, n_152);
  or g669 (n_622, wc33, n_153);
  not gc33 (wc33, n_154);
  or g670 (n_624, wc34, n_163);
  not gc34 (wc34, n_158);
  or g671 (n_627, wc35, n_159);
  not gc35 (wc35, n_160);
  or g672 (n_628, wc36, n_169);
  not gc36 (wc36, n_164);
  or g673 (n_631, wc37, n_165);
  not gc37 (wc37, n_166);
  or g674 (n_633, wc38, n_175);
  not gc38 (wc38, n_170);
  or g675 (n_636, wc39, n_171);
  not gc39 (wc39, n_172);
  or g676 (n_639, wc40, n_181);
  not gc40 (wc40, n_176);
  or g677 (n_642, wc41, n_177);
  not gc41 (wc41, n_178);
  or g678 (n_644, wc42, n_187);
  not gc42 (wc42, n_182);
  or g679 (n_647, wc43, n_183);
  not gc43 (wc43, n_184);
  or g680 (n_648, wc44, n_193);
  not gc44 (wc44, n_188);
  or g681 (n_651, wc45, n_189);
  not gc45 (wc45, n_190);
  or g682 (n_653, wc46, n_199);
  not gc46 (wc46, n_194);
  or g683 (n_656, wc47, n_195);
  not gc47 (wc47, n_196);
  or g684 (n_659, wc48, n_205);
  not gc48 (wc48, n_200);
  or g685 (n_662, wc49, n_201);
  not gc49 (wc49, n_202);
  or g686 (n_664, wc50, n_211);
  not gc50 (wc50, n_206);
  or g687 (n_667, wc51, n_207);
  not gc51 (wc51, n_208);
  or g688 (n_669, wc52, n_217);
  not gc52 (wc52, n_212);
  or g689 (n_672, wc53, n_213);
  not gc53 (wc53, n_214);
  or g690 (n_674, wc54, n_223);
  not gc54 (wc54, n_218);
  or g691 (n_677, wc55, n_219);
  not gc55 (wc55, n_220);
  or g692 (n_680, wc56, n_229);
  not gc56 (wc56, n_224);
  or g693 (n_683, wc57, n_225);
  not gc57 (wc57, n_226);
  or g694 (n_685, wc58, n_235);
  not gc58 (wc58, n_230);
  or g695 (n_688, wc59, n_231);
  not gc59 (wc59, n_232);
  or g696 (n_689, wc60, n_241);
  not gc60 (wc60, n_236);
  or g697 (n_692, wc61, n_237);
  not gc61 (wc61, n_238);
  or g698 (n_694, wc62, n_247);
  not gc62 (wc62, n_242);
  or g699 (n_697, wc63, n_243);
  not gc63 (wc63, n_244);
  or g700 (n_700, wc64, n_253);
  not gc64 (wc64, n_248);
  or g701 (n_703, wc65, n_249);
  not gc65 (wc65, n_250);
  or g702 (n_705, wc66, n_259);
  not gc66 (wc66, n_254);
  or g703 (n_708, wc67, n_255);
  not gc67 (wc67, n_256);
  or g704 (n_710, wc68, n_265);
  not gc68 (wc68, n_260);
  or g705 (n_713, wc69, n_261);
  not gc69 (wc69, n_262);
  or g706 (n_715, wc70, n_271);
  not gc70 (wc70, n_266);
  and g707 (n_356, wc71, n_353);
  not gc71 (wc71, n_348);
  and g708 (n_366, wc72, n_363);
  not gc72 (wc72, n_358);
  and g709 (n_375, n_268, wc73);
  not gc73 (wc73, n_269);
  and g710 (n_316, wc74, n_313);
  not gc74 (wc74, n_308);
  and g711 (n_326, wc75, n_323);
  not gc75 (wc75, n_318);
  and g712 (n_336, wc76, n_333);
  not gc76 (wc76, n_328);
  and g713 (n_346, wc77, n_343);
  not gc77 (wc77, n_338);
  and g714 (n_296, wc78, n_293);
  not gc78 (wc78, n_288);
  and g715 (n_306, wc79, n_303);
  not gc79 (wc79, n_298);
  and g716 (n_286, wc80, n_283);
  not gc80 (wc80, n_278);
  and g717 (n_463, wc81, n_301);
  not gc81 (wc81, n_393);
  and g718 (n_539, wc82, n_321);
  not gc82 (wc82, n_408);
  and g719 (n_493, wc83, n_341);
  not gc83 (wc83, n_423);
  and g720 (n_591, wc84, n_361);
  not gc84 (wc84, n_438);
  xor g721 (Z[1], n_138, n_614);
  or g722 (n_718, wc85, n_267);
  not gc85 (wc85, n_268);
  and g723 (n_435, wc86, n_355);
  not gc86 (wc86, n_356);
  and g724 (n_447, wc87, n_365);
  not gc87 (wc87, n_366);
  and g725 (n_376, wc88, n_373);
  not gc88 (wc88, n_368);
  and g726 (n_405, wc89, n_315);
  not gc89 (wc89, n_316);
  and g727 (n_417, wc90, n_325);
  not gc90 (wc90, n_326);
  and g728 (n_420, wc91, n_335);
  not gc91 (wc91, n_336);
  and g729 (n_432, wc92, n_345);
  not gc92 (wc92, n_346);
  and g730 (n_390, wc93, n_295);
  not gc93 (wc93, n_296);
  and g731 (n_402, wc94, n_305);
  not gc94 (wc94, n_306);
  and g732 (n_388, wc95, n_285);
  not gc95 (wc95, n_286);
  or g733 (n_274, wc96, n_151);
  not gc96 (wc96, n_272);
  and g734 (n_384, wc97, n_158);
  not gc97 (wc97, n_279);
  and g735 (n_456, wc98, n_170);
  not gc98 (wc98, n_289);
  and g736 (n_398, wc99, n_182);
  not gc99 (wc99, n_299);
  and g737 (n_532, wc100, n_194);
  not gc100 (wc100, n_309);
  and g738 (n_413, wc101, n_206);
  not gc101 (wc101, n_319);
  and g739 (n_481, wc102, n_218);
  not gc102 (wc102, n_329);
  and g740 (n_428, wc103, n_230);
  not gc103 (wc103, n_339);
  and g741 (n_584, wc104, n_242);
  not gc104 (wc104, n_349);
  and g742 (n_443, wc105, n_254);
  not gc105 (wc105, n_359);
  and g743 (n_517, wc106, n_266);
  not gc106 (wc106, n_369);
  or g744 (n_546, wc107, n_217);
  not gc107 (wc107, n_475);
  or g745 (n_554, n_480, wc108);
  not gc108 (wc108, n_475);
  or g746 (n_558, wc109, n_423);
  not gc109 (wc109, n_475);
  or g747 (n_598, wc110, n_265);
  not gc110 (wc110, n_511);
  or g748 (n_606, n_516, wc111);
  not gc111 (wc111, n_511);
  and g749 (n_522, wc112, n_375);
  not gc112 (wc112, n_376);
  or g750 (n_610, wc113, n_521);
  not gc113 (wc113, n_511);
  and g751 (n_395, wc114, n_301);
  not gc114 (wc114, n_390);
  and g752 (n_410, wc115, n_321);
  not gc115 (wc115, n_405);
  and g753 (n_425, wc116, n_341);
  not gc116 (wc116, n_420);
  and g754 (n_440, wc117, n_361);
  not gc117 (wc117, n_435);
  and g755 (n_508, n_447, wc118);
  not gc118 (wc118, n_448);
  and g756 (n_472, n_417, wc119);
  not gc119 (wc119, n_418);
  and g757 (n_505, n_432, wc120);
  not gc120 (wc120, n_433);
  and g758 (n_470, n_402, wc121);
  not gc121 (wc121, n_403);
  or g759 (n_389, n_386, wc122);
  not gc122 (wc122, n_378);
  or g760 (n_380, wc123, n_157);
  not gc123 (wc123, n_378);
  or g761 (n_385, n_382, wc124);
  not gc124 (wc124, n_378);
  and g762 (n_461, wc125, n_176);
  not gc125 (wc125, n_391);
  and g763 (n_464, wc126, n_298);
  not gc126 (wc126, n_395);
  and g764 (n_467, n_398, wc127);
  not gc127 (wc127, n_399);
  and g765 (n_537, wc128, n_200);
  not gc128 (wc128, n_406);
  and g766 (n_540, wc129, n_318);
  not gc129 (wc129, n_410);
  and g767 (n_543, n_413, wc130);
  not gc130 (wc130, n_414);
  and g768 (n_490, wc131, n_224);
  not gc131 (wc131, n_421);
  and g769 (n_495, wc132, n_338);
  not gc132 (wc132, n_425);
  and g770 (n_500, n_428, wc133);
  not gc133 (wc133, n_429);
  and g771 (n_589, wc134, n_248);
  not gc134 (wc134, n_436);
  and g772 (n_592, wc135, n_358);
  not gc135 (wc135, n_440);
  and g773 (n_595, n_443, wc136);
  not gc136 (wc136, n_444);
  and g774 (n_506, wc137, n_503);
  not gc137 (wc137, n_472);
  and g775 (n_478, wc138, n_331);
  not gc138 (wc138, n_472);
  and g776 (n_491, wc139, n_488);
  not gc139 (wc139, n_472);
  and g777 (n_496, wc140, n_493);
  not gc140 (wc140, n_472);
  and g778 (n_501, wc141, n_498);
  not gc141 (wc141, n_472);
  and g779 (n_514, wc142, n_371);
  not gc142 (wc142, n_508);
  and g780 (n_612, n_522, wc143);
  not gc143 (wc143, n_523);
  and g781 (n_576, wc144, n_505);
  not gc144 (wc144, n_506);
  or g782 (n_452, wc145, n_169);
  not gc145 (wc145, n_450);
  or g783 (n_457, n_454, wc146);
  not gc146 (wc146, n_450);
  or g784 (n_459, wc147, n_393);
  not gc147 (wc147, n_450);
  and g785 (n_548, wc148, n_212);
  not gc148 (wc148, n_473);
  and g786 (n_552, wc149, n_328);
  not gc149 (wc149, n_478);
  and g787 (n_556, n_481, wc150);
  not gc150 (wc150, n_482);
  and g788 (n_560, n_420, wc151);
  not gc151 (wc151, n_485);
  and g789 (n_564, wc152, n_490);
  not gc152 (wc152, n_491);
  and g790 (n_568, wc153, n_495);
  not gc153 (wc153, n_496);
  and g791 (n_572, wc154, n_500);
  not gc154 (wc154, n_501);
  and g792 (n_600, wc155, n_260);
  not gc155 (wc155, n_509);
  and g793 (n_604, wc156, n_368);
  not gc156 (wc156, n_514);
  and g794 (n_608, n_517, wc157);
  not gc157 (wc157, n_518);
  or g795 (n_577, n_574, wc158);
  not gc158 (wc158, n_526);
  or g796 (n_528, wc159, n_193);
  not gc159 (wc159, n_526);
  or g797 (n_533, n_530, wc160);
  not gc160 (wc160, n_526);
  or g798 (n_535, wc161, n_408);
  not gc161 (wc161, n_526);
  or g799 (n_549, n_546, wc162);
  not gc162 (wc162, n_526);
  or g800 (n_553, n_550, wc163);
  not gc163 (wc163, n_526);
  or g801 (n_557, n_554, wc164);
  not gc164 (wc164, n_526);
  or g802 (n_561, n_558, wc165);
  not gc165 (wc165, n_526);
  or g803 (n_565, n_562, wc166);
  not gc166 (wc166, n_526);
  or g804 (n_569, n_566, wc167);
  not gc167 (wc167, n_526);
  or g805 (n_573, n_570, wc168);
  not gc168 (wc168, n_526);
  or g806 (n_613, n_610, wc169);
  not gc169 (wc169, n_578);
  or g807 (n_580, wc170, n_241);
  not gc170 (wc170, n_578);
  or g808 (n_585, n_582, wc171);
  not gc171 (wc171, n_578);
  or g809 (n_587, wc172, n_438);
  not gc172 (wc172, n_578);
  or g810 (n_601, n_598, wc173);
  not gc173 (wc173, n_578);
  or g811 (n_605, wc174, n_602);
  not gc174 (wc174, n_578);
  or g812 (n_609, n_606, wc175);
  not gc175 (wc175, n_578);
endmodule

module add_signed_398_GENERIC(A, B, Z);
  input [43:0] A, B;
  output [44:0] Z;
  wire [43:0] A, B;
  wire [44:0] Z;
  add_signed_398_GENERIC_REAL g1(.A ({A[42], A[42:0]}), .B ({B[42],
       B[42:0]}), .Z (Z));
endmodule

module add_signed_412_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [42:0] A, B;
  output [43:0] Z;
  wire [42:0] A, B;
  wire [43:0] Z;
  wire n_134, n_135, n_138, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_148, n_149, n_150, n_151, n_152, n_154, n_155;
  wire n_156, n_157, n_158, n_160, n_161, n_162, n_163, n_164;
  wire n_166, n_167, n_168, n_169, n_170, n_172, n_173, n_174;
  wire n_175, n_176, n_178, n_179, n_180, n_181, n_182, n_184;
  wire n_185, n_186, n_187, n_188, n_190, n_191, n_192, n_193;
  wire n_194, n_196, n_197, n_198, n_199, n_200, n_202, n_203;
  wire n_204, n_205, n_206, n_208, n_209, n_210, n_211, n_212;
  wire n_214, n_215, n_216, n_217, n_218, n_220, n_221, n_222;
  wire n_223, n_224, n_226, n_227, n_228, n_229, n_230, n_232;
  wire n_233, n_234, n_235, n_236, n_238, n_239, n_240, n_241;
  wire n_242, n_244, n_245, n_246, n_247, n_248, n_250, n_251;
  wire n_252, n_253, n_254, n_256, n_257, n_258, n_259, n_260;
  wire n_262, n_263, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_272, n_274, n_276, n_277, n_279, n_280, n_282, n_284;
  wire n_286, n_287, n_289, n_290, n_292, n_294, n_296, n_297;
  wire n_299, n_300, n_302, n_304, n_306, n_307, n_309, n_310;
  wire n_312, n_314, n_316, n_317, n_319, n_320, n_322, n_324;
  wire n_326, n_327, n_329, n_330, n_332, n_334, n_336, n_337;
  wire n_339, n_340, n_342, n_344, n_346, n_347, n_349, n_350;
  wire n_352, n_354, n_356, n_357, n_359, n_360, n_361, n_362;
  wire n_364, n_366, n_368, n_369, n_370, n_372, n_373, n_374;
  wire n_376, n_377, n_378, n_379, n_381, n_383, n_385, n_386;
  wire n_387, n_389, n_390, n_391, n_393, n_394, n_396, n_398;
  wire n_400, n_401, n_402, n_404, n_405, n_406, n_408, n_409;
  wire n_411, n_413, n_415, n_416, n_417, n_419, n_420, n_421;
  wire n_423, n_424, n_426, n_428, n_430, n_431, n_432, n_434;
  wire n_435, n_436, n_438, n_440, n_441, n_442, n_444, n_445;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_463;
  wire n_466, n_468, n_469, n_470, n_473, n_476, n_478, n_479;
  wire n_481, n_483, n_484, n_486, n_488, n_489, n_491, n_493;
  wire n_494, n_496, n_497, n_499, n_502, n_504, n_505, n_506;
  wire n_509, n_511, n_512, n_513, n_515, n_516, n_518, n_519;
  wire n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_531, n_532, n_533, n_535, n_536, n_537;
  wire n_539, n_540, n_541, n_543, n_544, n_545, n_547, n_548;
  wire n_549, n_551, n_552, n_553, n_555, n_556, n_557, n_559;
  wire n_560, n_561, n_563, n_564, n_565, n_567, n_568, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578;
  wire n_579, n_580, n_581, n_583, n_584, n_585, n_587, n_588;
  wire n_589, n_591, n_592, n_593, n_594, n_596, n_597, n_598;
  wire n_600, n_601, n_602, n_603, n_605, n_606, n_607, n_609;
  wire n_610, n_611, n_612, n_614, n_615, n_617, n_618, n_620;
  wire n_621, n_622, n_623, n_625, n_626, n_627, n_629, n_630;
  wire n_631, n_632, n_634, n_635, n_637, n_638, n_640, n_641;
  wire n_642, n_643, n_645, n_646, n_647, n_648, n_650, n_651;
  wire n_652, n_653, n_655, n_656, n_658, n_659, n_661, n_662;
  wire n_663, n_664, n_666, n_667, n_668, n_670, n_671, n_672;
  wire n_673, n_675, n_676, n_678, n_679, n_681, n_682, n_683;
  wire n_684, n_686, n_687, n_688, n_689, n_691, n_692, n_693;
  wire n_694;
  not g3 (Z[43], n_134);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_135, A[0], B[0]);
  nor g9 (n_138, A[1], B[1]);
  nand g10 (n_141, A[1], B[1]);
  nor g11 (n_148, A[2], B[2]);
  nand g12 (n_143, A[2], B[2]);
  nor g13 (n_144, A[3], B[3]);
  nand g14 (n_145, A[3], B[3]);
  nor g15 (n_154, A[4], B[4]);
  nand g16 (n_149, A[4], B[4]);
  nor g17 (n_150, A[5], B[5]);
  nand g18 (n_151, A[5], B[5]);
  nor g19 (n_160, A[6], B[6]);
  nand g20 (n_155, A[6], B[6]);
  nor g21 (n_156, A[7], B[7]);
  nand g22 (n_157, A[7], B[7]);
  nor g23 (n_166, A[8], B[8]);
  nand g24 (n_161, A[8], B[8]);
  nor g25 (n_162, A[9], B[9]);
  nand g26 (n_163, A[9], B[9]);
  nor g27 (n_172, A[10], B[10]);
  nand g28 (n_167, A[10], B[10]);
  nor g29 (n_168, A[11], B[11]);
  nand g30 (n_169, A[11], B[11]);
  nor g31 (n_178, A[12], B[12]);
  nand g32 (n_173, A[12], B[12]);
  nor g33 (n_174, A[13], B[13]);
  nand g34 (n_175, A[13], B[13]);
  nor g35 (n_184, A[14], B[14]);
  nand g36 (n_179, A[14], B[14]);
  nor g37 (n_180, A[15], B[15]);
  nand g38 (n_181, A[15], B[15]);
  nor g39 (n_190, A[16], B[16]);
  nand g40 (n_185, A[16], B[16]);
  nor g41 (n_186, A[17], B[17]);
  nand g42 (n_187, A[17], B[17]);
  nor g43 (n_196, A[18], B[18]);
  nand g44 (n_191, A[18], B[18]);
  nor g45 (n_192, A[19], B[19]);
  nand g46 (n_193, A[19], B[19]);
  nor g47 (n_202, A[20], B[20]);
  nand g48 (n_197, A[20], B[20]);
  nor g49 (n_198, A[21], B[21]);
  nand g50 (n_199, A[21], B[21]);
  nor g51 (n_208, A[22], B[22]);
  nand g52 (n_203, A[22], B[22]);
  nor g53 (n_204, A[23], B[23]);
  nand g54 (n_205, A[23], B[23]);
  nor g55 (n_214, A[24], B[24]);
  nand g56 (n_209, A[24], B[24]);
  nor g57 (n_210, A[25], B[25]);
  nand g58 (n_211, A[25], B[25]);
  nor g59 (n_220, A[26], B[26]);
  nand g60 (n_215, A[26], B[26]);
  nor g61 (n_216, A[27], B[27]);
  nand g62 (n_217, A[27], B[27]);
  nor g63 (n_226, A[28], B[28]);
  nand g64 (n_221, A[28], B[28]);
  nor g65 (n_222, A[29], B[29]);
  nand g66 (n_223, A[29], B[29]);
  nor g67 (n_232, A[30], B[30]);
  nand g68 (n_227, A[30], B[30]);
  nor g69 (n_228, A[31], B[31]);
  nand g70 (n_229, A[31], B[31]);
  nor g71 (n_238, A[32], B[32]);
  nand g72 (n_233, A[32], B[32]);
  nor g73 (n_234, A[33], B[33]);
  nand g74 (n_235, A[33], B[33]);
  nor g75 (n_244, A[34], B[34]);
  nand g76 (n_239, A[34], B[34]);
  nor g77 (n_240, A[35], B[35]);
  nand g78 (n_241, A[35], B[35]);
  nor g79 (n_250, A[36], B[36]);
  nand g80 (n_245, A[36], B[36]);
  nor g81 (n_246, A[37], B[37]);
  nand g82 (n_247, A[37], B[37]);
  nor g83 (n_256, A[38], B[38]);
  nand g84 (n_251, A[38], B[38]);
  nor g85 (n_252, A[39], B[39]);
  nand g86 (n_253, A[39], B[39]);
  nor g87 (n_262, A[40], B[40]);
  nand g88 (n_257, A[40], B[40]);
  nor g89 (n_258, A[41], B[41]);
  nand g90 (n_259, A[41], B[41]);
  nand g95 (n_263, n_141, n_142);
  nor g96 (n_146, n_143, n_144);
  nor g99 (n_266, n_148, n_144);
  nor g100 (n_152, n_149, n_150);
  nor g103 (n_272, n_154, n_150);
  nor g104 (n_158, n_155, n_156);
  nor g107 (n_274, n_160, n_156);
  nor g108 (n_164, n_161, n_162);
  nor g111 (n_282, n_166, n_162);
  nor g112 (n_170, n_167, n_168);
  nor g115 (n_284, n_172, n_168);
  nor g116 (n_176, n_173, n_174);
  nor g119 (n_292, n_178, n_174);
  nor g120 (n_182, n_179, n_180);
  nor g123 (n_294, n_184, n_180);
  nor g124 (n_188, n_185, n_186);
  nor g127 (n_302, n_190, n_186);
  nor g128 (n_194, n_191, n_192);
  nor g131 (n_304, n_196, n_192);
  nor g132 (n_200, n_197, n_198);
  nor g135 (n_312, n_202, n_198);
  nor g136 (n_206, n_203, n_204);
  nor g139 (n_314, n_208, n_204);
  nor g140 (n_212, n_209, n_210);
  nor g143 (n_322, n_214, n_210);
  nor g144 (n_218, n_215, n_216);
  nor g147 (n_324, n_220, n_216);
  nor g148 (n_224, n_221, n_222);
  nor g151 (n_332, n_226, n_222);
  nor g152 (n_230, n_227, n_228);
  nor g155 (n_334, n_232, n_228);
  nor g156 (n_236, n_233, n_234);
  nor g159 (n_342, n_238, n_234);
  nor g160 (n_242, n_239, n_240);
  nor g163 (n_344, n_244, n_240);
  nor g164 (n_248, n_245, n_246);
  nor g167 (n_352, n_250, n_246);
  nor g168 (n_254, n_251, n_252);
  nor g171 (n_354, n_256, n_252);
  nor g172 (n_260, n_257, n_258);
  nor g175 (n_364, n_262, n_258);
  nand g178 (n_596, n_143, n_265);
  nand g179 (n_268, n_266, n_263);
  nand g180 (n_366, n_267, n_268);
  nor g181 (n_270, n_160, n_269);
  nand g190 (n_374, n_272, n_274);
  nor g191 (n_280, n_172, n_279);
  nand g200 (n_381, n_282, n_284);
  nor g201 (n_290, n_184, n_289);
  nand g210 (n_389, n_292, n_294);
  nor g211 (n_300, n_196, n_299);
  nand g220 (n_396, n_302, n_304);
  nor g221 (n_310, n_208, n_309);
  nand g230 (n_404, n_312, n_314);
  nor g231 (n_320, n_220, n_319);
  nand g240 (n_411, n_322, n_324);
  nor g241 (n_330, n_232, n_329);
  nand g250 (n_419, n_332, n_334);
  nor g251 (n_340, n_244, n_339);
  nand g260 (n_426, n_342, n_344);
  nor g261 (n_350, n_256, n_349);
  nand g270 (n_434, n_352, n_354);
  nor g271 (n_362, n_359, n_360);
  nand g278 (n_600, n_149, n_368);
  nand g279 (n_369, n_272, n_366);
  nand g280 (n_602, n_269, n_369);
  nand g283 (n_605, n_372, n_373);
  nand g286 (n_438, n_376, n_377);
  nor g287 (n_379, n_178, n_378);
  nor g290 (n_448, n_178, n_381);
  nor g296 (n_387, n_385, n_378);
  nor g299 (n_454, n_381, n_385);
  nor g300 (n_391, n_389, n_378);
  nor g303 (n_457, n_381, n_389);
  nor g304 (n_394, n_202, n_393);
  nor g307 (n_519, n_202, n_396);
  nor g313 (n_402, n_400, n_393);
  nor g316 (n_525, n_396, n_400);
  nor g317 (n_406, n_404, n_393);
  nor g320 (n_463, n_396, n_404);
  nor g321 (n_409, n_226, n_408);
  nor g324 (n_476, n_226, n_411);
  nor g330 (n_417, n_415, n_408);
  nor g333 (n_486, n_411, n_415);
  nor g334 (n_421, n_419, n_408);
  nor g337 (n_491, n_411, n_419);
  nor g338 (n_424, n_250, n_423);
  nor g341 (n_571, n_250, n_426);
  nor g347 (n_432, n_430, n_423);
  nor g350 (n_577, n_426, n_430);
  nor g351 (n_436, n_434, n_423);
  nor g354 (n_499, n_426, n_434);
  nand g357 (n_609, n_161, n_440);
  nand g358 (n_441, n_282, n_438);
  nand g359 (n_611, n_279, n_441);
  nand g362 (n_614, n_444, n_445);
  nand g365 (n_617, n_378, n_447);
  nand g366 (n_450, n_448, n_438);
  nand g367 (n_620, n_449, n_450);
  nand g368 (n_453, n_451, n_438);
  nand g369 (n_622, n_452, n_453);
  nand g370 (n_456, n_454, n_438);
  nand g371 (n_625, n_455, n_456);
  nand g372 (n_459, n_457, n_438);
  nand g373 (n_509, n_458, n_459);
  nor g374 (n_461, n_214, n_460);
  nand g383 (n_533, n_322, n_463);
  nor g384 (n_470, n_468, n_460);
  nor g389 (n_473, n_411, n_460);
  nand g398 (n_545, n_463, n_476);
  nand g403 (n_549, n_463, n_481);
  nand g408 (n_553, n_463, n_486);
  nand g413 (n_557, n_463, n_491);
  nor g414 (n_497, n_262, n_496);
  nand g423 (n_585, n_364, n_499);
  nor g424 (n_506, n_504, n_496);
  nand g431 (n_629, n_185, n_511);
  nand g432 (n_512, n_302, n_509);
  nand g433 (n_631, n_299, n_512);
  nand g436 (n_634, n_515, n_516);
  nand g439 (n_637, n_393, n_518);
  nand g440 (n_521, n_519, n_509);
  nand g441 (n_640, n_520, n_521);
  nand g442 (n_524, n_522, n_509);
  nand g443 (n_642, n_523, n_524);
  nand g444 (n_527, n_525, n_509);
  nand g445 (n_645, n_526, n_527);
  nand g446 (n_528, n_463, n_509);
  nand g447 (n_647, n_460, n_528);
  nand g450 (n_650, n_531, n_532);
  nand g453 (n_652, n_535, n_536);
  nand g456 (n_655, n_539, n_540);
  nand g459 (n_658, n_543, n_544);
  nand g462 (n_661, n_547, n_548);
  nand g465 (n_663, n_551, n_552);
  nand g468 (n_666, n_555, n_556);
  nand g471 (n_561, n_559, n_560);
  nand g474 (n_670, n_233, n_563);
  nand g475 (n_564, n_342, n_561);
  nand g476 (n_672, n_339, n_564);
  nand g479 (n_675, n_567, n_568);
  nand g482 (n_678, n_423, n_570);
  nand g483 (n_573, n_571, n_561);
  nand g484 (n_681, n_572, n_573);
  nand g485 (n_576, n_574, n_561);
  nand g486 (n_683, n_575, n_576);
  nand g487 (n_579, n_577, n_561);
  nand g488 (n_686, n_578, n_579);
  nand g489 (n_580, n_499, n_561);
  nand g490 (n_688, n_496, n_580);
  nand g493 (n_691, n_583, n_584);
  nand g496 (n_693, n_587, n_588);
  nand g499 (n_134, n_591, n_592);
  xnor g503 (Z[2], n_263, n_594);
  xnor g506 (Z[3], n_596, n_597);
  xnor g508 (Z[4], n_366, n_598);
  xnor g511 (Z[5], n_600, n_601);
  xnor g513 (Z[6], n_602, n_603);
  xnor g516 (Z[7], n_605, n_606);
  xnor g518 (Z[8], n_438, n_607);
  xnor g521 (Z[9], n_609, n_610);
  xnor g523 (Z[10], n_611, n_612);
  xnor g526 (Z[11], n_614, n_615);
  xnor g529 (Z[12], n_617, n_618);
  xnor g532 (Z[13], n_620, n_621);
  xnor g534 (Z[14], n_622, n_623);
  xnor g537 (Z[15], n_625, n_626);
  xnor g539 (Z[16], n_509, n_627);
  xnor g542 (Z[17], n_629, n_630);
  xnor g544 (Z[18], n_631, n_632);
  xnor g547 (Z[19], n_634, n_635);
  xnor g550 (Z[20], n_637, n_638);
  xnor g553 (Z[21], n_640, n_641);
  xnor g555 (Z[22], n_642, n_643);
  xnor g558 (Z[23], n_645, n_646);
  xnor g560 (Z[24], n_647, n_648);
  xnor g563 (Z[25], n_650, n_651);
  xnor g565 (Z[26], n_652, n_653);
  xnor g568 (Z[27], n_655, n_656);
  xnor g571 (Z[28], n_658, n_659);
  xnor g574 (Z[29], n_661, n_662);
  xnor g576 (Z[30], n_663, n_664);
  xnor g579 (Z[31], n_666, n_667);
  xnor g581 (Z[32], n_561, n_668);
  xnor g584 (Z[33], n_670, n_671);
  xnor g586 (Z[34], n_672, n_673);
  xnor g589 (Z[35], n_675, n_676);
  xnor g592 (Z[36], n_678, n_679);
  xnor g595 (Z[37], n_681, n_682);
  xnor g597 (Z[38], n_683, n_684);
  xnor g600 (Z[39], n_686, n_687);
  xnor g602 (Z[40], n_688, n_689);
  xnor g605 (Z[41], n_691, n_692);
  xnor g607 (Z[42], n_693, n_694);
  and g610 (n_359, A[42], B[42]);
  or g611 (n_361, A[42], B[42]);
  and g612 (n_339, wc, n_235);
  not gc (wc, n_236);
  and g613 (n_346, wc0, n_241);
  not gc0 (wc0, n_242);
  and g614 (n_349, wc1, n_247);
  not gc1 (wc1, n_248);
  and g615 (n_356, wc2, n_253);
  not gc2 (wc2, n_254);
  and g616 (n_360, wc3, n_259);
  not gc3 (wc3, n_260);
  and g617 (n_299, wc4, n_187);
  not gc4 (wc4, n_188);
  and g618 (n_306, wc5, n_193);
  not gc5 (wc5, n_194);
  and g619 (n_309, wc6, n_199);
  not gc6 (wc6, n_200);
  and g620 (n_316, wc7, n_205);
  not gc7 (wc7, n_206);
  and g621 (n_319, wc8, n_211);
  not gc8 (wc8, n_212);
  and g622 (n_326, wc9, n_217);
  not gc9 (wc9, n_218);
  and g623 (n_329, wc10, n_223);
  not gc10 (wc10, n_224);
  and g624 (n_336, wc11, n_229);
  not gc11 (wc11, n_230);
  and g625 (n_279, wc12, n_163);
  not gc12 (wc12, n_164);
  and g626 (n_286, wc13, n_169);
  not gc13 (wc13, n_170);
  and g627 (n_289, wc14, n_175);
  not gc14 (wc14, n_176);
  and g628 (n_296, wc15, n_181);
  not gc15 (wc15, n_182);
  and g629 (n_269, wc16, n_151);
  not gc16 (wc16, n_152);
  and g630 (n_276, wc17, n_157);
  not gc17 (wc17, n_158);
  and g631 (n_267, wc18, n_145);
  not gc18 (wc18, n_146);
  or g632 (n_142, n_135, n_138);
  or g633 (n_370, wc19, n_160);
  not gc19 (wc19, n_272);
  or g634 (n_442, wc20, n_172);
  not gc20 (wc20, n_282);
  or g635 (n_385, wc21, n_184);
  not gc21 (wc21, n_292);
  or g636 (n_513, wc22, n_196);
  not gc22 (wc22, n_302);
  or g637 (n_400, wc23, n_208);
  not gc23 (wc23, n_312);
  or g638 (n_468, wc24, n_220);
  not gc24 (wc24, n_322);
  or g639 (n_415, wc25, n_232);
  not gc25 (wc25, n_332);
  or g640 (n_565, wc26, n_244);
  not gc26 (wc26, n_342);
  or g641 (n_430, wc27, n_256);
  not gc27 (wc27, n_352);
  or g642 (n_593, wc28, n_138);
  not gc28 (wc28, n_141);
  or g643 (n_594, wc29, n_148);
  not gc29 (wc29, n_143);
  or g644 (n_597, wc30, n_144);
  not gc30 (wc30, n_145);
  or g645 (n_598, wc31, n_154);
  not gc31 (wc31, n_149);
  or g646 (n_601, wc32, n_150);
  not gc32 (wc32, n_151);
  or g647 (n_603, wc33, n_160);
  not gc33 (wc33, n_155);
  or g648 (n_606, wc34, n_156);
  not gc34 (wc34, n_157);
  or g649 (n_607, wc35, n_166);
  not gc35 (wc35, n_161);
  or g650 (n_610, wc36, n_162);
  not gc36 (wc36, n_163);
  or g651 (n_612, wc37, n_172);
  not gc37 (wc37, n_167);
  or g652 (n_615, wc38, n_168);
  not gc38 (wc38, n_169);
  or g653 (n_618, wc39, n_178);
  not gc39 (wc39, n_173);
  or g654 (n_621, wc40, n_174);
  not gc40 (wc40, n_175);
  or g655 (n_623, wc41, n_184);
  not gc41 (wc41, n_179);
  or g656 (n_626, wc42, n_180);
  not gc42 (wc42, n_181);
  or g657 (n_627, wc43, n_190);
  not gc43 (wc43, n_185);
  or g658 (n_630, wc44, n_186);
  not gc44 (wc44, n_187);
  or g659 (n_632, wc45, n_196);
  not gc45 (wc45, n_191);
  or g660 (n_635, wc46, n_192);
  not gc46 (wc46, n_193);
  or g661 (n_638, wc47, n_202);
  not gc47 (wc47, n_197);
  or g662 (n_641, wc48, n_198);
  not gc48 (wc48, n_199);
  or g663 (n_643, wc49, n_208);
  not gc49 (wc49, n_203);
  or g664 (n_646, wc50, n_204);
  not gc50 (wc50, n_205);
  or g665 (n_648, wc51, n_214);
  not gc51 (wc51, n_209);
  or g666 (n_651, wc52, n_210);
  not gc52 (wc52, n_211);
  or g667 (n_653, wc53, n_220);
  not gc53 (wc53, n_215);
  or g668 (n_656, wc54, n_216);
  not gc54 (wc54, n_217);
  or g669 (n_659, wc55, n_226);
  not gc55 (wc55, n_221);
  or g670 (n_662, wc56, n_222);
  not gc56 (wc56, n_223);
  or g671 (n_664, wc57, n_232);
  not gc57 (wc57, n_227);
  or g672 (n_667, wc58, n_228);
  not gc58 (wc58, n_229);
  or g673 (n_668, wc59, n_238);
  not gc59 (wc59, n_233);
  or g674 (n_671, wc60, n_234);
  not gc60 (wc60, n_235);
  or g675 (n_673, wc61, n_244);
  not gc61 (wc61, n_239);
  or g676 (n_676, wc62, n_240);
  not gc62 (wc62, n_241);
  or g677 (n_679, wc63, n_250);
  not gc63 (wc63, n_245);
  or g678 (n_682, wc64, n_246);
  not gc64 (wc64, n_247);
  or g679 (n_684, wc65, n_256);
  not gc65 (wc65, n_251);
  or g680 (n_687, wc66, n_252);
  not gc66 (wc66, n_253);
  or g681 (n_689, wc67, n_262);
  not gc67 (wc67, n_257);
  or g682 (n_692, wc68, n_258);
  not gc68 (wc68, n_259);
  or g683 (n_504, n_359, wc69);
  not gc69 (wc69, n_364);
  and g684 (n_347, wc70, n_344);
  not gc70 (wc70, n_339);
  and g685 (n_357, wc71, n_354);
  not gc71 (wc71, n_349);
  and g686 (n_307, wc72, n_304);
  not gc72 (wc72, n_299);
  and g687 (n_317, wc73, n_314);
  not gc73 (wc73, n_309);
  and g688 (n_327, wc74, n_324);
  not gc74 (wc74, n_319);
  and g689 (n_337, wc75, n_334);
  not gc75 (wc75, n_329);
  and g690 (n_287, wc76, n_284);
  not gc76 (wc76, n_279);
  and g691 (n_297, wc77, n_294);
  not gc77 (wc77, n_289);
  and g692 (n_277, wc78, n_274);
  not gc78 (wc78, n_269);
  and g693 (n_451, wc79, n_292);
  not gc79 (wc79, n_381);
  and g694 (n_522, wc80, n_312);
  not gc80 (wc80, n_396);
  and g695 (n_481, wc81, n_332);
  not gc81 (wc81, n_411);
  and g696 (n_574, wc82, n_352);
  not gc82 (wc82, n_426);
  xor g697 (Z[1], n_135, n_593);
  or g698 (n_694, wc83, n_359);
  not gc83 (wc83, n_361);
  and g699 (n_423, wc84, n_346);
  not gc84 (wc84, n_347);
  and g700 (n_435, wc85, n_356);
  not gc85 (wc85, n_357);
  and g701 (n_505, n_361, wc86);
  not gc86 (wc86, n_362);
  and g702 (n_393, wc87, n_306);
  not gc87 (wc87, n_307);
  and g703 (n_405, wc88, n_316);
  not gc88 (wc88, n_317);
  and g704 (n_408, wc89, n_326);
  not gc89 (wc89, n_327);
  and g705 (n_420, wc90, n_336);
  not gc90 (wc90, n_337);
  and g706 (n_378, wc91, n_286);
  not gc91 (wc91, n_287);
  and g707 (n_390, wc92, n_296);
  not gc92 (wc92, n_297);
  and g708 (n_376, wc93, n_276);
  not gc93 (wc93, n_277);
  or g709 (n_265, wc94, n_148);
  not gc94 (wc94, n_263);
  and g710 (n_372, wc95, n_155);
  not gc95 (wc95, n_270);
  and g711 (n_444, wc96, n_167);
  not gc96 (wc96, n_280);
  and g712 (n_386, wc97, n_179);
  not gc97 (wc97, n_290);
  and g713 (n_515, wc98, n_191);
  not gc98 (wc98, n_300);
  and g714 (n_401, wc99, n_203);
  not gc99 (wc99, n_310);
  and g715 (n_469, wc100, n_215);
  not gc100 (wc100, n_320);
  and g716 (n_416, wc101, n_227);
  not gc101 (wc101, n_330);
  and g717 (n_567, wc102, n_239);
  not gc102 (wc102, n_340);
  and g718 (n_431, wc103, n_251);
  not gc103 (wc103, n_350);
  or g719 (n_529, wc104, n_214);
  not gc104 (wc104, n_463);
  or g720 (n_537, n_468, wc105);
  not gc105 (wc105, n_463);
  or g721 (n_541, wc106, n_411);
  not gc106 (wc106, n_463);
  or g722 (n_581, wc107, n_262);
  not gc107 (wc107, n_499);
  or g723 (n_589, n_504, wc108);
  not gc108 (wc108, n_499);
  and g724 (n_383, wc109, n_292);
  not gc109 (wc109, n_378);
  and g725 (n_398, wc110, n_312);
  not gc110 (wc110, n_393);
  and g726 (n_413, wc111, n_332);
  not gc111 (wc111, n_408);
  and g727 (n_428, wc112, n_352);
  not gc112 (wc112, n_423);
  and g728 (n_496, n_435, wc113);
  not gc113 (wc113, n_436);
  and g729 (n_460, n_405, wc114);
  not gc114 (wc114, n_406);
  and g730 (n_493, n_420, wc115);
  not gc115 (wc115, n_421);
  and g731 (n_458, n_390, wc116);
  not gc116 (wc116, n_391);
  or g732 (n_377, n_374, wc117);
  not gc117 (wc117, n_366);
  or g733 (n_368, wc118, n_154);
  not gc118 (wc118, n_366);
  or g734 (n_373, n_370, wc119);
  not gc119 (wc119, n_366);
  and g735 (n_449, wc120, n_173);
  not gc120 (wc120, n_379);
  and g736 (n_452, wc121, n_289);
  not gc121 (wc121, n_383);
  and g737 (n_455, n_386, wc122);
  not gc122 (wc122, n_387);
  and g738 (n_520, wc123, n_197);
  not gc123 (wc123, n_394);
  and g739 (n_523, wc124, n_309);
  not gc124 (wc124, n_398);
  and g740 (n_526, n_401, wc125);
  not gc125 (wc125, n_402);
  and g741 (n_478, wc126, n_221);
  not gc126 (wc126, n_409);
  and g742 (n_483, wc127, n_329);
  not gc127 (wc127, n_413);
  and g743 (n_488, n_416, wc128);
  not gc128 (wc128, n_417);
  and g744 (n_572, wc129, n_245);
  not gc129 (wc129, n_424);
  and g745 (n_575, wc130, n_349);
  not gc130 (wc130, n_428);
  and g746 (n_578, n_431, wc131);
  not gc131 (wc131, n_432);
  and g747 (n_494, wc132, n_491);
  not gc132 (wc132, n_460);
  and g748 (n_466, wc133, n_322);
  not gc133 (wc133, n_460);
  and g749 (n_479, wc134, n_476);
  not gc134 (wc134, n_460);
  and g750 (n_484, wc135, n_481);
  not gc135 (wc135, n_460);
  and g751 (n_489, wc136, n_486);
  not gc136 (wc136, n_460);
  and g752 (n_502, wc137, n_364);
  not gc137 (wc137, n_496);
  and g753 (n_591, n_505, wc138);
  not gc138 (wc138, n_506);
  and g754 (n_559, wc139, n_493);
  not gc139 (wc139, n_494);
  or g755 (n_440, wc140, n_166);
  not gc140 (wc140, n_438);
  or g756 (n_445, n_442, wc141);
  not gc141 (wc141, n_438);
  or g757 (n_447, wc142, n_381);
  not gc142 (wc142, n_438);
  and g758 (n_531, wc143, n_209);
  not gc143 (wc143, n_461);
  and g759 (n_535, wc144, n_319);
  not gc144 (wc144, n_466);
  and g760 (n_539, n_469, wc145);
  not gc145 (wc145, n_470);
  and g761 (n_543, n_408, wc146);
  not gc146 (wc146, n_473);
  and g762 (n_547, wc147, n_478);
  not gc147 (wc147, n_479);
  and g763 (n_551, wc148, n_483);
  not gc148 (wc148, n_484);
  and g764 (n_555, wc149, n_488);
  not gc149 (wc149, n_489);
  and g765 (n_583, wc150, n_257);
  not gc150 (wc150, n_497);
  and g766 (n_587, wc151, n_360);
  not gc151 (wc151, n_502);
  or g767 (n_560, n_557, wc152);
  not gc152 (wc152, n_509);
  or g768 (n_511, wc153, n_190);
  not gc153 (wc153, n_509);
  or g769 (n_516, n_513, wc154);
  not gc154 (wc154, n_509);
  or g770 (n_518, wc155, n_396);
  not gc155 (wc155, n_509);
  or g771 (n_532, n_529, wc156);
  not gc156 (wc156, n_509);
  or g772 (n_536, n_533, wc157);
  not gc157 (wc157, n_509);
  or g773 (n_540, n_537, wc158);
  not gc158 (wc158, n_509);
  or g774 (n_544, n_541, wc159);
  not gc159 (wc159, n_509);
  or g775 (n_548, n_545, wc160);
  not gc160 (wc160, n_509);
  or g776 (n_552, n_549, wc161);
  not gc161 (wc161, n_509);
  or g777 (n_556, n_553, wc162);
  not gc162 (wc162, n_509);
  or g778 (n_592, n_589, wc163);
  not gc163 (wc163, n_561);
  or g779 (n_563, wc164, n_238);
  not gc164 (wc164, n_561);
  or g780 (n_568, n_565, wc165);
  not gc165 (wc165, n_561);
  or g781 (n_570, wc166, n_426);
  not gc166 (wc166, n_561);
  or g782 (n_584, n_581, wc167);
  not gc167 (wc167, n_561);
  or g783 (n_588, wc168, n_585);
  not gc168 (wc168, n_561);
endmodule

module add_signed_412_GENERIC(A, B, Z);
  input [42:0] A, B;
  output [43:0] Z;
  wire [42:0] A, B;
  wire [43:0] Z;
  add_signed_412_GENERIC_REAL g1(.A ({A[41], A[41:0]}), .B ({B[41],
       B[41:0]}), .Z (Z));
endmodule

module add_signed_412_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [42:0] A, B;
  output [43:0] Z;
  wire [42:0] A, B;
  wire [43:0] Z;
  wire n_134, n_135, n_138, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_148, n_149, n_150, n_151, n_152, n_154, n_155;
  wire n_156, n_157, n_158, n_160, n_161, n_162, n_163, n_164;
  wire n_166, n_167, n_168, n_169, n_170, n_172, n_173, n_174;
  wire n_175, n_176, n_178, n_179, n_180, n_181, n_182, n_184;
  wire n_185, n_186, n_187, n_188, n_190, n_191, n_192, n_193;
  wire n_194, n_196, n_197, n_198, n_199, n_200, n_202, n_203;
  wire n_204, n_205, n_206, n_208, n_209, n_210, n_211, n_212;
  wire n_214, n_215, n_216, n_217, n_218, n_220, n_221, n_222;
  wire n_223, n_224, n_226, n_227, n_228, n_229, n_230, n_232;
  wire n_233, n_234, n_235, n_236, n_238, n_239, n_240, n_241;
  wire n_242, n_244, n_245, n_246, n_247, n_248, n_250, n_251;
  wire n_252, n_253, n_254, n_256, n_257, n_258, n_259, n_260;
  wire n_262, n_263, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_272, n_274, n_276, n_277, n_279, n_280, n_282, n_284;
  wire n_286, n_287, n_289, n_290, n_292, n_294, n_296, n_297;
  wire n_299, n_300, n_302, n_304, n_306, n_307, n_309, n_310;
  wire n_312, n_314, n_316, n_317, n_319, n_320, n_322, n_324;
  wire n_326, n_327, n_329, n_330, n_332, n_334, n_336, n_337;
  wire n_339, n_340, n_342, n_344, n_346, n_347, n_349, n_350;
  wire n_352, n_354, n_356, n_357, n_359, n_360, n_361, n_362;
  wire n_364, n_366, n_368, n_369, n_370, n_372, n_373, n_374;
  wire n_376, n_377, n_378, n_379, n_381, n_383, n_385, n_386;
  wire n_387, n_389, n_390, n_391, n_393, n_394, n_396, n_398;
  wire n_400, n_401, n_402, n_404, n_405, n_406, n_408, n_409;
  wire n_411, n_413, n_415, n_416, n_417, n_419, n_420, n_421;
  wire n_423, n_424, n_426, n_428, n_430, n_431, n_432, n_434;
  wire n_435, n_436, n_438, n_440, n_441, n_442, n_444, n_445;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_463;
  wire n_466, n_468, n_469, n_470, n_473, n_476, n_478, n_479;
  wire n_481, n_483, n_484, n_486, n_488, n_489, n_491, n_493;
  wire n_494, n_496, n_497, n_499, n_502, n_504, n_505, n_506;
  wire n_509, n_511, n_512, n_513, n_515, n_516, n_518, n_519;
  wire n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_531, n_532, n_533, n_535, n_536, n_537;
  wire n_539, n_540, n_541, n_543, n_544, n_545, n_547, n_548;
  wire n_549, n_551, n_552, n_553, n_555, n_556, n_557, n_559;
  wire n_560, n_561, n_563, n_564, n_565, n_567, n_568, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578;
  wire n_579, n_580, n_581, n_583, n_584, n_585, n_587, n_588;
  wire n_589, n_591, n_592, n_593, n_594, n_596, n_597, n_598;
  wire n_600, n_601, n_602, n_603, n_605, n_606, n_607, n_609;
  wire n_610, n_611, n_612, n_614, n_615, n_617, n_618, n_620;
  wire n_621, n_622, n_623, n_625, n_626, n_627, n_629, n_630;
  wire n_631, n_632, n_634, n_635, n_637, n_638, n_640, n_641;
  wire n_642, n_643, n_645, n_646, n_647, n_648, n_650, n_651;
  wire n_652, n_653, n_655, n_656, n_658, n_659, n_661, n_662;
  wire n_663, n_664, n_666, n_667, n_668, n_670, n_671, n_672;
  wire n_673, n_675, n_676, n_678, n_679, n_681, n_682, n_683;
  wire n_684, n_686, n_687, n_688, n_689, n_691, n_692, n_693;
  wire n_694;
  not g3 (Z[43], n_134);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_135, A[0], B[0]);
  nor g9 (n_138, A[1], B[1]);
  nand g10 (n_141, A[1], B[1]);
  nor g11 (n_148, A[2], B[2]);
  nand g12 (n_143, A[2], B[2]);
  nor g13 (n_144, A[3], B[3]);
  nand g14 (n_145, A[3], B[3]);
  nor g15 (n_154, A[4], B[4]);
  nand g16 (n_149, A[4], B[4]);
  nor g17 (n_150, A[5], B[5]);
  nand g18 (n_151, A[5], B[5]);
  nor g19 (n_160, A[6], B[6]);
  nand g20 (n_155, A[6], B[6]);
  nor g21 (n_156, A[7], B[7]);
  nand g22 (n_157, A[7], B[7]);
  nor g23 (n_166, A[8], B[8]);
  nand g24 (n_161, A[8], B[8]);
  nor g25 (n_162, A[9], B[9]);
  nand g26 (n_163, A[9], B[9]);
  nor g27 (n_172, A[10], B[10]);
  nand g28 (n_167, A[10], B[10]);
  nor g29 (n_168, A[11], B[11]);
  nand g30 (n_169, A[11], B[11]);
  nor g31 (n_178, A[12], B[12]);
  nand g32 (n_173, A[12], B[12]);
  nor g33 (n_174, A[13], B[13]);
  nand g34 (n_175, A[13], B[13]);
  nor g35 (n_184, A[14], B[14]);
  nand g36 (n_179, A[14], B[14]);
  nor g37 (n_180, A[15], B[15]);
  nand g38 (n_181, A[15], B[15]);
  nor g39 (n_190, A[16], B[16]);
  nand g40 (n_185, A[16], B[16]);
  nor g41 (n_186, A[17], B[17]);
  nand g42 (n_187, A[17], B[17]);
  nor g43 (n_196, A[18], B[18]);
  nand g44 (n_191, A[18], B[18]);
  nor g45 (n_192, A[19], B[19]);
  nand g46 (n_193, A[19], B[19]);
  nor g47 (n_202, A[20], B[20]);
  nand g48 (n_197, A[20], B[20]);
  nor g49 (n_198, A[21], B[21]);
  nand g50 (n_199, A[21], B[21]);
  nor g51 (n_208, A[22], B[22]);
  nand g52 (n_203, A[22], B[22]);
  nor g53 (n_204, A[23], B[23]);
  nand g54 (n_205, A[23], B[23]);
  nor g55 (n_214, A[24], B[24]);
  nand g56 (n_209, A[24], B[24]);
  nor g57 (n_210, A[25], B[25]);
  nand g58 (n_211, A[25], B[25]);
  nor g59 (n_220, A[26], B[26]);
  nand g60 (n_215, A[26], B[26]);
  nor g61 (n_216, A[27], B[27]);
  nand g62 (n_217, A[27], B[27]);
  nor g63 (n_226, A[28], B[28]);
  nand g64 (n_221, A[28], B[28]);
  nor g65 (n_222, A[29], B[29]);
  nand g66 (n_223, A[29], B[29]);
  nor g67 (n_232, A[30], B[30]);
  nand g68 (n_227, A[30], B[30]);
  nor g69 (n_228, A[31], B[31]);
  nand g70 (n_229, A[31], B[31]);
  nor g71 (n_238, A[32], B[32]);
  nand g72 (n_233, A[32], B[32]);
  nor g73 (n_234, A[33], B[33]);
  nand g74 (n_235, A[33], B[33]);
  nor g75 (n_244, A[34], B[34]);
  nand g76 (n_239, A[34], B[34]);
  nor g77 (n_240, A[35], B[35]);
  nand g78 (n_241, A[35], B[35]);
  nor g79 (n_250, A[36], B[36]);
  nand g80 (n_245, A[36], B[36]);
  nor g81 (n_246, A[37], B[37]);
  nand g82 (n_247, A[37], B[37]);
  nor g83 (n_256, A[38], B[38]);
  nand g84 (n_251, A[38], B[38]);
  nor g85 (n_252, A[39], B[39]);
  nand g86 (n_253, A[39], B[39]);
  nor g87 (n_262, A[40], B[40]);
  nand g88 (n_257, A[40], B[40]);
  nor g89 (n_258, A[41], B[41]);
  nand g90 (n_259, A[41], B[41]);
  nand g95 (n_263, n_141, n_142);
  nor g96 (n_146, n_143, n_144);
  nor g99 (n_266, n_148, n_144);
  nor g100 (n_152, n_149, n_150);
  nor g103 (n_272, n_154, n_150);
  nor g104 (n_158, n_155, n_156);
  nor g107 (n_274, n_160, n_156);
  nor g108 (n_164, n_161, n_162);
  nor g111 (n_282, n_166, n_162);
  nor g112 (n_170, n_167, n_168);
  nor g115 (n_284, n_172, n_168);
  nor g116 (n_176, n_173, n_174);
  nor g119 (n_292, n_178, n_174);
  nor g120 (n_182, n_179, n_180);
  nor g123 (n_294, n_184, n_180);
  nor g124 (n_188, n_185, n_186);
  nor g127 (n_302, n_190, n_186);
  nor g128 (n_194, n_191, n_192);
  nor g131 (n_304, n_196, n_192);
  nor g132 (n_200, n_197, n_198);
  nor g135 (n_312, n_202, n_198);
  nor g136 (n_206, n_203, n_204);
  nor g139 (n_314, n_208, n_204);
  nor g140 (n_212, n_209, n_210);
  nor g143 (n_322, n_214, n_210);
  nor g144 (n_218, n_215, n_216);
  nor g147 (n_324, n_220, n_216);
  nor g148 (n_224, n_221, n_222);
  nor g151 (n_332, n_226, n_222);
  nor g152 (n_230, n_227, n_228);
  nor g155 (n_334, n_232, n_228);
  nor g156 (n_236, n_233, n_234);
  nor g159 (n_342, n_238, n_234);
  nor g160 (n_242, n_239, n_240);
  nor g163 (n_344, n_244, n_240);
  nor g164 (n_248, n_245, n_246);
  nor g167 (n_352, n_250, n_246);
  nor g168 (n_254, n_251, n_252);
  nor g171 (n_354, n_256, n_252);
  nor g172 (n_260, n_257, n_258);
  nor g175 (n_364, n_262, n_258);
  nand g178 (n_596, n_143, n_265);
  nand g179 (n_268, n_266, n_263);
  nand g180 (n_366, n_267, n_268);
  nor g181 (n_270, n_160, n_269);
  nand g190 (n_374, n_272, n_274);
  nor g191 (n_280, n_172, n_279);
  nand g200 (n_381, n_282, n_284);
  nor g201 (n_290, n_184, n_289);
  nand g210 (n_389, n_292, n_294);
  nor g211 (n_300, n_196, n_299);
  nand g220 (n_396, n_302, n_304);
  nor g221 (n_310, n_208, n_309);
  nand g230 (n_404, n_312, n_314);
  nor g231 (n_320, n_220, n_319);
  nand g240 (n_411, n_322, n_324);
  nor g241 (n_330, n_232, n_329);
  nand g250 (n_419, n_332, n_334);
  nor g251 (n_340, n_244, n_339);
  nand g260 (n_426, n_342, n_344);
  nor g261 (n_350, n_256, n_349);
  nand g270 (n_434, n_352, n_354);
  nor g271 (n_362, n_359, n_360);
  nand g278 (n_600, n_149, n_368);
  nand g279 (n_369, n_272, n_366);
  nand g280 (n_602, n_269, n_369);
  nand g283 (n_605, n_372, n_373);
  nand g286 (n_438, n_376, n_377);
  nor g287 (n_379, n_178, n_378);
  nor g290 (n_448, n_178, n_381);
  nor g296 (n_387, n_385, n_378);
  nor g299 (n_454, n_381, n_385);
  nor g300 (n_391, n_389, n_378);
  nor g303 (n_457, n_381, n_389);
  nor g304 (n_394, n_202, n_393);
  nor g307 (n_519, n_202, n_396);
  nor g313 (n_402, n_400, n_393);
  nor g316 (n_525, n_396, n_400);
  nor g317 (n_406, n_404, n_393);
  nor g320 (n_463, n_396, n_404);
  nor g321 (n_409, n_226, n_408);
  nor g324 (n_476, n_226, n_411);
  nor g330 (n_417, n_415, n_408);
  nor g333 (n_486, n_411, n_415);
  nor g334 (n_421, n_419, n_408);
  nor g337 (n_491, n_411, n_419);
  nor g338 (n_424, n_250, n_423);
  nor g341 (n_571, n_250, n_426);
  nor g347 (n_432, n_430, n_423);
  nor g350 (n_577, n_426, n_430);
  nor g351 (n_436, n_434, n_423);
  nor g354 (n_499, n_426, n_434);
  nand g357 (n_609, n_161, n_440);
  nand g358 (n_441, n_282, n_438);
  nand g359 (n_611, n_279, n_441);
  nand g362 (n_614, n_444, n_445);
  nand g365 (n_617, n_378, n_447);
  nand g366 (n_450, n_448, n_438);
  nand g367 (n_620, n_449, n_450);
  nand g368 (n_453, n_451, n_438);
  nand g369 (n_622, n_452, n_453);
  nand g370 (n_456, n_454, n_438);
  nand g371 (n_625, n_455, n_456);
  nand g372 (n_459, n_457, n_438);
  nand g373 (n_509, n_458, n_459);
  nor g374 (n_461, n_214, n_460);
  nand g383 (n_533, n_322, n_463);
  nor g384 (n_470, n_468, n_460);
  nor g389 (n_473, n_411, n_460);
  nand g398 (n_545, n_463, n_476);
  nand g403 (n_549, n_463, n_481);
  nand g408 (n_553, n_463, n_486);
  nand g413 (n_557, n_463, n_491);
  nor g414 (n_497, n_262, n_496);
  nand g423 (n_585, n_364, n_499);
  nor g424 (n_506, n_504, n_496);
  nand g431 (n_629, n_185, n_511);
  nand g432 (n_512, n_302, n_509);
  nand g433 (n_631, n_299, n_512);
  nand g436 (n_634, n_515, n_516);
  nand g439 (n_637, n_393, n_518);
  nand g440 (n_521, n_519, n_509);
  nand g441 (n_640, n_520, n_521);
  nand g442 (n_524, n_522, n_509);
  nand g443 (n_642, n_523, n_524);
  nand g444 (n_527, n_525, n_509);
  nand g445 (n_645, n_526, n_527);
  nand g446 (n_528, n_463, n_509);
  nand g447 (n_647, n_460, n_528);
  nand g450 (n_650, n_531, n_532);
  nand g453 (n_652, n_535, n_536);
  nand g456 (n_655, n_539, n_540);
  nand g459 (n_658, n_543, n_544);
  nand g462 (n_661, n_547, n_548);
  nand g465 (n_663, n_551, n_552);
  nand g468 (n_666, n_555, n_556);
  nand g471 (n_561, n_559, n_560);
  nand g474 (n_670, n_233, n_563);
  nand g475 (n_564, n_342, n_561);
  nand g476 (n_672, n_339, n_564);
  nand g479 (n_675, n_567, n_568);
  nand g482 (n_678, n_423, n_570);
  nand g483 (n_573, n_571, n_561);
  nand g484 (n_681, n_572, n_573);
  nand g485 (n_576, n_574, n_561);
  nand g486 (n_683, n_575, n_576);
  nand g487 (n_579, n_577, n_561);
  nand g488 (n_686, n_578, n_579);
  nand g489 (n_580, n_499, n_561);
  nand g490 (n_688, n_496, n_580);
  nand g493 (n_691, n_583, n_584);
  nand g496 (n_693, n_587, n_588);
  nand g499 (n_134, n_591, n_592);
  xnor g503 (Z[2], n_263, n_594);
  xnor g506 (Z[3], n_596, n_597);
  xnor g508 (Z[4], n_366, n_598);
  xnor g511 (Z[5], n_600, n_601);
  xnor g513 (Z[6], n_602, n_603);
  xnor g516 (Z[7], n_605, n_606);
  xnor g518 (Z[8], n_438, n_607);
  xnor g521 (Z[9], n_609, n_610);
  xnor g523 (Z[10], n_611, n_612);
  xnor g526 (Z[11], n_614, n_615);
  xnor g529 (Z[12], n_617, n_618);
  xnor g532 (Z[13], n_620, n_621);
  xnor g534 (Z[14], n_622, n_623);
  xnor g537 (Z[15], n_625, n_626);
  xnor g539 (Z[16], n_509, n_627);
  xnor g542 (Z[17], n_629, n_630);
  xnor g544 (Z[18], n_631, n_632);
  xnor g547 (Z[19], n_634, n_635);
  xnor g550 (Z[20], n_637, n_638);
  xnor g553 (Z[21], n_640, n_641);
  xnor g555 (Z[22], n_642, n_643);
  xnor g558 (Z[23], n_645, n_646);
  xnor g560 (Z[24], n_647, n_648);
  xnor g563 (Z[25], n_650, n_651);
  xnor g565 (Z[26], n_652, n_653);
  xnor g568 (Z[27], n_655, n_656);
  xnor g571 (Z[28], n_658, n_659);
  xnor g574 (Z[29], n_661, n_662);
  xnor g576 (Z[30], n_663, n_664);
  xnor g579 (Z[31], n_666, n_667);
  xnor g581 (Z[32], n_561, n_668);
  xnor g584 (Z[33], n_670, n_671);
  xnor g586 (Z[34], n_672, n_673);
  xnor g589 (Z[35], n_675, n_676);
  xnor g592 (Z[36], n_678, n_679);
  xnor g595 (Z[37], n_681, n_682);
  xnor g597 (Z[38], n_683, n_684);
  xnor g600 (Z[39], n_686, n_687);
  xnor g602 (Z[40], n_688, n_689);
  xnor g605 (Z[41], n_691, n_692);
  xnor g607 (Z[42], n_693, n_694);
  and g610 (n_359, A[42], B[42]);
  or g611 (n_361, A[42], B[42]);
  and g612 (n_339, wc, n_235);
  not gc (wc, n_236);
  and g613 (n_346, wc0, n_241);
  not gc0 (wc0, n_242);
  and g614 (n_349, wc1, n_247);
  not gc1 (wc1, n_248);
  and g615 (n_356, wc2, n_253);
  not gc2 (wc2, n_254);
  and g616 (n_360, wc3, n_259);
  not gc3 (wc3, n_260);
  and g617 (n_299, wc4, n_187);
  not gc4 (wc4, n_188);
  and g618 (n_306, wc5, n_193);
  not gc5 (wc5, n_194);
  and g619 (n_309, wc6, n_199);
  not gc6 (wc6, n_200);
  and g620 (n_316, wc7, n_205);
  not gc7 (wc7, n_206);
  and g621 (n_319, wc8, n_211);
  not gc8 (wc8, n_212);
  and g622 (n_326, wc9, n_217);
  not gc9 (wc9, n_218);
  and g623 (n_329, wc10, n_223);
  not gc10 (wc10, n_224);
  and g624 (n_336, wc11, n_229);
  not gc11 (wc11, n_230);
  and g625 (n_279, wc12, n_163);
  not gc12 (wc12, n_164);
  and g626 (n_286, wc13, n_169);
  not gc13 (wc13, n_170);
  and g627 (n_289, wc14, n_175);
  not gc14 (wc14, n_176);
  and g628 (n_296, wc15, n_181);
  not gc15 (wc15, n_182);
  and g629 (n_269, wc16, n_151);
  not gc16 (wc16, n_152);
  and g630 (n_276, wc17, n_157);
  not gc17 (wc17, n_158);
  and g631 (n_267, wc18, n_145);
  not gc18 (wc18, n_146);
  or g632 (n_142, n_135, n_138);
  or g633 (n_370, wc19, n_160);
  not gc19 (wc19, n_272);
  or g634 (n_442, wc20, n_172);
  not gc20 (wc20, n_282);
  or g635 (n_385, wc21, n_184);
  not gc21 (wc21, n_292);
  or g636 (n_513, wc22, n_196);
  not gc22 (wc22, n_302);
  or g637 (n_400, wc23, n_208);
  not gc23 (wc23, n_312);
  or g638 (n_468, wc24, n_220);
  not gc24 (wc24, n_322);
  or g639 (n_415, wc25, n_232);
  not gc25 (wc25, n_332);
  or g640 (n_565, wc26, n_244);
  not gc26 (wc26, n_342);
  or g641 (n_430, wc27, n_256);
  not gc27 (wc27, n_352);
  or g642 (n_593, wc28, n_138);
  not gc28 (wc28, n_141);
  or g643 (n_594, wc29, n_148);
  not gc29 (wc29, n_143);
  or g644 (n_597, wc30, n_144);
  not gc30 (wc30, n_145);
  or g645 (n_598, wc31, n_154);
  not gc31 (wc31, n_149);
  or g646 (n_601, wc32, n_150);
  not gc32 (wc32, n_151);
  or g647 (n_603, wc33, n_160);
  not gc33 (wc33, n_155);
  or g648 (n_606, wc34, n_156);
  not gc34 (wc34, n_157);
  or g649 (n_607, wc35, n_166);
  not gc35 (wc35, n_161);
  or g650 (n_610, wc36, n_162);
  not gc36 (wc36, n_163);
  or g651 (n_612, wc37, n_172);
  not gc37 (wc37, n_167);
  or g652 (n_615, wc38, n_168);
  not gc38 (wc38, n_169);
  or g653 (n_618, wc39, n_178);
  not gc39 (wc39, n_173);
  or g654 (n_621, wc40, n_174);
  not gc40 (wc40, n_175);
  or g655 (n_623, wc41, n_184);
  not gc41 (wc41, n_179);
  or g656 (n_626, wc42, n_180);
  not gc42 (wc42, n_181);
  or g657 (n_627, wc43, n_190);
  not gc43 (wc43, n_185);
  or g658 (n_630, wc44, n_186);
  not gc44 (wc44, n_187);
  or g659 (n_632, wc45, n_196);
  not gc45 (wc45, n_191);
  or g660 (n_635, wc46, n_192);
  not gc46 (wc46, n_193);
  or g661 (n_638, wc47, n_202);
  not gc47 (wc47, n_197);
  or g662 (n_641, wc48, n_198);
  not gc48 (wc48, n_199);
  or g663 (n_643, wc49, n_208);
  not gc49 (wc49, n_203);
  or g664 (n_646, wc50, n_204);
  not gc50 (wc50, n_205);
  or g665 (n_648, wc51, n_214);
  not gc51 (wc51, n_209);
  or g666 (n_651, wc52, n_210);
  not gc52 (wc52, n_211);
  or g667 (n_653, wc53, n_220);
  not gc53 (wc53, n_215);
  or g668 (n_656, wc54, n_216);
  not gc54 (wc54, n_217);
  or g669 (n_659, wc55, n_226);
  not gc55 (wc55, n_221);
  or g670 (n_662, wc56, n_222);
  not gc56 (wc56, n_223);
  or g671 (n_664, wc57, n_232);
  not gc57 (wc57, n_227);
  or g672 (n_667, wc58, n_228);
  not gc58 (wc58, n_229);
  or g673 (n_668, wc59, n_238);
  not gc59 (wc59, n_233);
  or g674 (n_671, wc60, n_234);
  not gc60 (wc60, n_235);
  or g675 (n_673, wc61, n_244);
  not gc61 (wc61, n_239);
  or g676 (n_676, wc62, n_240);
  not gc62 (wc62, n_241);
  or g677 (n_679, wc63, n_250);
  not gc63 (wc63, n_245);
  or g678 (n_682, wc64, n_246);
  not gc64 (wc64, n_247);
  or g679 (n_684, wc65, n_256);
  not gc65 (wc65, n_251);
  or g680 (n_687, wc66, n_252);
  not gc66 (wc66, n_253);
  or g681 (n_689, wc67, n_262);
  not gc67 (wc67, n_257);
  or g682 (n_692, wc68, n_258);
  not gc68 (wc68, n_259);
  or g683 (n_504, n_359, wc69);
  not gc69 (wc69, n_364);
  and g684 (n_347, wc70, n_344);
  not gc70 (wc70, n_339);
  and g685 (n_357, wc71, n_354);
  not gc71 (wc71, n_349);
  and g686 (n_307, wc72, n_304);
  not gc72 (wc72, n_299);
  and g687 (n_317, wc73, n_314);
  not gc73 (wc73, n_309);
  and g688 (n_327, wc74, n_324);
  not gc74 (wc74, n_319);
  and g689 (n_337, wc75, n_334);
  not gc75 (wc75, n_329);
  and g690 (n_287, wc76, n_284);
  not gc76 (wc76, n_279);
  and g691 (n_297, wc77, n_294);
  not gc77 (wc77, n_289);
  and g692 (n_277, wc78, n_274);
  not gc78 (wc78, n_269);
  and g693 (n_451, wc79, n_292);
  not gc79 (wc79, n_381);
  and g694 (n_522, wc80, n_312);
  not gc80 (wc80, n_396);
  and g695 (n_481, wc81, n_332);
  not gc81 (wc81, n_411);
  and g696 (n_574, wc82, n_352);
  not gc82 (wc82, n_426);
  xor g697 (Z[1], n_135, n_593);
  or g698 (n_694, wc83, n_359);
  not gc83 (wc83, n_361);
  and g699 (n_423, wc84, n_346);
  not gc84 (wc84, n_347);
  and g700 (n_435, wc85, n_356);
  not gc85 (wc85, n_357);
  and g701 (n_505, n_361, wc86);
  not gc86 (wc86, n_362);
  and g702 (n_393, wc87, n_306);
  not gc87 (wc87, n_307);
  and g703 (n_405, wc88, n_316);
  not gc88 (wc88, n_317);
  and g704 (n_408, wc89, n_326);
  not gc89 (wc89, n_327);
  and g705 (n_420, wc90, n_336);
  not gc90 (wc90, n_337);
  and g706 (n_378, wc91, n_286);
  not gc91 (wc91, n_287);
  and g707 (n_390, wc92, n_296);
  not gc92 (wc92, n_297);
  and g708 (n_376, wc93, n_276);
  not gc93 (wc93, n_277);
  or g709 (n_265, wc94, n_148);
  not gc94 (wc94, n_263);
  and g710 (n_372, wc95, n_155);
  not gc95 (wc95, n_270);
  and g711 (n_444, wc96, n_167);
  not gc96 (wc96, n_280);
  and g712 (n_386, wc97, n_179);
  not gc97 (wc97, n_290);
  and g713 (n_515, wc98, n_191);
  not gc98 (wc98, n_300);
  and g714 (n_401, wc99, n_203);
  not gc99 (wc99, n_310);
  and g715 (n_469, wc100, n_215);
  not gc100 (wc100, n_320);
  and g716 (n_416, wc101, n_227);
  not gc101 (wc101, n_330);
  and g717 (n_567, wc102, n_239);
  not gc102 (wc102, n_340);
  and g718 (n_431, wc103, n_251);
  not gc103 (wc103, n_350);
  or g719 (n_529, wc104, n_214);
  not gc104 (wc104, n_463);
  or g720 (n_537, n_468, wc105);
  not gc105 (wc105, n_463);
  or g721 (n_541, wc106, n_411);
  not gc106 (wc106, n_463);
  or g722 (n_581, wc107, n_262);
  not gc107 (wc107, n_499);
  or g723 (n_589, n_504, wc108);
  not gc108 (wc108, n_499);
  and g724 (n_383, wc109, n_292);
  not gc109 (wc109, n_378);
  and g725 (n_398, wc110, n_312);
  not gc110 (wc110, n_393);
  and g726 (n_413, wc111, n_332);
  not gc111 (wc111, n_408);
  and g727 (n_428, wc112, n_352);
  not gc112 (wc112, n_423);
  and g728 (n_496, n_435, wc113);
  not gc113 (wc113, n_436);
  and g729 (n_460, n_405, wc114);
  not gc114 (wc114, n_406);
  and g730 (n_493, n_420, wc115);
  not gc115 (wc115, n_421);
  and g731 (n_458, n_390, wc116);
  not gc116 (wc116, n_391);
  or g732 (n_377, n_374, wc117);
  not gc117 (wc117, n_366);
  or g733 (n_368, wc118, n_154);
  not gc118 (wc118, n_366);
  or g734 (n_373, n_370, wc119);
  not gc119 (wc119, n_366);
  and g735 (n_449, wc120, n_173);
  not gc120 (wc120, n_379);
  and g736 (n_452, wc121, n_289);
  not gc121 (wc121, n_383);
  and g737 (n_455, n_386, wc122);
  not gc122 (wc122, n_387);
  and g738 (n_520, wc123, n_197);
  not gc123 (wc123, n_394);
  and g739 (n_523, wc124, n_309);
  not gc124 (wc124, n_398);
  and g740 (n_526, n_401, wc125);
  not gc125 (wc125, n_402);
  and g741 (n_478, wc126, n_221);
  not gc126 (wc126, n_409);
  and g742 (n_483, wc127, n_329);
  not gc127 (wc127, n_413);
  and g743 (n_488, n_416, wc128);
  not gc128 (wc128, n_417);
  and g744 (n_572, wc129, n_245);
  not gc129 (wc129, n_424);
  and g745 (n_575, wc130, n_349);
  not gc130 (wc130, n_428);
  and g746 (n_578, n_431, wc131);
  not gc131 (wc131, n_432);
  and g747 (n_494, wc132, n_491);
  not gc132 (wc132, n_460);
  and g748 (n_466, wc133, n_322);
  not gc133 (wc133, n_460);
  and g749 (n_479, wc134, n_476);
  not gc134 (wc134, n_460);
  and g750 (n_484, wc135, n_481);
  not gc135 (wc135, n_460);
  and g751 (n_489, wc136, n_486);
  not gc136 (wc136, n_460);
  and g752 (n_502, wc137, n_364);
  not gc137 (wc137, n_496);
  and g753 (n_591, n_505, wc138);
  not gc138 (wc138, n_506);
  and g754 (n_559, wc139, n_493);
  not gc139 (wc139, n_494);
  or g755 (n_440, wc140, n_166);
  not gc140 (wc140, n_438);
  or g756 (n_445, n_442, wc141);
  not gc141 (wc141, n_438);
  or g757 (n_447, wc142, n_381);
  not gc142 (wc142, n_438);
  and g758 (n_531, wc143, n_209);
  not gc143 (wc143, n_461);
  and g759 (n_535, wc144, n_319);
  not gc144 (wc144, n_466);
  and g760 (n_539, n_469, wc145);
  not gc145 (wc145, n_470);
  and g761 (n_543, n_408, wc146);
  not gc146 (wc146, n_473);
  and g762 (n_547, wc147, n_478);
  not gc147 (wc147, n_479);
  and g763 (n_551, wc148, n_483);
  not gc148 (wc148, n_484);
  and g764 (n_555, wc149, n_488);
  not gc149 (wc149, n_489);
  and g765 (n_583, wc150, n_257);
  not gc150 (wc150, n_497);
  and g766 (n_587, wc151, n_360);
  not gc151 (wc151, n_502);
  or g767 (n_560, n_557, wc152);
  not gc152 (wc152, n_509);
  or g768 (n_511, wc153, n_190);
  not gc153 (wc153, n_509);
  or g769 (n_516, n_513, wc154);
  not gc154 (wc154, n_509);
  or g770 (n_518, wc155, n_396);
  not gc155 (wc155, n_509);
  or g771 (n_532, n_529, wc156);
  not gc156 (wc156, n_509);
  or g772 (n_536, n_533, wc157);
  not gc157 (wc157, n_509);
  or g773 (n_540, n_537, wc158);
  not gc158 (wc158, n_509);
  or g774 (n_544, n_541, wc159);
  not gc159 (wc159, n_509);
  or g775 (n_548, n_545, wc160);
  not gc160 (wc160, n_509);
  or g776 (n_552, n_549, wc161);
  not gc161 (wc161, n_509);
  or g777 (n_556, n_553, wc162);
  not gc162 (wc162, n_509);
  or g778 (n_592, n_589, wc163);
  not gc163 (wc163, n_561);
  or g779 (n_563, wc164, n_238);
  not gc164 (wc164, n_561);
  or g780 (n_568, n_565, wc165);
  not gc165 (wc165, n_561);
  or g781 (n_570, wc166, n_426);
  not gc166 (wc166, n_561);
  or g782 (n_584, n_581, wc167);
  not gc167 (wc167, n_561);
  or g783 (n_588, wc168, n_585);
  not gc168 (wc168, n_561);
endmodule

module add_signed_412_1_GENERIC(A, B, Z);
  input [42:0] A, B;
  output [43:0] Z;
  wire [42:0] A, B;
  wire [43:0] Z;
  add_signed_412_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_412_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [42:0] A, B;
  output [43:0] Z;
  wire [42:0] A, B;
  wire [43:0] Z;
  wire n_134, n_135, n_138, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_148, n_149, n_150, n_151, n_152, n_154, n_155;
  wire n_156, n_157, n_158, n_160, n_161, n_162, n_163, n_164;
  wire n_166, n_167, n_168, n_169, n_170, n_172, n_173, n_174;
  wire n_175, n_176, n_178, n_179, n_180, n_181, n_182, n_184;
  wire n_185, n_186, n_187, n_188, n_190, n_191, n_192, n_193;
  wire n_194, n_196, n_197, n_198, n_199, n_200, n_202, n_203;
  wire n_204, n_205, n_206, n_208, n_209, n_210, n_211, n_212;
  wire n_214, n_215, n_216, n_217, n_218, n_220, n_221, n_222;
  wire n_223, n_224, n_226, n_227, n_228, n_229, n_230, n_232;
  wire n_233, n_234, n_235, n_236, n_238, n_239, n_240, n_241;
  wire n_242, n_244, n_245, n_246, n_247, n_248, n_250, n_251;
  wire n_252, n_253, n_254, n_256, n_257, n_258, n_259, n_260;
  wire n_262, n_263, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_272, n_274, n_276, n_277, n_279, n_280, n_282, n_284;
  wire n_286, n_287, n_289, n_290, n_292, n_294, n_296, n_297;
  wire n_299, n_300, n_302, n_304, n_306, n_307, n_309, n_310;
  wire n_312, n_314, n_316, n_317, n_319, n_320, n_322, n_324;
  wire n_326, n_327, n_329, n_330, n_332, n_334, n_336, n_337;
  wire n_339, n_340, n_342, n_344, n_346, n_347, n_349, n_350;
  wire n_352, n_354, n_356, n_357, n_359, n_360, n_361, n_362;
  wire n_364, n_366, n_368, n_369, n_370, n_372, n_373, n_374;
  wire n_376, n_377, n_378, n_379, n_381, n_383, n_385, n_386;
  wire n_387, n_389, n_390, n_391, n_393, n_394, n_396, n_398;
  wire n_400, n_401, n_402, n_404, n_405, n_406, n_408, n_409;
  wire n_411, n_413, n_415, n_416, n_417, n_419, n_420, n_421;
  wire n_423, n_424, n_426, n_428, n_430, n_431, n_432, n_434;
  wire n_435, n_436, n_438, n_440, n_441, n_442, n_444, n_445;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_463;
  wire n_466, n_468, n_469, n_470, n_473, n_476, n_478, n_479;
  wire n_481, n_483, n_484, n_486, n_488, n_489, n_491, n_493;
  wire n_494, n_496, n_497, n_499, n_502, n_504, n_505, n_506;
  wire n_509, n_511, n_512, n_513, n_515, n_516, n_518, n_519;
  wire n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_531, n_532, n_533, n_535, n_536, n_537;
  wire n_539, n_540, n_541, n_543, n_544, n_545, n_547, n_548;
  wire n_549, n_551, n_552, n_553, n_555, n_556, n_557, n_559;
  wire n_560, n_561, n_563, n_564, n_565, n_567, n_568, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578;
  wire n_579, n_580, n_581, n_583, n_584, n_585, n_587, n_588;
  wire n_589, n_591, n_592, n_593, n_594, n_596, n_597, n_598;
  wire n_600, n_601, n_602, n_603, n_605, n_606, n_607, n_609;
  wire n_610, n_611, n_612, n_614, n_615, n_617, n_618, n_620;
  wire n_621, n_622, n_623, n_625, n_626, n_627, n_629, n_630;
  wire n_631, n_632, n_634, n_635, n_637, n_638, n_640, n_641;
  wire n_642, n_643, n_645, n_646, n_647, n_648, n_650, n_651;
  wire n_652, n_653, n_655, n_656, n_658, n_659, n_661, n_662;
  wire n_663, n_664, n_666, n_667, n_668, n_670, n_671, n_672;
  wire n_673, n_675, n_676, n_678, n_679, n_681, n_682, n_683;
  wire n_684, n_686, n_687, n_688, n_689, n_691, n_692, n_693;
  wire n_694;
  not g3 (Z[43], n_134);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_135, A[0], B[0]);
  nor g9 (n_138, A[1], B[1]);
  nand g10 (n_141, A[1], B[1]);
  nor g11 (n_148, A[2], B[2]);
  nand g12 (n_143, A[2], B[2]);
  nor g13 (n_144, A[3], B[3]);
  nand g14 (n_145, A[3], B[3]);
  nor g15 (n_154, A[4], B[4]);
  nand g16 (n_149, A[4], B[4]);
  nor g17 (n_150, A[5], B[5]);
  nand g18 (n_151, A[5], B[5]);
  nor g19 (n_160, A[6], B[6]);
  nand g20 (n_155, A[6], B[6]);
  nor g21 (n_156, A[7], B[7]);
  nand g22 (n_157, A[7], B[7]);
  nor g23 (n_166, A[8], B[8]);
  nand g24 (n_161, A[8], B[8]);
  nor g25 (n_162, A[9], B[9]);
  nand g26 (n_163, A[9], B[9]);
  nor g27 (n_172, A[10], B[10]);
  nand g28 (n_167, A[10], B[10]);
  nor g29 (n_168, A[11], B[11]);
  nand g30 (n_169, A[11], B[11]);
  nor g31 (n_178, A[12], B[12]);
  nand g32 (n_173, A[12], B[12]);
  nor g33 (n_174, A[13], B[13]);
  nand g34 (n_175, A[13], B[13]);
  nor g35 (n_184, A[14], B[14]);
  nand g36 (n_179, A[14], B[14]);
  nor g37 (n_180, A[15], B[15]);
  nand g38 (n_181, A[15], B[15]);
  nor g39 (n_190, A[16], B[16]);
  nand g40 (n_185, A[16], B[16]);
  nor g41 (n_186, A[17], B[17]);
  nand g42 (n_187, A[17], B[17]);
  nor g43 (n_196, A[18], B[18]);
  nand g44 (n_191, A[18], B[18]);
  nor g45 (n_192, A[19], B[19]);
  nand g46 (n_193, A[19], B[19]);
  nor g47 (n_202, A[20], B[20]);
  nand g48 (n_197, A[20], B[20]);
  nor g49 (n_198, A[21], B[21]);
  nand g50 (n_199, A[21], B[21]);
  nor g51 (n_208, A[22], B[22]);
  nand g52 (n_203, A[22], B[22]);
  nor g53 (n_204, A[23], B[23]);
  nand g54 (n_205, A[23], B[23]);
  nor g55 (n_214, A[24], B[24]);
  nand g56 (n_209, A[24], B[24]);
  nor g57 (n_210, A[25], B[25]);
  nand g58 (n_211, A[25], B[25]);
  nor g59 (n_220, A[26], B[26]);
  nand g60 (n_215, A[26], B[26]);
  nor g61 (n_216, A[27], B[27]);
  nand g62 (n_217, A[27], B[27]);
  nor g63 (n_226, A[28], B[28]);
  nand g64 (n_221, A[28], B[28]);
  nor g65 (n_222, A[29], B[29]);
  nand g66 (n_223, A[29], B[29]);
  nor g67 (n_232, A[30], B[30]);
  nand g68 (n_227, A[30], B[30]);
  nor g69 (n_228, A[31], B[31]);
  nand g70 (n_229, A[31], B[31]);
  nor g71 (n_238, A[32], B[32]);
  nand g72 (n_233, A[32], B[32]);
  nor g73 (n_234, A[33], B[33]);
  nand g74 (n_235, A[33], B[33]);
  nor g75 (n_244, A[34], B[34]);
  nand g76 (n_239, A[34], B[34]);
  nor g77 (n_240, A[35], B[35]);
  nand g78 (n_241, A[35], B[35]);
  nor g79 (n_250, A[36], B[36]);
  nand g80 (n_245, A[36], B[36]);
  nor g81 (n_246, A[37], B[37]);
  nand g82 (n_247, A[37], B[37]);
  nor g83 (n_256, A[38], B[38]);
  nand g84 (n_251, A[38], B[38]);
  nor g85 (n_252, A[39], B[39]);
  nand g86 (n_253, A[39], B[39]);
  nor g87 (n_262, A[40], B[40]);
  nand g88 (n_257, A[40], B[40]);
  nor g89 (n_258, A[41], B[41]);
  nand g90 (n_259, A[41], B[41]);
  nand g95 (n_263, n_141, n_142);
  nor g96 (n_146, n_143, n_144);
  nor g99 (n_266, n_148, n_144);
  nor g100 (n_152, n_149, n_150);
  nor g103 (n_272, n_154, n_150);
  nor g104 (n_158, n_155, n_156);
  nor g107 (n_274, n_160, n_156);
  nor g108 (n_164, n_161, n_162);
  nor g111 (n_282, n_166, n_162);
  nor g112 (n_170, n_167, n_168);
  nor g115 (n_284, n_172, n_168);
  nor g116 (n_176, n_173, n_174);
  nor g119 (n_292, n_178, n_174);
  nor g120 (n_182, n_179, n_180);
  nor g123 (n_294, n_184, n_180);
  nor g124 (n_188, n_185, n_186);
  nor g127 (n_302, n_190, n_186);
  nor g128 (n_194, n_191, n_192);
  nor g131 (n_304, n_196, n_192);
  nor g132 (n_200, n_197, n_198);
  nor g135 (n_312, n_202, n_198);
  nor g136 (n_206, n_203, n_204);
  nor g139 (n_314, n_208, n_204);
  nor g140 (n_212, n_209, n_210);
  nor g143 (n_322, n_214, n_210);
  nor g144 (n_218, n_215, n_216);
  nor g147 (n_324, n_220, n_216);
  nor g148 (n_224, n_221, n_222);
  nor g151 (n_332, n_226, n_222);
  nor g152 (n_230, n_227, n_228);
  nor g155 (n_334, n_232, n_228);
  nor g156 (n_236, n_233, n_234);
  nor g159 (n_342, n_238, n_234);
  nor g160 (n_242, n_239, n_240);
  nor g163 (n_344, n_244, n_240);
  nor g164 (n_248, n_245, n_246);
  nor g167 (n_352, n_250, n_246);
  nor g168 (n_254, n_251, n_252);
  nor g171 (n_354, n_256, n_252);
  nor g172 (n_260, n_257, n_258);
  nor g175 (n_364, n_262, n_258);
  nand g178 (n_596, n_143, n_265);
  nand g179 (n_268, n_266, n_263);
  nand g180 (n_366, n_267, n_268);
  nor g181 (n_270, n_160, n_269);
  nand g190 (n_374, n_272, n_274);
  nor g191 (n_280, n_172, n_279);
  nand g200 (n_381, n_282, n_284);
  nor g201 (n_290, n_184, n_289);
  nand g210 (n_389, n_292, n_294);
  nor g211 (n_300, n_196, n_299);
  nand g220 (n_396, n_302, n_304);
  nor g221 (n_310, n_208, n_309);
  nand g230 (n_404, n_312, n_314);
  nor g231 (n_320, n_220, n_319);
  nand g240 (n_411, n_322, n_324);
  nor g241 (n_330, n_232, n_329);
  nand g250 (n_419, n_332, n_334);
  nor g251 (n_340, n_244, n_339);
  nand g260 (n_426, n_342, n_344);
  nor g261 (n_350, n_256, n_349);
  nand g270 (n_434, n_352, n_354);
  nor g271 (n_362, n_359, n_360);
  nand g278 (n_600, n_149, n_368);
  nand g279 (n_369, n_272, n_366);
  nand g280 (n_602, n_269, n_369);
  nand g283 (n_605, n_372, n_373);
  nand g286 (n_438, n_376, n_377);
  nor g287 (n_379, n_178, n_378);
  nor g290 (n_448, n_178, n_381);
  nor g296 (n_387, n_385, n_378);
  nor g299 (n_454, n_381, n_385);
  nor g300 (n_391, n_389, n_378);
  nor g303 (n_457, n_381, n_389);
  nor g304 (n_394, n_202, n_393);
  nor g307 (n_519, n_202, n_396);
  nor g313 (n_402, n_400, n_393);
  nor g316 (n_525, n_396, n_400);
  nor g317 (n_406, n_404, n_393);
  nor g320 (n_463, n_396, n_404);
  nor g321 (n_409, n_226, n_408);
  nor g324 (n_476, n_226, n_411);
  nor g330 (n_417, n_415, n_408);
  nor g333 (n_486, n_411, n_415);
  nor g334 (n_421, n_419, n_408);
  nor g337 (n_491, n_411, n_419);
  nor g338 (n_424, n_250, n_423);
  nor g341 (n_571, n_250, n_426);
  nor g347 (n_432, n_430, n_423);
  nor g350 (n_577, n_426, n_430);
  nor g351 (n_436, n_434, n_423);
  nor g354 (n_499, n_426, n_434);
  nand g357 (n_609, n_161, n_440);
  nand g358 (n_441, n_282, n_438);
  nand g359 (n_611, n_279, n_441);
  nand g362 (n_614, n_444, n_445);
  nand g365 (n_617, n_378, n_447);
  nand g366 (n_450, n_448, n_438);
  nand g367 (n_620, n_449, n_450);
  nand g368 (n_453, n_451, n_438);
  nand g369 (n_622, n_452, n_453);
  nand g370 (n_456, n_454, n_438);
  nand g371 (n_625, n_455, n_456);
  nand g372 (n_459, n_457, n_438);
  nand g373 (n_509, n_458, n_459);
  nor g374 (n_461, n_214, n_460);
  nand g383 (n_533, n_322, n_463);
  nor g384 (n_470, n_468, n_460);
  nor g389 (n_473, n_411, n_460);
  nand g398 (n_545, n_463, n_476);
  nand g403 (n_549, n_463, n_481);
  nand g408 (n_553, n_463, n_486);
  nand g413 (n_557, n_463, n_491);
  nor g414 (n_497, n_262, n_496);
  nand g423 (n_585, n_364, n_499);
  nor g424 (n_506, n_504, n_496);
  nand g431 (n_629, n_185, n_511);
  nand g432 (n_512, n_302, n_509);
  nand g433 (n_631, n_299, n_512);
  nand g436 (n_634, n_515, n_516);
  nand g439 (n_637, n_393, n_518);
  nand g440 (n_521, n_519, n_509);
  nand g441 (n_640, n_520, n_521);
  nand g442 (n_524, n_522, n_509);
  nand g443 (n_642, n_523, n_524);
  nand g444 (n_527, n_525, n_509);
  nand g445 (n_645, n_526, n_527);
  nand g446 (n_528, n_463, n_509);
  nand g447 (n_647, n_460, n_528);
  nand g450 (n_650, n_531, n_532);
  nand g453 (n_652, n_535, n_536);
  nand g456 (n_655, n_539, n_540);
  nand g459 (n_658, n_543, n_544);
  nand g462 (n_661, n_547, n_548);
  nand g465 (n_663, n_551, n_552);
  nand g468 (n_666, n_555, n_556);
  nand g471 (n_561, n_559, n_560);
  nand g474 (n_670, n_233, n_563);
  nand g475 (n_564, n_342, n_561);
  nand g476 (n_672, n_339, n_564);
  nand g479 (n_675, n_567, n_568);
  nand g482 (n_678, n_423, n_570);
  nand g483 (n_573, n_571, n_561);
  nand g484 (n_681, n_572, n_573);
  nand g485 (n_576, n_574, n_561);
  nand g486 (n_683, n_575, n_576);
  nand g487 (n_579, n_577, n_561);
  nand g488 (n_686, n_578, n_579);
  nand g489 (n_580, n_499, n_561);
  nand g490 (n_688, n_496, n_580);
  nand g493 (n_691, n_583, n_584);
  nand g496 (n_693, n_587, n_588);
  nand g499 (n_134, n_591, n_592);
  xnor g503 (Z[2], n_263, n_594);
  xnor g506 (Z[3], n_596, n_597);
  xnor g508 (Z[4], n_366, n_598);
  xnor g511 (Z[5], n_600, n_601);
  xnor g513 (Z[6], n_602, n_603);
  xnor g516 (Z[7], n_605, n_606);
  xnor g518 (Z[8], n_438, n_607);
  xnor g521 (Z[9], n_609, n_610);
  xnor g523 (Z[10], n_611, n_612);
  xnor g526 (Z[11], n_614, n_615);
  xnor g529 (Z[12], n_617, n_618);
  xnor g532 (Z[13], n_620, n_621);
  xnor g534 (Z[14], n_622, n_623);
  xnor g537 (Z[15], n_625, n_626);
  xnor g539 (Z[16], n_509, n_627);
  xnor g542 (Z[17], n_629, n_630);
  xnor g544 (Z[18], n_631, n_632);
  xnor g547 (Z[19], n_634, n_635);
  xnor g550 (Z[20], n_637, n_638);
  xnor g553 (Z[21], n_640, n_641);
  xnor g555 (Z[22], n_642, n_643);
  xnor g558 (Z[23], n_645, n_646);
  xnor g560 (Z[24], n_647, n_648);
  xnor g563 (Z[25], n_650, n_651);
  xnor g565 (Z[26], n_652, n_653);
  xnor g568 (Z[27], n_655, n_656);
  xnor g571 (Z[28], n_658, n_659);
  xnor g574 (Z[29], n_661, n_662);
  xnor g576 (Z[30], n_663, n_664);
  xnor g579 (Z[31], n_666, n_667);
  xnor g581 (Z[32], n_561, n_668);
  xnor g584 (Z[33], n_670, n_671);
  xnor g586 (Z[34], n_672, n_673);
  xnor g589 (Z[35], n_675, n_676);
  xnor g592 (Z[36], n_678, n_679);
  xnor g595 (Z[37], n_681, n_682);
  xnor g597 (Z[38], n_683, n_684);
  xnor g600 (Z[39], n_686, n_687);
  xnor g602 (Z[40], n_688, n_689);
  xnor g605 (Z[41], n_691, n_692);
  xnor g607 (Z[42], n_693, n_694);
  and g610 (n_359, A[42], B[42]);
  or g611 (n_361, A[42], B[42]);
  and g612 (n_339, wc, n_235);
  not gc (wc, n_236);
  and g613 (n_346, wc0, n_241);
  not gc0 (wc0, n_242);
  and g614 (n_349, wc1, n_247);
  not gc1 (wc1, n_248);
  and g615 (n_356, wc2, n_253);
  not gc2 (wc2, n_254);
  and g616 (n_360, wc3, n_259);
  not gc3 (wc3, n_260);
  and g617 (n_299, wc4, n_187);
  not gc4 (wc4, n_188);
  and g618 (n_306, wc5, n_193);
  not gc5 (wc5, n_194);
  and g619 (n_309, wc6, n_199);
  not gc6 (wc6, n_200);
  and g620 (n_316, wc7, n_205);
  not gc7 (wc7, n_206);
  and g621 (n_319, wc8, n_211);
  not gc8 (wc8, n_212);
  and g622 (n_326, wc9, n_217);
  not gc9 (wc9, n_218);
  and g623 (n_329, wc10, n_223);
  not gc10 (wc10, n_224);
  and g624 (n_336, wc11, n_229);
  not gc11 (wc11, n_230);
  and g625 (n_279, wc12, n_163);
  not gc12 (wc12, n_164);
  and g626 (n_286, wc13, n_169);
  not gc13 (wc13, n_170);
  and g627 (n_289, wc14, n_175);
  not gc14 (wc14, n_176);
  and g628 (n_296, wc15, n_181);
  not gc15 (wc15, n_182);
  and g629 (n_269, wc16, n_151);
  not gc16 (wc16, n_152);
  and g630 (n_276, wc17, n_157);
  not gc17 (wc17, n_158);
  and g631 (n_267, wc18, n_145);
  not gc18 (wc18, n_146);
  or g632 (n_142, n_135, n_138);
  or g633 (n_370, wc19, n_160);
  not gc19 (wc19, n_272);
  or g634 (n_442, wc20, n_172);
  not gc20 (wc20, n_282);
  or g635 (n_385, wc21, n_184);
  not gc21 (wc21, n_292);
  or g636 (n_513, wc22, n_196);
  not gc22 (wc22, n_302);
  or g637 (n_400, wc23, n_208);
  not gc23 (wc23, n_312);
  or g638 (n_468, wc24, n_220);
  not gc24 (wc24, n_322);
  or g639 (n_415, wc25, n_232);
  not gc25 (wc25, n_332);
  or g640 (n_565, wc26, n_244);
  not gc26 (wc26, n_342);
  or g641 (n_430, wc27, n_256);
  not gc27 (wc27, n_352);
  or g642 (n_593, wc28, n_138);
  not gc28 (wc28, n_141);
  or g643 (n_594, wc29, n_148);
  not gc29 (wc29, n_143);
  or g644 (n_597, wc30, n_144);
  not gc30 (wc30, n_145);
  or g645 (n_598, wc31, n_154);
  not gc31 (wc31, n_149);
  or g646 (n_601, wc32, n_150);
  not gc32 (wc32, n_151);
  or g647 (n_603, wc33, n_160);
  not gc33 (wc33, n_155);
  or g648 (n_606, wc34, n_156);
  not gc34 (wc34, n_157);
  or g649 (n_607, wc35, n_166);
  not gc35 (wc35, n_161);
  or g650 (n_610, wc36, n_162);
  not gc36 (wc36, n_163);
  or g651 (n_612, wc37, n_172);
  not gc37 (wc37, n_167);
  or g652 (n_615, wc38, n_168);
  not gc38 (wc38, n_169);
  or g653 (n_618, wc39, n_178);
  not gc39 (wc39, n_173);
  or g654 (n_621, wc40, n_174);
  not gc40 (wc40, n_175);
  or g655 (n_623, wc41, n_184);
  not gc41 (wc41, n_179);
  or g656 (n_626, wc42, n_180);
  not gc42 (wc42, n_181);
  or g657 (n_627, wc43, n_190);
  not gc43 (wc43, n_185);
  or g658 (n_630, wc44, n_186);
  not gc44 (wc44, n_187);
  or g659 (n_632, wc45, n_196);
  not gc45 (wc45, n_191);
  or g660 (n_635, wc46, n_192);
  not gc46 (wc46, n_193);
  or g661 (n_638, wc47, n_202);
  not gc47 (wc47, n_197);
  or g662 (n_641, wc48, n_198);
  not gc48 (wc48, n_199);
  or g663 (n_643, wc49, n_208);
  not gc49 (wc49, n_203);
  or g664 (n_646, wc50, n_204);
  not gc50 (wc50, n_205);
  or g665 (n_648, wc51, n_214);
  not gc51 (wc51, n_209);
  or g666 (n_651, wc52, n_210);
  not gc52 (wc52, n_211);
  or g667 (n_653, wc53, n_220);
  not gc53 (wc53, n_215);
  or g668 (n_656, wc54, n_216);
  not gc54 (wc54, n_217);
  or g669 (n_659, wc55, n_226);
  not gc55 (wc55, n_221);
  or g670 (n_662, wc56, n_222);
  not gc56 (wc56, n_223);
  or g671 (n_664, wc57, n_232);
  not gc57 (wc57, n_227);
  or g672 (n_667, wc58, n_228);
  not gc58 (wc58, n_229);
  or g673 (n_668, wc59, n_238);
  not gc59 (wc59, n_233);
  or g674 (n_671, wc60, n_234);
  not gc60 (wc60, n_235);
  or g675 (n_673, wc61, n_244);
  not gc61 (wc61, n_239);
  or g676 (n_676, wc62, n_240);
  not gc62 (wc62, n_241);
  or g677 (n_679, wc63, n_250);
  not gc63 (wc63, n_245);
  or g678 (n_682, wc64, n_246);
  not gc64 (wc64, n_247);
  or g679 (n_684, wc65, n_256);
  not gc65 (wc65, n_251);
  or g680 (n_687, wc66, n_252);
  not gc66 (wc66, n_253);
  or g681 (n_689, wc67, n_262);
  not gc67 (wc67, n_257);
  or g682 (n_692, wc68, n_258);
  not gc68 (wc68, n_259);
  or g683 (n_504, n_359, wc69);
  not gc69 (wc69, n_364);
  and g684 (n_347, wc70, n_344);
  not gc70 (wc70, n_339);
  and g685 (n_357, wc71, n_354);
  not gc71 (wc71, n_349);
  and g686 (n_307, wc72, n_304);
  not gc72 (wc72, n_299);
  and g687 (n_317, wc73, n_314);
  not gc73 (wc73, n_309);
  and g688 (n_327, wc74, n_324);
  not gc74 (wc74, n_319);
  and g689 (n_337, wc75, n_334);
  not gc75 (wc75, n_329);
  and g690 (n_287, wc76, n_284);
  not gc76 (wc76, n_279);
  and g691 (n_297, wc77, n_294);
  not gc77 (wc77, n_289);
  and g692 (n_277, wc78, n_274);
  not gc78 (wc78, n_269);
  and g693 (n_451, wc79, n_292);
  not gc79 (wc79, n_381);
  and g694 (n_522, wc80, n_312);
  not gc80 (wc80, n_396);
  and g695 (n_481, wc81, n_332);
  not gc81 (wc81, n_411);
  and g696 (n_574, wc82, n_352);
  not gc82 (wc82, n_426);
  xor g697 (Z[1], n_135, n_593);
  or g698 (n_694, wc83, n_359);
  not gc83 (wc83, n_361);
  and g699 (n_423, wc84, n_346);
  not gc84 (wc84, n_347);
  and g700 (n_435, wc85, n_356);
  not gc85 (wc85, n_357);
  and g701 (n_505, n_361, wc86);
  not gc86 (wc86, n_362);
  and g702 (n_393, wc87, n_306);
  not gc87 (wc87, n_307);
  and g703 (n_405, wc88, n_316);
  not gc88 (wc88, n_317);
  and g704 (n_408, wc89, n_326);
  not gc89 (wc89, n_327);
  and g705 (n_420, wc90, n_336);
  not gc90 (wc90, n_337);
  and g706 (n_378, wc91, n_286);
  not gc91 (wc91, n_287);
  and g707 (n_390, wc92, n_296);
  not gc92 (wc92, n_297);
  and g708 (n_376, wc93, n_276);
  not gc93 (wc93, n_277);
  or g709 (n_265, wc94, n_148);
  not gc94 (wc94, n_263);
  and g710 (n_372, wc95, n_155);
  not gc95 (wc95, n_270);
  and g711 (n_444, wc96, n_167);
  not gc96 (wc96, n_280);
  and g712 (n_386, wc97, n_179);
  not gc97 (wc97, n_290);
  and g713 (n_515, wc98, n_191);
  not gc98 (wc98, n_300);
  and g714 (n_401, wc99, n_203);
  not gc99 (wc99, n_310);
  and g715 (n_469, wc100, n_215);
  not gc100 (wc100, n_320);
  and g716 (n_416, wc101, n_227);
  not gc101 (wc101, n_330);
  and g717 (n_567, wc102, n_239);
  not gc102 (wc102, n_340);
  and g718 (n_431, wc103, n_251);
  not gc103 (wc103, n_350);
  or g719 (n_529, wc104, n_214);
  not gc104 (wc104, n_463);
  or g720 (n_537, n_468, wc105);
  not gc105 (wc105, n_463);
  or g721 (n_541, wc106, n_411);
  not gc106 (wc106, n_463);
  or g722 (n_581, wc107, n_262);
  not gc107 (wc107, n_499);
  or g723 (n_589, n_504, wc108);
  not gc108 (wc108, n_499);
  and g724 (n_383, wc109, n_292);
  not gc109 (wc109, n_378);
  and g725 (n_398, wc110, n_312);
  not gc110 (wc110, n_393);
  and g726 (n_413, wc111, n_332);
  not gc111 (wc111, n_408);
  and g727 (n_428, wc112, n_352);
  not gc112 (wc112, n_423);
  and g728 (n_496, n_435, wc113);
  not gc113 (wc113, n_436);
  and g729 (n_460, n_405, wc114);
  not gc114 (wc114, n_406);
  and g730 (n_493, n_420, wc115);
  not gc115 (wc115, n_421);
  and g731 (n_458, n_390, wc116);
  not gc116 (wc116, n_391);
  or g732 (n_377, n_374, wc117);
  not gc117 (wc117, n_366);
  or g733 (n_368, wc118, n_154);
  not gc118 (wc118, n_366);
  or g734 (n_373, n_370, wc119);
  not gc119 (wc119, n_366);
  and g735 (n_449, wc120, n_173);
  not gc120 (wc120, n_379);
  and g736 (n_452, wc121, n_289);
  not gc121 (wc121, n_383);
  and g737 (n_455, n_386, wc122);
  not gc122 (wc122, n_387);
  and g738 (n_520, wc123, n_197);
  not gc123 (wc123, n_394);
  and g739 (n_523, wc124, n_309);
  not gc124 (wc124, n_398);
  and g740 (n_526, n_401, wc125);
  not gc125 (wc125, n_402);
  and g741 (n_478, wc126, n_221);
  not gc126 (wc126, n_409);
  and g742 (n_483, wc127, n_329);
  not gc127 (wc127, n_413);
  and g743 (n_488, n_416, wc128);
  not gc128 (wc128, n_417);
  and g744 (n_572, wc129, n_245);
  not gc129 (wc129, n_424);
  and g745 (n_575, wc130, n_349);
  not gc130 (wc130, n_428);
  and g746 (n_578, n_431, wc131);
  not gc131 (wc131, n_432);
  and g747 (n_494, wc132, n_491);
  not gc132 (wc132, n_460);
  and g748 (n_466, wc133, n_322);
  not gc133 (wc133, n_460);
  and g749 (n_479, wc134, n_476);
  not gc134 (wc134, n_460);
  and g750 (n_484, wc135, n_481);
  not gc135 (wc135, n_460);
  and g751 (n_489, wc136, n_486);
  not gc136 (wc136, n_460);
  and g752 (n_502, wc137, n_364);
  not gc137 (wc137, n_496);
  and g753 (n_591, n_505, wc138);
  not gc138 (wc138, n_506);
  and g754 (n_559, wc139, n_493);
  not gc139 (wc139, n_494);
  or g755 (n_440, wc140, n_166);
  not gc140 (wc140, n_438);
  or g756 (n_445, n_442, wc141);
  not gc141 (wc141, n_438);
  or g757 (n_447, wc142, n_381);
  not gc142 (wc142, n_438);
  and g758 (n_531, wc143, n_209);
  not gc143 (wc143, n_461);
  and g759 (n_535, wc144, n_319);
  not gc144 (wc144, n_466);
  and g760 (n_539, n_469, wc145);
  not gc145 (wc145, n_470);
  and g761 (n_543, n_408, wc146);
  not gc146 (wc146, n_473);
  and g762 (n_547, wc147, n_478);
  not gc147 (wc147, n_479);
  and g763 (n_551, wc148, n_483);
  not gc148 (wc148, n_484);
  and g764 (n_555, wc149, n_488);
  not gc149 (wc149, n_489);
  and g765 (n_583, wc150, n_257);
  not gc150 (wc150, n_497);
  and g766 (n_587, wc151, n_360);
  not gc151 (wc151, n_502);
  or g767 (n_560, n_557, wc152);
  not gc152 (wc152, n_509);
  or g768 (n_511, wc153, n_190);
  not gc153 (wc153, n_509);
  or g769 (n_516, n_513, wc154);
  not gc154 (wc154, n_509);
  or g770 (n_518, wc155, n_396);
  not gc155 (wc155, n_509);
  or g771 (n_532, n_529, wc156);
  not gc156 (wc156, n_509);
  or g772 (n_536, n_533, wc157);
  not gc157 (wc157, n_509);
  or g773 (n_540, n_537, wc158);
  not gc158 (wc158, n_509);
  or g774 (n_544, n_541, wc159);
  not gc159 (wc159, n_509);
  or g775 (n_548, n_545, wc160);
  not gc160 (wc160, n_509);
  or g776 (n_552, n_549, wc161);
  not gc161 (wc161, n_509);
  or g777 (n_556, n_553, wc162);
  not gc162 (wc162, n_509);
  or g778 (n_592, n_589, wc163);
  not gc163 (wc163, n_561);
  or g779 (n_563, wc164, n_238);
  not gc164 (wc164, n_561);
  or g780 (n_568, n_565, wc165);
  not gc165 (wc165, n_561);
  or g781 (n_570, wc166, n_426);
  not gc166 (wc166, n_561);
  or g782 (n_584, n_581, wc167);
  not gc167 (wc167, n_561);
  or g783 (n_588, wc168, n_585);
  not gc168 (wc168, n_561);
endmodule

module add_signed_412_2_GENERIC(A, B, Z);
  input [42:0] A, B;
  output [43:0] Z;
  wire [42:0] A, B;
  wire [43:0] Z;
  add_signed_412_2_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_4165_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [60:0] A, B;
  output [61:0] Z;
  wire [60:0] A, B;
  wire [61:0] Z;
  wire n_188, n_189, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367;
  wire n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431;
  wire n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439;
  wire n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447;
  wire n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455;
  wire n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463;
  wire n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492;
  not g3 (Z[61], n_188);
  nand g4 (n_189, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_194, A[1], B[1]);
  nand g13 (n_198, n_194, n_195, n_196);
  xor g14 (n_197, A[1], B[1]);
  nand g16 (n_199, A[2], B[2]);
  nand g17 (n_200, A[2], n_198);
  nand g18 (n_201, B[2], n_198);
  nand g19 (n_203, n_199, n_200, n_201);
  xor g20 (n_202, A[2], B[2]);
  xor g21 (Z[2], n_198, n_202);
  nand g22 (n_204, A[3], B[3]);
  nand g23 (n_205, A[3], n_203);
  nand g24 (n_206, B[3], n_203);
  nand g25 (n_208, n_204, n_205, n_206);
  xor g26 (n_207, A[3], B[3]);
  xor g27 (Z[3], n_203, n_207);
  nand g28 (n_209, A[4], B[4]);
  nand g29 (n_210, A[4], n_208);
  nand g30 (n_211, B[4], n_208);
  nand g31 (n_213, n_209, n_210, n_211);
  xor g32 (n_212, A[4], B[4]);
  xor g33 (Z[4], n_208, n_212);
  nand g34 (n_214, A[5], B[5]);
  nand g35 (n_215, A[5], n_213);
  nand g36 (n_216, B[5], n_213);
  nand g37 (n_218, n_214, n_215, n_216);
  xor g38 (n_217, A[5], B[5]);
  xor g39 (Z[5], n_213, n_217);
  nand g40 (n_219, A[6], B[6]);
  nand g41 (n_220, A[6], n_218);
  nand g42 (n_221, B[6], n_218);
  nand g43 (n_223, n_219, n_220, n_221);
  xor g44 (n_222, A[6], B[6]);
  xor g45 (Z[6], n_218, n_222);
  nand g46 (n_224, A[7], B[7]);
  nand g47 (n_225, A[7], n_223);
  nand g48 (n_226, B[7], n_223);
  nand g49 (n_228, n_224, n_225, n_226);
  xor g50 (n_227, A[7], B[7]);
  xor g51 (Z[7], n_223, n_227);
  nand g52 (n_229, A[8], B[8]);
  nand g53 (n_230, A[8], n_228);
  nand g54 (n_231, B[8], n_228);
  nand g55 (n_233, n_229, n_230, n_231);
  xor g56 (n_232, A[8], B[8]);
  xor g57 (Z[8], n_228, n_232);
  nand g58 (n_234, A[9], B[9]);
  nand g59 (n_235, A[9], n_233);
  nand g60 (n_236, B[9], n_233);
  nand g61 (n_238, n_234, n_235, n_236);
  xor g62 (n_237, A[9], B[9]);
  xor g63 (Z[9], n_233, n_237);
  nand g64 (n_239, A[10], B[10]);
  nand g65 (n_240, A[10], n_238);
  nand g66 (n_241, B[10], n_238);
  nand g67 (n_243, n_239, n_240, n_241);
  xor g68 (n_242, A[10], B[10]);
  xor g69 (Z[10], n_238, n_242);
  nand g70 (n_244, A[11], B[11]);
  nand g71 (n_245, A[11], n_243);
  nand g72 (n_246, B[11], n_243);
  nand g73 (n_248, n_244, n_245, n_246);
  xor g74 (n_247, A[11], B[11]);
  xor g75 (Z[11], n_243, n_247);
  nand g76 (n_249, A[12], B[12]);
  nand g77 (n_250, A[12], n_248);
  nand g78 (n_251, B[12], n_248);
  nand g79 (n_253, n_249, n_250, n_251);
  xor g80 (n_252, A[12], B[12]);
  xor g81 (Z[12], n_248, n_252);
  nand g82 (n_254, A[13], B[13]);
  nand g83 (n_255, A[13], n_253);
  nand g84 (n_256, B[13], n_253);
  nand g85 (n_258, n_254, n_255, n_256);
  xor g86 (n_257, A[13], B[13]);
  xor g87 (Z[13], n_253, n_257);
  nand g88 (n_259, A[14], B[14]);
  nand g89 (n_260, A[14], n_258);
  nand g90 (n_261, B[14], n_258);
  nand g91 (n_263, n_259, n_260, n_261);
  xor g92 (n_262, A[14], B[14]);
  xor g93 (Z[14], n_258, n_262);
  nand g94 (n_264, A[15], B[15]);
  nand g95 (n_265, A[15], n_263);
  nand g96 (n_266, B[15], n_263);
  nand g97 (n_268, n_264, n_265, n_266);
  xor g98 (n_267, A[15], B[15]);
  xor g99 (Z[15], n_263, n_267);
  nand g100 (n_269, A[16], B[16]);
  nand g101 (n_270, A[16], n_268);
  nand g102 (n_271, B[16], n_268);
  nand g103 (n_273, n_269, n_270, n_271);
  xor g104 (n_272, A[16], B[16]);
  xor g105 (Z[16], n_268, n_272);
  nand g106 (n_274, A[17], B[17]);
  nand g107 (n_275, A[17], n_273);
  nand g108 (n_276, B[17], n_273);
  nand g109 (n_278, n_274, n_275, n_276);
  xor g110 (n_277, A[17], B[17]);
  xor g111 (Z[17], n_273, n_277);
  nand g112 (n_279, A[18], B[18]);
  nand g113 (n_280, A[18], n_278);
  nand g114 (n_281, B[18], n_278);
  nand g115 (n_283, n_279, n_280, n_281);
  xor g116 (n_282, A[18], B[18]);
  xor g117 (Z[18], n_278, n_282);
  nand g118 (n_284, A[19], B[19]);
  nand g119 (n_285, A[19], n_283);
  nand g120 (n_286, B[19], n_283);
  nand g121 (n_288, n_284, n_285, n_286);
  xor g122 (n_287, A[19], B[19]);
  xor g123 (Z[19], n_283, n_287);
  nand g124 (n_289, A[20], B[20]);
  nand g125 (n_290, A[20], n_288);
  nand g126 (n_291, B[20], n_288);
  nand g127 (n_293, n_289, n_290, n_291);
  xor g128 (n_292, A[20], B[20]);
  xor g129 (Z[20], n_288, n_292);
  nand g130 (n_294, A[21], B[21]);
  nand g131 (n_295, A[21], n_293);
  nand g132 (n_296, B[21], n_293);
  nand g133 (n_298, n_294, n_295, n_296);
  xor g134 (n_297, A[21], B[21]);
  xor g135 (Z[21], n_293, n_297);
  nand g136 (n_299, A[22], B[22]);
  nand g137 (n_300, A[22], n_298);
  nand g138 (n_301, B[22], n_298);
  nand g139 (n_303, n_299, n_300, n_301);
  xor g140 (n_302, A[22], B[22]);
  xor g141 (Z[22], n_298, n_302);
  nand g142 (n_304, A[23], B[23]);
  nand g143 (n_305, A[23], n_303);
  nand g144 (n_306, B[23], n_303);
  nand g145 (n_308, n_304, n_305, n_306);
  xor g146 (n_307, A[23], B[23]);
  xor g147 (Z[23], n_303, n_307);
  nand g148 (n_309, A[24], B[24]);
  nand g149 (n_310, A[24], n_308);
  nand g150 (n_311, B[24], n_308);
  nand g151 (n_313, n_309, n_310, n_311);
  xor g152 (n_312, A[24], B[24]);
  xor g153 (Z[24], n_308, n_312);
  nand g154 (n_314, A[25], B[25]);
  nand g155 (n_315, A[25], n_313);
  nand g156 (n_316, B[25], n_313);
  nand g157 (n_318, n_314, n_315, n_316);
  xor g158 (n_317, A[25], B[25]);
  xor g159 (Z[25], n_313, n_317);
  nand g160 (n_319, A[26], B[26]);
  nand g161 (n_320, A[26], n_318);
  nand g162 (n_321, B[26], n_318);
  nand g163 (n_323, n_319, n_320, n_321);
  xor g164 (n_322, A[26], B[26]);
  xor g165 (Z[26], n_318, n_322);
  nand g166 (n_324, A[27], B[27]);
  nand g167 (n_325, A[27], n_323);
  nand g168 (n_326, B[27], n_323);
  nand g169 (n_328, n_324, n_325, n_326);
  xor g170 (n_327, A[27], B[27]);
  xor g171 (Z[27], n_323, n_327);
  nand g172 (n_329, A[28], B[28]);
  nand g173 (n_330, A[28], n_328);
  nand g174 (n_331, B[28], n_328);
  nand g175 (n_333, n_329, n_330, n_331);
  xor g176 (n_332, A[28], B[28]);
  xor g177 (Z[28], n_328, n_332);
  nand g178 (n_334, A[29], B[29]);
  nand g179 (n_335, A[29], n_333);
  nand g180 (n_336, B[29], n_333);
  nand g181 (n_338, n_334, n_335, n_336);
  xor g182 (n_337, A[29], B[29]);
  xor g183 (Z[29], n_333, n_337);
  nand g184 (n_339, A[30], B[30]);
  nand g185 (n_340, A[30], n_338);
  nand g186 (n_341, B[30], n_338);
  nand g187 (n_343, n_339, n_340, n_341);
  xor g188 (n_342, A[30], B[30]);
  xor g189 (Z[30], n_338, n_342);
  nand g190 (n_344, A[31], B[31]);
  nand g191 (n_345, A[31], n_343);
  nand g192 (n_346, B[31], n_343);
  nand g193 (n_348, n_344, n_345, n_346);
  xor g194 (n_347, A[31], B[31]);
  xor g195 (Z[31], n_343, n_347);
  nand g196 (n_349, A[32], B[32]);
  nand g197 (n_350, A[32], n_348);
  nand g198 (n_351, B[32], n_348);
  nand g199 (n_353, n_349, n_350, n_351);
  xor g200 (n_352, A[32], B[32]);
  xor g201 (Z[32], n_348, n_352);
  nand g202 (n_354, A[33], B[33]);
  nand g203 (n_355, A[33], n_353);
  nand g204 (n_356, B[33], n_353);
  nand g205 (n_358, n_354, n_355, n_356);
  xor g206 (n_357, A[33], B[33]);
  xor g207 (Z[33], n_353, n_357);
  nand g208 (n_359, A[34], B[34]);
  nand g209 (n_360, A[34], n_358);
  nand g210 (n_361, B[34], n_358);
  nand g211 (n_363, n_359, n_360, n_361);
  xor g212 (n_362, A[34], B[34]);
  xor g213 (Z[34], n_358, n_362);
  nand g214 (n_364, A[35], B[35]);
  nand g215 (n_365, A[35], n_363);
  nand g216 (n_366, B[35], n_363);
  nand g217 (n_368, n_364, n_365, n_366);
  xor g218 (n_367, A[35], B[35]);
  xor g219 (Z[35], n_363, n_367);
  nand g220 (n_369, A[36], B[36]);
  nand g221 (n_370, A[36], n_368);
  nand g222 (n_371, B[36], n_368);
  nand g223 (n_373, n_369, n_370, n_371);
  xor g224 (n_372, A[36], B[36]);
  xor g225 (Z[36], n_368, n_372);
  nand g226 (n_374, A[37], B[37]);
  nand g227 (n_375, A[37], n_373);
  nand g228 (n_376, B[37], n_373);
  nand g229 (n_378, n_374, n_375, n_376);
  xor g230 (n_377, A[37], B[37]);
  xor g231 (Z[37], n_373, n_377);
  nand g232 (n_379, A[38], B[38]);
  nand g233 (n_380, A[38], n_378);
  nand g234 (n_381, B[38], n_378);
  nand g235 (n_383, n_379, n_380, n_381);
  xor g236 (n_382, A[38], B[38]);
  xor g237 (Z[38], n_378, n_382);
  nand g238 (n_384, A[39], B[39]);
  nand g239 (n_385, A[39], n_383);
  nand g240 (n_386, B[39], n_383);
  nand g241 (n_388, n_384, n_385, n_386);
  xor g242 (n_387, A[39], B[39]);
  xor g243 (Z[39], n_383, n_387);
  nand g244 (n_389, A[40], B[40]);
  nand g245 (n_390, A[40], n_388);
  nand g246 (n_391, B[40], n_388);
  nand g247 (n_393, n_389, n_390, n_391);
  xor g248 (n_392, A[40], B[40]);
  xor g249 (Z[40], n_388, n_392);
  nand g250 (n_394, A[41], B[41]);
  nand g251 (n_395, A[41], n_393);
  nand g252 (n_396, B[41], n_393);
  nand g253 (n_398, n_394, n_395, n_396);
  xor g254 (n_397, A[41], B[41]);
  xor g255 (Z[41], n_393, n_397);
  nand g256 (n_399, A[42], B[42]);
  nand g257 (n_400, A[42], n_398);
  nand g258 (n_401, B[42], n_398);
  nand g259 (n_403, n_399, n_400, n_401);
  xor g260 (n_402, A[42], B[42]);
  xor g261 (Z[42], n_398, n_402);
  nand g262 (n_404, A[43], B[43]);
  nand g263 (n_405, A[43], n_403);
  nand g264 (n_406, B[43], n_403);
  nand g265 (n_408, n_404, n_405, n_406);
  xor g266 (n_407, A[43], B[43]);
  xor g267 (Z[43], n_403, n_407);
  nand g268 (n_409, A[44], B[44]);
  nand g269 (n_410, A[44], n_408);
  nand g270 (n_411, B[44], n_408);
  nand g271 (n_413, n_409, n_410, n_411);
  xor g272 (n_412, A[44], B[44]);
  xor g273 (Z[44], n_408, n_412);
  nand g274 (n_414, A[45], B[45]);
  nand g275 (n_415, A[45], n_413);
  nand g276 (n_416, B[45], n_413);
  nand g277 (n_418, n_414, n_415, n_416);
  xor g278 (n_417, A[45], B[45]);
  xor g279 (Z[45], n_413, n_417);
  nand g280 (n_419, A[46], B[46]);
  nand g281 (n_420, A[46], n_418);
  nand g282 (n_421, B[46], n_418);
  nand g283 (n_423, n_419, n_420, n_421);
  xor g284 (n_422, A[46], B[46]);
  xor g285 (Z[46], n_418, n_422);
  nand g286 (n_424, A[47], B[47]);
  nand g287 (n_425, A[47], n_423);
  nand g288 (n_426, B[47], n_423);
  nand g289 (n_428, n_424, n_425, n_426);
  xor g290 (n_427, A[47], B[47]);
  xor g291 (Z[47], n_423, n_427);
  nand g292 (n_429, A[48], B[48]);
  nand g293 (n_430, A[48], n_428);
  nand g294 (n_431, B[48], n_428);
  nand g295 (n_433, n_429, n_430, n_431);
  xor g296 (n_432, A[48], B[48]);
  xor g297 (Z[48], n_428, n_432);
  nand g298 (n_434, A[49], B[49]);
  nand g299 (n_435, A[49], n_433);
  nand g300 (n_436, B[49], n_433);
  nand g301 (n_438, n_434, n_435, n_436);
  xor g302 (n_437, A[49], B[49]);
  xor g303 (Z[49], n_433, n_437);
  nand g304 (n_439, A[50], B[50]);
  nand g305 (n_440, A[50], n_438);
  nand g306 (n_441, B[50], n_438);
  nand g307 (n_443, n_439, n_440, n_441);
  xor g308 (n_442, A[50], B[50]);
  xor g309 (Z[50], n_438, n_442);
  nand g310 (n_444, A[51], B[51]);
  nand g311 (n_445, A[51], n_443);
  nand g312 (n_446, B[51], n_443);
  nand g313 (n_448, n_444, n_445, n_446);
  xor g314 (n_447, A[51], B[51]);
  xor g315 (Z[51], n_443, n_447);
  nand g316 (n_449, A[52], B[52]);
  nand g317 (n_450, A[52], n_448);
  nand g318 (n_451, B[52], n_448);
  nand g319 (n_453, n_449, n_450, n_451);
  xor g320 (n_452, A[52], B[52]);
  xor g321 (Z[52], n_448, n_452);
  nand g322 (n_454, A[53], B[53]);
  nand g323 (n_455, A[53], n_453);
  nand g324 (n_456, B[53], n_453);
  nand g325 (n_458, n_454, n_455, n_456);
  xor g326 (n_457, A[53], B[53]);
  xor g327 (Z[53], n_453, n_457);
  nand g328 (n_459, A[54], B[54]);
  nand g329 (n_460, A[54], n_458);
  nand g330 (n_461, B[54], n_458);
  nand g331 (n_463, n_459, n_460, n_461);
  xor g332 (n_462, A[54], B[54]);
  xor g333 (Z[54], n_458, n_462);
  nand g334 (n_464, A[55], B[55]);
  nand g335 (n_465, A[55], n_463);
  nand g336 (n_466, B[55], n_463);
  nand g337 (n_468, n_464, n_465, n_466);
  xor g338 (n_467, A[55], B[55]);
  xor g339 (Z[55], n_463, n_467);
  nand g340 (n_469, A[56], B[56]);
  nand g341 (n_470, A[56], n_468);
  nand g342 (n_471, B[56], n_468);
  nand g343 (n_473, n_469, n_470, n_471);
  xor g344 (n_472, A[56], B[56]);
  xor g345 (Z[56], n_468, n_472);
  nand g346 (n_474, A[57], B[57]);
  nand g347 (n_475, A[57], n_473);
  nand g348 (n_476, B[57], n_473);
  nand g349 (n_478, n_474, n_475, n_476);
  xor g350 (n_477, A[57], B[57]);
  xor g351 (Z[57], n_473, n_477);
  nand g352 (n_479, A[58], B[58]);
  nand g353 (n_480, A[58], n_478);
  nand g354 (n_481, B[58], n_478);
  nand g355 (n_483, n_479, n_480, n_481);
  xor g356 (n_482, A[58], B[58]);
  xor g357 (Z[58], n_478, n_482);
  nand g358 (n_484, A[59], B[59]);
  nand g359 (n_485, A[59], n_483);
  nand g360 (n_486, B[59], n_483);
  nand g361 (n_488, n_484, n_485, n_486);
  xor g362 (n_487, A[59], B[59]);
  xor g363 (Z[59], n_483, n_487);
  nand g367 (n_188, n_489, n_490, n_491);
  xor g369 (Z[60], n_488, n_492);
  or g371 (n_489, A[60], B[60]);
  xor g372 (n_492, A[60], B[60]);
  or g373 (n_195, wc, n_189);
  not gc (wc, A[1]);
  or g374 (n_196, wc0, n_189);
  not gc0 (wc0, B[1]);
  xnor g375 (Z[1], n_189, n_197);
  or g376 (n_490, A[60], wc1);
  not gc1 (wc1, n_488);
  or g377 (n_491, B[60], wc2);
  not gc2 (wc2, n_488);
endmodule

module add_signed_4165_GENERIC(A, B, Z);
  input [60:0] A, B;
  output [61:0] Z;
  wire [60:0] A, B;
  wire [61:0] Z;
  add_signed_4165_GENERIC_REAL g1(.A ({A[60:2], A[0], A[0]}), .B (B),
       .Z (Z));
endmodule

module add_signed_4165_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [60:0] A, B;
  output [61:0] Z;
  wire [60:0] A, B;
  wire [61:0] Z;
  wire n_188, n_189, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367;
  wire n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431;
  wire n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439;
  wire n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447;
  wire n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455;
  wire n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463;
  wire n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492;
  not g3 (Z[61], n_188);
  nand g4 (n_189, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_194, A[1], B[1]);
  nand g13 (n_198, n_194, n_195, n_196);
  xor g14 (n_197, A[1], B[1]);
  nand g16 (n_199, A[2], B[2]);
  nand g17 (n_200, A[2], n_198);
  nand g18 (n_201, B[2], n_198);
  nand g19 (n_203, n_199, n_200, n_201);
  xor g20 (n_202, A[2], B[2]);
  xor g21 (Z[2], n_198, n_202);
  nand g22 (n_204, A[3], B[3]);
  nand g23 (n_205, A[3], n_203);
  nand g24 (n_206, B[3], n_203);
  nand g25 (n_208, n_204, n_205, n_206);
  xor g26 (n_207, A[3], B[3]);
  xor g27 (Z[3], n_203, n_207);
  nand g28 (n_209, A[4], B[4]);
  nand g29 (n_210, A[4], n_208);
  nand g30 (n_211, B[4], n_208);
  nand g31 (n_213, n_209, n_210, n_211);
  xor g32 (n_212, A[4], B[4]);
  xor g33 (Z[4], n_208, n_212);
  nand g34 (n_214, A[5], B[5]);
  nand g35 (n_215, A[5], n_213);
  nand g36 (n_216, B[5], n_213);
  nand g37 (n_218, n_214, n_215, n_216);
  xor g38 (n_217, A[5], B[5]);
  xor g39 (Z[5], n_213, n_217);
  nand g40 (n_219, A[6], B[6]);
  nand g41 (n_220, A[6], n_218);
  nand g42 (n_221, B[6], n_218);
  nand g43 (n_223, n_219, n_220, n_221);
  xor g44 (n_222, A[6], B[6]);
  xor g45 (Z[6], n_218, n_222);
  nand g46 (n_224, A[7], B[7]);
  nand g47 (n_225, A[7], n_223);
  nand g48 (n_226, B[7], n_223);
  nand g49 (n_228, n_224, n_225, n_226);
  xor g50 (n_227, A[7], B[7]);
  xor g51 (Z[7], n_223, n_227);
  nand g52 (n_229, A[8], B[8]);
  nand g53 (n_230, A[8], n_228);
  nand g54 (n_231, B[8], n_228);
  nand g55 (n_233, n_229, n_230, n_231);
  xor g56 (n_232, A[8], B[8]);
  xor g57 (Z[8], n_228, n_232);
  nand g58 (n_234, A[9], B[9]);
  nand g59 (n_235, A[9], n_233);
  nand g60 (n_236, B[9], n_233);
  nand g61 (n_238, n_234, n_235, n_236);
  xor g62 (n_237, A[9], B[9]);
  xor g63 (Z[9], n_233, n_237);
  nand g64 (n_239, A[10], B[10]);
  nand g65 (n_240, A[10], n_238);
  nand g66 (n_241, B[10], n_238);
  nand g67 (n_243, n_239, n_240, n_241);
  xor g68 (n_242, A[10], B[10]);
  xor g69 (Z[10], n_238, n_242);
  nand g70 (n_244, A[11], B[11]);
  nand g71 (n_245, A[11], n_243);
  nand g72 (n_246, B[11], n_243);
  nand g73 (n_248, n_244, n_245, n_246);
  xor g74 (n_247, A[11], B[11]);
  xor g75 (Z[11], n_243, n_247);
  nand g76 (n_249, A[12], B[12]);
  nand g77 (n_250, A[12], n_248);
  nand g78 (n_251, B[12], n_248);
  nand g79 (n_253, n_249, n_250, n_251);
  xor g80 (n_252, A[12], B[12]);
  xor g81 (Z[12], n_248, n_252);
  nand g82 (n_254, A[13], B[13]);
  nand g83 (n_255, A[13], n_253);
  nand g84 (n_256, B[13], n_253);
  nand g85 (n_258, n_254, n_255, n_256);
  xor g86 (n_257, A[13], B[13]);
  xor g87 (Z[13], n_253, n_257);
  nand g88 (n_259, A[14], B[14]);
  nand g89 (n_260, A[14], n_258);
  nand g90 (n_261, B[14], n_258);
  nand g91 (n_263, n_259, n_260, n_261);
  xor g92 (n_262, A[14], B[14]);
  xor g93 (Z[14], n_258, n_262);
  nand g94 (n_264, A[15], B[15]);
  nand g95 (n_265, A[15], n_263);
  nand g96 (n_266, B[15], n_263);
  nand g97 (n_268, n_264, n_265, n_266);
  xor g98 (n_267, A[15], B[15]);
  xor g99 (Z[15], n_263, n_267);
  nand g100 (n_269, A[16], B[16]);
  nand g101 (n_270, A[16], n_268);
  nand g102 (n_271, B[16], n_268);
  nand g103 (n_273, n_269, n_270, n_271);
  xor g104 (n_272, A[16], B[16]);
  xor g105 (Z[16], n_268, n_272);
  nand g106 (n_274, A[17], B[17]);
  nand g107 (n_275, A[17], n_273);
  nand g108 (n_276, B[17], n_273);
  nand g109 (n_278, n_274, n_275, n_276);
  xor g110 (n_277, A[17], B[17]);
  xor g111 (Z[17], n_273, n_277);
  nand g112 (n_279, A[18], B[18]);
  nand g113 (n_280, A[18], n_278);
  nand g114 (n_281, B[18], n_278);
  nand g115 (n_283, n_279, n_280, n_281);
  xor g116 (n_282, A[18], B[18]);
  xor g117 (Z[18], n_278, n_282);
  nand g118 (n_284, A[19], B[19]);
  nand g119 (n_285, A[19], n_283);
  nand g120 (n_286, B[19], n_283);
  nand g121 (n_288, n_284, n_285, n_286);
  xor g122 (n_287, A[19], B[19]);
  xor g123 (Z[19], n_283, n_287);
  nand g124 (n_289, A[20], B[20]);
  nand g125 (n_290, A[20], n_288);
  nand g126 (n_291, B[20], n_288);
  nand g127 (n_293, n_289, n_290, n_291);
  xor g128 (n_292, A[20], B[20]);
  xor g129 (Z[20], n_288, n_292);
  nand g130 (n_294, A[21], B[21]);
  nand g131 (n_295, A[21], n_293);
  nand g132 (n_296, B[21], n_293);
  nand g133 (n_298, n_294, n_295, n_296);
  xor g134 (n_297, A[21], B[21]);
  xor g135 (Z[21], n_293, n_297);
  nand g136 (n_299, A[22], B[22]);
  nand g137 (n_300, A[22], n_298);
  nand g138 (n_301, B[22], n_298);
  nand g139 (n_303, n_299, n_300, n_301);
  xor g140 (n_302, A[22], B[22]);
  xor g141 (Z[22], n_298, n_302);
  nand g142 (n_304, A[23], B[23]);
  nand g143 (n_305, A[23], n_303);
  nand g144 (n_306, B[23], n_303);
  nand g145 (n_308, n_304, n_305, n_306);
  xor g146 (n_307, A[23], B[23]);
  xor g147 (Z[23], n_303, n_307);
  nand g148 (n_309, A[24], B[24]);
  nand g149 (n_310, A[24], n_308);
  nand g150 (n_311, B[24], n_308);
  nand g151 (n_313, n_309, n_310, n_311);
  xor g152 (n_312, A[24], B[24]);
  xor g153 (Z[24], n_308, n_312);
  nand g154 (n_314, A[25], B[25]);
  nand g155 (n_315, A[25], n_313);
  nand g156 (n_316, B[25], n_313);
  nand g157 (n_318, n_314, n_315, n_316);
  xor g158 (n_317, A[25], B[25]);
  xor g159 (Z[25], n_313, n_317);
  nand g160 (n_319, A[26], B[26]);
  nand g161 (n_320, A[26], n_318);
  nand g162 (n_321, B[26], n_318);
  nand g163 (n_323, n_319, n_320, n_321);
  xor g164 (n_322, A[26], B[26]);
  xor g165 (Z[26], n_318, n_322);
  nand g166 (n_324, A[27], B[27]);
  nand g167 (n_325, A[27], n_323);
  nand g168 (n_326, B[27], n_323);
  nand g169 (n_328, n_324, n_325, n_326);
  xor g170 (n_327, A[27], B[27]);
  xor g171 (Z[27], n_323, n_327);
  nand g172 (n_329, A[28], B[28]);
  nand g173 (n_330, A[28], n_328);
  nand g174 (n_331, B[28], n_328);
  nand g175 (n_333, n_329, n_330, n_331);
  xor g176 (n_332, A[28], B[28]);
  xor g177 (Z[28], n_328, n_332);
  nand g178 (n_334, A[29], B[29]);
  nand g179 (n_335, A[29], n_333);
  nand g180 (n_336, B[29], n_333);
  nand g181 (n_338, n_334, n_335, n_336);
  xor g182 (n_337, A[29], B[29]);
  xor g183 (Z[29], n_333, n_337);
  nand g184 (n_339, A[30], B[30]);
  nand g185 (n_340, A[30], n_338);
  nand g186 (n_341, B[30], n_338);
  nand g187 (n_343, n_339, n_340, n_341);
  xor g188 (n_342, A[30], B[30]);
  xor g189 (Z[30], n_338, n_342);
  nand g190 (n_344, A[31], B[31]);
  nand g191 (n_345, A[31], n_343);
  nand g192 (n_346, B[31], n_343);
  nand g193 (n_348, n_344, n_345, n_346);
  xor g194 (n_347, A[31], B[31]);
  xor g195 (Z[31], n_343, n_347);
  nand g196 (n_349, A[32], B[32]);
  nand g197 (n_350, A[32], n_348);
  nand g198 (n_351, B[32], n_348);
  nand g199 (n_353, n_349, n_350, n_351);
  xor g200 (n_352, A[32], B[32]);
  xor g201 (Z[32], n_348, n_352);
  nand g202 (n_354, A[33], B[33]);
  nand g203 (n_355, A[33], n_353);
  nand g204 (n_356, B[33], n_353);
  nand g205 (n_358, n_354, n_355, n_356);
  xor g206 (n_357, A[33], B[33]);
  xor g207 (Z[33], n_353, n_357);
  nand g208 (n_359, A[34], B[34]);
  nand g209 (n_360, A[34], n_358);
  nand g210 (n_361, B[34], n_358);
  nand g211 (n_363, n_359, n_360, n_361);
  xor g212 (n_362, A[34], B[34]);
  xor g213 (Z[34], n_358, n_362);
  nand g214 (n_364, A[35], B[35]);
  nand g215 (n_365, A[35], n_363);
  nand g216 (n_366, B[35], n_363);
  nand g217 (n_368, n_364, n_365, n_366);
  xor g218 (n_367, A[35], B[35]);
  xor g219 (Z[35], n_363, n_367);
  nand g220 (n_369, A[36], B[36]);
  nand g221 (n_370, A[36], n_368);
  nand g222 (n_371, B[36], n_368);
  nand g223 (n_373, n_369, n_370, n_371);
  xor g224 (n_372, A[36], B[36]);
  xor g225 (Z[36], n_368, n_372);
  nand g226 (n_374, A[37], B[37]);
  nand g227 (n_375, A[37], n_373);
  nand g228 (n_376, B[37], n_373);
  nand g229 (n_378, n_374, n_375, n_376);
  xor g230 (n_377, A[37], B[37]);
  xor g231 (Z[37], n_373, n_377);
  nand g232 (n_379, A[38], B[38]);
  nand g233 (n_380, A[38], n_378);
  nand g234 (n_381, B[38], n_378);
  nand g235 (n_383, n_379, n_380, n_381);
  xor g236 (n_382, A[38], B[38]);
  xor g237 (Z[38], n_378, n_382);
  nand g238 (n_384, A[39], B[39]);
  nand g239 (n_385, A[39], n_383);
  nand g240 (n_386, B[39], n_383);
  nand g241 (n_388, n_384, n_385, n_386);
  xor g242 (n_387, A[39], B[39]);
  xor g243 (Z[39], n_383, n_387);
  nand g244 (n_389, A[40], B[40]);
  nand g245 (n_390, A[40], n_388);
  nand g246 (n_391, B[40], n_388);
  nand g247 (n_393, n_389, n_390, n_391);
  xor g248 (n_392, A[40], B[40]);
  xor g249 (Z[40], n_388, n_392);
  nand g250 (n_394, A[41], B[41]);
  nand g251 (n_395, A[41], n_393);
  nand g252 (n_396, B[41], n_393);
  nand g253 (n_398, n_394, n_395, n_396);
  xor g254 (n_397, A[41], B[41]);
  xor g255 (Z[41], n_393, n_397);
  nand g256 (n_399, A[42], B[42]);
  nand g257 (n_400, A[42], n_398);
  nand g258 (n_401, B[42], n_398);
  nand g259 (n_403, n_399, n_400, n_401);
  xor g260 (n_402, A[42], B[42]);
  xor g261 (Z[42], n_398, n_402);
  nand g262 (n_404, A[43], B[43]);
  nand g263 (n_405, A[43], n_403);
  nand g264 (n_406, B[43], n_403);
  nand g265 (n_408, n_404, n_405, n_406);
  xor g266 (n_407, A[43], B[43]);
  xor g267 (Z[43], n_403, n_407);
  nand g268 (n_409, A[44], B[44]);
  nand g269 (n_410, A[44], n_408);
  nand g270 (n_411, B[44], n_408);
  nand g271 (n_413, n_409, n_410, n_411);
  xor g272 (n_412, A[44], B[44]);
  xor g273 (Z[44], n_408, n_412);
  nand g274 (n_414, A[45], B[45]);
  nand g275 (n_415, A[45], n_413);
  nand g276 (n_416, B[45], n_413);
  nand g277 (n_418, n_414, n_415, n_416);
  xor g278 (n_417, A[45], B[45]);
  xor g279 (Z[45], n_413, n_417);
  nand g280 (n_419, A[46], B[46]);
  nand g281 (n_420, A[46], n_418);
  nand g282 (n_421, B[46], n_418);
  nand g283 (n_423, n_419, n_420, n_421);
  xor g284 (n_422, A[46], B[46]);
  xor g285 (Z[46], n_418, n_422);
  nand g286 (n_424, A[47], B[47]);
  nand g287 (n_425, A[47], n_423);
  nand g288 (n_426, B[47], n_423);
  nand g289 (n_428, n_424, n_425, n_426);
  xor g290 (n_427, A[47], B[47]);
  xor g291 (Z[47], n_423, n_427);
  nand g292 (n_429, A[48], B[48]);
  nand g293 (n_430, A[48], n_428);
  nand g294 (n_431, B[48], n_428);
  nand g295 (n_433, n_429, n_430, n_431);
  xor g296 (n_432, A[48], B[48]);
  xor g297 (Z[48], n_428, n_432);
  nand g298 (n_434, A[49], B[49]);
  nand g299 (n_435, A[49], n_433);
  nand g300 (n_436, B[49], n_433);
  nand g301 (n_438, n_434, n_435, n_436);
  xor g302 (n_437, A[49], B[49]);
  xor g303 (Z[49], n_433, n_437);
  nand g304 (n_439, A[50], B[50]);
  nand g305 (n_440, A[50], n_438);
  nand g306 (n_441, B[50], n_438);
  nand g307 (n_443, n_439, n_440, n_441);
  xor g308 (n_442, A[50], B[50]);
  xor g309 (Z[50], n_438, n_442);
  nand g310 (n_444, A[51], B[51]);
  nand g311 (n_445, A[51], n_443);
  nand g312 (n_446, B[51], n_443);
  nand g313 (n_448, n_444, n_445, n_446);
  xor g314 (n_447, A[51], B[51]);
  xor g315 (Z[51], n_443, n_447);
  nand g316 (n_449, A[52], B[52]);
  nand g317 (n_450, A[52], n_448);
  nand g318 (n_451, B[52], n_448);
  nand g319 (n_453, n_449, n_450, n_451);
  xor g320 (n_452, A[52], B[52]);
  xor g321 (Z[52], n_448, n_452);
  nand g322 (n_454, A[53], B[53]);
  nand g323 (n_455, A[53], n_453);
  nand g324 (n_456, B[53], n_453);
  nand g325 (n_458, n_454, n_455, n_456);
  xor g326 (n_457, A[53], B[53]);
  xor g327 (Z[53], n_453, n_457);
  nand g328 (n_459, A[54], B[54]);
  nand g329 (n_460, A[54], n_458);
  nand g330 (n_461, B[54], n_458);
  nand g331 (n_463, n_459, n_460, n_461);
  xor g332 (n_462, A[54], B[54]);
  xor g333 (Z[54], n_458, n_462);
  nand g334 (n_464, A[55], B[55]);
  nand g335 (n_465, A[55], n_463);
  nand g336 (n_466, B[55], n_463);
  nand g337 (n_468, n_464, n_465, n_466);
  xor g338 (n_467, A[55], B[55]);
  xor g339 (Z[55], n_463, n_467);
  nand g340 (n_469, A[56], B[56]);
  nand g341 (n_470, A[56], n_468);
  nand g342 (n_471, B[56], n_468);
  nand g343 (n_473, n_469, n_470, n_471);
  xor g344 (n_472, A[56], B[56]);
  xor g345 (Z[56], n_468, n_472);
  nand g346 (n_474, A[57], B[57]);
  nand g347 (n_475, A[57], n_473);
  nand g348 (n_476, B[57], n_473);
  nand g349 (n_478, n_474, n_475, n_476);
  xor g350 (n_477, A[57], B[57]);
  xor g351 (Z[57], n_473, n_477);
  nand g352 (n_479, A[58], B[58]);
  nand g353 (n_480, A[58], n_478);
  nand g354 (n_481, B[58], n_478);
  nand g355 (n_483, n_479, n_480, n_481);
  xor g356 (n_482, A[58], B[58]);
  xor g357 (Z[58], n_478, n_482);
  nand g358 (n_484, A[59], B[59]);
  nand g359 (n_485, A[59], n_483);
  nand g360 (n_486, B[59], n_483);
  nand g361 (n_488, n_484, n_485, n_486);
  xor g362 (n_487, A[59], B[59]);
  xor g363 (Z[59], n_483, n_487);
  nand g367 (n_188, n_489, n_490, n_491);
  xor g369 (Z[60], n_488, n_492);
  or g371 (n_489, A[60], B[60]);
  xor g372 (n_492, A[60], B[60]);
  or g373 (n_195, wc, n_189);
  not gc (wc, A[1]);
  or g374 (n_196, wc0, n_189);
  not gc0 (wc0, B[1]);
  xnor g375 (Z[1], n_189, n_197);
  or g376 (n_490, A[60], wc1);
  not gc1 (wc1, n_488);
  or g377 (n_491, B[60], wc2);
  not gc2 (wc2, n_488);
endmodule

module add_signed_4165_1_GENERIC(A, B, Z);
  input [60:0] A, B;
  output [61:0] Z;
  wire [60:0] A, B;
  wire [61:0] Z;
  add_signed_4165_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_426_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [41:0] A, B;
  output [42:0] Z;
  wire [41:0] A, B;
  wire [42:0] Z;
  wire n_131, n_132, n_135, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_145, n_146, n_147, n_148, n_149, n_151, n_152;
  wire n_153, n_154, n_155, n_157, n_158, n_159, n_160, n_161;
  wire n_163, n_164, n_165, n_166, n_167, n_169, n_170, n_171;
  wire n_172, n_173, n_175, n_176, n_177, n_178, n_179, n_181;
  wire n_182, n_183, n_184, n_185, n_187, n_188, n_189, n_190;
  wire n_191, n_193, n_194, n_195, n_196, n_197, n_199, n_200;
  wire n_201, n_202, n_203, n_205, n_206, n_207, n_208, n_209;
  wire n_211, n_212, n_213, n_214, n_215, n_217, n_218, n_219;
  wire n_220, n_221, n_223, n_224, n_225, n_226, n_227, n_229;
  wire n_230, n_231, n_232, n_233, n_235, n_236, n_237, n_238;
  wire n_239, n_241, n_242, n_243, n_244, n_245, n_247, n_248;
  wire n_249, n_250, n_251, n_253, n_254, n_255, n_256, n_257;
  wire n_259, n_260, n_262, n_263, n_264, n_265, n_266, n_267;
  wire n_269, n_271, n_273, n_274, n_276, n_277, n_279, n_281;
  wire n_283, n_284, n_286, n_287, n_289, n_291, n_293, n_294;
  wire n_296, n_297, n_299, n_301, n_303, n_304, n_306, n_307;
  wire n_309, n_311, n_313, n_314, n_316, n_317, n_319, n_321;
  wire n_323, n_324, n_326, n_327, n_329, n_331, n_333, n_334;
  wire n_336, n_337, n_339, n_341, n_343, n_344, n_346, n_347;
  wire n_349, n_351, n_353, n_354, n_356, n_358, n_359, n_360;
  wire n_362, n_363, n_364, n_366, n_367, n_368, n_369, n_371;
  wire n_373, n_375, n_376, n_377, n_379, n_380, n_381, n_383;
  wire n_384, n_386, n_388, n_390, n_391, n_392, n_394, n_395;
  wire n_396, n_398, n_399, n_401, n_403, n_405, n_406, n_407;
  wire n_409, n_410, n_411, n_413, n_414, n_416, n_418, n_420;
  wire n_421, n_422, n_424, n_425, n_426, n_428, n_430, n_431;
  wire n_432, n_434, n_435, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_453, n_456, n_458, n_459, n_460, n_463;
  wire n_466, n_468, n_469, n_471, n_473, n_474, n_476, n_478;
  wire n_479, n_481, n_483, n_484, n_486, n_487, n_489, n_491;
  wire n_493, n_494, n_496, n_498, n_499, n_500, n_502, n_503;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_518, n_519, n_520, n_522;
  wire n_523, n_524, n_526, n_527, n_528, n_530, n_531, n_532;
  wire n_534, n_535, n_536, n_538, n_539, n_540, n_542, n_543;
  wire n_544, n_546, n_547, n_548, n_550, n_551, n_552, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_562, n_563;
  wire n_564, n_565, n_566, n_567, n_568, n_570, n_571, n_572;
  wire n_574, n_575, n_576, n_577, n_579, n_580, n_581, n_583;
  wire n_584, n_585, n_586, n_588, n_589, n_590, n_592, n_593;
  wire n_594, n_595, n_597, n_598, n_600, n_601, n_603, n_604;
  wire n_605, n_606, n_608, n_609, n_610, n_612, n_613, n_614;
  wire n_615, n_617, n_618, n_620, n_621, n_623, n_624, n_625;
  wire n_626, n_628, n_629, n_630, n_631, n_633, n_634, n_635;
  wire n_636, n_638, n_639, n_641, n_642, n_644, n_645, n_646;
  wire n_647, n_649, n_650, n_651, n_653, n_654, n_655, n_656;
  wire n_658, n_659, n_661, n_662, n_664, n_665, n_666, n_667;
  wire n_669, n_670, n_671, n_672, n_674, n_675;
  not g3 (Z[42], n_131);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_132, A[0], B[0]);
  nor g9 (n_135, A[1], B[1]);
  nand g10 (n_138, A[1], B[1]);
  nor g11 (n_145, A[2], B[2]);
  nand g12 (n_140, A[2], B[2]);
  nor g13 (n_141, A[3], B[3]);
  nand g14 (n_142, A[3], B[3]);
  nor g15 (n_151, A[4], B[4]);
  nand g16 (n_146, A[4], B[4]);
  nor g17 (n_147, A[5], B[5]);
  nand g18 (n_148, A[5], B[5]);
  nor g19 (n_157, A[6], B[6]);
  nand g20 (n_152, A[6], B[6]);
  nor g21 (n_153, A[7], B[7]);
  nand g22 (n_154, A[7], B[7]);
  nor g23 (n_163, A[8], B[8]);
  nand g24 (n_158, A[8], B[8]);
  nor g25 (n_159, A[9], B[9]);
  nand g26 (n_160, A[9], B[9]);
  nor g27 (n_169, A[10], B[10]);
  nand g28 (n_164, A[10], B[10]);
  nor g29 (n_165, A[11], B[11]);
  nand g30 (n_166, A[11], B[11]);
  nor g31 (n_175, A[12], B[12]);
  nand g32 (n_170, A[12], B[12]);
  nor g33 (n_171, A[13], B[13]);
  nand g34 (n_172, A[13], B[13]);
  nor g35 (n_181, A[14], B[14]);
  nand g36 (n_176, A[14], B[14]);
  nor g37 (n_177, A[15], B[15]);
  nand g38 (n_178, A[15], B[15]);
  nor g39 (n_187, A[16], B[16]);
  nand g40 (n_182, A[16], B[16]);
  nor g41 (n_183, A[17], B[17]);
  nand g42 (n_184, A[17], B[17]);
  nor g43 (n_193, A[18], B[18]);
  nand g44 (n_188, A[18], B[18]);
  nor g45 (n_189, A[19], B[19]);
  nand g46 (n_190, A[19], B[19]);
  nor g47 (n_199, A[20], B[20]);
  nand g48 (n_194, A[20], B[20]);
  nor g49 (n_195, A[21], B[21]);
  nand g50 (n_196, A[21], B[21]);
  nor g51 (n_205, A[22], B[22]);
  nand g52 (n_200, A[22], B[22]);
  nor g53 (n_201, A[23], B[23]);
  nand g54 (n_202, A[23], B[23]);
  nor g55 (n_211, A[24], B[24]);
  nand g56 (n_206, A[24], B[24]);
  nor g57 (n_207, A[25], B[25]);
  nand g58 (n_208, A[25], B[25]);
  nor g59 (n_217, A[26], B[26]);
  nand g60 (n_212, A[26], B[26]);
  nor g61 (n_213, A[27], B[27]);
  nand g62 (n_214, A[27], B[27]);
  nor g63 (n_223, A[28], B[28]);
  nand g64 (n_218, A[28], B[28]);
  nor g65 (n_219, A[29], B[29]);
  nand g66 (n_220, A[29], B[29]);
  nor g67 (n_229, A[30], B[30]);
  nand g68 (n_224, A[30], B[30]);
  nor g69 (n_225, A[31], B[31]);
  nand g70 (n_226, A[31], B[31]);
  nor g71 (n_235, A[32], B[32]);
  nand g72 (n_230, A[32], B[32]);
  nor g73 (n_231, A[33], B[33]);
  nand g74 (n_232, A[33], B[33]);
  nor g75 (n_241, A[34], B[34]);
  nand g76 (n_236, A[34], B[34]);
  nor g77 (n_237, A[35], B[35]);
  nand g78 (n_238, A[35], B[35]);
  nor g79 (n_247, A[36], B[36]);
  nand g80 (n_242, A[36], B[36]);
  nor g81 (n_243, A[37], B[37]);
  nand g82 (n_244, A[37], B[37]);
  nor g83 (n_253, A[38], B[38]);
  nand g84 (n_248, A[38], B[38]);
  nor g85 (n_249, A[39], B[39]);
  nand g86 (n_250, A[39], B[39]);
  nor g87 (n_259, A[40], B[40]);
  nand g88 (n_254, A[40], B[40]);
  nand g93 (n_260, n_138, n_139);
  nor g94 (n_143, n_140, n_141);
  nor g97 (n_263, n_145, n_141);
  nor g98 (n_149, n_146, n_147);
  nor g101 (n_269, n_151, n_147);
  nor g102 (n_155, n_152, n_153);
  nor g105 (n_271, n_157, n_153);
  nor g106 (n_161, n_158, n_159);
  nor g109 (n_279, n_163, n_159);
  nor g110 (n_167, n_164, n_165);
  nor g113 (n_281, n_169, n_165);
  nor g114 (n_173, n_170, n_171);
  nor g117 (n_289, n_175, n_171);
  nor g118 (n_179, n_176, n_177);
  nor g121 (n_291, n_181, n_177);
  nor g122 (n_185, n_182, n_183);
  nor g125 (n_299, n_187, n_183);
  nor g126 (n_191, n_188, n_189);
  nor g129 (n_301, n_193, n_189);
  nor g130 (n_197, n_194, n_195);
  nor g133 (n_309, n_199, n_195);
  nor g134 (n_203, n_200, n_201);
  nor g137 (n_311, n_205, n_201);
  nor g138 (n_209, n_206, n_207);
  nor g141 (n_319, n_211, n_207);
  nor g142 (n_215, n_212, n_213);
  nor g145 (n_321, n_217, n_213);
  nor g146 (n_221, n_218, n_219);
  nor g149 (n_329, n_223, n_219);
  nor g150 (n_227, n_224, n_225);
  nor g153 (n_331, n_229, n_225);
  nor g154 (n_233, n_230, n_231);
  nor g157 (n_339, n_235, n_231);
  nor g158 (n_239, n_236, n_237);
  nor g161 (n_341, n_241, n_237);
  nor g162 (n_245, n_242, n_243);
  nor g165 (n_349, n_247, n_243);
  nor g166 (n_251, n_248, n_249);
  nor g169 (n_351, n_253, n_249);
  nor g170 (n_257, n_254, n_255);
  nor g173 (n_491, n_259, n_255);
  nand g176 (n_579, n_140, n_262);
  nand g177 (n_265, n_263, n_260);
  nand g178 (n_356, n_264, n_265);
  nor g179 (n_267, n_157, n_266);
  nand g188 (n_364, n_269, n_271);
  nor g189 (n_277, n_169, n_276);
  nand g198 (n_371, n_279, n_281);
  nor g199 (n_287, n_181, n_286);
  nand g208 (n_379, n_289, n_291);
  nor g209 (n_297, n_193, n_296);
  nand g218 (n_386, n_299, n_301);
  nor g219 (n_307, n_205, n_306);
  nand g228 (n_394, n_309, n_311);
  nor g229 (n_317, n_217, n_316);
  nand g238 (n_401, n_319, n_321);
  nor g239 (n_327, n_229, n_326);
  nand g248 (n_409, n_329, n_331);
  nor g249 (n_337, n_241, n_336);
  nand g258 (n_416, n_339, n_341);
  nor g259 (n_347, n_253, n_346);
  nand g268 (n_424, n_349, n_351);
  nand g271 (n_583, n_146, n_358);
  nand g272 (n_359, n_269, n_356);
  nand g273 (n_585, n_266, n_359);
  nand g276 (n_588, n_362, n_363);
  nand g279 (n_428, n_366, n_367);
  nor g280 (n_369, n_175, n_368);
  nor g283 (n_438, n_175, n_371);
  nor g289 (n_377, n_375, n_368);
  nor g292 (n_444, n_371, n_375);
  nor g293 (n_381, n_379, n_368);
  nor g296 (n_447, n_371, n_379);
  nor g297 (n_384, n_199, n_383);
  nor g300 (n_506, n_199, n_386);
  nor g306 (n_392, n_390, n_383);
  nor g309 (n_512, n_386, n_390);
  nor g310 (n_396, n_394, n_383);
  nor g313 (n_453, n_386, n_394);
  nor g314 (n_399, n_223, n_398);
  nor g317 (n_466, n_223, n_401);
  nor g323 (n_407, n_405, n_398);
  nor g326 (n_476, n_401, n_405);
  nor g327 (n_411, n_409, n_398);
  nor g330 (n_481, n_401, n_409);
  nor g331 (n_414, n_247, n_413);
  nor g334 (n_558, n_247, n_416);
  nor g340 (n_422, n_420, n_413);
  nor g343 (n_564, n_416, n_420);
  nor g344 (n_426, n_424, n_413);
  nor g347 (n_489, n_416, n_424);
  nand g350 (n_592, n_158, n_430);
  nand g351 (n_431, n_279, n_428);
  nand g352 (n_594, n_276, n_431);
  nand g355 (n_597, n_434, n_435);
  nand g358 (n_600, n_368, n_437);
  nand g359 (n_440, n_438, n_428);
  nand g360 (n_603, n_439, n_440);
  nand g361 (n_443, n_441, n_428);
  nand g362 (n_605, n_442, n_443);
  nand g363 (n_446, n_444, n_428);
  nand g364 (n_608, n_445, n_446);
  nand g365 (n_449, n_447, n_428);
  nand g366 (n_496, n_448, n_449);
  nor g367 (n_451, n_211, n_450);
  nand g376 (n_520, n_319, n_453);
  nor g377 (n_460, n_458, n_450);
  nor g382 (n_463, n_401, n_450);
  nand g391 (n_532, n_453, n_466);
  nand g396 (n_536, n_453, n_471);
  nand g401 (n_540, n_453, n_476);
  nand g406 (n_544, n_453, n_481);
  nor g407 (n_487, n_259, n_486);
  nand g416 (n_572, n_491, n_489);
  nand g419 (n_612, n_182, n_498);
  nand g420 (n_499, n_299, n_496);
  nand g421 (n_614, n_296, n_499);
  nand g424 (n_617, n_502, n_503);
  nand g427 (n_620, n_383, n_505);
  nand g428 (n_508, n_506, n_496);
  nand g429 (n_623, n_507, n_508);
  nand g430 (n_511, n_509, n_496);
  nand g431 (n_625, n_510, n_511);
  nand g432 (n_514, n_512, n_496);
  nand g433 (n_628, n_513, n_514);
  nand g434 (n_515, n_453, n_496);
  nand g435 (n_630, n_450, n_515);
  nand g438 (n_633, n_518, n_519);
  nand g441 (n_635, n_522, n_523);
  nand g444 (n_638, n_526, n_527);
  nand g447 (n_641, n_530, n_531);
  nand g450 (n_644, n_534, n_535);
  nand g453 (n_646, n_538, n_539);
  nand g456 (n_649, n_542, n_543);
  nand g459 (n_548, n_546, n_547);
  nand g462 (n_653, n_230, n_550);
  nand g463 (n_551, n_339, n_548);
  nand g464 (n_655, n_336, n_551);
  nand g467 (n_658, n_554, n_555);
  nand g470 (n_661, n_413, n_557);
  nand g471 (n_560, n_558, n_548);
  nand g472 (n_664, n_559, n_560);
  nand g473 (n_563, n_561, n_548);
  nand g474 (n_666, n_562, n_563);
  nand g475 (n_566, n_564, n_548);
  nand g476 (n_669, n_565, n_566);
  nand g477 (n_567, n_489, n_548);
  nand g478 (n_671, n_486, n_567);
  nand g481 (n_674, n_570, n_571);
  nand g484 (n_131, n_574, n_575);
  xnor g488 (Z[2], n_260, n_577);
  xnor g491 (Z[3], n_579, n_580);
  xnor g493 (Z[4], n_356, n_581);
  xnor g496 (Z[5], n_583, n_584);
  xnor g498 (Z[6], n_585, n_586);
  xnor g501 (Z[7], n_588, n_589);
  xnor g503 (Z[8], n_428, n_590);
  xnor g506 (Z[9], n_592, n_593);
  xnor g508 (Z[10], n_594, n_595);
  xnor g511 (Z[11], n_597, n_598);
  xnor g514 (Z[12], n_600, n_601);
  xnor g517 (Z[13], n_603, n_604);
  xnor g519 (Z[14], n_605, n_606);
  xnor g522 (Z[15], n_608, n_609);
  xnor g524 (Z[16], n_496, n_610);
  xnor g527 (Z[17], n_612, n_613);
  xnor g529 (Z[18], n_614, n_615);
  xnor g532 (Z[19], n_617, n_618);
  xnor g535 (Z[20], n_620, n_621);
  xnor g538 (Z[21], n_623, n_624);
  xnor g540 (Z[22], n_625, n_626);
  xnor g543 (Z[23], n_628, n_629);
  xnor g545 (Z[24], n_630, n_631);
  xnor g548 (Z[25], n_633, n_634);
  xnor g550 (Z[26], n_635, n_636);
  xnor g553 (Z[27], n_638, n_639);
  xnor g556 (Z[28], n_641, n_642);
  xnor g559 (Z[29], n_644, n_645);
  xnor g561 (Z[30], n_646, n_647);
  xnor g564 (Z[31], n_649, n_650);
  xnor g566 (Z[32], n_548, n_651);
  xnor g569 (Z[33], n_653, n_654);
  xnor g571 (Z[34], n_655, n_656);
  xnor g574 (Z[35], n_658, n_659);
  xnor g577 (Z[36], n_661, n_662);
  xnor g580 (Z[37], n_664, n_665);
  xnor g582 (Z[38], n_666, n_667);
  xnor g585 (Z[39], n_669, n_670);
  xnor g587 (Z[40], n_671, n_672);
  xnor g590 (Z[41], n_674, n_675);
  and g593 (n_255, A[41], B[41]);
  or g594 (n_256, A[41], B[41]);
  and g595 (n_336, wc, n_232);
  not gc (wc, n_233);
  and g596 (n_343, wc0, n_238);
  not gc0 (wc0, n_239);
  and g597 (n_346, wc1, n_244);
  not gc1 (wc1, n_245);
  and g598 (n_353, wc2, n_250);
  not gc2 (wc2, n_251);
  and g599 (n_296, wc3, n_184);
  not gc3 (wc3, n_185);
  and g600 (n_303, wc4, n_190);
  not gc4 (wc4, n_191);
  and g601 (n_306, wc5, n_196);
  not gc5 (wc5, n_197);
  and g602 (n_313, wc6, n_202);
  not gc6 (wc6, n_203);
  and g603 (n_316, wc7, n_208);
  not gc7 (wc7, n_209);
  and g604 (n_323, wc8, n_214);
  not gc8 (wc8, n_215);
  and g605 (n_326, wc9, n_220);
  not gc9 (wc9, n_221);
  and g606 (n_333, wc10, n_226);
  not gc10 (wc10, n_227);
  and g607 (n_276, wc11, n_160);
  not gc11 (wc11, n_161);
  and g608 (n_283, wc12, n_166);
  not gc12 (wc12, n_167);
  and g609 (n_286, wc13, n_172);
  not gc13 (wc13, n_173);
  and g610 (n_293, wc14, n_178);
  not gc14 (wc14, n_179);
  and g611 (n_266, wc15, n_148);
  not gc15 (wc15, n_149);
  and g612 (n_273, wc16, n_154);
  not gc16 (wc16, n_155);
  and g613 (n_264, wc17, n_142);
  not gc17 (wc17, n_143);
  or g614 (n_139, n_132, n_135);
  or g615 (n_360, wc18, n_157);
  not gc18 (wc18, n_269);
  or g616 (n_432, wc19, n_169);
  not gc19 (wc19, n_279);
  or g617 (n_375, wc20, n_181);
  not gc20 (wc20, n_289);
  or g618 (n_500, wc21, n_193);
  not gc21 (wc21, n_299);
  or g619 (n_390, wc22, n_205);
  not gc22 (wc22, n_309);
  or g620 (n_458, wc23, n_217);
  not gc23 (wc23, n_319);
  or g621 (n_405, wc24, n_229);
  not gc24 (wc24, n_329);
  or g622 (n_552, wc25, n_241);
  not gc25 (wc25, n_339);
  or g623 (n_420, wc26, n_253);
  not gc26 (wc26, n_349);
  or g624 (n_576, wc27, n_135);
  not gc27 (wc27, n_138);
  or g625 (n_577, wc28, n_145);
  not gc28 (wc28, n_140);
  or g626 (n_580, wc29, n_141);
  not gc29 (wc29, n_142);
  or g627 (n_581, wc30, n_151);
  not gc30 (wc30, n_146);
  or g628 (n_584, wc31, n_147);
  not gc31 (wc31, n_148);
  or g629 (n_586, wc32, n_157);
  not gc32 (wc32, n_152);
  or g630 (n_589, wc33, n_153);
  not gc33 (wc33, n_154);
  or g631 (n_590, wc34, n_163);
  not gc34 (wc34, n_158);
  or g632 (n_593, wc35, n_159);
  not gc35 (wc35, n_160);
  or g633 (n_595, wc36, n_169);
  not gc36 (wc36, n_164);
  or g634 (n_598, wc37, n_165);
  not gc37 (wc37, n_166);
  or g635 (n_601, wc38, n_175);
  not gc38 (wc38, n_170);
  or g636 (n_604, wc39, n_171);
  not gc39 (wc39, n_172);
  or g637 (n_606, wc40, n_181);
  not gc40 (wc40, n_176);
  or g638 (n_609, wc41, n_177);
  not gc41 (wc41, n_178);
  or g639 (n_610, wc42, n_187);
  not gc42 (wc42, n_182);
  or g640 (n_613, wc43, n_183);
  not gc43 (wc43, n_184);
  or g641 (n_615, wc44, n_193);
  not gc44 (wc44, n_188);
  or g642 (n_618, wc45, n_189);
  not gc45 (wc45, n_190);
  or g643 (n_621, wc46, n_199);
  not gc46 (wc46, n_194);
  or g644 (n_624, wc47, n_195);
  not gc47 (wc47, n_196);
  or g645 (n_626, wc48, n_205);
  not gc48 (wc48, n_200);
  or g646 (n_629, wc49, n_201);
  not gc49 (wc49, n_202);
  or g647 (n_631, wc50, n_211);
  not gc50 (wc50, n_206);
  or g648 (n_634, wc51, n_207);
  not gc51 (wc51, n_208);
  or g649 (n_636, wc52, n_217);
  not gc52 (wc52, n_212);
  or g650 (n_639, wc53, n_213);
  not gc53 (wc53, n_214);
  or g651 (n_642, wc54, n_223);
  not gc54 (wc54, n_218);
  or g652 (n_645, wc55, n_219);
  not gc55 (wc55, n_220);
  or g653 (n_647, wc56, n_229);
  not gc56 (wc56, n_224);
  or g654 (n_650, wc57, n_225);
  not gc57 (wc57, n_226);
  or g655 (n_651, wc58, n_235);
  not gc58 (wc58, n_230);
  or g656 (n_654, wc59, n_231);
  not gc59 (wc59, n_232);
  or g657 (n_656, wc60, n_241);
  not gc60 (wc60, n_236);
  or g658 (n_659, wc61, n_237);
  not gc61 (wc61, n_238);
  or g659 (n_662, wc62, n_247);
  not gc62 (wc62, n_242);
  or g660 (n_665, wc63, n_243);
  not gc63 (wc63, n_244);
  or g661 (n_667, wc64, n_253);
  not gc64 (wc64, n_248);
  or g662 (n_670, wc65, n_249);
  not gc65 (wc65, n_250);
  or g663 (n_672, wc66, n_259);
  not gc66 (wc66, n_254);
  and g664 (n_344, wc67, n_341);
  not gc67 (wc67, n_336);
  and g665 (n_354, wc68, n_351);
  not gc68 (wc68, n_346);
  and g666 (n_493, n_256, wc69);
  not gc69 (wc69, n_257);
  and g667 (n_304, wc70, n_301);
  not gc70 (wc70, n_296);
  and g668 (n_314, wc71, n_311);
  not gc71 (wc71, n_306);
  and g669 (n_324, wc72, n_321);
  not gc72 (wc72, n_316);
  and g670 (n_334, wc73, n_331);
  not gc73 (wc73, n_326);
  and g671 (n_284, wc74, n_281);
  not gc74 (wc74, n_276);
  and g672 (n_294, wc75, n_291);
  not gc75 (wc75, n_286);
  and g673 (n_274, wc76, n_271);
  not gc76 (wc76, n_266);
  and g674 (n_441, wc77, n_289);
  not gc77 (wc77, n_371);
  and g675 (n_509, wc78, n_309);
  not gc78 (wc78, n_386);
  and g676 (n_471, wc79, n_329);
  not gc79 (wc79, n_401);
  and g677 (n_561, wc80, n_349);
  not gc80 (wc80, n_416);
  xor g678 (Z[1], n_132, n_576);
  or g679 (n_675, wc81, n_255);
  not gc81 (wc81, n_256);
  and g680 (n_413, wc82, n_343);
  not gc82 (wc82, n_344);
  and g681 (n_425, wc83, n_353);
  not gc83 (wc83, n_354);
  and g682 (n_383, wc84, n_303);
  not gc84 (wc84, n_304);
  and g683 (n_395, wc85, n_313);
  not gc85 (wc85, n_314);
  and g684 (n_398, wc86, n_323);
  not gc86 (wc86, n_324);
  and g685 (n_410, wc87, n_333);
  not gc87 (wc87, n_334);
  and g686 (n_368, wc88, n_283);
  not gc88 (wc88, n_284);
  and g687 (n_380, wc89, n_293);
  not gc89 (wc89, n_294);
  and g688 (n_366, wc90, n_273);
  not gc90 (wc90, n_274);
  or g689 (n_262, wc91, n_145);
  not gc91 (wc91, n_260);
  and g690 (n_362, wc92, n_152);
  not gc92 (wc92, n_267);
  and g691 (n_434, wc93, n_164);
  not gc93 (wc93, n_277);
  and g692 (n_376, wc94, n_176);
  not gc94 (wc94, n_287);
  and g693 (n_502, wc95, n_188);
  not gc95 (wc95, n_297);
  and g694 (n_391, wc96, n_200);
  not gc96 (wc96, n_307);
  and g695 (n_459, wc97, n_212);
  not gc97 (wc97, n_317);
  and g696 (n_406, wc98, n_224);
  not gc98 (wc98, n_327);
  and g697 (n_554, wc99, n_236);
  not gc99 (wc99, n_337);
  and g698 (n_421, wc100, n_248);
  not gc100 (wc100, n_347);
  or g699 (n_516, wc101, n_211);
  not gc101 (wc101, n_453);
  or g700 (n_524, n_458, wc102);
  not gc102 (wc102, n_453);
  or g701 (n_528, wc103, n_401);
  not gc103 (wc103, n_453);
  or g702 (n_568, wc104, n_259);
  not gc104 (wc104, n_489);
  and g703 (n_373, wc105, n_289);
  not gc105 (wc105, n_368);
  and g704 (n_388, wc106, n_309);
  not gc106 (wc106, n_383);
  and g705 (n_403, wc107, n_329);
  not gc107 (wc107, n_398);
  and g706 (n_418, wc108, n_349);
  not gc108 (wc108, n_413);
  and g707 (n_486, n_425, wc109);
  not gc109 (wc109, n_426);
  and g708 (n_450, n_395, wc110);
  not gc110 (wc110, n_396);
  and g709 (n_483, n_410, wc111);
  not gc111 (wc111, n_411);
  and g710 (n_448, n_380, wc112);
  not gc112 (wc112, n_381);
  or g711 (n_367, n_364, wc113);
  not gc113 (wc113, n_356);
  or g712 (n_358, wc114, n_151);
  not gc114 (wc114, n_356);
  or g713 (n_363, n_360, wc115);
  not gc115 (wc115, n_356);
  and g714 (n_439, wc116, n_170);
  not gc116 (wc116, n_369);
  and g715 (n_442, wc117, n_286);
  not gc117 (wc117, n_373);
  and g716 (n_445, n_376, wc118);
  not gc118 (wc118, n_377);
  and g717 (n_507, wc119, n_194);
  not gc119 (wc119, n_384);
  and g718 (n_510, wc120, n_306);
  not gc120 (wc120, n_388);
  and g719 (n_513, n_391, wc121);
  not gc121 (wc121, n_392);
  and g720 (n_468, wc122, n_218);
  not gc122 (wc122, n_399);
  and g721 (n_473, wc123, n_326);
  not gc123 (wc123, n_403);
  and g722 (n_478, n_406, wc124);
  not gc124 (wc124, n_407);
  and g723 (n_559, wc125, n_242);
  not gc125 (wc125, n_414);
  and g724 (n_562, wc126, n_346);
  not gc126 (wc126, n_418);
  and g725 (n_565, n_421, wc127);
  not gc127 (wc127, n_422);
  and g726 (n_494, wc128, n_491);
  not gc128 (wc128, n_486);
  and g727 (n_484, wc129, n_481);
  not gc129 (wc129, n_450);
  and g728 (n_456, wc130, n_319);
  not gc130 (wc130, n_450);
  and g729 (n_469, wc131, n_466);
  not gc131 (wc131, n_450);
  and g730 (n_474, wc132, n_471);
  not gc132 (wc132, n_450);
  and g731 (n_479, wc133, n_476);
  not gc133 (wc133, n_450);
  and g732 (n_574, wc134, n_493);
  not gc134 (wc134, n_494);
  and g733 (n_546, wc135, n_483);
  not gc135 (wc135, n_484);
  or g734 (n_430, wc136, n_163);
  not gc136 (wc136, n_428);
  or g735 (n_435, n_432, wc137);
  not gc137 (wc137, n_428);
  or g736 (n_437, wc138, n_371);
  not gc138 (wc138, n_428);
  and g737 (n_518, wc139, n_206);
  not gc139 (wc139, n_451);
  and g738 (n_522, wc140, n_316);
  not gc140 (wc140, n_456);
  and g739 (n_526, n_459, wc141);
  not gc141 (wc141, n_460);
  and g740 (n_530, n_398, wc142);
  not gc142 (wc142, n_463);
  and g741 (n_534, wc143, n_468);
  not gc143 (wc143, n_469);
  and g742 (n_538, wc144, n_473);
  not gc144 (wc144, n_474);
  and g743 (n_542, wc145, n_478);
  not gc145 (wc145, n_479);
  and g744 (n_570, wc146, n_254);
  not gc146 (wc146, n_487);
  or g745 (n_547, n_544, wc147);
  not gc147 (wc147, n_496);
  or g746 (n_498, wc148, n_187);
  not gc148 (wc148, n_496);
  or g747 (n_503, n_500, wc149);
  not gc149 (wc149, n_496);
  or g748 (n_505, wc150, n_386);
  not gc150 (wc150, n_496);
  or g749 (n_519, n_516, wc151);
  not gc151 (wc151, n_496);
  or g750 (n_523, n_520, wc152);
  not gc152 (wc152, n_496);
  or g751 (n_527, n_524, wc153);
  not gc153 (wc153, n_496);
  or g752 (n_531, n_528, wc154);
  not gc154 (wc154, n_496);
  or g753 (n_535, n_532, wc155);
  not gc155 (wc155, n_496);
  or g754 (n_539, n_536, wc156);
  not gc156 (wc156, n_496);
  or g755 (n_543, n_540, wc157);
  not gc157 (wc157, n_496);
  or g756 (n_575, wc158, n_572);
  not gc158 (wc158, n_548);
  or g757 (n_550, wc159, n_235);
  not gc159 (wc159, n_548);
  or g758 (n_555, n_552, wc160);
  not gc160 (wc160, n_548);
  or g759 (n_557, wc161, n_416);
  not gc161 (wc161, n_548);
  or g760 (n_571, n_568, wc162);
  not gc162 (wc162, n_548);
endmodule

module add_signed_426_GENERIC(A, B, Z);
  input [41:0] A, B;
  output [42:0] Z;
  wire [41:0] A, B;
  wire [42:0] Z;
  add_signed_426_GENERIC_REAL g1(.A ({A[40], A[40:0]}), .B ({B[40],
       B[40:0]}), .Z (Z));
endmodule

module add_signed_440_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [40:0] A, B;
  output [41:0] Z;
  wire [40:0] A, B;
  wire [41:0] Z;
  wire n_128, n_129, n_132, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_142, n_143, n_144, n_145, n_146, n_148, n_149;
  wire n_150, n_151, n_152, n_154, n_155, n_156, n_157, n_158;
  wire n_160, n_161, n_162, n_163, n_164, n_166, n_167, n_168;
  wire n_169, n_170, n_172, n_173, n_174, n_175, n_176, n_178;
  wire n_179, n_180, n_181, n_182, n_184, n_185, n_186, n_187;
  wire n_188, n_190, n_191, n_192, n_193, n_194, n_196, n_197;
  wire n_198, n_199, n_200, n_202, n_203, n_204, n_205, n_206;
  wire n_208, n_209, n_210, n_211, n_212, n_214, n_215, n_216;
  wire n_217, n_218, n_220, n_221, n_222, n_223, n_224, n_226;
  wire n_227, n_228, n_229, n_230, n_232, n_233, n_234, n_235;
  wire n_236, n_238, n_239, n_240, n_241, n_242, n_244, n_245;
  wire n_246, n_247, n_248, n_250, n_251, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_260, n_262, n_264, n_265, n_267;
  wire n_268, n_270, n_272, n_274, n_275, n_277, n_278, n_280;
  wire n_282, n_284, n_285, n_287, n_288, n_290, n_292, n_294;
  wire n_295, n_297, n_298, n_300, n_302, n_304, n_305, n_307;
  wire n_308, n_310, n_312, n_314, n_315, n_317, n_318, n_320;
  wire n_322, n_324, n_325, n_327, n_328, n_330, n_332, n_334;
  wire n_335, n_337, n_338, n_340, n_342, n_344, n_345, n_347;
  wire n_349, n_350, n_351, n_353, n_354, n_355, n_357, n_358;
  wire n_359, n_360, n_362, n_364, n_366, n_367, n_368, n_370;
  wire n_371, n_372, n_374, n_375, n_377, n_379, n_381, n_382;
  wire n_383, n_385, n_386, n_387, n_389, n_390, n_392, n_394;
  wire n_396, n_397, n_398, n_400, n_401, n_402, n_404, n_405;
  wire n_407, n_409, n_411, n_412, n_413, n_415, n_416, n_417;
  wire n_419, n_421, n_422, n_423, n_425, n_426, n_428, n_429;
  wire n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437;
  wire n_438, n_439, n_440, n_441, n_442, n_444, n_447, n_449;
  wire n_450, n_451, n_454, n_457, n_459, n_460, n_462, n_464;
  wire n_465, n_467, n_469, n_470, n_472, n_474, n_475, n_477;
  wire n_478, n_479, n_480, n_482, n_484, n_486, n_487, n_488;
  wire n_490, n_491, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_506, n_507;
  wire n_508, n_510, n_511, n_512, n_514, n_515, n_516, n_518;
  wire n_519, n_520, n_522, n_523, n_524, n_526, n_527, n_528;
  wire n_530, n_531, n_532, n_534, n_535, n_536, n_538, n_539;
  wire n_540, n_542, n_543, n_545, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_558;
  wire n_559, n_560, n_561, n_563, n_564, n_565, n_567, n_568;
  wire n_569, n_570, n_572, n_573, n_574, n_576, n_577, n_578;
  wire n_579, n_581, n_582, n_584, n_585, n_587, n_588, n_589;
  wire n_590, n_592, n_593, n_594, n_596, n_597, n_598, n_599;
  wire n_601, n_602, n_604, n_605, n_607, n_608, n_609, n_610;
  wire n_612, n_613, n_614, n_615, n_617, n_618, n_619, n_620;
  wire n_622, n_623, n_625, n_626, n_628, n_629, n_630, n_631;
  wire n_633, n_634, n_635, n_637, n_638, n_639, n_640, n_642;
  wire n_643, n_645, n_646, n_648, n_649, n_650, n_651, n_653;
  wire n_654, n_655, n_656;
  not g3 (Z[41], n_128);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_129, A[0], B[0]);
  nor g9 (n_132, A[1], B[1]);
  nand g10 (n_135, A[1], B[1]);
  nor g11 (n_142, A[2], B[2]);
  nand g12 (n_137, A[2], B[2]);
  nor g13 (n_138, A[3], B[3]);
  nand g14 (n_139, A[3], B[3]);
  nor g15 (n_148, A[4], B[4]);
  nand g16 (n_143, A[4], B[4]);
  nor g17 (n_144, A[5], B[5]);
  nand g18 (n_145, A[5], B[5]);
  nor g19 (n_154, A[6], B[6]);
  nand g20 (n_149, A[6], B[6]);
  nor g21 (n_150, A[7], B[7]);
  nand g22 (n_151, A[7], B[7]);
  nor g23 (n_160, A[8], B[8]);
  nand g24 (n_155, A[8], B[8]);
  nor g25 (n_156, A[9], B[9]);
  nand g26 (n_157, A[9], B[9]);
  nor g27 (n_166, A[10], B[10]);
  nand g28 (n_161, A[10], B[10]);
  nor g29 (n_162, A[11], B[11]);
  nand g30 (n_163, A[11], B[11]);
  nor g31 (n_172, A[12], B[12]);
  nand g32 (n_167, A[12], B[12]);
  nor g33 (n_168, A[13], B[13]);
  nand g34 (n_169, A[13], B[13]);
  nor g35 (n_178, A[14], B[14]);
  nand g36 (n_173, A[14], B[14]);
  nor g37 (n_174, A[15], B[15]);
  nand g38 (n_175, A[15], B[15]);
  nor g39 (n_184, A[16], B[16]);
  nand g40 (n_179, A[16], B[16]);
  nor g41 (n_180, A[17], B[17]);
  nand g42 (n_181, A[17], B[17]);
  nor g43 (n_190, A[18], B[18]);
  nand g44 (n_185, A[18], B[18]);
  nor g45 (n_186, A[19], B[19]);
  nand g46 (n_187, A[19], B[19]);
  nor g47 (n_196, A[20], B[20]);
  nand g48 (n_191, A[20], B[20]);
  nor g49 (n_192, A[21], B[21]);
  nand g50 (n_193, A[21], B[21]);
  nor g51 (n_202, A[22], B[22]);
  nand g52 (n_197, A[22], B[22]);
  nor g53 (n_198, A[23], B[23]);
  nand g54 (n_199, A[23], B[23]);
  nor g55 (n_208, A[24], B[24]);
  nand g56 (n_203, A[24], B[24]);
  nor g57 (n_204, A[25], B[25]);
  nand g58 (n_205, A[25], B[25]);
  nor g59 (n_214, A[26], B[26]);
  nand g60 (n_209, A[26], B[26]);
  nor g61 (n_210, A[27], B[27]);
  nand g62 (n_211, A[27], B[27]);
  nor g63 (n_220, A[28], B[28]);
  nand g64 (n_215, A[28], B[28]);
  nor g65 (n_216, A[29], B[29]);
  nand g66 (n_217, A[29], B[29]);
  nor g67 (n_226, A[30], B[30]);
  nand g68 (n_221, A[30], B[30]);
  nor g69 (n_222, A[31], B[31]);
  nand g70 (n_223, A[31], B[31]);
  nor g71 (n_232, A[32], B[32]);
  nand g72 (n_227, A[32], B[32]);
  nor g73 (n_228, A[33], B[33]);
  nand g74 (n_229, A[33], B[33]);
  nor g75 (n_238, A[34], B[34]);
  nand g76 (n_233, A[34], B[34]);
  nor g77 (n_234, A[35], B[35]);
  nand g78 (n_235, A[35], B[35]);
  nor g79 (n_244, A[36], B[36]);
  nand g80 (n_239, A[36], B[36]);
  nor g81 (n_240, A[37], B[37]);
  nand g82 (n_241, A[37], B[37]);
  nor g83 (n_250, A[38], B[38]);
  nand g84 (n_245, A[38], B[38]);
  nor g85 (n_246, A[39], B[39]);
  nand g86 (n_247, A[39], B[39]);
  nand g91 (n_251, n_135, n_136);
  nor g92 (n_140, n_137, n_138);
  nor g95 (n_254, n_142, n_138);
  nor g96 (n_146, n_143, n_144);
  nor g99 (n_260, n_148, n_144);
  nor g100 (n_152, n_149, n_150);
  nor g103 (n_262, n_154, n_150);
  nor g104 (n_158, n_155, n_156);
  nor g107 (n_270, n_160, n_156);
  nor g108 (n_164, n_161, n_162);
  nor g111 (n_272, n_166, n_162);
  nor g112 (n_170, n_167, n_168);
  nor g115 (n_280, n_172, n_168);
  nor g116 (n_176, n_173, n_174);
  nor g119 (n_282, n_178, n_174);
  nor g120 (n_182, n_179, n_180);
  nor g123 (n_290, n_184, n_180);
  nor g124 (n_188, n_185, n_186);
  nor g127 (n_292, n_190, n_186);
  nor g128 (n_194, n_191, n_192);
  nor g131 (n_300, n_196, n_192);
  nor g132 (n_200, n_197, n_198);
  nor g135 (n_302, n_202, n_198);
  nor g136 (n_206, n_203, n_204);
  nor g139 (n_310, n_208, n_204);
  nor g140 (n_212, n_209, n_210);
  nor g143 (n_312, n_214, n_210);
  nor g144 (n_218, n_215, n_216);
  nor g147 (n_320, n_220, n_216);
  nor g148 (n_224, n_221, n_222);
  nor g151 (n_322, n_226, n_222);
  nor g152 (n_230, n_227, n_228);
  nor g155 (n_330, n_232, n_228);
  nor g156 (n_236, n_233, n_234);
  nor g159 (n_332, n_238, n_234);
  nor g160 (n_242, n_239, n_240);
  nor g163 (n_340, n_244, n_240);
  nor g164 (n_248, n_245, n_246);
  nor g167 (n_342, n_250, n_246);
  nand g170 (n_563, n_137, n_253);
  nand g171 (n_256, n_254, n_251);
  nand g172 (n_347, n_255, n_256);
  nor g173 (n_258, n_154, n_257);
  nand g182 (n_355, n_260, n_262);
  nor g183 (n_268, n_166, n_267);
  nand g192 (n_362, n_270, n_272);
  nor g193 (n_278, n_178, n_277);
  nand g202 (n_370, n_280, n_282);
  nor g203 (n_288, n_190, n_287);
  nand g212 (n_377, n_290, n_292);
  nor g213 (n_298, n_202, n_297);
  nand g222 (n_385, n_300, n_302);
  nor g223 (n_308, n_214, n_307);
  nand g232 (n_392, n_310, n_312);
  nor g233 (n_318, n_226, n_317);
  nand g242 (n_400, n_320, n_322);
  nor g243 (n_328, n_238, n_327);
  nand g252 (n_407, n_330, n_332);
  nor g253 (n_338, n_250, n_337);
  nand g262 (n_415, n_340, n_342);
  nand g265 (n_567, n_143, n_349);
  nand g266 (n_350, n_260, n_347);
  nand g267 (n_569, n_257, n_350);
  nand g270 (n_572, n_353, n_354);
  nand g273 (n_419, n_357, n_358);
  nor g274 (n_360, n_172, n_359);
  nor g277 (n_429, n_172, n_362);
  nor g283 (n_368, n_366, n_359);
  nor g286 (n_435, n_362, n_366);
  nor g287 (n_372, n_370, n_359);
  nor g290 (n_438, n_362, n_370);
  nor g291 (n_375, n_196, n_374);
  nor g294 (n_494, n_196, n_377);
  nor g300 (n_383, n_381, n_374);
  nor g303 (n_500, n_377, n_381);
  nor g304 (n_387, n_385, n_374);
  nor g307 (n_444, n_377, n_385);
  nor g308 (n_390, n_220, n_389);
  nor g311 (n_457, n_220, n_392);
  nor g317 (n_398, n_396, n_389);
  nor g320 (n_467, n_392, n_396);
  nor g321 (n_402, n_400, n_389);
  nor g324 (n_472, n_392, n_400);
  nor g325 (n_405, n_244, n_404);
  nor g328 (n_546, n_244, n_407);
  nor g334 (n_413, n_411, n_404);
  nor g337 (n_552, n_407, n_411);
  nor g338 (n_417, n_415, n_404);
  nor g341 (n_482, n_407, n_415);
  nand g344 (n_576, n_155, n_421);
  nand g345 (n_422, n_270, n_419);
  nand g346 (n_578, n_267, n_422);
  nand g349 (n_581, n_425, n_426);
  nand g352 (n_584, n_359, n_428);
  nand g353 (n_431, n_429, n_419);
  nand g354 (n_587, n_430, n_431);
  nand g355 (n_434, n_432, n_419);
  nand g356 (n_589, n_433, n_434);
  nand g357 (n_437, n_435, n_419);
  nand g358 (n_592, n_436, n_437);
  nand g359 (n_440, n_438, n_419);
  nand g360 (n_484, n_439, n_440);
  nor g361 (n_442, n_208, n_441);
  nand g370 (n_508, n_310, n_444);
  nor g371 (n_451, n_449, n_441);
  nor g376 (n_454, n_392, n_441);
  nand g385 (n_520, n_444, n_457);
  nand g390 (n_524, n_444, n_462);
  nand g395 (n_528, n_444, n_467);
  nand g400 (n_532, n_444, n_472);
  nor g401 (n_480, n_477, n_478);
  nand g408 (n_596, n_179, n_486);
  nand g409 (n_487, n_290, n_484);
  nand g410 (n_598, n_287, n_487);
  nand g413 (n_601, n_490, n_491);
  nand g416 (n_604, n_374, n_493);
  nand g417 (n_496, n_494, n_484);
  nand g418 (n_607, n_495, n_496);
  nand g419 (n_499, n_497, n_484);
  nand g420 (n_609, n_498, n_499);
  nand g421 (n_502, n_500, n_484);
  nand g422 (n_612, n_501, n_502);
  nand g423 (n_503, n_444, n_484);
  nand g424 (n_614, n_441, n_503);
  nand g427 (n_617, n_506, n_507);
  nand g430 (n_619, n_510, n_511);
  nand g433 (n_622, n_514, n_515);
  nand g436 (n_625, n_518, n_519);
  nand g439 (n_628, n_522, n_523);
  nand g442 (n_630, n_526, n_527);
  nand g445 (n_633, n_530, n_531);
  nand g448 (n_536, n_534, n_535);
  nand g451 (n_637, n_227, n_538);
  nand g452 (n_539, n_330, n_536);
  nand g453 (n_639, n_327, n_539);
  nand g456 (n_642, n_542, n_543);
  nand g459 (n_645, n_404, n_545);
  nand g460 (n_548, n_546, n_536);
  nand g461 (n_648, n_547, n_548);
  nand g462 (n_551, n_549, n_536);
  nand g463 (n_650, n_550, n_551);
  nand g464 (n_554, n_552, n_536);
  nand g465 (n_653, n_553, n_554);
  nand g466 (n_555, n_482, n_536);
  nand g467 (n_655, n_478, n_555);
  nand g470 (n_128, n_558, n_559);
  xnor g474 (Z[2], n_251, n_561);
  xnor g477 (Z[3], n_563, n_564);
  xnor g479 (Z[4], n_347, n_565);
  xnor g482 (Z[5], n_567, n_568);
  xnor g484 (Z[6], n_569, n_570);
  xnor g487 (Z[7], n_572, n_573);
  xnor g489 (Z[8], n_419, n_574);
  xnor g492 (Z[9], n_576, n_577);
  xnor g494 (Z[10], n_578, n_579);
  xnor g497 (Z[11], n_581, n_582);
  xnor g500 (Z[12], n_584, n_585);
  xnor g503 (Z[13], n_587, n_588);
  xnor g505 (Z[14], n_589, n_590);
  xnor g508 (Z[15], n_592, n_593);
  xnor g510 (Z[16], n_484, n_594);
  xnor g513 (Z[17], n_596, n_597);
  xnor g515 (Z[18], n_598, n_599);
  xnor g518 (Z[19], n_601, n_602);
  xnor g521 (Z[20], n_604, n_605);
  xnor g524 (Z[21], n_607, n_608);
  xnor g526 (Z[22], n_609, n_610);
  xnor g529 (Z[23], n_612, n_613);
  xnor g531 (Z[24], n_614, n_615);
  xnor g534 (Z[25], n_617, n_618);
  xnor g536 (Z[26], n_619, n_620);
  xnor g539 (Z[27], n_622, n_623);
  xnor g542 (Z[28], n_625, n_626);
  xnor g545 (Z[29], n_628, n_629);
  xnor g547 (Z[30], n_630, n_631);
  xnor g550 (Z[31], n_633, n_634);
  xnor g552 (Z[32], n_536, n_635);
  xnor g555 (Z[33], n_637, n_638);
  xnor g557 (Z[34], n_639, n_640);
  xnor g560 (Z[35], n_642, n_643);
  xnor g563 (Z[36], n_645, n_646);
  xnor g566 (Z[37], n_648, n_649);
  xnor g568 (Z[38], n_650, n_651);
  xnor g571 (Z[39], n_653, n_654);
  xnor g573 (Z[40], n_655, n_656);
  and g576 (n_477, A[40], B[40]);
  or g577 (n_479, A[40], B[40]);
  and g578 (n_327, wc, n_229);
  not gc (wc, n_230);
  and g579 (n_334, wc0, n_235);
  not gc0 (wc0, n_236);
  and g580 (n_337, wc1, n_241);
  not gc1 (wc1, n_242);
  and g581 (n_344, wc2, n_247);
  not gc2 (wc2, n_248);
  and g582 (n_287, wc3, n_181);
  not gc3 (wc3, n_182);
  and g583 (n_294, wc4, n_187);
  not gc4 (wc4, n_188);
  and g584 (n_297, wc5, n_193);
  not gc5 (wc5, n_194);
  and g585 (n_304, wc6, n_199);
  not gc6 (wc6, n_200);
  and g586 (n_307, wc7, n_205);
  not gc7 (wc7, n_206);
  and g587 (n_314, wc8, n_211);
  not gc8 (wc8, n_212);
  and g588 (n_317, wc9, n_217);
  not gc9 (wc9, n_218);
  and g589 (n_324, wc10, n_223);
  not gc10 (wc10, n_224);
  and g590 (n_267, wc11, n_157);
  not gc11 (wc11, n_158);
  and g591 (n_274, wc12, n_163);
  not gc12 (wc12, n_164);
  and g592 (n_277, wc13, n_169);
  not gc13 (wc13, n_170);
  and g593 (n_284, wc14, n_175);
  not gc14 (wc14, n_176);
  and g594 (n_257, wc15, n_145);
  not gc15 (wc15, n_146);
  and g595 (n_264, wc16, n_151);
  not gc16 (wc16, n_152);
  and g596 (n_255, wc17, n_139);
  not gc17 (wc17, n_140);
  or g597 (n_136, n_129, n_132);
  or g598 (n_351, wc18, n_154);
  not gc18 (wc18, n_260);
  or g599 (n_423, wc19, n_166);
  not gc19 (wc19, n_270);
  or g600 (n_366, wc20, n_178);
  not gc20 (wc20, n_280);
  or g601 (n_488, wc21, n_190);
  not gc21 (wc21, n_290);
  or g602 (n_381, wc22, n_202);
  not gc22 (wc22, n_300);
  or g603 (n_449, wc23, n_214);
  not gc23 (wc23, n_310);
  or g604 (n_396, wc24, n_226);
  not gc24 (wc24, n_320);
  or g605 (n_540, wc25, n_238);
  not gc25 (wc25, n_330);
  or g606 (n_411, wc26, n_250);
  not gc26 (wc26, n_340);
  or g607 (n_560, wc27, n_132);
  not gc27 (wc27, n_135);
  or g608 (n_561, wc28, n_142);
  not gc28 (wc28, n_137);
  or g609 (n_564, wc29, n_138);
  not gc29 (wc29, n_139);
  or g610 (n_565, wc30, n_148);
  not gc30 (wc30, n_143);
  or g611 (n_568, wc31, n_144);
  not gc31 (wc31, n_145);
  or g612 (n_570, wc32, n_154);
  not gc32 (wc32, n_149);
  or g613 (n_573, wc33, n_150);
  not gc33 (wc33, n_151);
  or g614 (n_574, wc34, n_160);
  not gc34 (wc34, n_155);
  or g615 (n_577, wc35, n_156);
  not gc35 (wc35, n_157);
  or g616 (n_579, wc36, n_166);
  not gc36 (wc36, n_161);
  or g617 (n_582, wc37, n_162);
  not gc37 (wc37, n_163);
  or g618 (n_585, wc38, n_172);
  not gc38 (wc38, n_167);
  or g619 (n_588, wc39, n_168);
  not gc39 (wc39, n_169);
  or g620 (n_590, wc40, n_178);
  not gc40 (wc40, n_173);
  or g621 (n_593, wc41, n_174);
  not gc41 (wc41, n_175);
  or g622 (n_594, wc42, n_184);
  not gc42 (wc42, n_179);
  or g623 (n_597, wc43, n_180);
  not gc43 (wc43, n_181);
  or g624 (n_599, wc44, n_190);
  not gc44 (wc44, n_185);
  or g625 (n_602, wc45, n_186);
  not gc45 (wc45, n_187);
  or g626 (n_605, wc46, n_196);
  not gc46 (wc46, n_191);
  or g627 (n_608, wc47, n_192);
  not gc47 (wc47, n_193);
  or g628 (n_610, wc48, n_202);
  not gc48 (wc48, n_197);
  or g629 (n_613, wc49, n_198);
  not gc49 (wc49, n_199);
  or g630 (n_615, wc50, n_208);
  not gc50 (wc50, n_203);
  or g631 (n_618, wc51, n_204);
  not gc51 (wc51, n_205);
  or g632 (n_620, wc52, n_214);
  not gc52 (wc52, n_209);
  or g633 (n_623, wc53, n_210);
  not gc53 (wc53, n_211);
  or g634 (n_626, wc54, n_220);
  not gc54 (wc54, n_215);
  or g635 (n_629, wc55, n_216);
  not gc55 (wc55, n_217);
  or g636 (n_631, wc56, n_226);
  not gc56 (wc56, n_221);
  or g637 (n_634, wc57, n_222);
  not gc57 (wc57, n_223);
  or g638 (n_635, wc58, n_232);
  not gc58 (wc58, n_227);
  or g639 (n_638, wc59, n_228);
  not gc59 (wc59, n_229);
  or g640 (n_640, wc60, n_238);
  not gc60 (wc60, n_233);
  or g641 (n_643, wc61, n_234);
  not gc61 (wc61, n_235);
  or g642 (n_646, wc62, n_244);
  not gc62 (wc62, n_239);
  or g643 (n_649, wc63, n_240);
  not gc63 (wc63, n_241);
  or g644 (n_651, wc64, n_250);
  not gc64 (wc64, n_245);
  or g645 (n_654, wc65, n_246);
  not gc65 (wc65, n_247);
  and g646 (n_335, wc66, n_332);
  not gc66 (wc66, n_327);
  and g647 (n_345, wc67, n_342);
  not gc67 (wc67, n_337);
  and g648 (n_295, wc68, n_292);
  not gc68 (wc68, n_287);
  and g649 (n_305, wc69, n_302);
  not gc69 (wc69, n_297);
  and g650 (n_315, wc70, n_312);
  not gc70 (wc70, n_307);
  and g651 (n_325, wc71, n_322);
  not gc71 (wc71, n_317);
  and g652 (n_275, wc72, n_272);
  not gc72 (wc72, n_267);
  and g653 (n_285, wc73, n_282);
  not gc73 (wc73, n_277);
  and g654 (n_265, wc74, n_262);
  not gc74 (wc74, n_257);
  and g655 (n_432, wc75, n_280);
  not gc75 (wc75, n_362);
  and g656 (n_497, wc76, n_300);
  not gc76 (wc76, n_377);
  and g657 (n_462, wc77, n_320);
  not gc77 (wc77, n_392);
  and g658 (n_549, wc78, n_340);
  not gc78 (wc78, n_407);
  xor g659 (Z[1], n_129, n_560);
  or g660 (n_656, wc79, n_477);
  not gc79 (wc79, n_479);
  and g661 (n_404, wc80, n_334);
  not gc80 (wc80, n_335);
  and g662 (n_416, wc81, n_344);
  not gc81 (wc81, n_345);
  and g663 (n_374, wc82, n_294);
  not gc82 (wc82, n_295);
  and g664 (n_386, wc83, n_304);
  not gc83 (wc83, n_305);
  and g665 (n_389, wc84, n_314);
  not gc84 (wc84, n_315);
  and g666 (n_401, wc85, n_324);
  not gc85 (wc85, n_325);
  and g667 (n_359, wc86, n_274);
  not gc86 (wc86, n_275);
  and g668 (n_371, wc87, n_284);
  not gc87 (wc87, n_285);
  and g669 (n_357, wc88, n_264);
  not gc88 (wc88, n_265);
  or g670 (n_556, n_477, wc89);
  not gc89 (wc89, n_482);
  or g671 (n_253, wc90, n_142);
  not gc90 (wc90, n_251);
  and g672 (n_353, wc91, n_149);
  not gc91 (wc91, n_258);
  and g673 (n_425, wc92, n_161);
  not gc92 (wc92, n_268);
  and g674 (n_367, wc93, n_173);
  not gc93 (wc93, n_278);
  and g675 (n_490, wc94, n_185);
  not gc94 (wc94, n_288);
  and g676 (n_382, wc95, n_197);
  not gc95 (wc95, n_298);
  and g677 (n_450, wc96, n_209);
  not gc96 (wc96, n_308);
  and g678 (n_397, wc97, n_221);
  not gc97 (wc97, n_318);
  and g679 (n_542, wc98, n_233);
  not gc98 (wc98, n_328);
  and g680 (n_412, wc99, n_245);
  not gc99 (wc99, n_338);
  or g681 (n_504, wc100, n_208);
  not gc100 (wc100, n_444);
  or g682 (n_512, n_449, wc101);
  not gc101 (wc101, n_444);
  or g683 (n_516, wc102, n_392);
  not gc102 (wc102, n_444);
  and g684 (n_364, wc103, n_280);
  not gc103 (wc103, n_359);
  and g685 (n_379, wc104, n_300);
  not gc104 (wc104, n_374);
  and g686 (n_394, wc105, n_320);
  not gc105 (wc105, n_389);
  and g687 (n_409, wc106, n_340);
  not gc106 (wc106, n_404);
  and g688 (n_478, n_416, wc107);
  not gc107 (wc107, n_417);
  and g689 (n_441, n_386, wc108);
  not gc108 (wc108, n_387);
  and g690 (n_474, n_401, wc109);
  not gc109 (wc109, n_402);
  and g691 (n_439, n_371, wc110);
  not gc110 (wc110, n_372);
  or g692 (n_358, n_355, wc111);
  not gc111 (wc111, n_347);
  or g693 (n_349, wc112, n_148);
  not gc112 (wc112, n_347);
  or g694 (n_354, n_351, wc113);
  not gc113 (wc113, n_347);
  and g695 (n_430, wc114, n_167);
  not gc114 (wc114, n_360);
  and g696 (n_433, wc115, n_277);
  not gc115 (wc115, n_364);
  and g697 (n_436, n_367, wc116);
  not gc116 (wc116, n_368);
  and g698 (n_495, wc117, n_191);
  not gc117 (wc117, n_375);
  and g699 (n_498, wc118, n_297);
  not gc118 (wc118, n_379);
  and g700 (n_501, n_382, wc119);
  not gc119 (wc119, n_383);
  and g701 (n_459, wc120, n_215);
  not gc120 (wc120, n_390);
  and g702 (n_464, wc121, n_317);
  not gc121 (wc121, n_394);
  and g703 (n_469, n_397, wc122);
  not gc122 (wc122, n_398);
  and g704 (n_547, wc123, n_239);
  not gc123 (wc123, n_405);
  and g705 (n_550, wc124, n_337);
  not gc124 (wc124, n_409);
  and g706 (n_553, n_412, wc125);
  not gc125 (wc125, n_413);
  and g707 (n_475, wc126, n_472);
  not gc126 (wc126, n_441);
  and g708 (n_447, wc127, n_310);
  not gc127 (wc127, n_441);
  and g709 (n_460, wc128, n_457);
  not gc128 (wc128, n_441);
  and g710 (n_465, wc129, n_462);
  not gc129 (wc129, n_441);
  and g711 (n_470, wc130, n_467);
  not gc130 (wc130, n_441);
  and g712 (n_558, n_479, wc131);
  not gc131 (wc131, n_480);
  and g713 (n_534, wc132, n_474);
  not gc132 (wc132, n_475);
  or g714 (n_421, wc133, n_160);
  not gc133 (wc133, n_419);
  or g715 (n_426, n_423, wc134);
  not gc134 (wc134, n_419);
  or g716 (n_428, wc135, n_362);
  not gc135 (wc135, n_419);
  and g717 (n_506, wc136, n_203);
  not gc136 (wc136, n_442);
  and g718 (n_510, wc137, n_307);
  not gc137 (wc137, n_447);
  and g719 (n_514, n_450, wc138);
  not gc138 (wc138, n_451);
  and g720 (n_518, n_389, wc139);
  not gc139 (wc139, n_454);
  and g721 (n_522, wc140, n_459);
  not gc140 (wc140, n_460);
  and g722 (n_526, wc141, n_464);
  not gc141 (wc141, n_465);
  and g723 (n_530, wc142, n_469);
  not gc142 (wc142, n_470);
  or g724 (n_535, n_532, wc143);
  not gc143 (wc143, n_484);
  or g725 (n_486, wc144, n_184);
  not gc144 (wc144, n_484);
  or g726 (n_491, n_488, wc145);
  not gc145 (wc145, n_484);
  or g727 (n_493, wc146, n_377);
  not gc146 (wc146, n_484);
  or g728 (n_507, n_504, wc147);
  not gc147 (wc147, n_484);
  or g729 (n_511, n_508, wc148);
  not gc148 (wc148, n_484);
  or g730 (n_515, n_512, wc149);
  not gc149 (wc149, n_484);
  or g731 (n_519, n_516, wc150);
  not gc150 (wc150, n_484);
  or g732 (n_523, n_520, wc151);
  not gc151 (wc151, n_484);
  or g733 (n_527, n_524, wc152);
  not gc152 (wc152, n_484);
  or g734 (n_531, n_528, wc153);
  not gc153 (wc153, n_484);
  or g735 (n_559, n_556, wc154);
  not gc154 (wc154, n_536);
  or g736 (n_538, wc155, n_232);
  not gc155 (wc155, n_536);
  or g737 (n_543, n_540, wc156);
  not gc156 (wc156, n_536);
  or g738 (n_545, wc157, n_407);
  not gc157 (wc157, n_536);
endmodule

module add_signed_440_GENERIC(A, B, Z);
  input [40:0] A, B;
  output [41:0] Z;
  wire [40:0] A, B;
  wire [41:0] Z;
  add_signed_440_GENERIC_REAL g1(.A ({A[39], A[39:0]}), .B ({B[39],
       B[39:0]}), .Z (Z));
endmodule

module add_signed_454_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [39:0] A, B;
  output [40:0] Z;
  wire [39:0] A, B;
  wire [40:0] Z;
  wire n_125, n_126, n_129, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_139, n_140, n_141, n_142, n_143, n_145, n_146;
  wire n_147, n_148, n_149, n_151, n_152, n_153, n_154, n_155;
  wire n_157, n_158, n_159, n_160, n_161, n_163, n_164, n_165;
  wire n_166, n_167, n_169, n_170, n_171, n_172, n_173, n_175;
  wire n_176, n_177, n_178, n_179, n_181, n_182, n_183, n_184;
  wire n_185, n_187, n_188, n_189, n_190, n_191, n_193, n_194;
  wire n_195, n_196, n_197, n_199, n_200, n_201, n_202, n_203;
  wire n_205, n_206, n_207, n_208, n_209, n_211, n_212, n_213;
  wire n_214, n_215, n_217, n_218, n_219, n_220, n_221, n_223;
  wire n_224, n_225, n_226, n_227, n_229, n_230, n_231, n_232;
  wire n_233, n_235, n_236, n_237, n_238, n_239, n_241, n_242;
  wire n_243, n_244, n_245, n_247, n_248, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_257, n_259, n_261, n_262, n_264;
  wire n_265, n_267, n_269, n_271, n_272, n_274, n_275, n_277;
  wire n_279, n_281, n_282, n_284, n_285, n_287, n_289, n_291;
  wire n_292, n_294, n_295, n_297, n_299, n_301, n_302, n_304;
  wire n_305, n_307, n_309, n_311, n_312, n_314, n_315, n_317;
  wire n_319, n_321, n_322, n_324, n_325, n_327, n_329, n_331;
  wire n_332, n_334, n_335, n_337, n_339, n_341, n_342, n_344;
  wire n_346, n_347, n_348, n_350, n_351, n_352, n_354, n_355;
  wire n_356, n_357, n_359, n_361, n_363, n_364, n_365, n_367;
  wire n_368, n_369, n_371, n_372, n_374, n_376, n_378, n_379;
  wire n_380, n_382, n_383, n_384, n_386, n_387, n_389, n_391;
  wire n_393, n_394, n_395, n_397, n_398, n_399, n_401, n_402;
  wire n_404, n_406, n_408, n_409, n_410, n_412, n_413, n_414;
  wire n_416, n_418, n_419, n_420, n_422, n_423, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_441, n_444, n_446;
  wire n_447, n_448, n_451, n_454, n_456, n_457, n_459, n_461;
  wire n_462, n_464, n_466, n_467, n_469, n_471, n_472, n_474;
  wire n_476, n_477, n_478, n_480, n_481, n_483, n_484, n_485;
  wire n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_494, n_496, n_497, n_498, n_500, n_501, n_502, n_504;
  wire n_505, n_506, n_508, n_509, n_510, n_512, n_513, n_514;
  wire n_516, n_517, n_518, n_520, n_521, n_522, n_524, n_525;
  wire n_526, n_528, n_529, n_530, n_532, n_533, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_551, n_552, n_553;
  wire n_555, n_556, n_557, n_558, n_560, n_561, n_562, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_572, n_573, n_575;
  wire n_576, n_577, n_578, n_580, n_581, n_582, n_584, n_585;
  wire n_586, n_587, n_589, n_590, n_592, n_593, n_595, n_596;
  wire n_597, n_598, n_600, n_601, n_602, n_603, n_605, n_606;
  wire n_607, n_608, n_610, n_611, n_613, n_614, n_616, n_617;
  wire n_618, n_619, n_621, n_622, n_623, n_625, n_626, n_627;
  wire n_628, n_630, n_631, n_633, n_634, n_636, n_637, n_638;
  wire n_639, n_641, n_642;
  not g3 (Z[40], n_125);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_126, A[0], B[0]);
  nor g9 (n_129, A[1], B[1]);
  nand g10 (n_132, A[1], B[1]);
  nor g11 (n_139, A[2], B[2]);
  nand g12 (n_134, A[2], B[2]);
  nor g13 (n_135, A[3], B[3]);
  nand g14 (n_136, A[3], B[3]);
  nor g15 (n_145, A[4], B[4]);
  nand g16 (n_140, A[4], B[4]);
  nor g17 (n_141, A[5], B[5]);
  nand g18 (n_142, A[5], B[5]);
  nor g19 (n_151, A[6], B[6]);
  nand g20 (n_146, A[6], B[6]);
  nor g21 (n_147, A[7], B[7]);
  nand g22 (n_148, A[7], B[7]);
  nor g23 (n_157, A[8], B[8]);
  nand g24 (n_152, A[8], B[8]);
  nor g25 (n_153, A[9], B[9]);
  nand g26 (n_154, A[9], B[9]);
  nor g27 (n_163, A[10], B[10]);
  nand g28 (n_158, A[10], B[10]);
  nor g29 (n_159, A[11], B[11]);
  nand g30 (n_160, A[11], B[11]);
  nor g31 (n_169, A[12], B[12]);
  nand g32 (n_164, A[12], B[12]);
  nor g33 (n_165, A[13], B[13]);
  nand g34 (n_166, A[13], B[13]);
  nor g35 (n_175, A[14], B[14]);
  nand g36 (n_170, A[14], B[14]);
  nor g37 (n_171, A[15], B[15]);
  nand g38 (n_172, A[15], B[15]);
  nor g39 (n_181, A[16], B[16]);
  nand g40 (n_176, A[16], B[16]);
  nor g41 (n_177, A[17], B[17]);
  nand g42 (n_178, A[17], B[17]);
  nor g43 (n_187, A[18], B[18]);
  nand g44 (n_182, A[18], B[18]);
  nor g45 (n_183, A[19], B[19]);
  nand g46 (n_184, A[19], B[19]);
  nor g47 (n_193, A[20], B[20]);
  nand g48 (n_188, A[20], B[20]);
  nor g49 (n_189, A[21], B[21]);
  nand g50 (n_190, A[21], B[21]);
  nor g51 (n_199, A[22], B[22]);
  nand g52 (n_194, A[22], B[22]);
  nor g53 (n_195, A[23], B[23]);
  nand g54 (n_196, A[23], B[23]);
  nor g55 (n_205, A[24], B[24]);
  nand g56 (n_200, A[24], B[24]);
  nor g57 (n_201, A[25], B[25]);
  nand g58 (n_202, A[25], B[25]);
  nor g59 (n_211, A[26], B[26]);
  nand g60 (n_206, A[26], B[26]);
  nor g61 (n_207, A[27], B[27]);
  nand g62 (n_208, A[27], B[27]);
  nor g63 (n_217, A[28], B[28]);
  nand g64 (n_212, A[28], B[28]);
  nor g65 (n_213, A[29], B[29]);
  nand g66 (n_214, A[29], B[29]);
  nor g67 (n_223, A[30], B[30]);
  nand g68 (n_218, A[30], B[30]);
  nor g69 (n_219, A[31], B[31]);
  nand g70 (n_220, A[31], B[31]);
  nor g71 (n_229, A[32], B[32]);
  nand g72 (n_224, A[32], B[32]);
  nor g73 (n_225, A[33], B[33]);
  nand g74 (n_226, A[33], B[33]);
  nor g75 (n_235, A[34], B[34]);
  nand g76 (n_230, A[34], B[34]);
  nor g77 (n_231, A[35], B[35]);
  nand g78 (n_232, A[35], B[35]);
  nor g79 (n_241, A[36], B[36]);
  nand g80 (n_236, A[36], B[36]);
  nor g81 (n_237, A[37], B[37]);
  nand g82 (n_238, A[37], B[37]);
  nor g83 (n_247, A[38], B[38]);
  nand g84 (n_242, A[38], B[38]);
  nand g89 (n_248, n_132, n_133);
  nor g90 (n_137, n_134, n_135);
  nor g93 (n_251, n_139, n_135);
  nor g94 (n_143, n_140, n_141);
  nor g97 (n_257, n_145, n_141);
  nor g98 (n_149, n_146, n_147);
  nor g101 (n_259, n_151, n_147);
  nor g102 (n_155, n_152, n_153);
  nor g105 (n_267, n_157, n_153);
  nor g106 (n_161, n_158, n_159);
  nor g109 (n_269, n_163, n_159);
  nor g110 (n_167, n_164, n_165);
  nor g113 (n_277, n_169, n_165);
  nor g114 (n_173, n_170, n_171);
  nor g117 (n_279, n_175, n_171);
  nor g118 (n_179, n_176, n_177);
  nor g121 (n_287, n_181, n_177);
  nor g122 (n_185, n_182, n_183);
  nor g125 (n_289, n_187, n_183);
  nor g126 (n_191, n_188, n_189);
  nor g129 (n_297, n_193, n_189);
  nor g130 (n_197, n_194, n_195);
  nor g133 (n_299, n_199, n_195);
  nor g134 (n_203, n_200, n_201);
  nor g137 (n_307, n_205, n_201);
  nor g138 (n_209, n_206, n_207);
  nor g141 (n_309, n_211, n_207);
  nor g142 (n_215, n_212, n_213);
  nor g145 (n_317, n_217, n_213);
  nor g146 (n_221, n_218, n_219);
  nor g149 (n_319, n_223, n_219);
  nor g150 (n_227, n_224, n_225);
  nor g153 (n_327, n_229, n_225);
  nor g154 (n_233, n_230, n_231);
  nor g157 (n_329, n_235, n_231);
  nor g158 (n_239, n_236, n_237);
  nor g161 (n_337, n_241, n_237);
  nor g162 (n_245, n_242, n_243);
  nor g165 (n_339, n_247, n_243);
  nand g168 (n_551, n_134, n_250);
  nand g169 (n_253, n_251, n_248);
  nand g170 (n_344, n_252, n_253);
  nor g171 (n_255, n_151, n_254);
  nand g180 (n_352, n_257, n_259);
  nor g181 (n_265, n_163, n_264);
  nand g190 (n_359, n_267, n_269);
  nor g191 (n_275, n_175, n_274);
  nand g200 (n_367, n_277, n_279);
  nor g201 (n_285, n_187, n_284);
  nand g210 (n_374, n_287, n_289);
  nor g211 (n_295, n_199, n_294);
  nand g220 (n_382, n_297, n_299);
  nor g221 (n_305, n_211, n_304);
  nand g230 (n_389, n_307, n_309);
  nor g231 (n_315, n_223, n_314);
  nand g240 (n_397, n_317, n_319);
  nor g241 (n_325, n_235, n_324);
  nand g250 (n_404, n_327, n_329);
  nor g251 (n_335, n_247, n_334);
  nand g260 (n_412, n_337, n_339);
  nand g263 (n_555, n_140, n_346);
  nand g264 (n_347, n_257, n_344);
  nand g265 (n_557, n_254, n_347);
  nand g268 (n_560, n_350, n_351);
  nand g271 (n_416, n_354, n_355);
  nor g272 (n_357, n_169, n_356);
  nor g275 (n_426, n_169, n_359);
  nor g281 (n_365, n_363, n_356);
  nor g284 (n_432, n_359, n_363);
  nor g285 (n_369, n_367, n_356);
  nor g288 (n_435, n_359, n_367);
  nor g289 (n_372, n_193, n_371);
  nor g292 (n_484, n_193, n_374);
  nor g298 (n_380, n_378, n_371);
  nor g301 (n_490, n_374, n_378);
  nor g302 (n_384, n_382, n_371);
  nor g305 (n_441, n_374, n_382);
  nor g306 (n_387, n_217, n_386);
  nor g309 (n_454, n_217, n_389);
  nor g315 (n_395, n_393, n_386);
  nor g318 (n_464, n_389, n_393);
  nor g319 (n_399, n_397, n_386);
  nor g322 (n_469, n_389, n_397);
  nor g323 (n_402, n_241, n_401);
  nor g326 (n_536, n_241, n_404);
  nor g332 (n_410, n_408, n_401);
  nor g335 (n_542, n_404, n_408);
  nor g336 (n_414, n_412, n_401);
  nor g339 (n_545, n_404, n_412);
  nand g342 (n_564, n_152, n_418);
  nand g343 (n_419, n_267, n_416);
  nand g344 (n_566, n_264, n_419);
  nand g347 (n_569, n_422, n_423);
  nand g350 (n_572, n_356, n_425);
  nand g351 (n_428, n_426, n_416);
  nand g352 (n_575, n_427, n_428);
  nand g353 (n_431, n_429, n_416);
  nand g354 (n_577, n_430, n_431);
  nand g355 (n_434, n_432, n_416);
  nand g356 (n_580, n_433, n_434);
  nand g357 (n_437, n_435, n_416);
  nand g358 (n_474, n_436, n_437);
  nor g359 (n_439, n_205, n_438);
  nand g368 (n_498, n_307, n_441);
  nor g369 (n_448, n_446, n_438);
  nor g374 (n_451, n_389, n_438);
  nand g383 (n_510, n_441, n_454);
  nand g388 (n_514, n_441, n_459);
  nand g393 (n_518, n_441, n_464);
  nand g398 (n_522, n_441, n_469);
  nand g401 (n_584, n_176, n_476);
  nand g402 (n_477, n_287, n_474);
  nand g403 (n_586, n_284, n_477);
  nand g406 (n_589, n_480, n_481);
  nand g409 (n_592, n_371, n_483);
  nand g410 (n_486, n_484, n_474);
  nand g411 (n_595, n_485, n_486);
  nand g412 (n_489, n_487, n_474);
  nand g413 (n_597, n_488, n_489);
  nand g414 (n_492, n_490, n_474);
  nand g415 (n_600, n_491, n_492);
  nand g416 (n_493, n_441, n_474);
  nand g417 (n_602, n_438, n_493);
  nand g420 (n_605, n_496, n_497);
  nand g423 (n_607, n_500, n_501);
  nand g426 (n_610, n_504, n_505);
  nand g429 (n_613, n_508, n_509);
  nand g432 (n_616, n_512, n_513);
  nand g435 (n_618, n_516, n_517);
  nand g438 (n_621, n_520, n_521);
  nand g441 (n_526, n_524, n_525);
  nand g444 (n_625, n_224, n_528);
  nand g445 (n_529, n_327, n_526);
  nand g446 (n_627, n_324, n_529);
  nand g449 (n_630, n_532, n_533);
  nand g452 (n_633, n_401, n_535);
  nand g453 (n_538, n_536, n_526);
  nand g454 (n_636, n_537, n_538);
  nand g455 (n_541, n_539, n_526);
  nand g456 (n_638, n_540, n_541);
  nand g457 (n_544, n_542, n_526);
  nand g458 (n_641, n_543, n_544);
  nand g459 (n_547, n_545, n_526);
  nand g460 (n_125, n_546, n_547);
  xnor g464 (Z[2], n_248, n_549);
  xnor g467 (Z[3], n_551, n_552);
  xnor g469 (Z[4], n_344, n_553);
  xnor g472 (Z[5], n_555, n_556);
  xnor g474 (Z[6], n_557, n_558);
  xnor g477 (Z[7], n_560, n_561);
  xnor g479 (Z[8], n_416, n_562);
  xnor g482 (Z[9], n_564, n_565);
  xnor g484 (Z[10], n_566, n_567);
  xnor g487 (Z[11], n_569, n_570);
  xnor g490 (Z[12], n_572, n_573);
  xnor g493 (Z[13], n_575, n_576);
  xnor g495 (Z[14], n_577, n_578);
  xnor g498 (Z[15], n_580, n_581);
  xnor g500 (Z[16], n_474, n_582);
  xnor g503 (Z[17], n_584, n_585);
  xnor g505 (Z[18], n_586, n_587);
  xnor g508 (Z[19], n_589, n_590);
  xnor g511 (Z[20], n_592, n_593);
  xnor g514 (Z[21], n_595, n_596);
  xnor g516 (Z[22], n_597, n_598);
  xnor g519 (Z[23], n_600, n_601);
  xnor g521 (Z[24], n_602, n_603);
  xnor g524 (Z[25], n_605, n_606);
  xnor g526 (Z[26], n_607, n_608);
  xnor g529 (Z[27], n_610, n_611);
  xnor g532 (Z[28], n_613, n_614);
  xnor g535 (Z[29], n_616, n_617);
  xnor g537 (Z[30], n_618, n_619);
  xnor g540 (Z[31], n_621, n_622);
  xnor g542 (Z[32], n_526, n_623);
  xnor g545 (Z[33], n_625, n_626);
  xnor g547 (Z[34], n_627, n_628);
  xnor g550 (Z[35], n_630, n_631);
  xnor g553 (Z[36], n_633, n_634);
  xnor g556 (Z[37], n_636, n_637);
  xnor g558 (Z[38], n_638, n_639);
  xnor g561 (Z[39], n_641, n_642);
  and g564 (n_243, A[39], B[39]);
  or g565 (n_244, A[39], B[39]);
  and g566 (n_324, wc, n_226);
  not gc (wc, n_227);
  and g567 (n_331, wc0, n_232);
  not gc0 (wc0, n_233);
  and g568 (n_334, wc1, n_238);
  not gc1 (wc1, n_239);
  and g569 (n_284, wc2, n_178);
  not gc2 (wc2, n_179);
  and g570 (n_291, wc3, n_184);
  not gc3 (wc3, n_185);
  and g571 (n_294, wc4, n_190);
  not gc4 (wc4, n_191);
  and g572 (n_301, wc5, n_196);
  not gc5 (wc5, n_197);
  and g573 (n_304, wc6, n_202);
  not gc6 (wc6, n_203);
  and g574 (n_311, wc7, n_208);
  not gc7 (wc7, n_209);
  and g575 (n_314, wc8, n_214);
  not gc8 (wc8, n_215);
  and g576 (n_321, wc9, n_220);
  not gc9 (wc9, n_221);
  and g577 (n_264, wc10, n_154);
  not gc10 (wc10, n_155);
  and g578 (n_271, wc11, n_160);
  not gc11 (wc11, n_161);
  and g579 (n_274, wc12, n_166);
  not gc12 (wc12, n_167);
  and g580 (n_281, wc13, n_172);
  not gc13 (wc13, n_173);
  and g581 (n_254, wc14, n_142);
  not gc14 (wc14, n_143);
  and g582 (n_261, wc15, n_148);
  not gc15 (wc15, n_149);
  and g583 (n_252, wc16, n_136);
  not gc16 (wc16, n_137);
  or g584 (n_133, n_126, n_129);
  or g585 (n_348, wc17, n_151);
  not gc17 (wc17, n_257);
  or g586 (n_420, wc18, n_163);
  not gc18 (wc18, n_267);
  or g587 (n_363, wc19, n_175);
  not gc19 (wc19, n_277);
  or g588 (n_478, wc20, n_187);
  not gc20 (wc20, n_287);
  or g589 (n_378, wc21, n_199);
  not gc21 (wc21, n_297);
  or g590 (n_446, wc22, n_211);
  not gc22 (wc22, n_307);
  or g591 (n_393, wc23, n_223);
  not gc23 (wc23, n_317);
  or g592 (n_530, wc24, n_235);
  not gc24 (wc24, n_327);
  or g593 (n_408, wc25, n_247);
  not gc25 (wc25, n_337);
  or g594 (n_548, wc26, n_129);
  not gc26 (wc26, n_132);
  or g595 (n_549, wc27, n_139);
  not gc27 (wc27, n_134);
  or g596 (n_552, wc28, n_135);
  not gc28 (wc28, n_136);
  or g597 (n_553, wc29, n_145);
  not gc29 (wc29, n_140);
  or g598 (n_556, wc30, n_141);
  not gc30 (wc30, n_142);
  or g599 (n_558, wc31, n_151);
  not gc31 (wc31, n_146);
  or g600 (n_561, wc32, n_147);
  not gc32 (wc32, n_148);
  or g601 (n_562, wc33, n_157);
  not gc33 (wc33, n_152);
  or g602 (n_565, wc34, n_153);
  not gc34 (wc34, n_154);
  or g603 (n_567, wc35, n_163);
  not gc35 (wc35, n_158);
  or g604 (n_570, wc36, n_159);
  not gc36 (wc36, n_160);
  or g605 (n_573, wc37, n_169);
  not gc37 (wc37, n_164);
  or g606 (n_576, wc38, n_165);
  not gc38 (wc38, n_166);
  or g607 (n_578, wc39, n_175);
  not gc39 (wc39, n_170);
  or g608 (n_581, wc40, n_171);
  not gc40 (wc40, n_172);
  or g609 (n_582, wc41, n_181);
  not gc41 (wc41, n_176);
  or g610 (n_585, wc42, n_177);
  not gc42 (wc42, n_178);
  or g611 (n_587, wc43, n_187);
  not gc43 (wc43, n_182);
  or g612 (n_590, wc44, n_183);
  not gc44 (wc44, n_184);
  or g613 (n_593, wc45, n_193);
  not gc45 (wc45, n_188);
  or g614 (n_596, wc46, n_189);
  not gc46 (wc46, n_190);
  or g615 (n_598, wc47, n_199);
  not gc47 (wc47, n_194);
  or g616 (n_601, wc48, n_195);
  not gc48 (wc48, n_196);
  or g617 (n_603, wc49, n_205);
  not gc49 (wc49, n_200);
  or g618 (n_606, wc50, n_201);
  not gc50 (wc50, n_202);
  or g619 (n_608, wc51, n_211);
  not gc51 (wc51, n_206);
  or g620 (n_611, wc52, n_207);
  not gc52 (wc52, n_208);
  or g621 (n_614, wc53, n_217);
  not gc53 (wc53, n_212);
  or g622 (n_617, wc54, n_213);
  not gc54 (wc54, n_214);
  or g623 (n_619, wc55, n_223);
  not gc55 (wc55, n_218);
  or g624 (n_622, wc56, n_219);
  not gc56 (wc56, n_220);
  or g625 (n_623, wc57, n_229);
  not gc57 (wc57, n_224);
  or g626 (n_626, wc58, n_225);
  not gc58 (wc58, n_226);
  or g627 (n_628, wc59, n_235);
  not gc59 (wc59, n_230);
  or g628 (n_631, wc60, n_231);
  not gc60 (wc60, n_232);
  or g629 (n_634, wc61, n_241);
  not gc61 (wc61, n_236);
  or g630 (n_637, wc62, n_237);
  not gc62 (wc62, n_238);
  or g631 (n_639, wc63, n_247);
  not gc63 (wc63, n_242);
  and g632 (n_332, wc64, n_329);
  not gc64 (wc64, n_324);
  and g633 (n_341, n_244, wc65);
  not gc65 (wc65, n_245);
  and g634 (n_292, wc66, n_289);
  not gc66 (wc66, n_284);
  and g635 (n_302, wc67, n_299);
  not gc67 (wc67, n_294);
  and g636 (n_312, wc68, n_309);
  not gc68 (wc68, n_304);
  and g637 (n_322, wc69, n_319);
  not gc69 (wc69, n_314);
  and g638 (n_272, wc70, n_269);
  not gc70 (wc70, n_264);
  and g639 (n_282, wc71, n_279);
  not gc71 (wc71, n_274);
  and g640 (n_262, wc72, n_259);
  not gc72 (wc72, n_254);
  and g641 (n_429, wc73, n_277);
  not gc73 (wc73, n_359);
  and g642 (n_487, wc74, n_297);
  not gc74 (wc74, n_374);
  and g643 (n_459, wc75, n_317);
  not gc75 (wc75, n_389);
  and g644 (n_539, wc76, n_337);
  not gc76 (wc76, n_404);
  xor g645 (Z[1], n_126, n_548);
  or g646 (n_642, wc77, n_243);
  not gc77 (wc77, n_244);
  and g647 (n_401, wc78, n_331);
  not gc78 (wc78, n_332);
  and g648 (n_342, wc79, n_339);
  not gc79 (wc79, n_334);
  and g649 (n_371, wc80, n_291);
  not gc80 (wc80, n_292);
  and g650 (n_383, wc81, n_301);
  not gc81 (wc81, n_302);
  and g651 (n_386, wc82, n_311);
  not gc82 (wc82, n_312);
  and g652 (n_398, wc83, n_321);
  not gc83 (wc83, n_322);
  and g653 (n_356, wc84, n_271);
  not gc84 (wc84, n_272);
  and g654 (n_368, wc85, n_281);
  not gc85 (wc85, n_282);
  and g655 (n_354, wc86, n_261);
  not gc86 (wc86, n_262);
  or g656 (n_250, wc87, n_139);
  not gc87 (wc87, n_248);
  and g657 (n_350, wc88, n_146);
  not gc88 (wc88, n_255);
  and g658 (n_422, wc89, n_158);
  not gc89 (wc89, n_265);
  and g659 (n_364, wc90, n_170);
  not gc90 (wc90, n_275);
  and g660 (n_480, wc91, n_182);
  not gc91 (wc91, n_285);
  and g661 (n_379, wc92, n_194);
  not gc92 (wc92, n_295);
  and g662 (n_447, wc93, n_206);
  not gc93 (wc93, n_305);
  and g663 (n_394, wc94, n_218);
  not gc94 (wc94, n_315);
  and g664 (n_532, wc95, n_230);
  not gc95 (wc95, n_325);
  and g665 (n_409, wc96, n_242);
  not gc96 (wc96, n_335);
  or g666 (n_494, wc97, n_205);
  not gc97 (wc97, n_441);
  or g667 (n_502, n_446, wc98);
  not gc98 (wc98, n_441);
  or g668 (n_506, wc99, n_389);
  not gc99 (wc99, n_441);
  and g669 (n_413, wc100, n_341);
  not gc100 (wc100, n_342);
  and g670 (n_361, wc101, n_277);
  not gc101 (wc101, n_356);
  and g671 (n_376, wc102, n_297);
  not gc102 (wc102, n_371);
  and g672 (n_391, wc103, n_317);
  not gc103 (wc103, n_386);
  and g673 (n_406, wc104, n_337);
  not gc104 (wc104, n_401);
  and g674 (n_438, n_383, wc105);
  not gc105 (wc105, n_384);
  and g675 (n_471, n_398, wc106);
  not gc106 (wc106, n_399);
  and g676 (n_436, n_368, wc107);
  not gc107 (wc107, n_369);
  or g677 (n_355, n_352, wc108);
  not gc108 (wc108, n_344);
  or g678 (n_346, wc109, n_145);
  not gc109 (wc109, n_344);
  or g679 (n_351, n_348, wc110);
  not gc110 (wc110, n_344);
  and g680 (n_427, wc111, n_164);
  not gc111 (wc111, n_357);
  and g681 (n_430, wc112, n_274);
  not gc112 (wc112, n_361);
  and g682 (n_433, n_364, wc113);
  not gc113 (wc113, n_365);
  and g683 (n_485, wc114, n_188);
  not gc114 (wc114, n_372);
  and g684 (n_488, wc115, n_294);
  not gc115 (wc115, n_376);
  and g685 (n_491, n_379, wc116);
  not gc116 (wc116, n_380);
  and g686 (n_456, wc117, n_212);
  not gc117 (wc117, n_387);
  and g687 (n_461, wc118, n_314);
  not gc118 (wc118, n_391);
  and g688 (n_466, n_394, wc119);
  not gc119 (wc119, n_395);
  and g689 (n_537, wc120, n_236);
  not gc120 (wc120, n_402);
  and g690 (n_540, wc121, n_334);
  not gc121 (wc121, n_406);
  and g691 (n_543, n_409, wc122);
  not gc122 (wc122, n_410);
  and g692 (n_546, n_413, wc123);
  not gc123 (wc123, n_414);
  and g693 (n_472, wc124, n_469);
  not gc124 (wc124, n_438);
  and g694 (n_444, wc125, n_307);
  not gc125 (wc125, n_438);
  and g695 (n_457, wc126, n_454);
  not gc126 (wc126, n_438);
  and g696 (n_462, wc127, n_459);
  not gc127 (wc127, n_438);
  and g697 (n_467, wc128, n_464);
  not gc128 (wc128, n_438);
  and g698 (n_524, wc129, n_471);
  not gc129 (wc129, n_472);
  or g699 (n_418, wc130, n_157);
  not gc130 (wc130, n_416);
  or g700 (n_423, n_420, wc131);
  not gc131 (wc131, n_416);
  or g701 (n_425, wc132, n_359);
  not gc132 (wc132, n_416);
  and g702 (n_496, wc133, n_200);
  not gc133 (wc133, n_439);
  and g703 (n_500, wc134, n_304);
  not gc134 (wc134, n_444);
  and g704 (n_504, n_447, wc135);
  not gc135 (wc135, n_448);
  and g705 (n_508, n_386, wc136);
  not gc136 (wc136, n_451);
  and g706 (n_512, wc137, n_456);
  not gc137 (wc137, n_457);
  and g707 (n_516, wc138, n_461);
  not gc138 (wc138, n_462);
  and g708 (n_520, wc139, n_466);
  not gc139 (wc139, n_467);
  or g709 (n_525, n_522, wc140);
  not gc140 (wc140, n_474);
  or g710 (n_476, wc141, n_181);
  not gc141 (wc141, n_474);
  or g711 (n_481, n_478, wc142);
  not gc142 (wc142, n_474);
  or g712 (n_483, wc143, n_374);
  not gc143 (wc143, n_474);
  or g713 (n_497, n_494, wc144);
  not gc144 (wc144, n_474);
  or g714 (n_501, n_498, wc145);
  not gc145 (wc145, n_474);
  or g715 (n_505, n_502, wc146);
  not gc146 (wc146, n_474);
  or g716 (n_509, n_506, wc147);
  not gc147 (wc147, n_474);
  or g717 (n_513, n_510, wc148);
  not gc148 (wc148, n_474);
  or g718 (n_517, n_514, wc149);
  not gc149 (wc149, n_474);
  or g719 (n_521, n_518, wc150);
  not gc150 (wc150, n_474);
  or g720 (n_528, wc151, n_229);
  not gc151 (wc151, n_526);
  or g721 (n_533, n_530, wc152);
  not gc152 (wc152, n_526);
  or g722 (n_535, wc153, n_404);
  not gc153 (wc153, n_526);
endmodule

module add_signed_454_GENERIC(A, B, Z);
  input [39:0] A, B;
  output [40:0] Z;
  wire [39:0] A, B;
  wire [40:0] Z;
  add_signed_454_GENERIC_REAL g1(.A ({A[38], A[38:0]}), .B ({B[38],
       B[38:0]}), .Z (Z));
endmodule

module add_signed_468_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [38:0] A, B;
  output [39:0] Z;
  wire [38:0] A, B;
  wire [39:0] Z;
  wire n_122, n_123, n_126, n_129, n_130, n_131, n_132, n_133;
  wire n_134, n_136, n_137, n_138, n_139, n_140, n_142, n_143;
  wire n_144, n_145, n_146, n_148, n_149, n_150, n_151, n_152;
  wire n_154, n_155, n_156, n_157, n_158, n_160, n_161, n_162;
  wire n_163, n_164, n_166, n_167, n_168, n_169, n_170, n_172;
  wire n_173, n_174, n_175, n_176, n_178, n_179, n_180, n_181;
  wire n_182, n_184, n_185, n_186, n_187, n_188, n_190, n_191;
  wire n_192, n_193, n_194, n_196, n_197, n_198, n_199, n_200;
  wire n_202, n_203, n_204, n_205, n_206, n_208, n_209, n_210;
  wire n_211, n_212, n_214, n_215, n_216, n_217, n_218, n_220;
  wire n_221, n_222, n_223, n_224, n_226, n_227, n_228, n_229;
  wire n_230, n_232, n_233, n_234, n_235, n_236, n_238, n_239;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_248, n_250;
  wire n_252, n_253, n_255, n_256, n_258, n_260, n_262, n_263;
  wire n_265, n_266, n_268, n_270, n_272, n_273, n_275, n_276;
  wire n_278, n_280, n_282, n_283, n_285, n_286, n_288, n_290;
  wire n_292, n_293, n_295, n_296, n_298, n_300, n_302, n_303;
  wire n_305, n_306, n_308, n_310, n_312, n_313, n_315, n_316;
  wire n_318, n_320, n_322, n_323, n_325, n_326, n_327, n_328;
  wire n_330, n_332, n_334, n_335, n_336, n_338, n_339, n_340;
  wire n_342, n_343, n_344, n_345, n_347, n_349, n_351, n_352;
  wire n_353, n_355, n_356, n_357, n_359, n_360, n_362, n_364;
  wire n_366, n_367, n_368, n_370, n_371, n_372, n_374, n_375;
  wire n_377, n_379, n_381, n_382, n_383, n_385, n_386, n_387;
  wire n_389, n_390, n_392, n_394, n_396, n_397, n_398, n_400;
  wire n_402, n_403, n_404, n_406, n_407, n_409, n_410, n_411;
  wire n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419;
  wire n_420, n_421, n_422, n_423, n_425, n_428, n_430, n_431;
  wire n_432, n_435, n_438, n_440, n_441, n_443, n_445, n_446;
  wire n_448, n_450, n_451, n_453, n_455, n_456, n_458, n_460;
  wire n_461, n_462, n_464, n_465, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_480, n_481, n_482, n_484, n_485, n_486, n_488, n_489;
  wire n_490, n_492, n_493, n_494, n_496, n_497, n_498, n_500;
  wire n_501, n_502, n_504, n_505, n_506, n_508, n_509, n_510;
  wire n_512, n_513, n_514, n_516, n_517, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_532, n_533, n_534, n_536, n_537, n_538, n_539;
  wire n_541, n_542, n_543, n_545, n_546, n_547, n_548, n_550;
  wire n_551, n_553, n_554, n_556, n_557, n_558, n_559, n_561;
  wire n_562, n_563, n_565, n_566, n_567, n_568, n_570, n_571;
  wire n_573, n_574, n_576, n_577, n_578, n_579, n_581, n_582;
  wire n_583, n_584, n_586, n_587, n_588, n_589, n_591, n_592;
  wire n_594, n_595, n_597, n_598, n_599, n_600, n_602, n_603;
  wire n_604, n_606, n_607, n_608, n_609, n_611, n_612, n_614;
  wire n_615, n_617, n_618, n_619, n_620;
  not g3 (Z[39], n_122);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_123, A[0], B[0]);
  nor g9 (n_126, A[1], B[1]);
  nand g10 (n_129, A[1], B[1]);
  nor g11 (n_136, A[2], B[2]);
  nand g12 (n_131, A[2], B[2]);
  nor g13 (n_132, A[3], B[3]);
  nand g14 (n_133, A[3], B[3]);
  nor g15 (n_142, A[4], B[4]);
  nand g16 (n_137, A[4], B[4]);
  nor g17 (n_138, A[5], B[5]);
  nand g18 (n_139, A[5], B[5]);
  nor g19 (n_148, A[6], B[6]);
  nand g20 (n_143, A[6], B[6]);
  nor g21 (n_144, A[7], B[7]);
  nand g22 (n_145, A[7], B[7]);
  nor g23 (n_154, A[8], B[8]);
  nand g24 (n_149, A[8], B[8]);
  nor g25 (n_150, A[9], B[9]);
  nand g26 (n_151, A[9], B[9]);
  nor g27 (n_160, A[10], B[10]);
  nand g28 (n_155, A[10], B[10]);
  nor g29 (n_156, A[11], B[11]);
  nand g30 (n_157, A[11], B[11]);
  nor g31 (n_166, A[12], B[12]);
  nand g32 (n_161, A[12], B[12]);
  nor g33 (n_162, A[13], B[13]);
  nand g34 (n_163, A[13], B[13]);
  nor g35 (n_172, A[14], B[14]);
  nand g36 (n_167, A[14], B[14]);
  nor g37 (n_168, A[15], B[15]);
  nand g38 (n_169, A[15], B[15]);
  nor g39 (n_178, A[16], B[16]);
  nand g40 (n_173, A[16], B[16]);
  nor g41 (n_174, A[17], B[17]);
  nand g42 (n_175, A[17], B[17]);
  nor g43 (n_184, A[18], B[18]);
  nand g44 (n_179, A[18], B[18]);
  nor g45 (n_180, A[19], B[19]);
  nand g46 (n_181, A[19], B[19]);
  nor g47 (n_190, A[20], B[20]);
  nand g48 (n_185, A[20], B[20]);
  nor g49 (n_186, A[21], B[21]);
  nand g50 (n_187, A[21], B[21]);
  nor g51 (n_196, A[22], B[22]);
  nand g52 (n_191, A[22], B[22]);
  nor g53 (n_192, A[23], B[23]);
  nand g54 (n_193, A[23], B[23]);
  nor g55 (n_202, A[24], B[24]);
  nand g56 (n_197, A[24], B[24]);
  nor g57 (n_198, A[25], B[25]);
  nand g58 (n_199, A[25], B[25]);
  nor g59 (n_208, A[26], B[26]);
  nand g60 (n_203, A[26], B[26]);
  nor g61 (n_204, A[27], B[27]);
  nand g62 (n_205, A[27], B[27]);
  nor g63 (n_214, A[28], B[28]);
  nand g64 (n_209, A[28], B[28]);
  nor g65 (n_210, A[29], B[29]);
  nand g66 (n_211, A[29], B[29]);
  nor g67 (n_220, A[30], B[30]);
  nand g68 (n_215, A[30], B[30]);
  nor g69 (n_216, A[31], B[31]);
  nand g70 (n_217, A[31], B[31]);
  nor g71 (n_226, A[32], B[32]);
  nand g72 (n_221, A[32], B[32]);
  nor g73 (n_222, A[33], B[33]);
  nand g74 (n_223, A[33], B[33]);
  nor g75 (n_232, A[34], B[34]);
  nand g76 (n_227, A[34], B[34]);
  nor g77 (n_228, A[35], B[35]);
  nand g78 (n_229, A[35], B[35]);
  nor g79 (n_238, A[36], B[36]);
  nand g80 (n_233, A[36], B[36]);
  nor g81 (n_234, A[37], B[37]);
  nand g82 (n_235, A[37], B[37]);
  nand g87 (n_239, n_129, n_130);
  nor g88 (n_134, n_131, n_132);
  nor g91 (n_242, n_136, n_132);
  nor g92 (n_140, n_137, n_138);
  nor g95 (n_248, n_142, n_138);
  nor g96 (n_146, n_143, n_144);
  nor g99 (n_250, n_148, n_144);
  nor g100 (n_152, n_149, n_150);
  nor g103 (n_258, n_154, n_150);
  nor g104 (n_158, n_155, n_156);
  nor g107 (n_260, n_160, n_156);
  nor g108 (n_164, n_161, n_162);
  nor g111 (n_268, n_166, n_162);
  nor g112 (n_170, n_167, n_168);
  nor g115 (n_270, n_172, n_168);
  nor g116 (n_176, n_173, n_174);
  nor g119 (n_278, n_178, n_174);
  nor g120 (n_182, n_179, n_180);
  nor g123 (n_280, n_184, n_180);
  nor g124 (n_188, n_185, n_186);
  nor g127 (n_288, n_190, n_186);
  nor g128 (n_194, n_191, n_192);
  nor g131 (n_290, n_196, n_192);
  nor g132 (n_200, n_197, n_198);
  nor g135 (n_298, n_202, n_198);
  nor g136 (n_206, n_203, n_204);
  nor g139 (n_300, n_208, n_204);
  nor g140 (n_212, n_209, n_210);
  nor g143 (n_308, n_214, n_210);
  nor g144 (n_218, n_215, n_216);
  nor g147 (n_310, n_220, n_216);
  nor g148 (n_224, n_221, n_222);
  nor g151 (n_318, n_226, n_222);
  nor g152 (n_230, n_227, n_228);
  nor g155 (n_320, n_232, n_228);
  nor g156 (n_236, n_233, n_234);
  nor g159 (n_330, n_238, n_234);
  nand g162 (n_532, n_131, n_241);
  nand g163 (n_244, n_242, n_239);
  nand g164 (n_332, n_243, n_244);
  nor g165 (n_246, n_148, n_245);
  nand g174 (n_340, n_248, n_250);
  nor g175 (n_256, n_160, n_255);
  nand g184 (n_347, n_258, n_260);
  nor g185 (n_266, n_172, n_265);
  nand g194 (n_355, n_268, n_270);
  nor g195 (n_276, n_184, n_275);
  nand g204 (n_362, n_278, n_280);
  nor g205 (n_286, n_196, n_285);
  nand g214 (n_370, n_288, n_290);
  nor g215 (n_296, n_208, n_295);
  nand g224 (n_377, n_298, n_300);
  nor g225 (n_306, n_220, n_305);
  nand g234 (n_385, n_308, n_310);
  nor g235 (n_316, n_232, n_315);
  nand g244 (n_392, n_318, n_320);
  nor g245 (n_328, n_325, n_326);
  nand g252 (n_536, n_137, n_334);
  nand g253 (n_335, n_248, n_332);
  nand g254 (n_538, n_245, n_335);
  nand g257 (n_541, n_338, n_339);
  nand g260 (n_400, n_342, n_343);
  nor g261 (n_345, n_166, n_344);
  nor g264 (n_410, n_166, n_347);
  nor g270 (n_353, n_351, n_344);
  nor g273 (n_416, n_347, n_351);
  nor g274 (n_357, n_355, n_344);
  nor g277 (n_419, n_347, n_355);
  nor g278 (n_360, n_190, n_359);
  nor g281 (n_468, n_190, n_362);
  nor g287 (n_368, n_366, n_359);
  nor g290 (n_474, n_362, n_366);
  nor g291 (n_372, n_370, n_359);
  nor g294 (n_425, n_362, n_370);
  nor g295 (n_375, n_214, n_374);
  nor g298 (n_438, n_214, n_377);
  nor g304 (n_383, n_381, n_374);
  nor g307 (n_448, n_377, n_381);
  nor g308 (n_387, n_385, n_374);
  nor g311 (n_453, n_377, n_385);
  nor g312 (n_390, n_238, n_389);
  nor g315 (n_520, n_238, n_392);
  nor g321 (n_398, n_396, n_389);
  nor g324 (n_526, n_392, n_396);
  nand g327 (n_545, n_149, n_402);
  nand g328 (n_403, n_258, n_400);
  nand g329 (n_547, n_255, n_403);
  nand g332 (n_550, n_406, n_407);
  nand g335 (n_553, n_344, n_409);
  nand g336 (n_412, n_410, n_400);
  nand g337 (n_556, n_411, n_412);
  nand g338 (n_415, n_413, n_400);
  nand g339 (n_558, n_414, n_415);
  nand g340 (n_418, n_416, n_400);
  nand g341 (n_561, n_417, n_418);
  nand g342 (n_421, n_419, n_400);
  nand g343 (n_458, n_420, n_421);
  nor g344 (n_423, n_202, n_422);
  nand g353 (n_482, n_298, n_425);
  nor g354 (n_432, n_430, n_422);
  nor g359 (n_435, n_377, n_422);
  nand g368 (n_494, n_425, n_438);
  nand g373 (n_498, n_425, n_443);
  nand g378 (n_502, n_425, n_448);
  nand g383 (n_506, n_425, n_453);
  nand g386 (n_565, n_173, n_460);
  nand g387 (n_461, n_278, n_458);
  nand g388 (n_567, n_275, n_461);
  nand g391 (n_570, n_464, n_465);
  nand g394 (n_573, n_359, n_467);
  nand g395 (n_470, n_468, n_458);
  nand g396 (n_576, n_469, n_470);
  nand g397 (n_473, n_471, n_458);
  nand g398 (n_578, n_472, n_473);
  nand g399 (n_476, n_474, n_458);
  nand g400 (n_581, n_475, n_476);
  nand g401 (n_477, n_425, n_458);
  nand g402 (n_583, n_422, n_477);
  nand g405 (n_586, n_480, n_481);
  nand g408 (n_588, n_484, n_485);
  nand g411 (n_591, n_488, n_489);
  nand g414 (n_594, n_492, n_493);
  nand g417 (n_597, n_496, n_497);
  nand g420 (n_599, n_500, n_501);
  nand g423 (n_602, n_504, n_505);
  nand g426 (n_510, n_508, n_509);
  nand g429 (n_606, n_221, n_512);
  nand g430 (n_513, n_318, n_510);
  nand g431 (n_608, n_315, n_513);
  nand g434 (n_611, n_516, n_517);
  nand g437 (n_614, n_389, n_519);
  nand g438 (n_522, n_520, n_510);
  nand g439 (n_617, n_521, n_522);
  nand g440 (n_525, n_523, n_510);
  nand g441 (n_619, n_524, n_525);
  nand g442 (n_528, n_526, n_510);
  nand g443 (n_122, n_527, n_528);
  xnor g447 (Z[2], n_239, n_530);
  xnor g450 (Z[3], n_532, n_533);
  xnor g452 (Z[4], n_332, n_534);
  xnor g455 (Z[5], n_536, n_537);
  xnor g457 (Z[6], n_538, n_539);
  xnor g460 (Z[7], n_541, n_542);
  xnor g462 (Z[8], n_400, n_543);
  xnor g465 (Z[9], n_545, n_546);
  xnor g467 (Z[10], n_547, n_548);
  xnor g470 (Z[11], n_550, n_551);
  xnor g473 (Z[12], n_553, n_554);
  xnor g476 (Z[13], n_556, n_557);
  xnor g478 (Z[14], n_558, n_559);
  xnor g481 (Z[15], n_561, n_562);
  xnor g483 (Z[16], n_458, n_563);
  xnor g486 (Z[17], n_565, n_566);
  xnor g488 (Z[18], n_567, n_568);
  xnor g491 (Z[19], n_570, n_571);
  xnor g494 (Z[20], n_573, n_574);
  xnor g497 (Z[21], n_576, n_577);
  xnor g499 (Z[22], n_578, n_579);
  xnor g502 (Z[23], n_581, n_582);
  xnor g504 (Z[24], n_583, n_584);
  xnor g507 (Z[25], n_586, n_587);
  xnor g509 (Z[26], n_588, n_589);
  xnor g512 (Z[27], n_591, n_592);
  xnor g515 (Z[28], n_594, n_595);
  xnor g518 (Z[29], n_597, n_598);
  xnor g520 (Z[30], n_599, n_600);
  xnor g523 (Z[31], n_602, n_603);
  xnor g525 (Z[32], n_510, n_604);
  xnor g528 (Z[33], n_606, n_607);
  xnor g530 (Z[34], n_608, n_609);
  xnor g533 (Z[35], n_611, n_612);
  xnor g536 (Z[36], n_614, n_615);
  xnor g539 (Z[37], n_617, n_618);
  xnor g541 (Z[38], n_619, n_620);
  and g544 (n_325, A[38], B[38]);
  or g545 (n_327, A[38], B[38]);
  and g546 (n_315, wc, n_223);
  not gc (wc, n_224);
  and g547 (n_322, wc0, n_229);
  not gc0 (wc0, n_230);
  and g548 (n_326, wc1, n_235);
  not gc1 (wc1, n_236);
  and g549 (n_275, wc2, n_175);
  not gc2 (wc2, n_176);
  and g550 (n_282, wc3, n_181);
  not gc3 (wc3, n_182);
  and g551 (n_285, wc4, n_187);
  not gc4 (wc4, n_188);
  and g552 (n_292, wc5, n_193);
  not gc5 (wc5, n_194);
  and g553 (n_295, wc6, n_199);
  not gc6 (wc6, n_200);
  and g554 (n_302, wc7, n_205);
  not gc7 (wc7, n_206);
  and g555 (n_305, wc8, n_211);
  not gc8 (wc8, n_212);
  and g556 (n_312, wc9, n_217);
  not gc9 (wc9, n_218);
  and g557 (n_255, wc10, n_151);
  not gc10 (wc10, n_152);
  and g558 (n_262, wc11, n_157);
  not gc11 (wc11, n_158);
  and g559 (n_265, wc12, n_163);
  not gc12 (wc12, n_164);
  and g560 (n_272, wc13, n_169);
  not gc13 (wc13, n_170);
  and g561 (n_245, wc14, n_139);
  not gc14 (wc14, n_140);
  and g562 (n_252, wc15, n_145);
  not gc15 (wc15, n_146);
  and g563 (n_243, wc16, n_133);
  not gc16 (wc16, n_134);
  or g564 (n_130, n_123, n_126);
  or g565 (n_336, wc17, n_148);
  not gc17 (wc17, n_248);
  or g566 (n_404, wc18, n_160);
  not gc18 (wc18, n_258);
  or g567 (n_351, wc19, n_172);
  not gc19 (wc19, n_268);
  or g568 (n_462, wc20, n_184);
  not gc20 (wc20, n_278);
  or g569 (n_366, wc21, n_196);
  not gc21 (wc21, n_288);
  or g570 (n_430, wc22, n_208);
  not gc22 (wc22, n_298);
  or g571 (n_381, wc23, n_220);
  not gc23 (wc23, n_308);
  or g572 (n_514, wc24, n_232);
  not gc24 (wc24, n_318);
  or g573 (n_529, wc25, n_126);
  not gc25 (wc25, n_129);
  or g574 (n_530, wc26, n_136);
  not gc26 (wc26, n_131);
  or g575 (n_533, wc27, n_132);
  not gc27 (wc27, n_133);
  or g576 (n_534, wc28, n_142);
  not gc28 (wc28, n_137);
  or g577 (n_537, wc29, n_138);
  not gc29 (wc29, n_139);
  or g578 (n_539, wc30, n_148);
  not gc30 (wc30, n_143);
  or g579 (n_542, wc31, n_144);
  not gc31 (wc31, n_145);
  or g580 (n_543, wc32, n_154);
  not gc32 (wc32, n_149);
  or g581 (n_546, wc33, n_150);
  not gc33 (wc33, n_151);
  or g582 (n_548, wc34, n_160);
  not gc34 (wc34, n_155);
  or g583 (n_551, wc35, n_156);
  not gc35 (wc35, n_157);
  or g584 (n_554, wc36, n_166);
  not gc36 (wc36, n_161);
  or g585 (n_557, wc37, n_162);
  not gc37 (wc37, n_163);
  or g586 (n_559, wc38, n_172);
  not gc38 (wc38, n_167);
  or g587 (n_562, wc39, n_168);
  not gc39 (wc39, n_169);
  or g588 (n_563, wc40, n_178);
  not gc40 (wc40, n_173);
  or g589 (n_566, wc41, n_174);
  not gc41 (wc41, n_175);
  or g590 (n_568, wc42, n_184);
  not gc42 (wc42, n_179);
  or g591 (n_571, wc43, n_180);
  not gc43 (wc43, n_181);
  or g592 (n_574, wc44, n_190);
  not gc44 (wc44, n_185);
  or g593 (n_577, wc45, n_186);
  not gc45 (wc45, n_187);
  or g594 (n_579, wc46, n_196);
  not gc46 (wc46, n_191);
  or g595 (n_582, wc47, n_192);
  not gc47 (wc47, n_193);
  or g596 (n_584, wc48, n_202);
  not gc48 (wc48, n_197);
  or g597 (n_587, wc49, n_198);
  not gc49 (wc49, n_199);
  or g598 (n_589, wc50, n_208);
  not gc50 (wc50, n_203);
  or g599 (n_592, wc51, n_204);
  not gc51 (wc51, n_205);
  or g600 (n_595, wc52, n_214);
  not gc52 (wc52, n_209);
  or g601 (n_598, wc53, n_210);
  not gc53 (wc53, n_211);
  or g602 (n_600, wc54, n_220);
  not gc54 (wc54, n_215);
  or g603 (n_603, wc55, n_216);
  not gc55 (wc55, n_217);
  or g604 (n_604, wc56, n_226);
  not gc56 (wc56, n_221);
  or g605 (n_607, wc57, n_222);
  not gc57 (wc57, n_223);
  or g606 (n_609, wc58, n_232);
  not gc58 (wc58, n_227);
  or g607 (n_612, wc59, n_228);
  not gc59 (wc59, n_229);
  or g608 (n_615, wc60, n_238);
  not gc60 (wc60, n_233);
  or g609 (n_618, wc61, n_234);
  not gc61 (wc61, n_235);
  or g610 (n_396, n_325, wc62);
  not gc62 (wc62, n_330);
  and g611 (n_323, wc63, n_320);
  not gc63 (wc63, n_315);
  and g612 (n_283, wc64, n_280);
  not gc64 (wc64, n_275);
  and g613 (n_293, wc65, n_290);
  not gc65 (wc65, n_285);
  and g614 (n_303, wc66, n_300);
  not gc66 (wc66, n_295);
  and g615 (n_313, wc67, n_310);
  not gc67 (wc67, n_305);
  and g616 (n_263, wc68, n_260);
  not gc68 (wc68, n_255);
  and g617 (n_273, wc69, n_270);
  not gc69 (wc69, n_265);
  and g618 (n_253, wc70, n_250);
  not gc70 (wc70, n_245);
  and g619 (n_413, wc71, n_268);
  not gc71 (wc71, n_347);
  and g620 (n_471, wc72, n_288);
  not gc72 (wc72, n_362);
  and g621 (n_443, wc73, n_308);
  not gc73 (wc73, n_377);
  and g622 (n_523, wc74, n_330);
  not gc74 (wc74, n_392);
  xor g623 (Z[1], n_123, n_529);
  or g624 (n_620, wc75, n_325);
  not gc75 (wc75, n_327);
  and g625 (n_389, wc76, n_322);
  not gc76 (wc76, n_323);
  and g626 (n_397, n_327, wc77);
  not gc77 (wc77, n_328);
  and g627 (n_359, wc78, n_282);
  not gc78 (wc78, n_283);
  and g628 (n_371, wc79, n_292);
  not gc79 (wc79, n_293);
  and g629 (n_374, wc80, n_302);
  not gc80 (wc80, n_303);
  and g630 (n_386, wc81, n_312);
  not gc81 (wc81, n_313);
  and g631 (n_344, wc82, n_262);
  not gc82 (wc82, n_263);
  and g632 (n_356, wc83, n_272);
  not gc83 (wc83, n_273);
  and g633 (n_342, wc84, n_252);
  not gc84 (wc84, n_253);
  or g634 (n_241, wc85, n_136);
  not gc85 (wc85, n_239);
  and g635 (n_338, wc86, n_143);
  not gc86 (wc86, n_246);
  and g636 (n_406, wc87, n_155);
  not gc87 (wc87, n_256);
  and g637 (n_352, wc88, n_167);
  not gc88 (wc88, n_266);
  and g638 (n_464, wc89, n_179);
  not gc89 (wc89, n_276);
  and g639 (n_367, wc90, n_191);
  not gc90 (wc90, n_286);
  and g640 (n_431, wc91, n_203);
  not gc91 (wc91, n_296);
  and g641 (n_382, wc92, n_215);
  not gc92 (wc92, n_306);
  and g642 (n_516, wc93, n_227);
  not gc93 (wc93, n_316);
  or g643 (n_478, wc94, n_202);
  not gc94 (wc94, n_425);
  or g644 (n_486, n_430, wc95);
  not gc95 (wc95, n_425);
  or g645 (n_490, wc96, n_377);
  not gc96 (wc96, n_425);
  and g646 (n_349, wc97, n_268);
  not gc97 (wc97, n_344);
  and g647 (n_364, wc98, n_288);
  not gc98 (wc98, n_359);
  and g648 (n_379, wc99, n_308);
  not gc99 (wc99, n_374);
  and g649 (n_394, wc100, n_330);
  not gc100 (wc100, n_389);
  and g650 (n_527, n_397, wc101);
  not gc101 (wc101, n_398);
  and g651 (n_422, n_371, wc102);
  not gc102 (wc102, n_372);
  and g652 (n_455, n_386, wc103);
  not gc103 (wc103, n_387);
  and g653 (n_420, n_356, wc104);
  not gc104 (wc104, n_357);
  or g654 (n_343, n_340, wc105);
  not gc105 (wc105, n_332);
  or g655 (n_334, wc106, n_142);
  not gc106 (wc106, n_332);
  or g656 (n_339, n_336, wc107);
  not gc107 (wc107, n_332);
  and g657 (n_411, wc108, n_161);
  not gc108 (wc108, n_345);
  and g658 (n_414, wc109, n_265);
  not gc109 (wc109, n_349);
  and g659 (n_417, n_352, wc110);
  not gc110 (wc110, n_353);
  and g660 (n_469, wc111, n_185);
  not gc111 (wc111, n_360);
  and g661 (n_472, wc112, n_285);
  not gc112 (wc112, n_364);
  and g662 (n_475, n_367, wc113);
  not gc113 (wc113, n_368);
  and g663 (n_440, wc114, n_209);
  not gc114 (wc114, n_375);
  and g664 (n_445, wc115, n_305);
  not gc115 (wc115, n_379);
  and g665 (n_450, n_382, wc116);
  not gc116 (wc116, n_383);
  and g666 (n_521, wc117, n_233);
  not gc117 (wc117, n_390);
  and g667 (n_524, wc118, n_326);
  not gc118 (wc118, n_394);
  and g668 (n_456, wc119, n_453);
  not gc119 (wc119, n_422);
  and g669 (n_428, wc120, n_298);
  not gc120 (wc120, n_422);
  and g670 (n_441, wc121, n_438);
  not gc121 (wc121, n_422);
  and g671 (n_446, wc122, n_443);
  not gc122 (wc122, n_422);
  and g672 (n_451, wc123, n_448);
  not gc123 (wc123, n_422);
  and g673 (n_508, wc124, n_455);
  not gc124 (wc124, n_456);
  or g674 (n_402, wc125, n_154);
  not gc125 (wc125, n_400);
  or g675 (n_407, n_404, wc126);
  not gc126 (wc126, n_400);
  or g676 (n_409, wc127, n_347);
  not gc127 (wc127, n_400);
  and g677 (n_480, wc128, n_197);
  not gc128 (wc128, n_423);
  and g678 (n_484, wc129, n_295);
  not gc129 (wc129, n_428);
  and g679 (n_488, n_431, wc130);
  not gc130 (wc130, n_432);
  and g680 (n_492, n_374, wc131);
  not gc131 (wc131, n_435);
  and g681 (n_496, wc132, n_440);
  not gc132 (wc132, n_441);
  and g682 (n_500, wc133, n_445);
  not gc133 (wc133, n_446);
  and g683 (n_504, wc134, n_450);
  not gc134 (wc134, n_451);
  or g684 (n_509, n_506, wc135);
  not gc135 (wc135, n_458);
  or g685 (n_460, wc136, n_178);
  not gc136 (wc136, n_458);
  or g686 (n_465, n_462, wc137);
  not gc137 (wc137, n_458);
  or g687 (n_467, wc138, n_362);
  not gc138 (wc138, n_458);
  or g688 (n_481, n_478, wc139);
  not gc139 (wc139, n_458);
  or g689 (n_485, n_482, wc140);
  not gc140 (wc140, n_458);
  or g690 (n_489, n_486, wc141);
  not gc141 (wc141, n_458);
  or g691 (n_493, n_490, wc142);
  not gc142 (wc142, n_458);
  or g692 (n_497, n_494, wc143);
  not gc143 (wc143, n_458);
  or g693 (n_501, n_498, wc144);
  not gc144 (wc144, n_458);
  or g694 (n_505, n_502, wc145);
  not gc145 (wc145, n_458);
  or g695 (n_512, wc146, n_226);
  not gc146 (wc146, n_510);
  or g696 (n_517, n_514, wc147);
  not gc147 (wc147, n_510);
  or g697 (n_519, wc148, n_392);
  not gc148 (wc148, n_510);
endmodule

module add_signed_468_GENERIC(A, B, Z);
  input [38:0] A, B;
  output [39:0] Z;
  wire [38:0] A, B;
  wire [39:0] Z;
  add_signed_468_GENERIC_REAL g1(.A ({A[37], A[37:0]}), .B ({B[37],
       B[37:0]}), .Z (Z));
endmodule

module add_signed_4709_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [58:0] A, B;
  output [59:0] Z;
  wire [58:0] A, B;
  wire [59:0] Z;
  wire n_182, n_183, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476;
  not g3 (Z[59], n_182);
  nand g4 (n_183, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_188, A[1], B[1]);
  nand g13 (n_192, n_188, n_189, n_190);
  xor g14 (n_191, A[1], B[1]);
  nand g16 (n_193, A[2], B[2]);
  nand g17 (n_194, A[2], n_192);
  nand g18 (n_195, B[2], n_192);
  nand g19 (n_197, n_193, n_194, n_195);
  xor g20 (n_196, A[2], B[2]);
  xor g21 (Z[2], n_192, n_196);
  nand g22 (n_198, A[3], B[3]);
  nand g23 (n_199, A[3], n_197);
  nand g24 (n_200, B[3], n_197);
  nand g25 (n_202, n_198, n_199, n_200);
  xor g26 (n_201, A[3], B[3]);
  xor g27 (Z[3], n_197, n_201);
  nand g28 (n_203, A[4], B[4]);
  nand g29 (n_204, A[4], n_202);
  nand g30 (n_205, B[4], n_202);
  nand g31 (n_207, n_203, n_204, n_205);
  xor g32 (n_206, A[4], B[4]);
  xor g33 (Z[4], n_202, n_206);
  nand g34 (n_208, A[5], B[5]);
  nand g35 (n_209, A[5], n_207);
  nand g36 (n_210, B[5], n_207);
  nand g37 (n_212, n_208, n_209, n_210);
  xor g38 (n_211, A[5], B[5]);
  xor g39 (Z[5], n_207, n_211);
  nand g40 (n_213, A[6], B[6]);
  nand g41 (n_214, A[6], n_212);
  nand g42 (n_215, B[6], n_212);
  nand g43 (n_217, n_213, n_214, n_215);
  xor g44 (n_216, A[6], B[6]);
  xor g45 (Z[6], n_212, n_216);
  nand g46 (n_218, A[7], B[7]);
  nand g47 (n_219, A[7], n_217);
  nand g48 (n_220, B[7], n_217);
  nand g49 (n_222, n_218, n_219, n_220);
  xor g50 (n_221, A[7], B[7]);
  xor g51 (Z[7], n_217, n_221);
  nand g52 (n_223, A[8], B[8]);
  nand g53 (n_224, A[8], n_222);
  nand g54 (n_225, B[8], n_222);
  nand g55 (n_227, n_223, n_224, n_225);
  xor g56 (n_226, A[8], B[8]);
  xor g57 (Z[8], n_222, n_226);
  nand g58 (n_228, A[9], B[9]);
  nand g59 (n_229, A[9], n_227);
  nand g60 (n_230, B[9], n_227);
  nand g61 (n_232, n_228, n_229, n_230);
  xor g62 (n_231, A[9], B[9]);
  xor g63 (Z[9], n_227, n_231);
  nand g64 (n_233, A[10], B[10]);
  nand g65 (n_234, A[10], n_232);
  nand g66 (n_235, B[10], n_232);
  nand g67 (n_237, n_233, n_234, n_235);
  xor g68 (n_236, A[10], B[10]);
  xor g69 (Z[10], n_232, n_236);
  nand g70 (n_238, A[11], B[11]);
  nand g71 (n_239, A[11], n_237);
  nand g72 (n_240, B[11], n_237);
  nand g73 (n_242, n_238, n_239, n_240);
  xor g74 (n_241, A[11], B[11]);
  xor g75 (Z[11], n_237, n_241);
  nand g76 (n_243, A[12], B[12]);
  nand g77 (n_244, A[12], n_242);
  nand g78 (n_245, B[12], n_242);
  nand g79 (n_247, n_243, n_244, n_245);
  xor g80 (n_246, A[12], B[12]);
  xor g81 (Z[12], n_242, n_246);
  nand g82 (n_248, A[13], B[13]);
  nand g83 (n_249, A[13], n_247);
  nand g84 (n_250, B[13], n_247);
  nand g85 (n_252, n_248, n_249, n_250);
  xor g86 (n_251, A[13], B[13]);
  xor g87 (Z[13], n_247, n_251);
  nand g88 (n_253, A[14], B[14]);
  nand g89 (n_254, A[14], n_252);
  nand g90 (n_255, B[14], n_252);
  nand g91 (n_257, n_253, n_254, n_255);
  xor g92 (n_256, A[14], B[14]);
  xor g93 (Z[14], n_252, n_256);
  nand g94 (n_258, A[15], B[15]);
  nand g95 (n_259, A[15], n_257);
  nand g96 (n_260, B[15], n_257);
  nand g97 (n_262, n_258, n_259, n_260);
  xor g98 (n_261, A[15], B[15]);
  xor g99 (Z[15], n_257, n_261);
  nand g100 (n_263, A[16], B[16]);
  nand g101 (n_264, A[16], n_262);
  nand g102 (n_265, B[16], n_262);
  nand g103 (n_267, n_263, n_264, n_265);
  xor g104 (n_266, A[16], B[16]);
  xor g105 (Z[16], n_262, n_266);
  nand g106 (n_268, A[17], B[17]);
  nand g107 (n_269, A[17], n_267);
  nand g108 (n_270, B[17], n_267);
  nand g109 (n_272, n_268, n_269, n_270);
  xor g110 (n_271, A[17], B[17]);
  xor g111 (Z[17], n_267, n_271);
  nand g112 (n_273, A[18], B[18]);
  nand g113 (n_274, A[18], n_272);
  nand g114 (n_275, B[18], n_272);
  nand g115 (n_277, n_273, n_274, n_275);
  xor g116 (n_276, A[18], B[18]);
  xor g117 (Z[18], n_272, n_276);
  nand g118 (n_278, A[19], B[19]);
  nand g119 (n_279, A[19], n_277);
  nand g120 (n_280, B[19], n_277);
  nand g121 (n_282, n_278, n_279, n_280);
  xor g122 (n_281, A[19], B[19]);
  xor g123 (Z[19], n_277, n_281);
  nand g124 (n_283, A[20], B[20]);
  nand g125 (n_284, A[20], n_282);
  nand g126 (n_285, B[20], n_282);
  nand g127 (n_287, n_283, n_284, n_285);
  xor g128 (n_286, A[20], B[20]);
  xor g129 (Z[20], n_282, n_286);
  nand g130 (n_288, A[21], B[21]);
  nand g131 (n_289, A[21], n_287);
  nand g132 (n_290, B[21], n_287);
  nand g133 (n_292, n_288, n_289, n_290);
  xor g134 (n_291, A[21], B[21]);
  xor g135 (Z[21], n_287, n_291);
  nand g136 (n_293, A[22], B[22]);
  nand g137 (n_294, A[22], n_292);
  nand g138 (n_295, B[22], n_292);
  nand g139 (n_297, n_293, n_294, n_295);
  xor g140 (n_296, A[22], B[22]);
  xor g141 (Z[22], n_292, n_296);
  nand g142 (n_298, A[23], B[23]);
  nand g143 (n_299, A[23], n_297);
  nand g144 (n_300, B[23], n_297);
  nand g145 (n_302, n_298, n_299, n_300);
  xor g146 (n_301, A[23], B[23]);
  xor g147 (Z[23], n_297, n_301);
  nand g148 (n_303, A[24], B[24]);
  nand g149 (n_304, A[24], n_302);
  nand g150 (n_305, B[24], n_302);
  nand g151 (n_307, n_303, n_304, n_305);
  xor g152 (n_306, A[24], B[24]);
  xor g153 (Z[24], n_302, n_306);
  nand g154 (n_308, A[25], B[25]);
  nand g155 (n_309, A[25], n_307);
  nand g156 (n_310, B[25], n_307);
  nand g157 (n_312, n_308, n_309, n_310);
  xor g158 (n_311, A[25], B[25]);
  xor g159 (Z[25], n_307, n_311);
  nand g160 (n_313, A[26], B[26]);
  nand g161 (n_314, A[26], n_312);
  nand g162 (n_315, B[26], n_312);
  nand g163 (n_317, n_313, n_314, n_315);
  xor g164 (n_316, A[26], B[26]);
  xor g165 (Z[26], n_312, n_316);
  nand g166 (n_318, A[27], B[27]);
  nand g167 (n_319, A[27], n_317);
  nand g168 (n_320, B[27], n_317);
  nand g169 (n_322, n_318, n_319, n_320);
  xor g170 (n_321, A[27], B[27]);
  xor g171 (Z[27], n_317, n_321);
  nand g172 (n_323, A[28], B[28]);
  nand g173 (n_324, A[28], n_322);
  nand g174 (n_325, B[28], n_322);
  nand g175 (n_327, n_323, n_324, n_325);
  xor g176 (n_326, A[28], B[28]);
  xor g177 (Z[28], n_322, n_326);
  nand g178 (n_328, A[29], B[29]);
  nand g179 (n_329, A[29], n_327);
  nand g180 (n_330, B[29], n_327);
  nand g181 (n_332, n_328, n_329, n_330);
  xor g182 (n_331, A[29], B[29]);
  xor g183 (Z[29], n_327, n_331);
  nand g184 (n_333, A[30], B[30]);
  nand g185 (n_334, A[30], n_332);
  nand g186 (n_335, B[30], n_332);
  nand g187 (n_337, n_333, n_334, n_335);
  xor g188 (n_336, A[30], B[30]);
  xor g189 (Z[30], n_332, n_336);
  nand g190 (n_338, A[31], B[31]);
  nand g191 (n_339, A[31], n_337);
  nand g192 (n_340, B[31], n_337);
  nand g193 (n_342, n_338, n_339, n_340);
  xor g194 (n_341, A[31], B[31]);
  xor g195 (Z[31], n_337, n_341);
  nand g196 (n_343, A[32], B[32]);
  nand g197 (n_344, A[32], n_342);
  nand g198 (n_345, B[32], n_342);
  nand g199 (n_347, n_343, n_344, n_345);
  xor g200 (n_346, A[32], B[32]);
  xor g201 (Z[32], n_342, n_346);
  nand g202 (n_348, A[33], B[33]);
  nand g203 (n_349, A[33], n_347);
  nand g204 (n_350, B[33], n_347);
  nand g205 (n_352, n_348, n_349, n_350);
  xor g206 (n_351, A[33], B[33]);
  xor g207 (Z[33], n_347, n_351);
  nand g208 (n_353, A[34], B[34]);
  nand g209 (n_354, A[34], n_352);
  nand g210 (n_355, B[34], n_352);
  nand g211 (n_357, n_353, n_354, n_355);
  xor g212 (n_356, A[34], B[34]);
  xor g213 (Z[34], n_352, n_356);
  nand g214 (n_358, A[35], B[35]);
  nand g215 (n_359, A[35], n_357);
  nand g216 (n_360, B[35], n_357);
  nand g217 (n_362, n_358, n_359, n_360);
  xor g218 (n_361, A[35], B[35]);
  xor g219 (Z[35], n_357, n_361);
  nand g220 (n_363, A[36], B[36]);
  nand g221 (n_364, A[36], n_362);
  nand g222 (n_365, B[36], n_362);
  nand g223 (n_367, n_363, n_364, n_365);
  xor g224 (n_366, A[36], B[36]);
  xor g225 (Z[36], n_362, n_366);
  nand g226 (n_368, A[37], B[37]);
  nand g227 (n_369, A[37], n_367);
  nand g228 (n_370, B[37], n_367);
  nand g229 (n_372, n_368, n_369, n_370);
  xor g230 (n_371, A[37], B[37]);
  xor g231 (Z[37], n_367, n_371);
  nand g232 (n_373, A[38], B[38]);
  nand g233 (n_374, A[38], n_372);
  nand g234 (n_375, B[38], n_372);
  nand g235 (n_377, n_373, n_374, n_375);
  xor g236 (n_376, A[38], B[38]);
  xor g237 (Z[38], n_372, n_376);
  nand g238 (n_378, A[39], B[39]);
  nand g239 (n_379, A[39], n_377);
  nand g240 (n_380, B[39], n_377);
  nand g241 (n_382, n_378, n_379, n_380);
  xor g242 (n_381, A[39], B[39]);
  xor g243 (Z[39], n_377, n_381);
  nand g244 (n_383, A[40], B[40]);
  nand g245 (n_384, A[40], n_382);
  nand g246 (n_385, B[40], n_382);
  nand g247 (n_387, n_383, n_384, n_385);
  xor g248 (n_386, A[40], B[40]);
  xor g249 (Z[40], n_382, n_386);
  nand g250 (n_388, A[41], B[41]);
  nand g251 (n_389, A[41], n_387);
  nand g252 (n_390, B[41], n_387);
  nand g253 (n_392, n_388, n_389, n_390);
  xor g254 (n_391, A[41], B[41]);
  xor g255 (Z[41], n_387, n_391);
  nand g256 (n_393, A[42], B[42]);
  nand g257 (n_394, A[42], n_392);
  nand g258 (n_395, B[42], n_392);
  nand g259 (n_397, n_393, n_394, n_395);
  xor g260 (n_396, A[42], B[42]);
  xor g261 (Z[42], n_392, n_396);
  nand g262 (n_398, A[43], B[43]);
  nand g263 (n_399, A[43], n_397);
  nand g264 (n_400, B[43], n_397);
  nand g265 (n_402, n_398, n_399, n_400);
  xor g266 (n_401, A[43], B[43]);
  xor g267 (Z[43], n_397, n_401);
  nand g268 (n_403, A[44], B[44]);
  nand g269 (n_404, A[44], n_402);
  nand g270 (n_405, B[44], n_402);
  nand g271 (n_407, n_403, n_404, n_405);
  xor g272 (n_406, A[44], B[44]);
  xor g273 (Z[44], n_402, n_406);
  nand g274 (n_408, A[45], B[45]);
  nand g275 (n_409, A[45], n_407);
  nand g276 (n_410, B[45], n_407);
  nand g277 (n_412, n_408, n_409, n_410);
  xor g278 (n_411, A[45], B[45]);
  xor g279 (Z[45], n_407, n_411);
  nand g280 (n_413, A[46], B[46]);
  nand g281 (n_414, A[46], n_412);
  nand g282 (n_415, B[46], n_412);
  nand g283 (n_417, n_413, n_414, n_415);
  xor g284 (n_416, A[46], B[46]);
  xor g285 (Z[46], n_412, n_416);
  nand g286 (n_418, A[47], B[47]);
  nand g287 (n_419, A[47], n_417);
  nand g288 (n_420, B[47], n_417);
  nand g289 (n_422, n_418, n_419, n_420);
  xor g290 (n_421, A[47], B[47]);
  xor g291 (Z[47], n_417, n_421);
  nand g292 (n_423, A[48], B[48]);
  nand g293 (n_424, A[48], n_422);
  nand g294 (n_425, B[48], n_422);
  nand g295 (n_427, n_423, n_424, n_425);
  xor g296 (n_426, A[48], B[48]);
  xor g297 (Z[48], n_422, n_426);
  nand g298 (n_428, A[49], B[49]);
  nand g299 (n_429, A[49], n_427);
  nand g300 (n_430, B[49], n_427);
  nand g301 (n_432, n_428, n_429, n_430);
  xor g302 (n_431, A[49], B[49]);
  xor g303 (Z[49], n_427, n_431);
  nand g304 (n_433, A[50], B[50]);
  nand g305 (n_434, A[50], n_432);
  nand g306 (n_435, B[50], n_432);
  nand g307 (n_437, n_433, n_434, n_435);
  xor g308 (n_436, A[50], B[50]);
  xor g309 (Z[50], n_432, n_436);
  nand g310 (n_438, A[51], B[51]);
  nand g311 (n_439, A[51], n_437);
  nand g312 (n_440, B[51], n_437);
  nand g313 (n_442, n_438, n_439, n_440);
  xor g314 (n_441, A[51], B[51]);
  xor g315 (Z[51], n_437, n_441);
  nand g316 (n_443, A[52], B[52]);
  nand g317 (n_444, A[52], n_442);
  nand g318 (n_445, B[52], n_442);
  nand g319 (n_447, n_443, n_444, n_445);
  xor g320 (n_446, A[52], B[52]);
  xor g321 (Z[52], n_442, n_446);
  nand g322 (n_448, A[53], B[53]);
  nand g323 (n_449, A[53], n_447);
  nand g324 (n_450, B[53], n_447);
  nand g325 (n_452, n_448, n_449, n_450);
  xor g326 (n_451, A[53], B[53]);
  xor g327 (Z[53], n_447, n_451);
  nand g328 (n_453, A[54], B[54]);
  nand g329 (n_454, A[54], n_452);
  nand g330 (n_455, B[54], n_452);
  nand g331 (n_457, n_453, n_454, n_455);
  xor g332 (n_456, A[54], B[54]);
  xor g333 (Z[54], n_452, n_456);
  nand g334 (n_458, A[55], B[55]);
  nand g335 (n_459, A[55], n_457);
  nand g336 (n_460, B[55], n_457);
  nand g337 (n_462, n_458, n_459, n_460);
  xor g338 (n_461, A[55], B[55]);
  xor g339 (Z[55], n_457, n_461);
  nand g340 (n_463, A[56], B[56]);
  nand g341 (n_464, A[56], n_462);
  nand g342 (n_465, B[56], n_462);
  nand g343 (n_467, n_463, n_464, n_465);
  xor g344 (n_466, A[56], B[56]);
  xor g345 (Z[56], n_462, n_466);
  nand g346 (n_468, A[57], B[57]);
  nand g347 (n_469, A[57], n_467);
  nand g348 (n_470, B[57], n_467);
  nand g349 (n_472, n_468, n_469, n_470);
  xor g350 (n_471, A[57], B[57]);
  xor g351 (Z[57], n_467, n_471);
  nand g355 (n_182, n_473, n_474, n_475);
  xor g357 (Z[58], n_472, n_476);
  or g359 (n_473, A[58], B[58]);
  xor g360 (n_476, A[58], B[58]);
  or g361 (n_189, wc, n_183);
  not gc (wc, A[1]);
  or g362 (n_190, wc0, n_183);
  not gc0 (wc0, B[1]);
  xnor g363 (Z[1], n_183, n_191);
  or g364 (n_474, A[58], wc1);
  not gc1 (wc1, n_472);
  or g365 (n_475, B[58], wc2);
  not gc2 (wc2, n_472);
endmodule

module add_signed_4709_GENERIC(A, B, Z);
  input [58:0] A, B;
  output [59:0] Z;
  wire [58:0] A, B;
  wire [59:0] Z;
  add_signed_4709_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_4709_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [58:0] A, B;
  output [59:0] Z;
  wire [58:0] A, B;
  wire [59:0] Z;
  wire n_182, n_183, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476;
  not g3 (Z[59], n_182);
  nand g4 (n_183, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_188, A[1], B[1]);
  nand g13 (n_192, n_188, n_189, n_190);
  xor g14 (n_191, A[1], B[1]);
  nand g16 (n_193, A[2], B[2]);
  nand g17 (n_194, A[2], n_192);
  nand g18 (n_195, B[2], n_192);
  nand g19 (n_197, n_193, n_194, n_195);
  xor g20 (n_196, A[2], B[2]);
  xor g21 (Z[2], n_192, n_196);
  nand g22 (n_198, A[3], B[3]);
  nand g23 (n_199, A[3], n_197);
  nand g24 (n_200, B[3], n_197);
  nand g25 (n_202, n_198, n_199, n_200);
  xor g26 (n_201, A[3], B[3]);
  xor g27 (Z[3], n_197, n_201);
  nand g28 (n_203, A[4], B[4]);
  nand g29 (n_204, A[4], n_202);
  nand g30 (n_205, B[4], n_202);
  nand g31 (n_207, n_203, n_204, n_205);
  xor g32 (n_206, A[4], B[4]);
  xor g33 (Z[4], n_202, n_206);
  nand g34 (n_208, A[5], B[5]);
  nand g35 (n_209, A[5], n_207);
  nand g36 (n_210, B[5], n_207);
  nand g37 (n_212, n_208, n_209, n_210);
  xor g38 (n_211, A[5], B[5]);
  xor g39 (Z[5], n_207, n_211);
  nand g40 (n_213, A[6], B[6]);
  nand g41 (n_214, A[6], n_212);
  nand g42 (n_215, B[6], n_212);
  nand g43 (n_217, n_213, n_214, n_215);
  xor g44 (n_216, A[6], B[6]);
  xor g45 (Z[6], n_212, n_216);
  nand g46 (n_218, A[7], B[7]);
  nand g47 (n_219, A[7], n_217);
  nand g48 (n_220, B[7], n_217);
  nand g49 (n_222, n_218, n_219, n_220);
  xor g50 (n_221, A[7], B[7]);
  xor g51 (Z[7], n_217, n_221);
  nand g52 (n_223, A[8], B[8]);
  nand g53 (n_224, A[8], n_222);
  nand g54 (n_225, B[8], n_222);
  nand g55 (n_227, n_223, n_224, n_225);
  xor g56 (n_226, A[8], B[8]);
  xor g57 (Z[8], n_222, n_226);
  nand g58 (n_228, A[9], B[9]);
  nand g59 (n_229, A[9], n_227);
  nand g60 (n_230, B[9], n_227);
  nand g61 (n_232, n_228, n_229, n_230);
  xor g62 (n_231, A[9], B[9]);
  xor g63 (Z[9], n_227, n_231);
  nand g64 (n_233, A[10], B[10]);
  nand g65 (n_234, A[10], n_232);
  nand g66 (n_235, B[10], n_232);
  nand g67 (n_237, n_233, n_234, n_235);
  xor g68 (n_236, A[10], B[10]);
  xor g69 (Z[10], n_232, n_236);
  nand g70 (n_238, A[11], B[11]);
  nand g71 (n_239, A[11], n_237);
  nand g72 (n_240, B[11], n_237);
  nand g73 (n_242, n_238, n_239, n_240);
  xor g74 (n_241, A[11], B[11]);
  xor g75 (Z[11], n_237, n_241);
  nand g76 (n_243, A[12], B[12]);
  nand g77 (n_244, A[12], n_242);
  nand g78 (n_245, B[12], n_242);
  nand g79 (n_247, n_243, n_244, n_245);
  xor g80 (n_246, A[12], B[12]);
  xor g81 (Z[12], n_242, n_246);
  nand g82 (n_248, A[13], B[13]);
  nand g83 (n_249, A[13], n_247);
  nand g84 (n_250, B[13], n_247);
  nand g85 (n_252, n_248, n_249, n_250);
  xor g86 (n_251, A[13], B[13]);
  xor g87 (Z[13], n_247, n_251);
  nand g88 (n_253, A[14], B[14]);
  nand g89 (n_254, A[14], n_252);
  nand g90 (n_255, B[14], n_252);
  nand g91 (n_257, n_253, n_254, n_255);
  xor g92 (n_256, A[14], B[14]);
  xor g93 (Z[14], n_252, n_256);
  nand g94 (n_258, A[15], B[15]);
  nand g95 (n_259, A[15], n_257);
  nand g96 (n_260, B[15], n_257);
  nand g97 (n_262, n_258, n_259, n_260);
  xor g98 (n_261, A[15], B[15]);
  xor g99 (Z[15], n_257, n_261);
  nand g100 (n_263, A[16], B[16]);
  nand g101 (n_264, A[16], n_262);
  nand g102 (n_265, B[16], n_262);
  nand g103 (n_267, n_263, n_264, n_265);
  xor g104 (n_266, A[16], B[16]);
  xor g105 (Z[16], n_262, n_266);
  nand g106 (n_268, A[17], B[17]);
  nand g107 (n_269, A[17], n_267);
  nand g108 (n_270, B[17], n_267);
  nand g109 (n_272, n_268, n_269, n_270);
  xor g110 (n_271, A[17], B[17]);
  xor g111 (Z[17], n_267, n_271);
  nand g112 (n_273, A[18], B[18]);
  nand g113 (n_274, A[18], n_272);
  nand g114 (n_275, B[18], n_272);
  nand g115 (n_277, n_273, n_274, n_275);
  xor g116 (n_276, A[18], B[18]);
  xor g117 (Z[18], n_272, n_276);
  nand g118 (n_278, A[19], B[19]);
  nand g119 (n_279, A[19], n_277);
  nand g120 (n_280, B[19], n_277);
  nand g121 (n_282, n_278, n_279, n_280);
  xor g122 (n_281, A[19], B[19]);
  xor g123 (Z[19], n_277, n_281);
  nand g124 (n_283, A[20], B[20]);
  nand g125 (n_284, A[20], n_282);
  nand g126 (n_285, B[20], n_282);
  nand g127 (n_287, n_283, n_284, n_285);
  xor g128 (n_286, A[20], B[20]);
  xor g129 (Z[20], n_282, n_286);
  nand g130 (n_288, A[21], B[21]);
  nand g131 (n_289, A[21], n_287);
  nand g132 (n_290, B[21], n_287);
  nand g133 (n_292, n_288, n_289, n_290);
  xor g134 (n_291, A[21], B[21]);
  xor g135 (Z[21], n_287, n_291);
  nand g136 (n_293, A[22], B[22]);
  nand g137 (n_294, A[22], n_292);
  nand g138 (n_295, B[22], n_292);
  nand g139 (n_297, n_293, n_294, n_295);
  xor g140 (n_296, A[22], B[22]);
  xor g141 (Z[22], n_292, n_296);
  nand g142 (n_298, A[23], B[23]);
  nand g143 (n_299, A[23], n_297);
  nand g144 (n_300, B[23], n_297);
  nand g145 (n_302, n_298, n_299, n_300);
  xor g146 (n_301, A[23], B[23]);
  xor g147 (Z[23], n_297, n_301);
  nand g148 (n_303, A[24], B[24]);
  nand g149 (n_304, A[24], n_302);
  nand g150 (n_305, B[24], n_302);
  nand g151 (n_307, n_303, n_304, n_305);
  xor g152 (n_306, A[24], B[24]);
  xor g153 (Z[24], n_302, n_306);
  nand g154 (n_308, A[25], B[25]);
  nand g155 (n_309, A[25], n_307);
  nand g156 (n_310, B[25], n_307);
  nand g157 (n_312, n_308, n_309, n_310);
  xor g158 (n_311, A[25], B[25]);
  xor g159 (Z[25], n_307, n_311);
  nand g160 (n_313, A[26], B[26]);
  nand g161 (n_314, A[26], n_312);
  nand g162 (n_315, B[26], n_312);
  nand g163 (n_317, n_313, n_314, n_315);
  xor g164 (n_316, A[26], B[26]);
  xor g165 (Z[26], n_312, n_316);
  nand g166 (n_318, A[27], B[27]);
  nand g167 (n_319, A[27], n_317);
  nand g168 (n_320, B[27], n_317);
  nand g169 (n_322, n_318, n_319, n_320);
  xor g170 (n_321, A[27], B[27]);
  xor g171 (Z[27], n_317, n_321);
  nand g172 (n_323, A[28], B[28]);
  nand g173 (n_324, A[28], n_322);
  nand g174 (n_325, B[28], n_322);
  nand g175 (n_327, n_323, n_324, n_325);
  xor g176 (n_326, A[28], B[28]);
  xor g177 (Z[28], n_322, n_326);
  nand g178 (n_328, A[29], B[29]);
  nand g179 (n_329, A[29], n_327);
  nand g180 (n_330, B[29], n_327);
  nand g181 (n_332, n_328, n_329, n_330);
  xor g182 (n_331, A[29], B[29]);
  xor g183 (Z[29], n_327, n_331);
  nand g184 (n_333, A[30], B[30]);
  nand g185 (n_334, A[30], n_332);
  nand g186 (n_335, B[30], n_332);
  nand g187 (n_337, n_333, n_334, n_335);
  xor g188 (n_336, A[30], B[30]);
  xor g189 (Z[30], n_332, n_336);
  nand g190 (n_338, A[31], B[31]);
  nand g191 (n_339, A[31], n_337);
  nand g192 (n_340, B[31], n_337);
  nand g193 (n_342, n_338, n_339, n_340);
  xor g194 (n_341, A[31], B[31]);
  xor g195 (Z[31], n_337, n_341);
  nand g196 (n_343, A[32], B[32]);
  nand g197 (n_344, A[32], n_342);
  nand g198 (n_345, B[32], n_342);
  nand g199 (n_347, n_343, n_344, n_345);
  xor g200 (n_346, A[32], B[32]);
  xor g201 (Z[32], n_342, n_346);
  nand g202 (n_348, A[33], B[33]);
  nand g203 (n_349, A[33], n_347);
  nand g204 (n_350, B[33], n_347);
  nand g205 (n_352, n_348, n_349, n_350);
  xor g206 (n_351, A[33], B[33]);
  xor g207 (Z[33], n_347, n_351);
  nand g208 (n_353, A[34], B[34]);
  nand g209 (n_354, A[34], n_352);
  nand g210 (n_355, B[34], n_352);
  nand g211 (n_357, n_353, n_354, n_355);
  xor g212 (n_356, A[34], B[34]);
  xor g213 (Z[34], n_352, n_356);
  nand g214 (n_358, A[35], B[35]);
  nand g215 (n_359, A[35], n_357);
  nand g216 (n_360, B[35], n_357);
  nand g217 (n_362, n_358, n_359, n_360);
  xor g218 (n_361, A[35], B[35]);
  xor g219 (Z[35], n_357, n_361);
  nand g220 (n_363, A[36], B[36]);
  nand g221 (n_364, A[36], n_362);
  nand g222 (n_365, B[36], n_362);
  nand g223 (n_367, n_363, n_364, n_365);
  xor g224 (n_366, A[36], B[36]);
  xor g225 (Z[36], n_362, n_366);
  nand g226 (n_368, A[37], B[37]);
  nand g227 (n_369, A[37], n_367);
  nand g228 (n_370, B[37], n_367);
  nand g229 (n_372, n_368, n_369, n_370);
  xor g230 (n_371, A[37], B[37]);
  xor g231 (Z[37], n_367, n_371);
  nand g232 (n_373, A[38], B[38]);
  nand g233 (n_374, A[38], n_372);
  nand g234 (n_375, B[38], n_372);
  nand g235 (n_377, n_373, n_374, n_375);
  xor g236 (n_376, A[38], B[38]);
  xor g237 (Z[38], n_372, n_376);
  nand g238 (n_378, A[39], B[39]);
  nand g239 (n_379, A[39], n_377);
  nand g240 (n_380, B[39], n_377);
  nand g241 (n_382, n_378, n_379, n_380);
  xor g242 (n_381, A[39], B[39]);
  xor g243 (Z[39], n_377, n_381);
  nand g244 (n_383, A[40], B[40]);
  nand g245 (n_384, A[40], n_382);
  nand g246 (n_385, B[40], n_382);
  nand g247 (n_387, n_383, n_384, n_385);
  xor g248 (n_386, A[40], B[40]);
  xor g249 (Z[40], n_382, n_386);
  nand g250 (n_388, A[41], B[41]);
  nand g251 (n_389, A[41], n_387);
  nand g252 (n_390, B[41], n_387);
  nand g253 (n_392, n_388, n_389, n_390);
  xor g254 (n_391, A[41], B[41]);
  xor g255 (Z[41], n_387, n_391);
  nand g256 (n_393, A[42], B[42]);
  nand g257 (n_394, A[42], n_392);
  nand g258 (n_395, B[42], n_392);
  nand g259 (n_397, n_393, n_394, n_395);
  xor g260 (n_396, A[42], B[42]);
  xor g261 (Z[42], n_392, n_396);
  nand g262 (n_398, A[43], B[43]);
  nand g263 (n_399, A[43], n_397);
  nand g264 (n_400, B[43], n_397);
  nand g265 (n_402, n_398, n_399, n_400);
  xor g266 (n_401, A[43], B[43]);
  xor g267 (Z[43], n_397, n_401);
  nand g268 (n_403, A[44], B[44]);
  nand g269 (n_404, A[44], n_402);
  nand g270 (n_405, B[44], n_402);
  nand g271 (n_407, n_403, n_404, n_405);
  xor g272 (n_406, A[44], B[44]);
  xor g273 (Z[44], n_402, n_406);
  nand g274 (n_408, A[45], B[45]);
  nand g275 (n_409, A[45], n_407);
  nand g276 (n_410, B[45], n_407);
  nand g277 (n_412, n_408, n_409, n_410);
  xor g278 (n_411, A[45], B[45]);
  xor g279 (Z[45], n_407, n_411);
  nand g280 (n_413, A[46], B[46]);
  nand g281 (n_414, A[46], n_412);
  nand g282 (n_415, B[46], n_412);
  nand g283 (n_417, n_413, n_414, n_415);
  xor g284 (n_416, A[46], B[46]);
  xor g285 (Z[46], n_412, n_416);
  nand g286 (n_418, A[47], B[47]);
  nand g287 (n_419, A[47], n_417);
  nand g288 (n_420, B[47], n_417);
  nand g289 (n_422, n_418, n_419, n_420);
  xor g290 (n_421, A[47], B[47]);
  xor g291 (Z[47], n_417, n_421);
  nand g292 (n_423, A[48], B[48]);
  nand g293 (n_424, A[48], n_422);
  nand g294 (n_425, B[48], n_422);
  nand g295 (n_427, n_423, n_424, n_425);
  xor g296 (n_426, A[48], B[48]);
  xor g297 (Z[48], n_422, n_426);
  nand g298 (n_428, A[49], B[49]);
  nand g299 (n_429, A[49], n_427);
  nand g300 (n_430, B[49], n_427);
  nand g301 (n_432, n_428, n_429, n_430);
  xor g302 (n_431, A[49], B[49]);
  xor g303 (Z[49], n_427, n_431);
  nand g304 (n_433, A[50], B[50]);
  nand g305 (n_434, A[50], n_432);
  nand g306 (n_435, B[50], n_432);
  nand g307 (n_437, n_433, n_434, n_435);
  xor g308 (n_436, A[50], B[50]);
  xor g309 (Z[50], n_432, n_436);
  nand g310 (n_438, A[51], B[51]);
  nand g311 (n_439, A[51], n_437);
  nand g312 (n_440, B[51], n_437);
  nand g313 (n_442, n_438, n_439, n_440);
  xor g314 (n_441, A[51], B[51]);
  xor g315 (Z[51], n_437, n_441);
  nand g316 (n_443, A[52], B[52]);
  nand g317 (n_444, A[52], n_442);
  nand g318 (n_445, B[52], n_442);
  nand g319 (n_447, n_443, n_444, n_445);
  xor g320 (n_446, A[52], B[52]);
  xor g321 (Z[52], n_442, n_446);
  nand g322 (n_448, A[53], B[53]);
  nand g323 (n_449, A[53], n_447);
  nand g324 (n_450, B[53], n_447);
  nand g325 (n_452, n_448, n_449, n_450);
  xor g326 (n_451, A[53], B[53]);
  xor g327 (Z[53], n_447, n_451);
  nand g328 (n_453, A[54], B[54]);
  nand g329 (n_454, A[54], n_452);
  nand g330 (n_455, B[54], n_452);
  nand g331 (n_457, n_453, n_454, n_455);
  xor g332 (n_456, A[54], B[54]);
  xor g333 (Z[54], n_452, n_456);
  nand g334 (n_458, A[55], B[55]);
  nand g335 (n_459, A[55], n_457);
  nand g336 (n_460, B[55], n_457);
  nand g337 (n_462, n_458, n_459, n_460);
  xor g338 (n_461, A[55], B[55]);
  xor g339 (Z[55], n_457, n_461);
  nand g340 (n_463, A[56], B[56]);
  nand g341 (n_464, A[56], n_462);
  nand g342 (n_465, B[56], n_462);
  nand g343 (n_467, n_463, n_464, n_465);
  xor g344 (n_466, A[56], B[56]);
  xor g345 (Z[56], n_462, n_466);
  nand g346 (n_468, A[57], B[57]);
  nand g347 (n_469, A[57], n_467);
  nand g348 (n_470, B[57], n_467);
  nand g349 (n_472, n_468, n_469, n_470);
  xor g350 (n_471, A[57], B[57]);
  xor g351 (Z[57], n_467, n_471);
  nand g355 (n_182, n_473, n_474, n_475);
  xor g357 (Z[58], n_472, n_476);
  or g359 (n_473, A[58], B[58]);
  xor g360 (n_476, A[58], B[58]);
  or g361 (n_189, wc, n_183);
  not gc (wc, A[1]);
  or g362 (n_190, wc0, n_183);
  not gc0 (wc0, B[1]);
  xnor g363 (Z[1], n_183, n_191);
  or g364 (n_474, A[58], wc1);
  not gc1 (wc1, n_472);
  or g365 (n_475, B[58], wc2);
  not gc2 (wc2, n_472);
endmodule

module add_signed_4709_1_GENERIC(A, B, Z);
  input [58:0] A, B;
  output [59:0] Z;
  wire [58:0] A, B;
  wire [59:0] Z;
  add_signed_4709_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_4709_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [58:0] A, B;
  output [59:0] Z;
  wire [58:0] A, B;
  wire [59:0] Z;
  wire n_182, n_183, n_186, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_196, n_197, n_198, n_199, n_200, n_202, n_203;
  wire n_204, n_205, n_206, n_208, n_209, n_210, n_211, n_212;
  wire n_214, n_215, n_216, n_217, n_218, n_220, n_221, n_222;
  wire n_223, n_224, n_226, n_227, n_228, n_229, n_230, n_232;
  wire n_233, n_234, n_235, n_236, n_238, n_239, n_240, n_241;
  wire n_242, n_244, n_245, n_246, n_247, n_248, n_250, n_251;
  wire n_252, n_253, n_254, n_256, n_257, n_258, n_259, n_260;
  wire n_262, n_263, n_264, n_265, n_266, n_268, n_269, n_270;
  wire n_271, n_272, n_274, n_275, n_276, n_277, n_278, n_280;
  wire n_281, n_282, n_283, n_284, n_286, n_287, n_288, n_289;
  wire n_290, n_292, n_293, n_294, n_295, n_296, n_298, n_299;
  wire n_300, n_301, n_302, n_304, n_305, n_306, n_307, n_308;
  wire n_310, n_311, n_312, n_313, n_314, n_316, n_317, n_318;
  wire n_319, n_320, n_322, n_323, n_324, n_325, n_326, n_328;
  wire n_329, n_330, n_331, n_332, n_334, n_335, n_336, n_337;
  wire n_338, n_340, n_341, n_342, n_343, n_344, n_346, n_347;
  wire n_348, n_349, n_350, n_352, n_353, n_354, n_355, n_356;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_366;
  wire n_367, n_369, n_370, n_371, n_373, n_374, n_376, n_377;
  wire n_378, n_380, n_381, n_383, n_384, n_385, n_387, n_388;
  wire n_390, n_391, n_392, n_394, n_395, n_397, n_398, n_399;
  wire n_401, n_402, n_404, n_405, n_406, n_408, n_409, n_411;
  wire n_412, n_413, n_415, n_416, n_418, n_419, n_420, n_422;
  wire n_423, n_425, n_426, n_427, n_429, n_430, n_432, n_433;
  wire n_434, n_436, n_437, n_439, n_440, n_441, n_443, n_444;
  wire n_446, n_447, n_448, n_450, n_451, n_453, n_454, n_455;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_464, n_465;
  wire n_466, n_467, n_468, n_470, n_471, n_472, n_473, n_474;
  wire n_476, n_477, n_478, n_479, n_480, n_482, n_483, n_484;
  wire n_485, n_486, n_488, n_489, n_490, n_491, n_492, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_502, n_503;
  wire n_505, n_506, n_507, n_509, n_510, n_512, n_513, n_514;
  wire n_516, n_517, n_518, n_519, n_521, n_522, n_523, n_524;
  wire n_525, n_526, n_527, n_528, n_530, n_532, n_533, n_535;
  wire n_537, n_538, n_540, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562;
  wire n_563, n_564, n_565, n_567, n_569, n_570, n_572, n_574;
  wire n_575, n_577, n_579, n_580, n_582, n_584, n_585, n_587;
  wire n_589, n_590, n_592, n_594, n_595, n_597, n_599, n_600;
  wire n_602, n_604, n_605, n_607, n_609, n_610, n_612, n_614;
  wire n_615, n_617, n_619, n_620, n_622, n_624, n_625, n_627;
  wire n_629, n_630, n_632, n_634, n_635, n_636, n_638, n_639;
  wire n_640, n_641, n_643, n_644, n_645, n_647, n_648, n_649;
  wire n_651, n_652, n_653, n_655, n_656, n_657, n_659, n_660;
  wire n_661, n_663, n_664, n_665, n_667, n_668, n_669, n_671;
  wire n_672, n_673, n_675, n_676, n_677, n_679, n_680, n_681;
  wire n_683, n_684, n_685, n_687, n_688, n_689, n_691, n_692;
  wire n_693, n_695, n_696, n_697, n_699, n_700, n_701, n_703;
  wire n_704, n_705, n_707, n_708, n_709, n_711, n_712, n_713;
  wire n_715, n_716, n_717, n_719, n_720, n_721, n_723, n_724;
  wire n_725, n_727, n_728, n_729, n_731, n_732, n_733, n_735;
  wire n_736, n_737, n_739, n_740, n_741, n_743, n_744, n_745;
  wire n_747, n_748, n_749, n_751, n_752, n_753;
  not g3 (Z[59], n_182);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_183, A[0], B[0]);
  nor g9 (n_186, A[1], B[1]);
  nand g10 (n_189, A[1], B[1]);
  nor g11 (n_196, A[2], B[2]);
  nand g12 (n_191, A[2], B[2]);
  nor g13 (n_192, A[3], B[3]);
  nand g14 (n_193, A[3], B[3]);
  nor g15 (n_202, A[4], B[4]);
  nand g16 (n_197, A[4], B[4]);
  nor g17 (n_198, A[5], B[5]);
  nand g18 (n_199, A[5], B[5]);
  nor g19 (n_208, A[6], B[6]);
  nand g20 (n_203, A[6], B[6]);
  nor g21 (n_204, A[7], B[7]);
  nand g22 (n_205, A[7], B[7]);
  nor g23 (n_214, A[8], B[8]);
  nand g24 (n_209, A[8], B[8]);
  nor g25 (n_210, A[9], B[9]);
  nand g26 (n_211, A[9], B[9]);
  nor g27 (n_220, A[10], B[10]);
  nand g28 (n_215, A[10], B[10]);
  nor g29 (n_216, A[11], B[11]);
  nand g30 (n_217, A[11], B[11]);
  nor g31 (n_226, A[12], B[12]);
  nand g32 (n_221, A[12], B[12]);
  nor g33 (n_222, A[13], B[13]);
  nand g34 (n_223, A[13], B[13]);
  nor g35 (n_232, A[14], B[14]);
  nand g36 (n_227, A[14], B[14]);
  nor g37 (n_228, A[15], B[15]);
  nand g38 (n_229, A[15], B[15]);
  nor g39 (n_238, A[16], B[16]);
  nand g40 (n_233, A[16], B[16]);
  nor g41 (n_234, A[17], B[17]);
  nand g42 (n_235, A[17], B[17]);
  nor g43 (n_244, A[18], B[18]);
  nand g44 (n_239, A[18], B[18]);
  nor g45 (n_240, A[19], B[19]);
  nand g46 (n_241, A[19], B[19]);
  nor g47 (n_250, A[20], B[20]);
  nand g48 (n_245, A[20], B[20]);
  nor g49 (n_246, A[21], B[21]);
  nand g50 (n_247, A[21], B[21]);
  nor g51 (n_256, A[22], B[22]);
  nand g52 (n_251, A[22], B[22]);
  nor g53 (n_252, A[23], B[23]);
  nand g54 (n_253, A[23], B[23]);
  nor g55 (n_262, A[24], B[24]);
  nand g56 (n_257, A[24], B[24]);
  nor g57 (n_258, A[25], B[25]);
  nand g58 (n_259, A[25], B[25]);
  nor g59 (n_268, A[26], B[26]);
  nand g60 (n_263, A[26], B[26]);
  nor g61 (n_264, A[27], B[27]);
  nand g62 (n_265, A[27], B[27]);
  nor g63 (n_274, A[28], B[28]);
  nand g64 (n_269, A[28], B[28]);
  nor g65 (n_270, A[29], B[29]);
  nand g66 (n_271, A[29], B[29]);
  nor g67 (n_280, A[30], B[30]);
  nand g68 (n_275, A[30], B[30]);
  nor g69 (n_276, A[31], B[31]);
  nand g70 (n_277, A[31], B[31]);
  nor g71 (n_286, A[32], B[32]);
  nand g72 (n_281, A[32], B[32]);
  nor g73 (n_282, A[33], B[33]);
  nand g74 (n_283, A[33], B[33]);
  nor g75 (n_292, A[34], B[34]);
  nand g76 (n_287, A[34], B[34]);
  nor g77 (n_288, A[35], B[35]);
  nand g78 (n_289, A[35], B[35]);
  nor g79 (n_298, A[36], B[36]);
  nand g80 (n_293, A[36], B[36]);
  nor g81 (n_294, A[37], B[37]);
  nand g82 (n_295, A[37], B[37]);
  nor g83 (n_304, A[38], B[38]);
  nand g84 (n_299, A[38], B[38]);
  nor g85 (n_300, A[39], B[39]);
  nand g86 (n_301, A[39], B[39]);
  nor g87 (n_310, A[40], B[40]);
  nand g88 (n_305, A[40], B[40]);
  nor g89 (n_306, A[41], B[41]);
  nand g90 (n_307, A[41], B[41]);
  nor g91 (n_316, A[42], B[42]);
  nand g92 (n_311, A[42], B[42]);
  nor g93 (n_312, A[43], B[43]);
  nand g94 (n_313, A[43], B[43]);
  nor g95 (n_322, A[44], B[44]);
  nand g96 (n_317, A[44], B[44]);
  nor g97 (n_318, A[45], B[45]);
  nand g98 (n_319, A[45], B[45]);
  nor g99 (n_328, A[46], B[46]);
  nand g100 (n_323, A[46], B[46]);
  nor g101 (n_324, A[47], B[47]);
  nand g102 (n_325, A[47], B[47]);
  nor g103 (n_334, A[48], B[48]);
  nand g104 (n_329, A[48], B[48]);
  nor g105 (n_330, A[49], B[49]);
  nand g106 (n_331, A[49], B[49]);
  nor g107 (n_340, A[50], B[50]);
  nand g108 (n_335, A[50], B[50]);
  nor g109 (n_336, A[51], B[51]);
  nand g110 (n_337, A[51], B[51]);
  nor g111 (n_346, A[52], B[52]);
  nand g112 (n_341, A[52], B[52]);
  nor g113 (n_342, A[53], B[53]);
  nand g114 (n_343, A[53], B[53]);
  nor g115 (n_352, A[54], B[54]);
  nand g116 (n_347, A[54], B[54]);
  nor g117 (n_348, A[55], B[55]);
  nand g118 (n_349, A[55], B[55]);
  nor g119 (n_358, A[56], B[56]);
  nand g120 (n_353, A[56], B[56]);
  nor g121 (n_354, A[57], B[57]);
  nand g122 (n_355, A[57], B[57]);
  nand g127 (n_360, n_189, n_190);
  nor g128 (n_194, n_191, n_192);
  nor g131 (n_359, n_196, n_192);
  nor g132 (n_200, n_197, n_198);
  nor g135 (n_369, n_202, n_198);
  nor g136 (n_206, n_203, n_204);
  nor g139 (n_363, n_208, n_204);
  nor g140 (n_212, n_209, n_210);
  nor g143 (n_376, n_214, n_210);
  nor g144 (n_218, n_215, n_216);
  nor g147 (n_370, n_220, n_216);
  nor g148 (n_224, n_221, n_222);
  nor g151 (n_383, n_226, n_222);
  nor g152 (n_230, n_227, n_228);
  nor g155 (n_377, n_232, n_228);
  nor g156 (n_236, n_233, n_234);
  nor g159 (n_390, n_238, n_234);
  nor g160 (n_242, n_239, n_240);
  nor g163 (n_384, n_244, n_240);
  nor g164 (n_248, n_245, n_246);
  nor g167 (n_397, n_250, n_246);
  nor g168 (n_254, n_251, n_252);
  nor g171 (n_391, n_256, n_252);
  nor g172 (n_260, n_257, n_258);
  nor g175 (n_404, n_262, n_258);
  nor g176 (n_266, n_263, n_264);
  nor g179 (n_398, n_268, n_264);
  nor g180 (n_272, n_269, n_270);
  nor g183 (n_411, n_274, n_270);
  nor g184 (n_278, n_275, n_276);
  nor g187 (n_405, n_280, n_276);
  nor g188 (n_284, n_281, n_282);
  nor g191 (n_418, n_286, n_282);
  nor g192 (n_290, n_287, n_288);
  nor g195 (n_412, n_292, n_288);
  nor g196 (n_296, n_293, n_294);
  nor g199 (n_425, n_298, n_294);
  nor g200 (n_302, n_299, n_300);
  nor g203 (n_419, n_304, n_300);
  nor g204 (n_308, n_305, n_306);
  nor g207 (n_432, n_310, n_306);
  nor g208 (n_314, n_311, n_312);
  nor g211 (n_426, n_316, n_312);
  nor g212 (n_320, n_317, n_318);
  nor g215 (n_439, n_322, n_318);
  nor g216 (n_326, n_323, n_324);
  nor g219 (n_433, n_328, n_324);
  nor g220 (n_332, n_329, n_330);
  nor g223 (n_446, n_334, n_330);
  nor g224 (n_338, n_335, n_336);
  nor g227 (n_440, n_340, n_336);
  nor g228 (n_344, n_341, n_342);
  nor g231 (n_453, n_346, n_342);
  nor g232 (n_350, n_347, n_348);
  nor g235 (n_447, n_352, n_348);
  nor g236 (n_356, n_353, n_354);
  nor g239 (n_562, n_358, n_354);
  nand g240 (n_362, n_359, n_360);
  nand g241 (n_455, n_361, n_362);
  nand g246 (n_454, n_369, n_363);
  nand g251 (n_464, n_376, n_370);
  nand g256 (n_459, n_383, n_377);
  nand g261 (n_470, n_390, n_384);
  nand g266 (n_465, n_397, n_391);
  nand g271 (n_476, n_404, n_398);
  nand g276 (n_471, n_411, n_405);
  nand g281 (n_482, n_418, n_412);
  nand g286 (n_477, n_425, n_419);
  nand g291 (n_488, n_432, n_426);
  nand g296 (n_483, n_439, n_433);
  nand g301 (n_494, n_446, n_440);
  nand g306 (n_489, n_453, n_447);
  nand g309 (n_496, n_457, n_458);
  nor g310 (n_462, n_459, n_460);
  nor g313 (n_495, n_464, n_459);
  nor g314 (n_468, n_465, n_466);
  nor g317 (n_505, n_470, n_465);
  nor g318 (n_474, n_471, n_472);
  nor g321 (n_499, n_476, n_471);
  nor g322 (n_480, n_477, n_478);
  nor g325 (n_512, n_482, n_477);
  nor g326 (n_486, n_483, n_484);
  nor g329 (n_506, n_488, n_483);
  nor g330 (n_492, n_489, n_490);
  nor g333 (n_525, n_494, n_489);
  nand g334 (n_498, n_495, n_496);
  nand g335 (n_514, n_497, n_498);
  nand g340 (n_513, n_505, n_499);
  nand g345 (n_518, n_512, n_506);
  nand g348 (n_519, n_516, n_517);
  nand g351 (n_526, n_521, n_522);
  nand g352 (n_523, n_505, n_514);
  nand g353 (n_533, n_500, n_523);
  nand g354 (n_524, n_512, n_519);
  nand g355 (n_538, n_507, n_524);
  nand g356 (n_528, n_525, n_526);
  nand g357 (n_563, n_527, n_528);
  nand g360 (n_545, n_460, n_530);
  nand g363 (n_548, n_466, n_532);
  nand g366 (n_551, n_472, n_535);
  nand g369 (n_554, n_478, n_537);
  nand g372 (n_557, n_484, n_540);
  nand g375 (n_560, n_490, n_542);
  nand g376 (n_543, n_369, n_455);
  nand g377 (n_570, n_364, n_543);
  nand g378 (n_544, n_376, n_496);
  nand g379 (n_575, n_371, n_544);
  nand g380 (n_546, n_383, n_545);
  nand g381 (n_580, n_378, n_546);
  nand g382 (n_547, n_390, n_514);
  nand g383 (n_585, n_385, n_547);
  nand g384 (n_549, n_397, n_548);
  nand g385 (n_590, n_392, n_549);
  nand g386 (n_550, n_404, n_533);
  nand g387 (n_595, n_399, n_550);
  nand g388 (n_552, n_411, n_551);
  nand g389 (n_600, n_406, n_552);
  nand g390 (n_553, n_418, n_519);
  nand g391 (n_605, n_413, n_553);
  nand g392 (n_555, n_425, n_554);
  nand g393 (n_610, n_420, n_555);
  nand g394 (n_556, n_432, n_538);
  nand g395 (n_615, n_427, n_556);
  nand g396 (n_558, n_439, n_557);
  nand g397 (n_620, n_434, n_558);
  nand g398 (n_559, n_446, n_526);
  nand g399 (n_625, n_441, n_559);
  nand g400 (n_561, n_453, n_560);
  nand g401 (n_630, n_448, n_561);
  nand g402 (n_565, n_562, n_563);
  nand g403 (n_636, n_564, n_565);
  nand g406 (n_643, n_191, n_567);
  nand g409 (n_647, n_197, n_569);
  nand g412 (n_651, n_203, n_572);
  nand g415 (n_655, n_209, n_574);
  nand g418 (n_659, n_215, n_577);
  nand g421 (n_663, n_221, n_579);
  nand g424 (n_667, n_227, n_582);
  nand g427 (n_671, n_233, n_584);
  nand g430 (n_675, n_239, n_587);
  nand g433 (n_679, n_245, n_589);
  nand g436 (n_683, n_251, n_592);
  nand g439 (n_687, n_257, n_594);
  nand g442 (n_691, n_263, n_597);
  nand g445 (n_695, n_269, n_599);
  nand g448 (n_699, n_275, n_602);
  nand g451 (n_703, n_281, n_604);
  nand g454 (n_707, n_287, n_607);
  nand g457 (n_711, n_293, n_609);
  nand g460 (n_715, n_299, n_612);
  nand g463 (n_719, n_305, n_614);
  nand g466 (n_723, n_311, n_617);
  nand g469 (n_727, n_317, n_619);
  nand g472 (n_731, n_323, n_622);
  nand g475 (n_735, n_329, n_624);
  nand g478 (n_739, n_335, n_627);
  nand g481 (n_743, n_341, n_629);
  nand g484 (n_747, n_347, n_632);
  nand g487 (n_751, n_353, n_634);
  nand g490 (n_182, n_638, n_639);
  xnor g494 (Z[2], n_360, n_641);
  xnor g497 (Z[3], n_643, n_644);
  xnor g499 (Z[4], n_455, n_645);
  xnor g502 (Z[5], n_647, n_648);
  xnor g504 (Z[6], n_570, n_649);
  xnor g507 (Z[7], n_651, n_652);
  xnor g509 (Z[8], n_496, n_653);
  xnor g512 (Z[9], n_655, n_656);
  xnor g514 (Z[10], n_575, n_657);
  xnor g517 (Z[11], n_659, n_660);
  xnor g519 (Z[12], n_545, n_661);
  xnor g522 (Z[13], n_663, n_664);
  xnor g524 (Z[14], n_580, n_665);
  xnor g527 (Z[15], n_667, n_668);
  xnor g529 (Z[16], n_514, n_669);
  xnor g532 (Z[17], n_671, n_672);
  xnor g534 (Z[18], n_585, n_673);
  xnor g537 (Z[19], n_675, n_676);
  xnor g539 (Z[20], n_548, n_677);
  xnor g542 (Z[21], n_679, n_680);
  xnor g544 (Z[22], n_590, n_681);
  xnor g547 (Z[23], n_683, n_684);
  xnor g549 (Z[24], n_533, n_685);
  xnor g552 (Z[25], n_687, n_688);
  xnor g554 (Z[26], n_595, n_689);
  xnor g557 (Z[27], n_691, n_692);
  xnor g559 (Z[28], n_551, n_693);
  xnor g562 (Z[29], n_695, n_696);
  xnor g564 (Z[30], n_600, n_697);
  xnor g567 (Z[31], n_699, n_700);
  xnor g569 (Z[32], n_519, n_701);
  xnor g572 (Z[33], n_703, n_704);
  xnor g574 (Z[34], n_605, n_705);
  xnor g577 (Z[35], n_707, n_708);
  xnor g579 (Z[36], n_554, n_709);
  xnor g582 (Z[37], n_711, n_712);
  xnor g584 (Z[38], n_610, n_713);
  xnor g587 (Z[39], n_715, n_716);
  xnor g589 (Z[40], n_538, n_717);
  xnor g592 (Z[41], n_719, n_720);
  xnor g594 (Z[42], n_615, n_721);
  xnor g597 (Z[43], n_723, n_724);
  xnor g599 (Z[44], n_557, n_725);
  xnor g602 (Z[45], n_727, n_728);
  xnor g604 (Z[46], n_620, n_729);
  xnor g607 (Z[47], n_731, n_732);
  xnor g609 (Z[48], n_526, n_733);
  xnor g612 (Z[49], n_735, n_736);
  xnor g614 (Z[50], n_625, n_737);
  xnor g617 (Z[51], n_739, n_740);
  xnor g619 (Z[52], n_560, n_741);
  xnor g622 (Z[53], n_743, n_744);
  xnor g624 (Z[54], n_630, n_745);
  xnor g627 (Z[55], n_747, n_748);
  xnor g629 (Z[56], n_563, n_749);
  xnor g632 (Z[57], n_751, n_752);
  xnor g634 (Z[58], n_636, n_753);
  or g637 (n_638, A[58], B[58]);
  and g638 (n_635, A[58], B[58]);
  and g639 (n_564, wc, n_355);
  not gc (wc, n_356);
  and g640 (n_441, wc0, n_331);
  not gc0 (wc0, n_332);
  and g641 (n_443, wc1, n_337);
  not gc1 (wc1, n_338);
  and g642 (n_448, wc2, n_343);
  not gc2 (wc2, n_344);
  and g643 (n_450, wc3, n_349);
  not gc3 (wc3, n_350);
  and g644 (n_413, wc4, n_283);
  not gc4 (wc4, n_284);
  and g645 (n_415, wc5, n_289);
  not gc5 (wc5, n_290);
  and g646 (n_420, wc6, n_295);
  not gc6 (wc6, n_296);
  and g647 (n_422, wc7, n_301);
  not gc7 (wc7, n_302);
  and g648 (n_427, wc8, n_307);
  not gc8 (wc8, n_308);
  and g649 (n_429, wc9, n_313);
  not gc9 (wc9, n_314);
  and g650 (n_434, wc10, n_319);
  not gc10 (wc10, n_320);
  and g651 (n_436, wc11, n_325);
  not gc11 (wc11, n_326);
  and g652 (n_385, wc12, n_235);
  not gc12 (wc12, n_236);
  and g653 (n_387, wc13, n_241);
  not gc13 (wc13, n_242);
  and g654 (n_392, wc14, n_247);
  not gc14 (wc14, n_248);
  and g655 (n_394, wc15, n_253);
  not gc15 (wc15, n_254);
  and g656 (n_399, wc16, n_259);
  not gc16 (wc16, n_260);
  and g657 (n_401, wc17, n_265);
  not gc17 (wc17, n_266);
  and g658 (n_406, wc18, n_271);
  not gc18 (wc18, n_272);
  and g659 (n_408, wc19, n_277);
  not gc19 (wc19, n_278);
  and g660 (n_371, wc20, n_211);
  not gc20 (wc20, n_212);
  and g661 (n_373, wc21, n_217);
  not gc21 (wc21, n_218);
  and g662 (n_378, wc22, n_223);
  not gc22 (wc22, n_224);
  and g663 (n_380, wc23, n_229);
  not gc23 (wc23, n_230);
  and g664 (n_364, wc24, n_199);
  not gc24 (wc24, n_200);
  and g665 (n_366, wc25, n_205);
  not gc25 (wc25, n_206);
  and g666 (n_361, wc26, n_193);
  not gc26 (wc26, n_194);
  or g667 (n_190, n_183, n_186);
  or g668 (n_640, wc27, n_186);
  not gc27 (wc27, n_189);
  or g669 (n_641, wc28, n_196);
  not gc28 (wc28, n_191);
  or g670 (n_644, wc29, n_192);
  not gc29 (wc29, n_193);
  or g671 (n_645, wc30, n_202);
  not gc30 (wc30, n_197);
  or g672 (n_648, wc31, n_198);
  not gc31 (wc31, n_199);
  or g673 (n_649, wc32, n_208);
  not gc32 (wc32, n_203);
  or g674 (n_652, wc33, n_204);
  not gc33 (wc33, n_205);
  or g675 (n_653, wc34, n_214);
  not gc34 (wc34, n_209);
  or g676 (n_656, wc35, n_210);
  not gc35 (wc35, n_211);
  or g677 (n_657, wc36, n_220);
  not gc36 (wc36, n_215);
  or g678 (n_660, wc37, n_216);
  not gc37 (wc37, n_217);
  or g679 (n_661, wc38, n_226);
  not gc38 (wc38, n_221);
  or g680 (n_664, wc39, n_222);
  not gc39 (wc39, n_223);
  or g681 (n_665, wc40, n_232);
  not gc40 (wc40, n_227);
  or g682 (n_668, wc41, n_228);
  not gc41 (wc41, n_229);
  or g683 (n_669, wc42, n_238);
  not gc42 (wc42, n_233);
  or g684 (n_672, wc43, n_234);
  not gc43 (wc43, n_235);
  or g685 (n_673, wc44, n_244);
  not gc44 (wc44, n_239);
  or g686 (n_676, wc45, n_240);
  not gc45 (wc45, n_241);
  or g687 (n_677, wc46, n_250);
  not gc46 (wc46, n_245);
  or g688 (n_680, wc47, n_246);
  not gc47 (wc47, n_247);
  or g689 (n_681, wc48, n_256);
  not gc48 (wc48, n_251);
  or g690 (n_684, wc49, n_252);
  not gc49 (wc49, n_253);
  or g691 (n_685, wc50, n_262);
  not gc50 (wc50, n_257);
  or g692 (n_688, wc51, n_258);
  not gc51 (wc51, n_259);
  or g693 (n_689, wc52, n_268);
  not gc52 (wc52, n_263);
  or g694 (n_692, wc53, n_264);
  not gc53 (wc53, n_265);
  or g695 (n_693, wc54, n_274);
  not gc54 (wc54, n_269);
  or g696 (n_696, wc55, n_270);
  not gc55 (wc55, n_271);
  or g697 (n_697, wc56, n_280);
  not gc56 (wc56, n_275);
  or g698 (n_700, wc57, n_276);
  not gc57 (wc57, n_277);
  or g699 (n_701, wc58, n_286);
  not gc58 (wc58, n_281);
  or g700 (n_704, wc59, n_282);
  not gc59 (wc59, n_283);
  or g701 (n_705, wc60, n_292);
  not gc60 (wc60, n_287);
  or g702 (n_708, wc61, n_288);
  not gc61 (wc61, n_289);
  or g703 (n_709, wc62, n_298);
  not gc62 (wc62, n_293);
  or g704 (n_712, wc63, n_294);
  not gc63 (wc63, n_295);
  or g705 (n_713, wc64, n_304);
  not gc64 (wc64, n_299);
  or g706 (n_716, wc65, n_300);
  not gc65 (wc65, n_301);
  or g707 (n_717, wc66, n_310);
  not gc66 (wc66, n_305);
  or g708 (n_720, wc67, n_306);
  not gc67 (wc67, n_307);
  or g709 (n_721, wc68, n_316);
  not gc68 (wc68, n_311);
  or g710 (n_724, wc69, n_312);
  not gc69 (wc69, n_313);
  or g711 (n_725, wc70, n_322);
  not gc70 (wc70, n_317);
  or g712 (n_728, wc71, n_318);
  not gc71 (wc71, n_319);
  or g713 (n_729, wc72, n_328);
  not gc72 (wc72, n_323);
  or g714 (n_732, wc73, n_324);
  not gc73 (wc73, n_325);
  or g715 (n_733, wc74, n_334);
  not gc74 (wc74, n_329);
  or g716 (n_736, wc75, n_330);
  not gc75 (wc75, n_331);
  or g717 (n_737, wc76, n_340);
  not gc76 (wc76, n_335);
  or g718 (n_740, wc77, n_336);
  not gc77 (wc77, n_337);
  or g719 (n_741, wc78, n_346);
  not gc78 (wc78, n_341);
  or g720 (n_744, wc79, n_342);
  not gc79 (wc79, n_343);
  or g721 (n_745, wc80, n_352);
  not gc80 (wc80, n_347);
  or g722 (n_748, wc81, n_348);
  not gc81 (wc81, n_349);
  or g723 (n_749, wc82, n_358);
  not gc82 (wc82, n_353);
  or g724 (n_752, wc83, n_354);
  not gc83 (wc83, n_355);
  and g725 (n_444, wc84, n_440);
  not gc84 (wc84, n_441);
  and g726 (n_451, wc85, n_447);
  not gc85 (wc85, n_448);
  and g727 (n_416, wc86, n_412);
  not gc86 (wc86, n_413);
  and g728 (n_423, wc87, n_419);
  not gc87 (wc87, n_420);
  and g729 (n_430, wc88, n_426);
  not gc88 (wc88, n_427);
  and g730 (n_437, wc89, n_433);
  not gc89 (wc89, n_434);
  and g731 (n_388, wc90, n_384);
  not gc90 (wc90, n_385);
  and g732 (n_395, wc91, n_391);
  not gc91 (wc91, n_392);
  and g733 (n_402, wc92, n_398);
  not gc92 (wc92, n_399);
  and g734 (n_409, wc93, n_405);
  not gc93 (wc93, n_406);
  and g735 (n_374, wc94, n_370);
  not gc94 (wc94, n_371);
  and g736 (n_381, wc95, n_377);
  not gc95 (wc95, n_378);
  and g737 (n_367, wc96, n_363);
  not gc96 (wc96, n_364);
  xor g738 (Z[1], n_183, n_640);
  or g739 (n_753, n_635, wc97);
  not gc97 (wc97, n_638);
  and g740 (n_490, wc98, n_443);
  not gc98 (wc98, n_444);
  and g741 (n_491, wc99, n_450);
  not gc99 (wc99, n_451);
  and g742 (n_478, wc100, n_415);
  not gc100 (wc100, n_416);
  and g743 (n_479, wc101, n_422);
  not gc101 (wc101, n_423);
  and g744 (n_484, wc102, n_429);
  not gc102 (wc102, n_430);
  and g745 (n_485, wc103, n_436);
  not gc103 (wc103, n_437);
  and g746 (n_466, wc104, n_387);
  not gc104 (wc104, n_388);
  and g747 (n_467, wc105, n_394);
  not gc105 (wc105, n_395);
  and g748 (n_472, wc106, n_401);
  not gc106 (wc106, n_402);
  and g749 (n_473, wc107, n_408);
  not gc107 (wc107, n_409);
  and g750 (n_460, wc108, n_373);
  not gc108 (wc108, n_374);
  and g751 (n_461, wc109, n_380);
  not gc109 (wc109, n_381);
  and g752 (n_457, wc110, n_366);
  not gc110 (wc110, n_367);
  or g753 (n_567, wc111, n_196);
  not gc111 (wc111, n_360);
  and g754 (n_527, n_491, wc112);
  not gc112 (wc112, n_492);
  and g755 (n_507, n_479, wc113);
  not gc113 (wc113, n_480);
  and g756 (n_509, n_485, wc114);
  not gc114 (wc114, n_486);
  and g757 (n_500, n_467, wc115);
  not gc115 (wc115, n_468);
  and g758 (n_502, n_473, wc116);
  not gc116 (wc116, n_474);
  and g759 (n_497, n_461, wc117);
  not gc117 (wc117, n_462);
  or g760 (n_458, n_454, wc118);
  not gc118 (wc118, n_455);
  or g761 (n_569, wc119, n_202);
  not gc119 (wc119, n_455);
  and g762 (n_510, wc120, n_506);
  not gc120 (wc120, n_507);
  and g763 (n_503, wc121, n_499);
  not gc121 (wc121, n_500);
  and g764 (n_521, wc122, n_509);
  not gc122 (wc122, n_510);
  and g765 (n_516, wc123, n_502);
  not gc123 (wc123, n_503);
  or g766 (n_530, wc124, n_464);
  not gc124 (wc124, n_496);
  or g767 (n_572, wc125, n_208);
  not gc125 (wc125, n_570);
  or g768 (n_574, wc126, n_214);
  not gc126 (wc126, n_496);
  or g769 (n_517, n_513, wc127);
  not gc127 (wc127, n_514);
  or g770 (n_532, wc128, n_470);
  not gc128 (wc128, n_514);
  or g771 (n_577, wc129, n_220);
  not gc129 (wc129, n_575);
  or g772 (n_579, wc130, n_226);
  not gc130 (wc130, n_545);
  or g773 (n_584, wc131, n_238);
  not gc131 (wc131, n_514);
  or g774 (n_522, wc132, n_518);
  not gc132 (wc132, n_519);
  or g775 (n_535, wc133, n_476);
  not gc133 (wc133, n_533);
  or g776 (n_537, wc134, n_482);
  not gc134 (wc134, n_519);
  or g777 (n_582, wc135, n_232);
  not gc135 (wc135, n_580);
  or g778 (n_587, wc136, n_244);
  not gc136 (wc136, n_585);
  or g779 (n_589, wc137, n_250);
  not gc137 (wc137, n_548);
  or g780 (n_594, wc138, n_262);
  not gc138 (wc138, n_533);
  or g781 (n_604, wc139, n_286);
  not gc139 (wc139, n_519);
  or g782 (n_540, wc140, n_488);
  not gc140 (wc140, n_538);
  or g783 (n_542, wc141, n_494);
  not gc141 (wc141, n_526);
  or g784 (n_592, wc142, n_256);
  not gc142 (wc142, n_590);
  or g785 (n_597, wc143, n_268);
  not gc143 (wc143, n_595);
  or g786 (n_599, wc144, n_274);
  not gc144 (wc144, n_551);
  or g787 (n_607, wc145, n_292);
  not gc145 (wc145, n_605);
  or g788 (n_609, wc146, n_298);
  not gc146 (wc146, n_554);
  or g789 (n_614, wc147, n_310);
  not gc147 (wc147, n_538);
  or g790 (n_624, wc148, n_334);
  not gc148 (wc148, n_526);
  or g791 (n_602, wc149, n_280);
  not gc149 (wc149, n_600);
  or g792 (n_612, wc150, n_304);
  not gc150 (wc150, n_610);
  or g793 (n_617, wc151, n_316);
  not gc151 (wc151, n_615);
  or g794 (n_619, wc152, n_322);
  not gc152 (wc152, n_557);
  or g795 (n_627, wc153, n_340);
  not gc153 (wc153, n_625);
  or g796 (n_629, wc154, n_346);
  not gc154 (wc154, n_560);
  or g797 (n_634, wc155, n_358);
  not gc155 (wc155, n_563);
  or g798 (n_639, n_635, wc156);
  not gc156 (wc156, n_636);
  or g799 (n_622, wc157, n_328);
  not gc157 (wc157, n_620);
  or g800 (n_632, wc158, n_352);
  not gc158 (wc158, n_630);
endmodule

module add_signed_4709_2_GENERIC(A, B, Z);
  input [58:0] A, B;
  output [59:0] Z;
  wire [58:0] A, B;
  wire [59:0] Z;
  add_signed_4709_2_GENERIC_REAL g1(.A ({A[58:2], A[0], A[0]}), .B (B),
       .Z (Z));
endmodule

module add_signed_4709_3_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [58:0] A, B;
  output [59:0] Z;
  wire [58:0] A, B;
  wire [59:0] Z;
  wire n_182, n_183, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476;
  not g3 (Z[59], n_182);
  nand g4 (n_183, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_188, A[1], B[1]);
  nand g13 (n_192, n_188, n_189, n_190);
  xor g14 (n_191, A[1], B[1]);
  nand g16 (n_193, A[2], B[2]);
  nand g17 (n_194, A[2], n_192);
  nand g18 (n_195, B[2], n_192);
  nand g19 (n_197, n_193, n_194, n_195);
  xor g20 (n_196, A[2], B[2]);
  xor g21 (Z[2], n_192, n_196);
  nand g22 (n_198, A[3], B[3]);
  nand g23 (n_199, A[3], n_197);
  nand g24 (n_200, B[3], n_197);
  nand g25 (n_202, n_198, n_199, n_200);
  xor g26 (n_201, A[3], B[3]);
  xor g27 (Z[3], n_197, n_201);
  nand g28 (n_203, A[4], B[4]);
  nand g29 (n_204, A[4], n_202);
  nand g30 (n_205, B[4], n_202);
  nand g31 (n_207, n_203, n_204, n_205);
  xor g32 (n_206, A[4], B[4]);
  xor g33 (Z[4], n_202, n_206);
  nand g34 (n_208, A[5], B[5]);
  nand g35 (n_209, A[5], n_207);
  nand g36 (n_210, B[5], n_207);
  nand g37 (n_212, n_208, n_209, n_210);
  xor g38 (n_211, A[5], B[5]);
  xor g39 (Z[5], n_207, n_211);
  nand g40 (n_213, A[6], B[6]);
  nand g41 (n_214, A[6], n_212);
  nand g42 (n_215, B[6], n_212);
  nand g43 (n_217, n_213, n_214, n_215);
  xor g44 (n_216, A[6], B[6]);
  xor g45 (Z[6], n_212, n_216);
  nand g46 (n_218, A[7], B[7]);
  nand g47 (n_219, A[7], n_217);
  nand g48 (n_220, B[7], n_217);
  nand g49 (n_222, n_218, n_219, n_220);
  xor g50 (n_221, A[7], B[7]);
  xor g51 (Z[7], n_217, n_221);
  nand g52 (n_223, A[8], B[8]);
  nand g53 (n_224, A[8], n_222);
  nand g54 (n_225, B[8], n_222);
  nand g55 (n_227, n_223, n_224, n_225);
  xor g56 (n_226, A[8], B[8]);
  xor g57 (Z[8], n_222, n_226);
  nand g58 (n_228, A[9], B[9]);
  nand g59 (n_229, A[9], n_227);
  nand g60 (n_230, B[9], n_227);
  nand g61 (n_232, n_228, n_229, n_230);
  xor g62 (n_231, A[9], B[9]);
  xor g63 (Z[9], n_227, n_231);
  nand g64 (n_233, A[10], B[10]);
  nand g65 (n_234, A[10], n_232);
  nand g66 (n_235, B[10], n_232);
  nand g67 (n_237, n_233, n_234, n_235);
  xor g68 (n_236, A[10], B[10]);
  xor g69 (Z[10], n_232, n_236);
  nand g70 (n_238, A[11], B[11]);
  nand g71 (n_239, A[11], n_237);
  nand g72 (n_240, B[11], n_237);
  nand g73 (n_242, n_238, n_239, n_240);
  xor g74 (n_241, A[11], B[11]);
  xor g75 (Z[11], n_237, n_241);
  nand g76 (n_243, A[12], B[12]);
  nand g77 (n_244, A[12], n_242);
  nand g78 (n_245, B[12], n_242);
  nand g79 (n_247, n_243, n_244, n_245);
  xor g80 (n_246, A[12], B[12]);
  xor g81 (Z[12], n_242, n_246);
  nand g82 (n_248, A[13], B[13]);
  nand g83 (n_249, A[13], n_247);
  nand g84 (n_250, B[13], n_247);
  nand g85 (n_252, n_248, n_249, n_250);
  xor g86 (n_251, A[13], B[13]);
  xor g87 (Z[13], n_247, n_251);
  nand g88 (n_253, A[14], B[14]);
  nand g89 (n_254, A[14], n_252);
  nand g90 (n_255, B[14], n_252);
  nand g91 (n_257, n_253, n_254, n_255);
  xor g92 (n_256, A[14], B[14]);
  xor g93 (Z[14], n_252, n_256);
  nand g94 (n_258, A[15], B[15]);
  nand g95 (n_259, A[15], n_257);
  nand g96 (n_260, B[15], n_257);
  nand g97 (n_262, n_258, n_259, n_260);
  xor g98 (n_261, A[15], B[15]);
  xor g99 (Z[15], n_257, n_261);
  nand g100 (n_263, A[16], B[16]);
  nand g101 (n_264, A[16], n_262);
  nand g102 (n_265, B[16], n_262);
  nand g103 (n_267, n_263, n_264, n_265);
  xor g104 (n_266, A[16], B[16]);
  xor g105 (Z[16], n_262, n_266);
  nand g106 (n_268, A[17], B[17]);
  nand g107 (n_269, A[17], n_267);
  nand g108 (n_270, B[17], n_267);
  nand g109 (n_272, n_268, n_269, n_270);
  xor g110 (n_271, A[17], B[17]);
  xor g111 (Z[17], n_267, n_271);
  nand g112 (n_273, A[18], B[18]);
  nand g113 (n_274, A[18], n_272);
  nand g114 (n_275, B[18], n_272);
  nand g115 (n_277, n_273, n_274, n_275);
  xor g116 (n_276, A[18], B[18]);
  xor g117 (Z[18], n_272, n_276);
  nand g118 (n_278, A[19], B[19]);
  nand g119 (n_279, A[19], n_277);
  nand g120 (n_280, B[19], n_277);
  nand g121 (n_282, n_278, n_279, n_280);
  xor g122 (n_281, A[19], B[19]);
  xor g123 (Z[19], n_277, n_281);
  nand g124 (n_283, A[20], B[20]);
  nand g125 (n_284, A[20], n_282);
  nand g126 (n_285, B[20], n_282);
  nand g127 (n_287, n_283, n_284, n_285);
  xor g128 (n_286, A[20], B[20]);
  xor g129 (Z[20], n_282, n_286);
  nand g130 (n_288, A[21], B[21]);
  nand g131 (n_289, A[21], n_287);
  nand g132 (n_290, B[21], n_287);
  nand g133 (n_292, n_288, n_289, n_290);
  xor g134 (n_291, A[21], B[21]);
  xor g135 (Z[21], n_287, n_291);
  nand g136 (n_293, A[22], B[22]);
  nand g137 (n_294, A[22], n_292);
  nand g138 (n_295, B[22], n_292);
  nand g139 (n_297, n_293, n_294, n_295);
  xor g140 (n_296, A[22], B[22]);
  xor g141 (Z[22], n_292, n_296);
  nand g142 (n_298, A[23], B[23]);
  nand g143 (n_299, A[23], n_297);
  nand g144 (n_300, B[23], n_297);
  nand g145 (n_302, n_298, n_299, n_300);
  xor g146 (n_301, A[23], B[23]);
  xor g147 (Z[23], n_297, n_301);
  nand g148 (n_303, A[24], B[24]);
  nand g149 (n_304, A[24], n_302);
  nand g150 (n_305, B[24], n_302);
  nand g151 (n_307, n_303, n_304, n_305);
  xor g152 (n_306, A[24], B[24]);
  xor g153 (Z[24], n_302, n_306);
  nand g154 (n_308, A[25], B[25]);
  nand g155 (n_309, A[25], n_307);
  nand g156 (n_310, B[25], n_307);
  nand g157 (n_312, n_308, n_309, n_310);
  xor g158 (n_311, A[25], B[25]);
  xor g159 (Z[25], n_307, n_311);
  nand g160 (n_313, A[26], B[26]);
  nand g161 (n_314, A[26], n_312);
  nand g162 (n_315, B[26], n_312);
  nand g163 (n_317, n_313, n_314, n_315);
  xor g164 (n_316, A[26], B[26]);
  xor g165 (Z[26], n_312, n_316);
  nand g166 (n_318, A[27], B[27]);
  nand g167 (n_319, A[27], n_317);
  nand g168 (n_320, B[27], n_317);
  nand g169 (n_322, n_318, n_319, n_320);
  xor g170 (n_321, A[27], B[27]);
  xor g171 (Z[27], n_317, n_321);
  nand g172 (n_323, A[28], B[28]);
  nand g173 (n_324, A[28], n_322);
  nand g174 (n_325, B[28], n_322);
  nand g175 (n_327, n_323, n_324, n_325);
  xor g176 (n_326, A[28], B[28]);
  xor g177 (Z[28], n_322, n_326);
  nand g178 (n_328, A[29], B[29]);
  nand g179 (n_329, A[29], n_327);
  nand g180 (n_330, B[29], n_327);
  nand g181 (n_332, n_328, n_329, n_330);
  xor g182 (n_331, A[29], B[29]);
  xor g183 (Z[29], n_327, n_331);
  nand g184 (n_333, A[30], B[30]);
  nand g185 (n_334, A[30], n_332);
  nand g186 (n_335, B[30], n_332);
  nand g187 (n_337, n_333, n_334, n_335);
  xor g188 (n_336, A[30], B[30]);
  xor g189 (Z[30], n_332, n_336);
  nand g190 (n_338, A[31], B[31]);
  nand g191 (n_339, A[31], n_337);
  nand g192 (n_340, B[31], n_337);
  nand g193 (n_342, n_338, n_339, n_340);
  xor g194 (n_341, A[31], B[31]);
  xor g195 (Z[31], n_337, n_341);
  nand g196 (n_343, A[32], B[32]);
  nand g197 (n_344, A[32], n_342);
  nand g198 (n_345, B[32], n_342);
  nand g199 (n_347, n_343, n_344, n_345);
  xor g200 (n_346, A[32], B[32]);
  xor g201 (Z[32], n_342, n_346);
  nand g202 (n_348, A[33], B[33]);
  nand g203 (n_349, A[33], n_347);
  nand g204 (n_350, B[33], n_347);
  nand g205 (n_352, n_348, n_349, n_350);
  xor g206 (n_351, A[33], B[33]);
  xor g207 (Z[33], n_347, n_351);
  nand g208 (n_353, A[34], B[34]);
  nand g209 (n_354, A[34], n_352);
  nand g210 (n_355, B[34], n_352);
  nand g211 (n_357, n_353, n_354, n_355);
  xor g212 (n_356, A[34], B[34]);
  xor g213 (Z[34], n_352, n_356);
  nand g214 (n_358, A[35], B[35]);
  nand g215 (n_359, A[35], n_357);
  nand g216 (n_360, B[35], n_357);
  nand g217 (n_362, n_358, n_359, n_360);
  xor g218 (n_361, A[35], B[35]);
  xor g219 (Z[35], n_357, n_361);
  nand g220 (n_363, A[36], B[36]);
  nand g221 (n_364, A[36], n_362);
  nand g222 (n_365, B[36], n_362);
  nand g223 (n_367, n_363, n_364, n_365);
  xor g224 (n_366, A[36], B[36]);
  xor g225 (Z[36], n_362, n_366);
  nand g226 (n_368, A[37], B[37]);
  nand g227 (n_369, A[37], n_367);
  nand g228 (n_370, B[37], n_367);
  nand g229 (n_372, n_368, n_369, n_370);
  xor g230 (n_371, A[37], B[37]);
  xor g231 (Z[37], n_367, n_371);
  nand g232 (n_373, A[38], B[38]);
  nand g233 (n_374, A[38], n_372);
  nand g234 (n_375, B[38], n_372);
  nand g235 (n_377, n_373, n_374, n_375);
  xor g236 (n_376, A[38], B[38]);
  xor g237 (Z[38], n_372, n_376);
  nand g238 (n_378, A[39], B[39]);
  nand g239 (n_379, A[39], n_377);
  nand g240 (n_380, B[39], n_377);
  nand g241 (n_382, n_378, n_379, n_380);
  xor g242 (n_381, A[39], B[39]);
  xor g243 (Z[39], n_377, n_381);
  nand g244 (n_383, A[40], B[40]);
  nand g245 (n_384, A[40], n_382);
  nand g246 (n_385, B[40], n_382);
  nand g247 (n_387, n_383, n_384, n_385);
  xor g248 (n_386, A[40], B[40]);
  xor g249 (Z[40], n_382, n_386);
  nand g250 (n_388, A[41], B[41]);
  nand g251 (n_389, A[41], n_387);
  nand g252 (n_390, B[41], n_387);
  nand g253 (n_392, n_388, n_389, n_390);
  xor g254 (n_391, A[41], B[41]);
  xor g255 (Z[41], n_387, n_391);
  nand g256 (n_393, A[42], B[42]);
  nand g257 (n_394, A[42], n_392);
  nand g258 (n_395, B[42], n_392);
  nand g259 (n_397, n_393, n_394, n_395);
  xor g260 (n_396, A[42], B[42]);
  xor g261 (Z[42], n_392, n_396);
  nand g262 (n_398, A[43], B[43]);
  nand g263 (n_399, A[43], n_397);
  nand g264 (n_400, B[43], n_397);
  nand g265 (n_402, n_398, n_399, n_400);
  xor g266 (n_401, A[43], B[43]);
  xor g267 (Z[43], n_397, n_401);
  nand g268 (n_403, A[44], B[44]);
  nand g269 (n_404, A[44], n_402);
  nand g270 (n_405, B[44], n_402);
  nand g271 (n_407, n_403, n_404, n_405);
  xor g272 (n_406, A[44], B[44]);
  xor g273 (Z[44], n_402, n_406);
  nand g274 (n_408, A[45], B[45]);
  nand g275 (n_409, A[45], n_407);
  nand g276 (n_410, B[45], n_407);
  nand g277 (n_412, n_408, n_409, n_410);
  xor g278 (n_411, A[45], B[45]);
  xor g279 (Z[45], n_407, n_411);
  nand g280 (n_413, A[46], B[46]);
  nand g281 (n_414, A[46], n_412);
  nand g282 (n_415, B[46], n_412);
  nand g283 (n_417, n_413, n_414, n_415);
  xor g284 (n_416, A[46], B[46]);
  xor g285 (Z[46], n_412, n_416);
  nand g286 (n_418, A[47], B[47]);
  nand g287 (n_419, A[47], n_417);
  nand g288 (n_420, B[47], n_417);
  nand g289 (n_422, n_418, n_419, n_420);
  xor g290 (n_421, A[47], B[47]);
  xor g291 (Z[47], n_417, n_421);
  nand g292 (n_423, A[48], B[48]);
  nand g293 (n_424, A[48], n_422);
  nand g294 (n_425, B[48], n_422);
  nand g295 (n_427, n_423, n_424, n_425);
  xor g296 (n_426, A[48], B[48]);
  xor g297 (Z[48], n_422, n_426);
  nand g298 (n_428, A[49], B[49]);
  nand g299 (n_429, A[49], n_427);
  nand g300 (n_430, B[49], n_427);
  nand g301 (n_432, n_428, n_429, n_430);
  xor g302 (n_431, A[49], B[49]);
  xor g303 (Z[49], n_427, n_431);
  nand g304 (n_433, A[50], B[50]);
  nand g305 (n_434, A[50], n_432);
  nand g306 (n_435, B[50], n_432);
  nand g307 (n_437, n_433, n_434, n_435);
  xor g308 (n_436, A[50], B[50]);
  xor g309 (Z[50], n_432, n_436);
  nand g310 (n_438, A[51], B[51]);
  nand g311 (n_439, A[51], n_437);
  nand g312 (n_440, B[51], n_437);
  nand g313 (n_442, n_438, n_439, n_440);
  xor g314 (n_441, A[51], B[51]);
  xor g315 (Z[51], n_437, n_441);
  nand g316 (n_443, A[52], B[52]);
  nand g317 (n_444, A[52], n_442);
  nand g318 (n_445, B[52], n_442);
  nand g319 (n_447, n_443, n_444, n_445);
  xor g320 (n_446, A[52], B[52]);
  xor g321 (Z[52], n_442, n_446);
  nand g322 (n_448, A[53], B[53]);
  nand g323 (n_449, A[53], n_447);
  nand g324 (n_450, B[53], n_447);
  nand g325 (n_452, n_448, n_449, n_450);
  xor g326 (n_451, A[53], B[53]);
  xor g327 (Z[53], n_447, n_451);
  nand g328 (n_453, A[54], B[54]);
  nand g329 (n_454, A[54], n_452);
  nand g330 (n_455, B[54], n_452);
  nand g331 (n_457, n_453, n_454, n_455);
  xor g332 (n_456, A[54], B[54]);
  xor g333 (Z[54], n_452, n_456);
  nand g334 (n_458, A[55], B[55]);
  nand g335 (n_459, A[55], n_457);
  nand g336 (n_460, B[55], n_457);
  nand g337 (n_462, n_458, n_459, n_460);
  xor g338 (n_461, A[55], B[55]);
  xor g339 (Z[55], n_457, n_461);
  nand g340 (n_463, A[56], B[56]);
  nand g341 (n_464, A[56], n_462);
  nand g342 (n_465, B[56], n_462);
  nand g343 (n_467, n_463, n_464, n_465);
  xor g344 (n_466, A[56], B[56]);
  xor g345 (Z[56], n_462, n_466);
  nand g346 (n_468, A[57], B[57]);
  nand g347 (n_469, A[57], n_467);
  nand g348 (n_470, B[57], n_467);
  nand g349 (n_472, n_468, n_469, n_470);
  xor g350 (n_471, A[57], B[57]);
  xor g351 (Z[57], n_467, n_471);
  nand g355 (n_182, n_473, n_474, n_475);
  xor g357 (Z[58], n_472, n_476);
  or g359 (n_473, A[58], B[58]);
  xor g360 (n_476, A[58], B[58]);
  or g361 (n_189, wc, n_183);
  not gc (wc, A[1]);
  or g362 (n_190, wc0, n_183);
  not gc0 (wc0, B[1]);
  xnor g363 (Z[1], n_183, n_191);
  or g364 (n_474, A[58], wc1);
  not gc1 (wc1, n_472);
  or g365 (n_475, B[58], wc2);
  not gc2 (wc2, n_472);
endmodule

module add_signed_4709_3_GENERIC(A, B, Z);
  input [58:0] A, B;
  output [59:0] Z;
  wire [58:0] A, B;
  wire [59:0] Z;
  add_signed_4709_3_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_508_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [36:0] A, B;
  output [37:0] Z;
  wire [36:0] A, B;
  wire [37:0] Z;
  wire n_116, n_117, n_120, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_130, n_131, n_132, n_133, n_134, n_136, n_137;
  wire n_138, n_139, n_140, n_142, n_143, n_144, n_145, n_146;
  wire n_148, n_149, n_150, n_151, n_152, n_154, n_155, n_156;
  wire n_157, n_158, n_160, n_161, n_162, n_163, n_164, n_166;
  wire n_167, n_168, n_169, n_170, n_172, n_173, n_174, n_175;
  wire n_176, n_178, n_179, n_180, n_181, n_182, n_184, n_185;
  wire n_186, n_187, n_188, n_190, n_191, n_192, n_193, n_194;
  wire n_196, n_197, n_198, n_199, n_200, n_202, n_203, n_204;
  wire n_205, n_206, n_208, n_209, n_210, n_211, n_212, n_214;
  wire n_215, n_216, n_217, n_218, n_220, n_221, n_222, n_223;
  wire n_224, n_226, n_227, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_236, n_238, n_240, n_241, n_243, n_244, n_246;
  wire n_248, n_250, n_251, n_253, n_254, n_256, n_258, n_260;
  wire n_261, n_263, n_264, n_266, n_268, n_270, n_271, n_273;
  wire n_274, n_276, n_278, n_280, n_281, n_283, n_284, n_286;
  wire n_288, n_290, n_291, n_293, n_294, n_296, n_298, n_300;
  wire n_301, n_303, n_304, n_306, n_308, n_310, n_311, n_313;
  wire n_315, n_316, n_317, n_319, n_320, n_321, n_323, n_324;
  wire n_325, n_326, n_328, n_330, n_332, n_333, n_334, n_336;
  wire n_337, n_338, n_340, n_341, n_343, n_345, n_347, n_348;
  wire n_349, n_351, n_352, n_353, n_355, n_356, n_358, n_360;
  wire n_362, n_363, n_364, n_366, n_367, n_368, n_370, n_371;
  wire n_372, n_373, n_375, n_376, n_378, n_379, n_380, n_382;
  wire n_383, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_401, n_404, n_406, n_407, n_408, n_411, n_414, n_416;
  wire n_417, n_419, n_421, n_422, n_424, n_426, n_427, n_429;
  wire n_431, n_432, n_434, n_436, n_437, n_438, n_440, n_441;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_456, n_457, n_458, n_460;
  wire n_461, n_462, n_464, n_465, n_466, n_468, n_469, n_470;
  wire n_472, n_473, n_474, n_476, n_477, n_478, n_480, n_481;
  wire n_482, n_484, n_485, n_486, n_488, n_489, n_490, n_492;
  wire n_493, n_495, n_496, n_497, n_498, n_499, n_500, n_502;
  wire n_503, n_504, n_506, n_507, n_508, n_509, n_511, n_512;
  wire n_513, n_515, n_516, n_517, n_518, n_520, n_521, n_523;
  wire n_524, n_526, n_527, n_528, n_529, n_531, n_532, n_533;
  wire n_535, n_536, n_537, n_538, n_540, n_541, n_543, n_544;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_556, n_557, n_558, n_559, n_561, n_562, n_564, n_565;
  wire n_567, n_568, n_569, n_570, n_572, n_573, n_574, n_576;
  wire n_577, n_578, n_579, n_581, n_582, n_584, n_585;
  not g3 (Z[37], n_116);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_117, A[0], B[0]);
  nor g9 (n_120, A[1], B[1]);
  nand g10 (n_123, A[1], B[1]);
  nor g11 (n_130, A[2], B[2]);
  nand g12 (n_125, A[2], B[2]);
  nor g13 (n_126, A[3], B[3]);
  nand g14 (n_127, A[3], B[3]);
  nor g15 (n_136, A[4], B[4]);
  nand g16 (n_131, A[4], B[4]);
  nor g17 (n_132, A[5], B[5]);
  nand g18 (n_133, A[5], B[5]);
  nor g19 (n_142, A[6], B[6]);
  nand g20 (n_137, A[6], B[6]);
  nor g21 (n_138, A[7], B[7]);
  nand g22 (n_139, A[7], B[7]);
  nor g23 (n_148, A[8], B[8]);
  nand g24 (n_143, A[8], B[8]);
  nor g25 (n_144, A[9], B[9]);
  nand g26 (n_145, A[9], B[9]);
  nor g27 (n_154, A[10], B[10]);
  nand g28 (n_149, A[10], B[10]);
  nor g29 (n_150, A[11], B[11]);
  nand g30 (n_151, A[11], B[11]);
  nor g31 (n_160, A[12], B[12]);
  nand g32 (n_155, A[12], B[12]);
  nor g33 (n_156, A[13], B[13]);
  nand g34 (n_157, A[13], B[13]);
  nor g35 (n_166, A[14], B[14]);
  nand g36 (n_161, A[14], B[14]);
  nor g37 (n_162, A[15], B[15]);
  nand g38 (n_163, A[15], B[15]);
  nor g39 (n_172, A[16], B[16]);
  nand g40 (n_167, A[16], B[16]);
  nor g41 (n_168, A[17], B[17]);
  nand g42 (n_169, A[17], B[17]);
  nor g43 (n_178, A[18], B[18]);
  nand g44 (n_173, A[18], B[18]);
  nor g45 (n_174, A[19], B[19]);
  nand g46 (n_175, A[19], B[19]);
  nor g47 (n_184, A[20], B[20]);
  nand g48 (n_179, A[20], B[20]);
  nor g49 (n_180, A[21], B[21]);
  nand g50 (n_181, A[21], B[21]);
  nor g51 (n_190, A[22], B[22]);
  nand g52 (n_185, A[22], B[22]);
  nor g53 (n_186, A[23], B[23]);
  nand g54 (n_187, A[23], B[23]);
  nor g55 (n_196, A[24], B[24]);
  nand g56 (n_191, A[24], B[24]);
  nor g57 (n_192, A[25], B[25]);
  nand g58 (n_193, A[25], B[25]);
  nor g59 (n_202, A[26], B[26]);
  nand g60 (n_197, A[26], B[26]);
  nor g61 (n_198, A[27], B[27]);
  nand g62 (n_199, A[27], B[27]);
  nor g63 (n_208, A[28], B[28]);
  nand g64 (n_203, A[28], B[28]);
  nor g65 (n_204, A[29], B[29]);
  nand g66 (n_205, A[29], B[29]);
  nor g67 (n_214, A[30], B[30]);
  nand g68 (n_209, A[30], B[30]);
  nor g69 (n_210, A[31], B[31]);
  nand g70 (n_211, A[31], B[31]);
  nor g71 (n_220, A[32], B[32]);
  nand g72 (n_215, A[32], B[32]);
  nor g73 (n_216, A[33], B[33]);
  nand g74 (n_217, A[33], B[33]);
  nor g75 (n_226, A[34], B[34]);
  nand g76 (n_221, A[34], B[34]);
  nor g77 (n_222, A[35], B[35]);
  nand g78 (n_223, A[35], B[35]);
  nand g83 (n_227, n_123, n_124);
  nor g84 (n_128, n_125, n_126);
  nor g87 (n_230, n_130, n_126);
  nor g88 (n_134, n_131, n_132);
  nor g91 (n_236, n_136, n_132);
  nor g92 (n_140, n_137, n_138);
  nor g95 (n_238, n_142, n_138);
  nor g96 (n_146, n_143, n_144);
  nor g99 (n_246, n_148, n_144);
  nor g100 (n_152, n_149, n_150);
  nor g103 (n_248, n_154, n_150);
  nor g104 (n_158, n_155, n_156);
  nor g107 (n_256, n_160, n_156);
  nor g108 (n_164, n_161, n_162);
  nor g111 (n_258, n_166, n_162);
  nor g112 (n_170, n_167, n_168);
  nor g115 (n_266, n_172, n_168);
  nor g116 (n_176, n_173, n_174);
  nor g119 (n_268, n_178, n_174);
  nor g120 (n_182, n_179, n_180);
  nor g123 (n_276, n_184, n_180);
  nor g124 (n_188, n_185, n_186);
  nor g127 (n_278, n_190, n_186);
  nor g128 (n_194, n_191, n_192);
  nor g131 (n_286, n_196, n_192);
  nor g132 (n_200, n_197, n_198);
  nor g135 (n_288, n_202, n_198);
  nor g136 (n_206, n_203, n_204);
  nor g139 (n_296, n_208, n_204);
  nor g140 (n_212, n_209, n_210);
  nor g143 (n_298, n_214, n_210);
  nor g144 (n_218, n_215, n_216);
  nor g147 (n_306, n_220, n_216);
  nor g148 (n_224, n_221, n_222);
  nor g151 (n_308, n_226, n_222);
  nand g154 (n_502, n_125, n_229);
  nand g155 (n_232, n_230, n_227);
  nand g156 (n_313, n_231, n_232);
  nor g157 (n_234, n_142, n_233);
  nand g166 (n_321, n_236, n_238);
  nor g167 (n_244, n_154, n_243);
  nand g176 (n_328, n_246, n_248);
  nor g177 (n_254, n_166, n_253);
  nand g186 (n_336, n_256, n_258);
  nor g187 (n_264, n_178, n_263);
  nand g196 (n_343, n_266, n_268);
  nor g197 (n_274, n_190, n_273);
  nand g206 (n_351, n_276, n_278);
  nor g207 (n_284, n_202, n_283);
  nand g216 (n_358, n_286, n_288);
  nor g217 (n_294, n_214, n_293);
  nand g226 (n_366, n_296, n_298);
  nor g227 (n_304, n_226, n_303);
  nand g236 (n_375, n_306, n_308);
  nand g239 (n_506, n_131, n_315);
  nand g240 (n_316, n_236, n_313);
  nand g241 (n_508, n_233, n_316);
  nand g244 (n_511, n_319, n_320);
  nand g247 (n_376, n_323, n_324);
  nor g248 (n_326, n_160, n_325);
  nor g251 (n_386, n_160, n_328);
  nor g257 (n_334, n_332, n_325);
  nor g260 (n_392, n_328, n_332);
  nor g261 (n_338, n_336, n_325);
  nor g264 (n_395, n_328, n_336);
  nor g265 (n_341, n_184, n_340);
  nor g268 (n_444, n_184, n_343);
  nor g274 (n_349, n_347, n_340);
  nor g277 (n_450, n_343, n_347);
  nor g278 (n_353, n_351, n_340);
  nor g281 (n_401, n_343, n_351);
  nor g282 (n_356, n_208, n_355);
  nor g285 (n_414, n_208, n_358);
  nor g291 (n_364, n_362, n_355);
  nor g294 (n_424, n_358, n_362);
  nor g295 (n_368, n_366, n_355);
  nor g298 (n_429, n_358, n_366);
  nor g299 (n_373, n_370, n_371);
  nor g302 (n_496, n_370, n_375);
  nand g305 (n_515, n_143, n_378);
  nand g306 (n_379, n_246, n_376);
  nand g307 (n_517, n_243, n_379);
  nand g310 (n_520, n_382, n_383);
  nand g313 (n_523, n_325, n_385);
  nand g314 (n_388, n_386, n_376);
  nand g315 (n_526, n_387, n_388);
  nand g316 (n_391, n_389, n_376);
  nand g317 (n_528, n_390, n_391);
  nand g318 (n_394, n_392, n_376);
  nand g319 (n_531, n_393, n_394);
  nand g320 (n_397, n_395, n_376);
  nand g321 (n_434, n_396, n_397);
  nor g322 (n_399, n_196, n_398);
  nand g331 (n_458, n_286, n_401);
  nor g332 (n_408, n_406, n_398);
  nor g337 (n_411, n_358, n_398);
  nand g346 (n_470, n_401, n_414);
  nand g351 (n_474, n_401, n_419);
  nand g356 (n_478, n_401, n_424);
  nand g361 (n_482, n_401, n_429);
  nand g364 (n_535, n_167, n_436);
  nand g365 (n_437, n_266, n_434);
  nand g366 (n_537, n_263, n_437);
  nand g369 (n_540, n_440, n_441);
  nand g372 (n_543, n_340, n_443);
  nand g373 (n_446, n_444, n_434);
  nand g374 (n_546, n_445, n_446);
  nand g375 (n_449, n_447, n_434);
  nand g376 (n_548, n_448, n_449);
  nand g377 (n_452, n_450, n_434);
  nand g378 (n_551, n_451, n_452);
  nand g379 (n_453, n_401, n_434);
  nand g380 (n_553, n_398, n_453);
  nand g383 (n_556, n_456, n_457);
  nand g386 (n_558, n_460, n_461);
  nand g389 (n_561, n_464, n_465);
  nand g392 (n_564, n_468, n_469);
  nand g395 (n_567, n_472, n_473);
  nand g398 (n_569, n_476, n_477);
  nand g401 (n_572, n_480, n_481);
  nand g404 (n_486, n_484, n_485);
  nand g407 (n_576, n_215, n_488);
  nand g408 (n_489, n_306, n_486);
  nand g409 (n_578, n_303, n_489);
  nand g412 (n_581, n_492, n_493);
  nand g415 (n_584, n_371, n_495);
  nand g416 (n_498, n_496, n_486);
  nand g417 (n_116, n_497, n_498);
  xnor g421 (Z[2], n_227, n_500);
  xnor g424 (Z[3], n_502, n_503);
  xnor g426 (Z[4], n_313, n_504);
  xnor g429 (Z[5], n_506, n_507);
  xnor g431 (Z[6], n_508, n_509);
  xnor g434 (Z[7], n_511, n_512);
  xnor g436 (Z[8], n_376, n_513);
  xnor g439 (Z[9], n_515, n_516);
  xnor g441 (Z[10], n_517, n_518);
  xnor g444 (Z[11], n_520, n_521);
  xnor g447 (Z[12], n_523, n_524);
  xnor g450 (Z[13], n_526, n_527);
  xnor g452 (Z[14], n_528, n_529);
  xnor g455 (Z[15], n_531, n_532);
  xnor g457 (Z[16], n_434, n_533);
  xnor g460 (Z[17], n_535, n_536);
  xnor g462 (Z[18], n_537, n_538);
  xnor g465 (Z[19], n_540, n_541);
  xnor g468 (Z[20], n_543, n_544);
  xnor g471 (Z[21], n_546, n_547);
  xnor g473 (Z[22], n_548, n_549);
  xnor g476 (Z[23], n_551, n_552);
  xnor g478 (Z[24], n_553, n_554);
  xnor g481 (Z[25], n_556, n_557);
  xnor g483 (Z[26], n_558, n_559);
  xnor g486 (Z[27], n_561, n_562);
  xnor g489 (Z[28], n_564, n_565);
  xnor g492 (Z[29], n_567, n_568);
  xnor g494 (Z[30], n_569, n_570);
  xnor g497 (Z[31], n_572, n_573);
  xnor g499 (Z[32], n_486, n_574);
  xnor g502 (Z[33], n_576, n_577);
  xnor g504 (Z[34], n_578, n_579);
  xnor g507 (Z[35], n_581, n_582);
  xnor g510 (Z[36], n_584, n_585);
  and g513 (n_370, A[36], B[36]);
  or g514 (n_372, A[36], B[36]);
  and g515 (n_303, wc, n_217);
  not gc (wc, n_218);
  and g516 (n_310, wc0, n_223);
  not gc0 (wc0, n_224);
  and g517 (n_263, wc1, n_169);
  not gc1 (wc1, n_170);
  and g518 (n_270, wc2, n_175);
  not gc2 (wc2, n_176);
  and g519 (n_273, wc3, n_181);
  not gc3 (wc3, n_182);
  and g520 (n_280, wc4, n_187);
  not gc4 (wc4, n_188);
  and g521 (n_283, wc5, n_193);
  not gc5 (wc5, n_194);
  and g522 (n_290, wc6, n_199);
  not gc6 (wc6, n_200);
  and g523 (n_293, wc7, n_205);
  not gc7 (wc7, n_206);
  and g524 (n_300, wc8, n_211);
  not gc8 (wc8, n_212);
  and g525 (n_243, wc9, n_145);
  not gc9 (wc9, n_146);
  and g526 (n_250, wc10, n_151);
  not gc10 (wc10, n_152);
  and g527 (n_253, wc11, n_157);
  not gc11 (wc11, n_158);
  and g528 (n_260, wc12, n_163);
  not gc12 (wc12, n_164);
  and g529 (n_233, wc13, n_133);
  not gc13 (wc13, n_134);
  and g530 (n_240, wc14, n_139);
  not gc14 (wc14, n_140);
  and g531 (n_231, wc15, n_127);
  not gc15 (wc15, n_128);
  or g532 (n_124, n_117, n_120);
  or g533 (n_317, wc16, n_142);
  not gc16 (wc16, n_236);
  or g534 (n_380, wc17, n_154);
  not gc17 (wc17, n_246);
  or g535 (n_332, wc18, n_166);
  not gc18 (wc18, n_256);
  or g536 (n_438, wc19, n_178);
  not gc19 (wc19, n_266);
  or g537 (n_347, wc20, n_190);
  not gc20 (wc20, n_276);
  or g538 (n_406, wc21, n_202);
  not gc21 (wc21, n_286);
  or g539 (n_362, wc22, n_214);
  not gc22 (wc22, n_296);
  or g540 (n_490, wc23, n_226);
  not gc23 (wc23, n_306);
  or g541 (n_499, wc24, n_120);
  not gc24 (wc24, n_123);
  or g542 (n_500, wc25, n_130);
  not gc25 (wc25, n_125);
  or g543 (n_503, wc26, n_126);
  not gc26 (wc26, n_127);
  or g544 (n_504, wc27, n_136);
  not gc27 (wc27, n_131);
  or g545 (n_507, wc28, n_132);
  not gc28 (wc28, n_133);
  or g546 (n_509, wc29, n_142);
  not gc29 (wc29, n_137);
  or g547 (n_512, wc30, n_138);
  not gc30 (wc30, n_139);
  or g548 (n_513, wc31, n_148);
  not gc31 (wc31, n_143);
  or g549 (n_516, wc32, n_144);
  not gc32 (wc32, n_145);
  or g550 (n_518, wc33, n_154);
  not gc33 (wc33, n_149);
  or g551 (n_521, wc34, n_150);
  not gc34 (wc34, n_151);
  or g552 (n_524, wc35, n_160);
  not gc35 (wc35, n_155);
  or g553 (n_527, wc36, n_156);
  not gc36 (wc36, n_157);
  or g554 (n_529, wc37, n_166);
  not gc37 (wc37, n_161);
  or g555 (n_532, wc38, n_162);
  not gc38 (wc38, n_163);
  or g556 (n_533, wc39, n_172);
  not gc39 (wc39, n_167);
  or g557 (n_536, wc40, n_168);
  not gc40 (wc40, n_169);
  or g558 (n_538, wc41, n_178);
  not gc41 (wc41, n_173);
  or g559 (n_541, wc42, n_174);
  not gc42 (wc42, n_175);
  or g560 (n_544, wc43, n_184);
  not gc43 (wc43, n_179);
  or g561 (n_547, wc44, n_180);
  not gc44 (wc44, n_181);
  or g562 (n_549, wc45, n_190);
  not gc45 (wc45, n_185);
  or g563 (n_552, wc46, n_186);
  not gc46 (wc46, n_187);
  or g564 (n_554, wc47, n_196);
  not gc47 (wc47, n_191);
  or g565 (n_557, wc48, n_192);
  not gc48 (wc48, n_193);
  or g566 (n_559, wc49, n_202);
  not gc49 (wc49, n_197);
  or g567 (n_562, wc50, n_198);
  not gc50 (wc50, n_199);
  or g568 (n_565, wc51, n_208);
  not gc51 (wc51, n_203);
  or g569 (n_568, wc52, n_204);
  not gc52 (wc52, n_205);
  or g570 (n_570, wc53, n_214);
  not gc53 (wc53, n_209);
  or g571 (n_573, wc54, n_210);
  not gc54 (wc54, n_211);
  or g572 (n_574, wc55, n_220);
  not gc55 (wc55, n_215);
  or g573 (n_577, wc56, n_216);
  not gc56 (wc56, n_217);
  or g574 (n_579, wc57, n_226);
  not gc57 (wc57, n_221);
  or g575 (n_582, wc58, n_222);
  not gc58 (wc58, n_223);
  and g576 (n_311, wc59, n_308);
  not gc59 (wc59, n_303);
  and g577 (n_271, wc60, n_268);
  not gc60 (wc60, n_263);
  and g578 (n_281, wc61, n_278);
  not gc61 (wc61, n_273);
  and g579 (n_291, wc62, n_288);
  not gc62 (wc62, n_283);
  and g580 (n_301, wc63, n_298);
  not gc63 (wc63, n_293);
  and g581 (n_251, wc64, n_248);
  not gc64 (wc64, n_243);
  and g582 (n_261, wc65, n_258);
  not gc65 (wc65, n_253);
  and g583 (n_241, wc66, n_238);
  not gc66 (wc66, n_233);
  and g584 (n_389, wc67, n_256);
  not gc67 (wc67, n_328);
  and g585 (n_447, wc68, n_276);
  not gc68 (wc68, n_343);
  and g586 (n_419, wc69, n_296);
  not gc69 (wc69, n_358);
  xor g587 (Z[1], n_117, n_499);
  or g588 (n_585, wc70, n_370);
  not gc70 (wc70, n_372);
  and g589 (n_371, wc71, n_310);
  not gc71 (wc71, n_311);
  and g590 (n_340, wc72, n_270);
  not gc72 (wc72, n_271);
  and g591 (n_352, wc73, n_280);
  not gc73 (wc73, n_281);
  and g592 (n_355, wc74, n_290);
  not gc74 (wc74, n_291);
  and g593 (n_367, wc75, n_300);
  not gc75 (wc75, n_301);
  and g594 (n_325, wc76, n_250);
  not gc76 (wc76, n_251);
  and g595 (n_337, wc77, n_260);
  not gc77 (wc77, n_261);
  and g596 (n_323, wc78, n_240);
  not gc78 (wc78, n_241);
  or g597 (n_229, wc79, n_130);
  not gc79 (wc79, n_227);
  and g598 (n_319, wc80, n_137);
  not gc80 (wc80, n_234);
  and g599 (n_382, wc81, n_149);
  not gc81 (wc81, n_244);
  and g600 (n_333, wc82, n_161);
  not gc82 (wc82, n_254);
  and g601 (n_440, wc83, n_173);
  not gc83 (wc83, n_264);
  and g602 (n_348, wc84, n_185);
  not gc84 (wc84, n_274);
  and g603 (n_407, wc85, n_197);
  not gc85 (wc85, n_284);
  and g604 (n_363, wc86, n_209);
  not gc86 (wc86, n_294);
  and g605 (n_492, wc87, n_221);
  not gc87 (wc87, n_304);
  or g606 (n_454, wc88, n_196);
  not gc88 (wc88, n_401);
  or g607 (n_462, n_406, wc89);
  not gc89 (wc89, n_401);
  or g608 (n_466, wc90, n_358);
  not gc90 (wc90, n_401);
  and g609 (n_330, wc91, n_256);
  not gc91 (wc91, n_325);
  and g610 (n_345, wc92, n_276);
  not gc92 (wc92, n_340);
  and g611 (n_360, wc93, n_296);
  not gc93 (wc93, n_355);
  and g612 (n_497, n_372, wc94);
  not gc94 (wc94, n_373);
  and g613 (n_398, n_352, wc95);
  not gc95 (wc95, n_353);
  and g614 (n_431, n_367, wc96);
  not gc96 (wc96, n_368);
  and g615 (n_396, n_337, wc97);
  not gc97 (wc97, n_338);
  or g616 (n_324, n_321, wc98);
  not gc98 (wc98, n_313);
  or g617 (n_315, wc99, n_136);
  not gc99 (wc99, n_313);
  or g618 (n_320, n_317, wc100);
  not gc100 (wc100, n_313);
  and g619 (n_387, wc101, n_155);
  not gc101 (wc101, n_326);
  and g620 (n_390, wc102, n_253);
  not gc102 (wc102, n_330);
  and g621 (n_393, n_333, wc103);
  not gc103 (wc103, n_334);
  and g622 (n_445, wc104, n_179);
  not gc104 (wc104, n_341);
  and g623 (n_448, wc105, n_273);
  not gc105 (wc105, n_345);
  and g624 (n_451, n_348, wc106);
  not gc106 (wc106, n_349);
  and g625 (n_416, wc107, n_203);
  not gc107 (wc107, n_356);
  and g626 (n_421, wc108, n_293);
  not gc108 (wc108, n_360);
  and g627 (n_426, n_363, wc109);
  not gc109 (wc109, n_364);
  and g628 (n_432, wc110, n_429);
  not gc110 (wc110, n_398);
  and g629 (n_404, wc111, n_286);
  not gc111 (wc111, n_398);
  and g630 (n_417, wc112, n_414);
  not gc112 (wc112, n_398);
  and g631 (n_422, wc113, n_419);
  not gc113 (wc113, n_398);
  and g632 (n_427, wc114, n_424);
  not gc114 (wc114, n_398);
  and g633 (n_484, wc115, n_431);
  not gc115 (wc115, n_432);
  or g634 (n_378, wc116, n_148);
  not gc116 (wc116, n_376);
  or g635 (n_383, n_380, wc117);
  not gc117 (wc117, n_376);
  or g636 (n_385, wc118, n_328);
  not gc118 (wc118, n_376);
  and g637 (n_456, wc119, n_191);
  not gc119 (wc119, n_399);
  and g638 (n_460, wc120, n_283);
  not gc120 (wc120, n_404);
  and g639 (n_464, n_407, wc121);
  not gc121 (wc121, n_408);
  and g640 (n_468, n_355, wc122);
  not gc122 (wc122, n_411);
  and g641 (n_472, wc123, n_416);
  not gc123 (wc123, n_417);
  and g642 (n_476, wc124, n_421);
  not gc124 (wc124, n_422);
  and g643 (n_480, wc125, n_426);
  not gc125 (wc125, n_427);
  or g644 (n_485, n_482, wc126);
  not gc126 (wc126, n_434);
  or g645 (n_436, wc127, n_172);
  not gc127 (wc127, n_434);
  or g646 (n_441, n_438, wc128);
  not gc128 (wc128, n_434);
  or g647 (n_443, wc129, n_343);
  not gc129 (wc129, n_434);
  or g648 (n_457, n_454, wc130);
  not gc130 (wc130, n_434);
  or g649 (n_461, n_458, wc131);
  not gc131 (wc131, n_434);
  or g650 (n_465, n_462, wc132);
  not gc132 (wc132, n_434);
  or g651 (n_469, n_466, wc133);
  not gc133 (wc133, n_434);
  or g652 (n_473, n_470, wc134);
  not gc134 (wc134, n_434);
  or g653 (n_477, n_474, wc135);
  not gc135 (wc135, n_434);
  or g654 (n_481, n_478, wc136);
  not gc136 (wc136, n_434);
  or g655 (n_488, wc137, n_220);
  not gc137 (wc137, n_486);
  or g656 (n_493, n_490, wc138);
  not gc138 (wc138, n_486);
  or g657 (n_495, wc139, n_375);
  not gc139 (wc139, n_486);
endmodule

module add_signed_508_GENERIC(A, B, Z);
  input [36:0] A, B;
  output [37:0] Z;
  wire [36:0] A, B;
  wire [37:0] Z;
  add_signed_508_GENERIC_REAL g1(.A ({A[35], A[35:0]}), .B ({B[35],
       B[35:0]}), .Z (Z));
endmodule

module add_signed_522_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [35:0] A, B;
  output [36:0] Z;
  wire [35:0] A, B;
  wire [36:0] Z;
  wire n_113, n_114, n_117, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_127, n_128, n_129, n_130, n_131, n_133, n_134;
  wire n_135, n_136, n_137, n_139, n_140, n_141, n_142, n_143;
  wire n_145, n_146, n_147, n_148, n_149, n_151, n_152, n_153;
  wire n_154, n_155, n_157, n_158, n_159, n_160, n_161, n_163;
  wire n_164, n_165, n_166, n_167, n_169, n_170, n_171, n_172;
  wire n_173, n_175, n_176, n_177, n_178, n_179, n_181, n_182;
  wire n_183, n_184, n_185, n_187, n_188, n_189, n_190, n_191;
  wire n_193, n_194, n_195, n_196, n_197, n_199, n_200, n_201;
  wire n_202, n_203, n_205, n_206, n_207, n_208, n_209, n_211;
  wire n_212, n_213, n_214, n_215, n_217, n_218, n_219, n_220;
  wire n_221, n_223, n_224, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_233, n_235, n_237, n_238, n_240, n_241, n_243;
  wire n_245, n_247, n_248, n_250, n_251, n_253, n_255, n_257;
  wire n_258, n_260, n_261, n_263, n_265, n_267, n_268, n_270;
  wire n_271, n_273, n_275, n_277, n_278, n_280, n_281, n_283;
  wire n_285, n_287, n_288, n_290, n_291, n_293, n_295, n_297;
  wire n_298, n_300, n_301, n_303, n_305, n_307, n_308, n_310;
  wire n_312, n_313, n_314, n_316, n_317, n_318, n_320, n_321;
  wire n_322, n_323, n_325, n_327, n_329, n_330, n_331, n_333;
  wire n_334, n_335, n_337, n_338, n_340, n_342, n_344, n_345;
  wire n_346, n_348, n_349, n_350, n_352, n_353, n_355, n_357;
  wire n_359, n_360, n_361, n_363, n_364, n_365, n_367, n_369;
  wire n_370, n_371, n_373, n_374, n_376, n_377, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_390, n_392, n_395, n_397, n_398, n_399;
  wire n_402, n_405, n_407, n_408, n_410, n_412, n_413, n_415;
  wire n_417, n_418, n_420, n_422, n_423, n_425, n_427, n_428;
  wire n_429, n_431, n_432, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_447;
  wire n_448, n_449, n_451, n_452, n_453, n_455, n_456, n_457;
  wire n_459, n_460, n_461, n_463, n_464, n_465, n_467, n_468;
  wire n_469, n_471, n_472, n_473, n_475, n_476, n_477, n_479;
  wire n_480, n_481, n_483, n_484, n_485, n_487, n_488, n_489;
  wire n_490, n_492, n_493, n_494, n_496, n_497, n_498, n_499;
  wire n_501, n_502, n_503, n_505, n_506, n_507, n_508, n_510;
  wire n_511, n_513, n_514, n_516, n_517, n_518, n_519, n_521;
  wire n_522, n_523, n_525, n_526, n_527, n_528, n_530, n_531;
  wire n_533, n_534, n_536, n_537, n_538, n_539, n_541, n_542;
  wire n_543, n_544, n_546, n_547, n_548, n_549, n_551, n_552;
  wire n_554, n_555, n_557, n_558, n_559, n_560, n_562, n_563;
  wire n_564, n_566, n_567, n_568, n_569, n_571, n_572;
  not g3 (Z[36], n_113);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_114, A[0], B[0]);
  nor g9 (n_117, A[1], B[1]);
  nand g10 (n_120, A[1], B[1]);
  nor g11 (n_127, A[2], B[2]);
  nand g12 (n_122, A[2], B[2]);
  nor g13 (n_123, A[3], B[3]);
  nand g14 (n_124, A[3], B[3]);
  nor g15 (n_133, A[4], B[4]);
  nand g16 (n_128, A[4], B[4]);
  nor g17 (n_129, A[5], B[5]);
  nand g18 (n_130, A[5], B[5]);
  nor g19 (n_139, A[6], B[6]);
  nand g20 (n_134, A[6], B[6]);
  nor g21 (n_135, A[7], B[7]);
  nand g22 (n_136, A[7], B[7]);
  nor g23 (n_145, A[8], B[8]);
  nand g24 (n_140, A[8], B[8]);
  nor g25 (n_141, A[9], B[9]);
  nand g26 (n_142, A[9], B[9]);
  nor g27 (n_151, A[10], B[10]);
  nand g28 (n_146, A[10], B[10]);
  nor g29 (n_147, A[11], B[11]);
  nand g30 (n_148, A[11], B[11]);
  nor g31 (n_157, A[12], B[12]);
  nand g32 (n_152, A[12], B[12]);
  nor g33 (n_153, A[13], B[13]);
  nand g34 (n_154, A[13], B[13]);
  nor g35 (n_163, A[14], B[14]);
  nand g36 (n_158, A[14], B[14]);
  nor g37 (n_159, A[15], B[15]);
  nand g38 (n_160, A[15], B[15]);
  nor g39 (n_169, A[16], B[16]);
  nand g40 (n_164, A[16], B[16]);
  nor g41 (n_165, A[17], B[17]);
  nand g42 (n_166, A[17], B[17]);
  nor g43 (n_175, A[18], B[18]);
  nand g44 (n_170, A[18], B[18]);
  nor g45 (n_171, A[19], B[19]);
  nand g46 (n_172, A[19], B[19]);
  nor g47 (n_181, A[20], B[20]);
  nand g48 (n_176, A[20], B[20]);
  nor g49 (n_177, A[21], B[21]);
  nand g50 (n_178, A[21], B[21]);
  nor g51 (n_187, A[22], B[22]);
  nand g52 (n_182, A[22], B[22]);
  nor g53 (n_183, A[23], B[23]);
  nand g54 (n_184, A[23], B[23]);
  nor g55 (n_193, A[24], B[24]);
  nand g56 (n_188, A[24], B[24]);
  nor g57 (n_189, A[25], B[25]);
  nand g58 (n_190, A[25], B[25]);
  nor g59 (n_199, A[26], B[26]);
  nand g60 (n_194, A[26], B[26]);
  nor g61 (n_195, A[27], B[27]);
  nand g62 (n_196, A[27], B[27]);
  nor g63 (n_205, A[28], B[28]);
  nand g64 (n_200, A[28], B[28]);
  nor g65 (n_201, A[29], B[29]);
  nand g66 (n_202, A[29], B[29]);
  nor g67 (n_211, A[30], B[30]);
  nand g68 (n_206, A[30], B[30]);
  nor g69 (n_207, A[31], B[31]);
  nand g70 (n_208, A[31], B[31]);
  nor g71 (n_217, A[32], B[32]);
  nand g72 (n_212, A[32], B[32]);
  nor g73 (n_213, A[33], B[33]);
  nand g74 (n_214, A[33], B[33]);
  nor g75 (n_223, A[34], B[34]);
  nand g76 (n_218, A[34], B[34]);
  nand g81 (n_224, n_120, n_121);
  nor g82 (n_125, n_122, n_123);
  nor g85 (n_227, n_127, n_123);
  nor g86 (n_131, n_128, n_129);
  nor g89 (n_233, n_133, n_129);
  nor g90 (n_137, n_134, n_135);
  nor g93 (n_235, n_139, n_135);
  nor g94 (n_143, n_140, n_141);
  nor g97 (n_243, n_145, n_141);
  nor g98 (n_149, n_146, n_147);
  nor g101 (n_245, n_151, n_147);
  nor g102 (n_155, n_152, n_153);
  nor g105 (n_253, n_157, n_153);
  nor g106 (n_161, n_158, n_159);
  nor g109 (n_255, n_163, n_159);
  nor g110 (n_167, n_164, n_165);
  nor g113 (n_263, n_169, n_165);
  nor g114 (n_173, n_170, n_171);
  nor g117 (n_265, n_175, n_171);
  nor g118 (n_179, n_176, n_177);
  nor g121 (n_273, n_181, n_177);
  nor g122 (n_185, n_182, n_183);
  nor g125 (n_275, n_187, n_183);
  nor g126 (n_191, n_188, n_189);
  nor g129 (n_283, n_193, n_189);
  nor g130 (n_197, n_194, n_195);
  nor g133 (n_285, n_199, n_195);
  nor g134 (n_203, n_200, n_201);
  nor g137 (n_293, n_205, n_201);
  nor g138 (n_209, n_206, n_207);
  nor g141 (n_295, n_211, n_207);
  nor g142 (n_215, n_212, n_213);
  nor g145 (n_303, n_217, n_213);
  nor g146 (n_221, n_218, n_219);
  nor g149 (n_305, n_223, n_219);
  nand g152 (n_492, n_122, n_226);
  nand g153 (n_229, n_227, n_224);
  nand g154 (n_310, n_228, n_229);
  nor g155 (n_231, n_139, n_230);
  nand g164 (n_318, n_233, n_235);
  nor g165 (n_241, n_151, n_240);
  nand g174 (n_325, n_243, n_245);
  nor g175 (n_251, n_163, n_250);
  nand g184 (n_333, n_253, n_255);
  nor g185 (n_261, n_175, n_260);
  nand g194 (n_340, n_263, n_265);
  nor g195 (n_271, n_187, n_270);
  nand g204 (n_348, n_273, n_275);
  nor g205 (n_281, n_199, n_280);
  nand g214 (n_355, n_283, n_285);
  nor g215 (n_291, n_211, n_290);
  nand g224 (n_363, n_293, n_295);
  nor g225 (n_301, n_223, n_300);
  nand g234 (n_485, n_303, n_305);
  nand g237 (n_496, n_128, n_312);
  nand g238 (n_313, n_233, n_310);
  nand g239 (n_498, n_230, n_313);
  nand g242 (n_501, n_316, n_317);
  nand g245 (n_367, n_320, n_321);
  nor g246 (n_323, n_157, n_322);
  nor g249 (n_377, n_157, n_325);
  nor g255 (n_331, n_329, n_322);
  nor g258 (n_383, n_325, n_329);
  nor g259 (n_335, n_333, n_322);
  nor g262 (n_386, n_325, n_333);
  nor g263 (n_338, n_181, n_337);
  nor g266 (n_435, n_181, n_340);
  nor g272 (n_346, n_344, n_337);
  nor g275 (n_441, n_340, n_344);
  nor g276 (n_350, n_348, n_337);
  nor g279 (n_392, n_340, n_348);
  nor g280 (n_353, n_205, n_352);
  nor g283 (n_405, n_205, n_355);
  nor g289 (n_361, n_359, n_352);
  nor g292 (n_415, n_355, n_359);
  nor g293 (n_365, n_363, n_352);
  nor g296 (n_420, n_355, n_363);
  nand g299 (n_505, n_140, n_369);
  nand g300 (n_370, n_243, n_367);
  nand g301 (n_507, n_240, n_370);
  nand g304 (n_510, n_373, n_374);
  nand g307 (n_513, n_322, n_376);
  nand g308 (n_379, n_377, n_367);
  nand g309 (n_516, n_378, n_379);
  nand g310 (n_382, n_380, n_367);
  nand g311 (n_518, n_381, n_382);
  nand g312 (n_385, n_383, n_367);
  nand g313 (n_521, n_384, n_385);
  nand g314 (n_388, n_386, n_367);
  nand g315 (n_425, n_387, n_388);
  nor g316 (n_390, n_193, n_389);
  nand g325 (n_449, n_283, n_392);
  nor g326 (n_399, n_397, n_389);
  nor g331 (n_402, n_355, n_389);
  nand g340 (n_461, n_392, n_405);
  nand g345 (n_465, n_392, n_410);
  nand g350 (n_469, n_392, n_415);
  nand g355 (n_473, n_392, n_420);
  nand g358 (n_525, n_164, n_427);
  nand g359 (n_428, n_263, n_425);
  nand g360 (n_527, n_260, n_428);
  nand g363 (n_530, n_431, n_432);
  nand g366 (n_533, n_337, n_434);
  nand g367 (n_437, n_435, n_425);
  nand g368 (n_536, n_436, n_437);
  nand g369 (n_440, n_438, n_425);
  nand g370 (n_538, n_439, n_440);
  nand g371 (n_443, n_441, n_425);
  nand g372 (n_541, n_442, n_443);
  nand g373 (n_444, n_392, n_425);
  nand g374 (n_543, n_389, n_444);
  nand g377 (n_546, n_447, n_448);
  nand g380 (n_548, n_451, n_452);
  nand g383 (n_551, n_455, n_456);
  nand g386 (n_554, n_459, n_460);
  nand g389 (n_557, n_463, n_464);
  nand g392 (n_559, n_467, n_468);
  nand g395 (n_562, n_471, n_472);
  nand g398 (n_477, n_475, n_476);
  nand g401 (n_566, n_212, n_479);
  nand g402 (n_480, n_303, n_477);
  nand g403 (n_568, n_300, n_480);
  nand g406 (n_571, n_483, n_484);
  nand g409 (n_113, n_487, n_488);
  xnor g413 (Z[2], n_224, n_490);
  xnor g416 (Z[3], n_492, n_493);
  xnor g418 (Z[4], n_310, n_494);
  xnor g421 (Z[5], n_496, n_497);
  xnor g423 (Z[6], n_498, n_499);
  xnor g426 (Z[7], n_501, n_502);
  xnor g428 (Z[8], n_367, n_503);
  xnor g431 (Z[9], n_505, n_506);
  xnor g433 (Z[10], n_507, n_508);
  xnor g436 (Z[11], n_510, n_511);
  xnor g439 (Z[12], n_513, n_514);
  xnor g442 (Z[13], n_516, n_517);
  xnor g444 (Z[14], n_518, n_519);
  xnor g447 (Z[15], n_521, n_522);
  xnor g449 (Z[16], n_425, n_523);
  xnor g452 (Z[17], n_525, n_526);
  xnor g454 (Z[18], n_527, n_528);
  xnor g457 (Z[19], n_530, n_531);
  xnor g460 (Z[20], n_533, n_534);
  xnor g463 (Z[21], n_536, n_537);
  xnor g465 (Z[22], n_538, n_539);
  xnor g468 (Z[23], n_541, n_542);
  xnor g470 (Z[24], n_543, n_544);
  xnor g473 (Z[25], n_546, n_547);
  xnor g475 (Z[26], n_548, n_549);
  xnor g478 (Z[27], n_551, n_552);
  xnor g481 (Z[28], n_554, n_555);
  xnor g484 (Z[29], n_557, n_558);
  xnor g486 (Z[30], n_559, n_560);
  xnor g489 (Z[31], n_562, n_563);
  xnor g491 (Z[32], n_477, n_564);
  xnor g494 (Z[33], n_566, n_567);
  xnor g496 (Z[34], n_568, n_569);
  xnor g499 (Z[35], n_571, n_572);
  and g502 (n_219, A[35], B[35]);
  or g503 (n_220, A[35], B[35]);
  and g504 (n_300, wc, n_214);
  not gc (wc, n_215);
  and g505 (n_260, wc0, n_166);
  not gc0 (wc0, n_167);
  and g506 (n_267, wc1, n_172);
  not gc1 (wc1, n_173);
  and g507 (n_270, wc2, n_178);
  not gc2 (wc2, n_179);
  and g508 (n_277, wc3, n_184);
  not gc3 (wc3, n_185);
  and g509 (n_280, wc4, n_190);
  not gc4 (wc4, n_191);
  and g510 (n_287, wc5, n_196);
  not gc5 (wc5, n_197);
  and g511 (n_290, wc6, n_202);
  not gc6 (wc6, n_203);
  and g512 (n_297, wc7, n_208);
  not gc7 (wc7, n_209);
  and g513 (n_240, wc8, n_142);
  not gc8 (wc8, n_143);
  and g514 (n_247, wc9, n_148);
  not gc9 (wc9, n_149);
  and g515 (n_250, wc10, n_154);
  not gc10 (wc10, n_155);
  and g516 (n_257, wc11, n_160);
  not gc11 (wc11, n_161);
  and g517 (n_230, wc12, n_130);
  not gc12 (wc12, n_131);
  and g518 (n_237, wc13, n_136);
  not gc13 (wc13, n_137);
  and g519 (n_228, wc14, n_124);
  not gc14 (wc14, n_125);
  or g520 (n_121, n_114, n_117);
  or g521 (n_314, wc15, n_139);
  not gc15 (wc15, n_233);
  or g522 (n_371, wc16, n_151);
  not gc16 (wc16, n_243);
  or g523 (n_329, wc17, n_163);
  not gc17 (wc17, n_253);
  or g524 (n_429, wc18, n_175);
  not gc18 (wc18, n_263);
  or g525 (n_344, wc19, n_187);
  not gc19 (wc19, n_273);
  or g526 (n_397, wc20, n_199);
  not gc20 (wc20, n_283);
  or g527 (n_359, wc21, n_211);
  not gc21 (wc21, n_293);
  or g528 (n_481, wc22, n_223);
  not gc22 (wc22, n_303);
  or g529 (n_489, wc23, n_117);
  not gc23 (wc23, n_120);
  or g530 (n_490, wc24, n_127);
  not gc24 (wc24, n_122);
  or g531 (n_493, wc25, n_123);
  not gc25 (wc25, n_124);
  or g532 (n_494, wc26, n_133);
  not gc26 (wc26, n_128);
  or g533 (n_497, wc27, n_129);
  not gc27 (wc27, n_130);
  or g534 (n_499, wc28, n_139);
  not gc28 (wc28, n_134);
  or g535 (n_502, wc29, n_135);
  not gc29 (wc29, n_136);
  or g536 (n_503, wc30, n_145);
  not gc30 (wc30, n_140);
  or g537 (n_506, wc31, n_141);
  not gc31 (wc31, n_142);
  or g538 (n_508, wc32, n_151);
  not gc32 (wc32, n_146);
  or g539 (n_511, wc33, n_147);
  not gc33 (wc33, n_148);
  or g540 (n_514, wc34, n_157);
  not gc34 (wc34, n_152);
  or g541 (n_517, wc35, n_153);
  not gc35 (wc35, n_154);
  or g542 (n_519, wc36, n_163);
  not gc36 (wc36, n_158);
  or g543 (n_522, wc37, n_159);
  not gc37 (wc37, n_160);
  or g544 (n_523, wc38, n_169);
  not gc38 (wc38, n_164);
  or g545 (n_526, wc39, n_165);
  not gc39 (wc39, n_166);
  or g546 (n_528, wc40, n_175);
  not gc40 (wc40, n_170);
  or g547 (n_531, wc41, n_171);
  not gc41 (wc41, n_172);
  or g548 (n_534, wc42, n_181);
  not gc42 (wc42, n_176);
  or g549 (n_537, wc43, n_177);
  not gc43 (wc43, n_178);
  or g550 (n_539, wc44, n_187);
  not gc44 (wc44, n_182);
  or g551 (n_542, wc45, n_183);
  not gc45 (wc45, n_184);
  or g552 (n_544, wc46, n_193);
  not gc46 (wc46, n_188);
  or g553 (n_547, wc47, n_189);
  not gc47 (wc47, n_190);
  or g554 (n_549, wc48, n_199);
  not gc48 (wc48, n_194);
  or g555 (n_552, wc49, n_195);
  not gc49 (wc49, n_196);
  or g556 (n_555, wc50, n_205);
  not gc50 (wc50, n_200);
  or g557 (n_558, wc51, n_201);
  not gc51 (wc51, n_202);
  or g558 (n_560, wc52, n_211);
  not gc52 (wc52, n_206);
  or g559 (n_563, wc53, n_207);
  not gc53 (wc53, n_208);
  or g560 (n_564, wc54, n_217);
  not gc54 (wc54, n_212);
  or g561 (n_567, wc55, n_213);
  not gc55 (wc55, n_214);
  or g562 (n_569, wc56, n_223);
  not gc56 (wc56, n_218);
  and g563 (n_307, n_220, wc57);
  not gc57 (wc57, n_221);
  and g564 (n_268, wc58, n_265);
  not gc58 (wc58, n_260);
  and g565 (n_278, wc59, n_275);
  not gc59 (wc59, n_270);
  and g566 (n_288, wc60, n_285);
  not gc60 (wc60, n_280);
  and g567 (n_298, wc61, n_295);
  not gc61 (wc61, n_290);
  and g568 (n_248, wc62, n_245);
  not gc62 (wc62, n_240);
  and g569 (n_258, wc63, n_255);
  not gc63 (wc63, n_250);
  and g570 (n_238, wc64, n_235);
  not gc64 (wc64, n_230);
  and g571 (n_380, wc65, n_253);
  not gc65 (wc65, n_325);
  and g572 (n_438, wc66, n_273);
  not gc66 (wc66, n_340);
  and g573 (n_410, wc67, n_293);
  not gc67 (wc67, n_355);
  xor g574 (Z[1], n_114, n_489);
  or g575 (n_572, wc68, n_219);
  not gc68 (wc68, n_220);
  and g576 (n_308, wc69, n_305);
  not gc69 (wc69, n_300);
  and g577 (n_337, wc70, n_267);
  not gc70 (wc70, n_268);
  and g578 (n_349, wc71, n_277);
  not gc71 (wc71, n_278);
  and g579 (n_352, wc72, n_287);
  not gc72 (wc72, n_288);
  and g580 (n_364, wc73, n_297);
  not gc73 (wc73, n_298);
  and g581 (n_322, wc74, n_247);
  not gc74 (wc74, n_248);
  and g582 (n_334, wc75, n_257);
  not gc75 (wc75, n_258);
  and g583 (n_320, wc76, n_237);
  not gc76 (wc76, n_238);
  or g584 (n_226, wc77, n_127);
  not gc77 (wc77, n_224);
  and g585 (n_316, wc78, n_134);
  not gc78 (wc78, n_231);
  and g586 (n_373, wc79, n_146);
  not gc79 (wc79, n_241);
  and g587 (n_330, wc80, n_158);
  not gc80 (wc80, n_251);
  and g588 (n_431, wc81, n_170);
  not gc81 (wc81, n_261);
  and g589 (n_345, wc82, n_182);
  not gc82 (wc82, n_271);
  and g590 (n_398, wc83, n_194);
  not gc83 (wc83, n_281);
  and g591 (n_360, wc84, n_206);
  not gc84 (wc84, n_291);
  and g592 (n_483, wc85, n_218);
  not gc85 (wc85, n_301);
  or g593 (n_445, wc86, n_193);
  not gc86 (wc86, n_392);
  or g594 (n_453, n_397, wc87);
  not gc87 (wc87, n_392);
  or g595 (n_457, wc88, n_355);
  not gc88 (wc88, n_392);
  and g596 (n_487, wc89, n_307);
  not gc89 (wc89, n_308);
  and g597 (n_327, wc90, n_253);
  not gc90 (wc90, n_322);
  and g598 (n_342, wc91, n_273);
  not gc91 (wc91, n_337);
  and g599 (n_357, wc92, n_293);
  not gc92 (wc92, n_352);
  and g600 (n_389, n_349, wc93);
  not gc93 (wc93, n_350);
  and g601 (n_422, n_364, wc94);
  not gc94 (wc94, n_365);
  and g602 (n_387, n_334, wc95);
  not gc95 (wc95, n_335);
  or g603 (n_321, n_318, wc96);
  not gc96 (wc96, n_310);
  or g604 (n_312, wc97, n_133);
  not gc97 (wc97, n_310);
  or g605 (n_317, n_314, wc98);
  not gc98 (wc98, n_310);
  and g606 (n_378, wc99, n_152);
  not gc99 (wc99, n_323);
  and g607 (n_381, wc100, n_250);
  not gc100 (wc100, n_327);
  and g608 (n_384, n_330, wc101);
  not gc101 (wc101, n_331);
  and g609 (n_436, wc102, n_176);
  not gc102 (wc102, n_338);
  and g610 (n_439, wc103, n_270);
  not gc103 (wc103, n_342);
  and g611 (n_442, n_345, wc104);
  not gc104 (wc104, n_346);
  and g612 (n_407, wc105, n_200);
  not gc105 (wc105, n_353);
  and g613 (n_412, wc106, n_290);
  not gc106 (wc106, n_357);
  and g614 (n_417, n_360, wc107);
  not gc107 (wc107, n_361);
  and g615 (n_423, wc108, n_420);
  not gc108 (wc108, n_389);
  and g616 (n_395, wc109, n_283);
  not gc109 (wc109, n_389);
  and g617 (n_408, wc110, n_405);
  not gc110 (wc110, n_389);
  and g618 (n_413, wc111, n_410);
  not gc111 (wc111, n_389);
  and g619 (n_418, wc112, n_415);
  not gc112 (wc112, n_389);
  and g620 (n_475, wc113, n_422);
  not gc113 (wc113, n_423);
  or g621 (n_369, wc114, n_145);
  not gc114 (wc114, n_367);
  or g622 (n_374, n_371, wc115);
  not gc115 (wc115, n_367);
  or g623 (n_376, wc116, n_325);
  not gc116 (wc116, n_367);
  and g624 (n_447, wc117, n_188);
  not gc117 (wc117, n_390);
  and g625 (n_451, wc118, n_280);
  not gc118 (wc118, n_395);
  and g626 (n_455, n_398, wc119);
  not gc119 (wc119, n_399);
  and g627 (n_459, n_352, wc120);
  not gc120 (wc120, n_402);
  and g628 (n_463, wc121, n_407);
  not gc121 (wc121, n_408);
  and g629 (n_467, wc122, n_412);
  not gc122 (wc122, n_413);
  and g630 (n_471, wc123, n_417);
  not gc123 (wc123, n_418);
  or g631 (n_476, n_473, wc124);
  not gc124 (wc124, n_425);
  or g632 (n_427, wc125, n_169);
  not gc125 (wc125, n_425);
  or g633 (n_432, n_429, wc126);
  not gc126 (wc126, n_425);
  or g634 (n_434, wc127, n_340);
  not gc127 (wc127, n_425);
  or g635 (n_448, n_445, wc128);
  not gc128 (wc128, n_425);
  or g636 (n_452, n_449, wc129);
  not gc129 (wc129, n_425);
  or g637 (n_456, n_453, wc130);
  not gc130 (wc130, n_425);
  or g638 (n_460, n_457, wc131);
  not gc131 (wc131, n_425);
  or g639 (n_464, n_461, wc132);
  not gc132 (wc132, n_425);
  or g640 (n_468, n_465, wc133);
  not gc133 (wc133, n_425);
  or g641 (n_472, n_469, wc134);
  not gc134 (wc134, n_425);
  or g642 (n_488, wc135, n_485);
  not gc135 (wc135, n_477);
  or g643 (n_479, wc136, n_217);
  not gc136 (wc136, n_477);
  or g644 (n_484, n_481, wc137);
  not gc137 (wc137, n_477);
endmodule

module add_signed_522_GENERIC(A, B, Z);
  input [35:0] A, B;
  output [36:0] Z;
  wire [35:0] A, B;
  wire [36:0] Z;
  add_signed_522_GENERIC_REAL g1(.A ({A[34], A[34:0]}), .B ({B[34],
       B[34:0]}), .Z (Z));
endmodule

module add_signed_533_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [37:0] A, B;
  output [37:0] Z;
  wire [37:0] A, B;
  wire [37:0] Z;
  wire n_120, n_123, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_133, n_134, n_135, n_136, n_137, n_139, n_140, n_141;
  wire n_142, n_143, n_145, n_146, n_147, n_148, n_149, n_151;
  wire n_152, n_153, n_154, n_155, n_157, n_158, n_159, n_160;
  wire n_161, n_163, n_164, n_165, n_166, n_167, n_169, n_170;
  wire n_171, n_172, n_173, n_175, n_176, n_177, n_178, n_179;
  wire n_181, n_182, n_183, n_184, n_185, n_187, n_188, n_189;
  wire n_190, n_191, n_193, n_194, n_195, n_196, n_197, n_199;
  wire n_200, n_201, n_202, n_203, n_205, n_206, n_207, n_208;
  wire n_209, n_211, n_212, n_213, n_214, n_215, n_217, n_218;
  wire n_219, n_220, n_221, n_223, n_224, n_225, n_226, n_227;
  wire n_229, n_230, n_231, n_232, n_235, n_236, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_245, n_247, n_249, n_250;
  wire n_252, n_253, n_255, n_257, n_259, n_260, n_262, n_263;
  wire n_265, n_267, n_269, n_270, n_272, n_273, n_275, n_277;
  wire n_279, n_280, n_282, n_283, n_285, n_287, n_289, n_290;
  wire n_292, n_293, n_295, n_297, n_299, n_300, n_302, n_303;
  wire n_305, n_307, n_309, n_310, n_312, n_313, n_315, n_317;
  wire n_319, n_320, n_322, n_324, n_325, n_326, n_328, n_329;
  wire n_330, n_332, n_333, n_334, n_335, n_337, n_339, n_341;
  wire n_342, n_343, n_345, n_346, n_347, n_349, n_350, n_352;
  wire n_354, n_356, n_357, n_358, n_360, n_361, n_362, n_364;
  wire n_365, n_367, n_369, n_371, n_372, n_373, n_375, n_376;
  wire n_377, n_379, n_380, n_382, n_388, n_390, n_391, n_392;
  wire n_394, n_395, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_413, n_416, n_418, n_419, n_420, n_423, n_426;
  wire n_428, n_429, n_431, n_433, n_434, n_436, n_438, n_439;
  wire n_441, n_443, n_444, n_446, n_448, n_449, n_450, n_452;
  wire n_453, n_455, n_456, n_457, n_458, n_459, n_460, n_461;
  wire n_462, n_463, n_464, n_465, n_466, n_468, n_469, n_470;
  wire n_472, n_473, n_474, n_476, n_477, n_478, n_480, n_481;
  wire n_482, n_484, n_485, n_486, n_488, n_489, n_490, n_492;
  wire n_493, n_494, n_496, n_497, n_498, n_500, n_501, n_502;
  wire n_504, n_505, n_507, n_508, n_509, n_510, n_514, n_515;
  wire n_517, n_518, n_519, n_521, n_522, n_523, n_524, n_526;
  wire n_527, n_528, n_530, n_531, n_532, n_533, n_535, n_536;
  wire n_538, n_539, n_541, n_542, n_543, n_544, n_546, n_547;
  wire n_548, n_550, n_551, n_552, n_553, n_555, n_556, n_558;
  wire n_559, n_561, n_562, n_563, n_564, n_566, n_567, n_568;
  wire n_569, n_571, n_572, n_573, n_574, n_576, n_577, n_579;
  wire n_580, n_582, n_583, n_584, n_585, n_587, n_588, n_589;
  wire n_591, n_592, n_593, n_594, n_596, n_597, n_599, n_600;
  wire n_602, n_603;
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_120, A[0], B[0]);
  nor g9 (n_123, A[1], B[1]);
  nand g10 (n_126, A[1], B[1]);
  nor g11 (n_133, A[2], B[2]);
  nand g12 (n_128, A[2], B[2]);
  nor g13 (n_129, A[3], B[3]);
  nand g14 (n_130, A[3], B[3]);
  nor g15 (n_139, A[4], B[4]);
  nand g16 (n_134, A[4], B[4]);
  nor g17 (n_135, A[5], B[5]);
  nand g18 (n_136, A[5], B[5]);
  nor g19 (n_145, A[6], B[6]);
  nand g20 (n_140, A[6], B[6]);
  nor g21 (n_141, A[7], B[7]);
  nand g22 (n_142, A[7], B[7]);
  nor g23 (n_151, A[8], B[8]);
  nand g24 (n_146, A[8], B[8]);
  nor g25 (n_147, A[9], B[9]);
  nand g26 (n_148, A[9], B[9]);
  nor g27 (n_157, A[10], B[10]);
  nand g28 (n_152, A[10], B[10]);
  nor g29 (n_153, A[11], B[11]);
  nand g30 (n_154, A[11], B[11]);
  nor g31 (n_163, A[12], B[12]);
  nand g32 (n_158, A[12], B[12]);
  nor g33 (n_159, A[13], B[13]);
  nand g34 (n_160, A[13], B[13]);
  nor g35 (n_169, A[14], B[14]);
  nand g36 (n_164, A[14], B[14]);
  nor g37 (n_165, A[15], B[15]);
  nand g38 (n_166, A[15], B[15]);
  nor g39 (n_175, A[16], B[16]);
  nand g40 (n_170, A[16], B[16]);
  nor g41 (n_171, A[17], B[17]);
  nand g42 (n_172, A[17], B[17]);
  nor g43 (n_181, A[18], B[18]);
  nand g44 (n_176, A[18], B[18]);
  nor g45 (n_177, A[19], B[19]);
  nand g46 (n_178, A[19], B[19]);
  nor g47 (n_187, A[20], B[20]);
  nand g48 (n_182, A[20], B[20]);
  nor g49 (n_183, A[21], B[21]);
  nand g50 (n_184, A[21], B[21]);
  nor g51 (n_193, A[22], B[22]);
  nand g52 (n_188, A[22], B[22]);
  nor g53 (n_189, A[23], B[23]);
  nand g54 (n_190, A[23], B[23]);
  nor g55 (n_199, A[24], B[24]);
  nand g56 (n_194, A[24], B[24]);
  nor g57 (n_195, A[25], B[25]);
  nand g58 (n_196, A[25], B[25]);
  nor g59 (n_205, A[26], B[26]);
  nand g60 (n_200, A[26], B[26]);
  nor g61 (n_201, A[27], B[27]);
  nand g62 (n_202, A[27], B[27]);
  nor g63 (n_211, A[28], B[28]);
  nand g64 (n_206, A[28], B[28]);
  nor g65 (n_207, A[29], B[29]);
  nand g66 (n_208, A[29], B[29]);
  nor g67 (n_217, A[30], B[30]);
  nand g68 (n_212, A[30], B[30]);
  nor g69 (n_213, A[31], B[31]);
  nand g70 (n_214, A[31], B[31]);
  nor g71 (n_223, A[32], B[32]);
  nand g72 (n_218, A[32], B[32]);
  nor g73 (n_219, A[33], B[33]);
  nand g74 (n_220, A[33], B[33]);
  nor g75 (n_229, A[34], B[34]);
  nand g76 (n_224, A[34], B[34]);
  nor g77 (n_225, A[35], B[35]);
  nand g78 (n_226, A[35], B[35]);
  nor g79 (n_235, A[36], B[36]);
  nand g80 (n_230, A[36], B[36]);
  nand g85 (n_236, n_126, n_127);
  nor g86 (n_131, n_128, n_129);
  nor g89 (n_239, n_133, n_129);
  nor g90 (n_137, n_134, n_135);
  nor g93 (n_245, n_139, n_135);
  nor g94 (n_143, n_140, n_141);
  nor g97 (n_247, n_145, n_141);
  nor g98 (n_149, n_146, n_147);
  nor g101 (n_255, n_151, n_147);
  nor g102 (n_155, n_152, n_153);
  nor g105 (n_257, n_157, n_153);
  nor g106 (n_161, n_158, n_159);
  nor g109 (n_265, n_163, n_159);
  nor g110 (n_167, n_164, n_165);
  nor g113 (n_267, n_169, n_165);
  nor g114 (n_173, n_170, n_171);
  nor g117 (n_275, n_175, n_171);
  nor g118 (n_179, n_176, n_177);
  nor g121 (n_277, n_181, n_177);
  nor g122 (n_185, n_182, n_183);
  nor g125 (n_285, n_187, n_183);
  nor g126 (n_191, n_188, n_189);
  nor g129 (n_287, n_193, n_189);
  nor g130 (n_197, n_194, n_195);
  nor g133 (n_295, n_199, n_195);
  nor g134 (n_203, n_200, n_201);
  nor g137 (n_297, n_205, n_201);
  nor g138 (n_209, n_206, n_207);
  nor g141 (n_305, n_211, n_207);
  nor g142 (n_215, n_212, n_213);
  nor g145 (n_307, n_217, n_213);
  nor g146 (n_221, n_218, n_219);
  nor g149 (n_315, n_223, n_219);
  nor g150 (n_227, n_224, n_225);
  nor g153 (n_317, n_229, n_225);
  nand g160 (n_517, n_128, n_238);
  nand g161 (n_241, n_239, n_236);
  nand g162 (n_322, n_240, n_241);
  nor g163 (n_243, n_145, n_242);
  nand g172 (n_330, n_245, n_247);
  nor g173 (n_253, n_157, n_252);
  nand g182 (n_337, n_255, n_257);
  nor g183 (n_263, n_169, n_262);
  nand g192 (n_345, n_265, n_267);
  nor g193 (n_273, n_181, n_272);
  nand g202 (n_352, n_275, n_277);
  nor g203 (n_283, n_193, n_282);
  nand g212 (n_360, n_285, n_287);
  nor g213 (n_293, n_205, n_292);
  nand g222 (n_367, n_295, n_297);
  nor g223 (n_303, n_217, n_302);
  nand g232 (n_375, n_305, n_307);
  nor g233 (n_313, n_229, n_312);
  nand g242 (n_382, n_315, n_317);
  nand g245 (n_521, n_134, n_324);
  nand g246 (n_325, n_245, n_322);
  nand g247 (n_523, n_242, n_325);
  nand g250 (n_526, n_328, n_329);
  nand g253 (n_388, n_332, n_333);
  nor g254 (n_335, n_163, n_334);
  nor g257 (n_398, n_163, n_337);
  nor g263 (n_343, n_341, n_334);
  nor g266 (n_404, n_337, n_341);
  nor g267 (n_347, n_345, n_334);
  nor g270 (n_407, n_337, n_345);
  nor g271 (n_350, n_187, n_349);
  nor g274 (n_456, n_187, n_352);
  nor g280 (n_358, n_356, n_349);
  nor g283 (n_462, n_352, n_356);
  nor g284 (n_362, n_360, n_349);
  nor g287 (n_413, n_352, n_360);
  nor g288 (n_365, n_211, n_364);
  nor g291 (n_426, n_211, n_367);
  nor g297 (n_373, n_371, n_364);
  nor g300 (n_436, n_367, n_371);
  nor g301 (n_377, n_375, n_364);
  nor g304 (n_441, n_367, n_375);
  nor g305 (n_380, n_235, n_379);
  nor g308 (n_508, n_235, n_382);
  nand g316 (n_530, n_146, n_390);
  nand g317 (n_391, n_255, n_388);
  nand g318 (n_532, n_252, n_391);
  nand g321 (n_535, n_394, n_395);
  nand g324 (n_538, n_334, n_397);
  nand g325 (n_400, n_398, n_388);
  nand g326 (n_541, n_399, n_400);
  nand g327 (n_403, n_401, n_388);
  nand g328 (n_543, n_402, n_403);
  nand g329 (n_406, n_404, n_388);
  nand g330 (n_546, n_405, n_406);
  nand g331 (n_409, n_407, n_388);
  nand g332 (n_446, n_408, n_409);
  nor g333 (n_411, n_199, n_410);
  nand g342 (n_470, n_295, n_413);
  nor g343 (n_420, n_418, n_410);
  nor g348 (n_423, n_367, n_410);
  nand g357 (n_482, n_413, n_426);
  nand g362 (n_486, n_413, n_431);
  nand g367 (n_490, n_413, n_436);
  nand g372 (n_494, n_413, n_441);
  nand g375 (n_550, n_170, n_448);
  nand g376 (n_449, n_275, n_446);
  nand g377 (n_552, n_272, n_449);
  nand g380 (n_555, n_452, n_453);
  nand g383 (n_558, n_349, n_455);
  nand g384 (n_458, n_456, n_446);
  nand g385 (n_561, n_457, n_458);
  nand g386 (n_461, n_459, n_446);
  nand g387 (n_563, n_460, n_461);
  nand g388 (n_464, n_462, n_446);
  nand g389 (n_566, n_463, n_464);
  nand g390 (n_465, n_413, n_446);
  nand g391 (n_568, n_410, n_465);
  nand g394 (n_571, n_468, n_469);
  nand g397 (n_573, n_472, n_473);
  nand g400 (n_576, n_476, n_477);
  nand g403 (n_579, n_480, n_481);
  nand g406 (n_582, n_484, n_485);
  nand g409 (n_584, n_488, n_489);
  nand g412 (n_587, n_492, n_493);
  nand g415 (n_498, n_496, n_497);
  nand g418 (n_591, n_218, n_500);
  nand g419 (n_501, n_315, n_498);
  nand g420 (n_593, n_312, n_501);
  nand g423 (n_596, n_504, n_505);
  nand g426 (n_599, n_379, n_507);
  nand g427 (n_510, n_508, n_498);
  nand g428 (n_602, n_509, n_510);
  xnor g434 (Z[2], n_236, n_515);
  xnor g437 (Z[3], n_517, n_518);
  xnor g439 (Z[4], n_322, n_519);
  xnor g442 (Z[5], n_521, n_522);
  xnor g444 (Z[6], n_523, n_524);
  xnor g447 (Z[7], n_526, n_527);
  xnor g449 (Z[8], n_388, n_528);
  xnor g452 (Z[9], n_530, n_531);
  xnor g454 (Z[10], n_532, n_533);
  xnor g457 (Z[11], n_535, n_536);
  xnor g460 (Z[12], n_538, n_539);
  xnor g463 (Z[13], n_541, n_542);
  xnor g465 (Z[14], n_543, n_544);
  xnor g468 (Z[15], n_546, n_547);
  xnor g470 (Z[16], n_446, n_548);
  xnor g473 (Z[17], n_550, n_551);
  xnor g475 (Z[18], n_552, n_553);
  xnor g478 (Z[19], n_555, n_556);
  xnor g481 (Z[20], n_558, n_559);
  xnor g484 (Z[21], n_561, n_562);
  xnor g486 (Z[22], n_563, n_564);
  xnor g489 (Z[23], n_566, n_567);
  xnor g491 (Z[24], n_568, n_569);
  xnor g494 (Z[25], n_571, n_572);
  xnor g496 (Z[26], n_573, n_574);
  xnor g499 (Z[27], n_576, n_577);
  xnor g502 (Z[28], n_579, n_580);
  xnor g505 (Z[29], n_582, n_583);
  xnor g507 (Z[30], n_584, n_585);
  xnor g510 (Z[31], n_587, n_588);
  xnor g512 (Z[32], n_498, n_589);
  xnor g515 (Z[33], n_591, n_592);
  xnor g517 (Z[34], n_593, n_594);
  xnor g520 (Z[35], n_596, n_597);
  xnor g523 (Z[36], n_599, n_600);
  xnor g526 (Z[37], n_602, n_603);
  and g529 (n_231, A[37], B[37]);
  or g530 (n_232, A[37], B[37]);
  or g531 (n_127, n_120, n_123);
  and g532 (n_240, wc, n_130);
  not gc (wc, n_131);
  and g533 (n_242, wc0, n_136);
  not gc0 (wc0, n_137);
  and g534 (n_249, wc1, n_142);
  not gc1 (wc1, n_143);
  and g535 (n_252, wc2, n_148);
  not gc2 (wc2, n_149);
  and g536 (n_259, wc3, n_154);
  not gc3 (wc3, n_155);
  and g537 (n_262, wc4, n_160);
  not gc4 (wc4, n_161);
  and g538 (n_269, wc5, n_166);
  not gc5 (wc5, n_167);
  and g539 (n_272, wc6, n_172);
  not gc6 (wc6, n_173);
  and g540 (n_279, wc7, n_178);
  not gc7 (wc7, n_179);
  and g541 (n_282, wc8, n_184);
  not gc8 (wc8, n_185);
  and g542 (n_289, wc9, n_190);
  not gc9 (wc9, n_191);
  and g543 (n_292, wc10, n_196);
  not gc10 (wc10, n_197);
  and g544 (n_299, wc11, n_202);
  not gc11 (wc11, n_203);
  and g545 (n_302, wc12, n_208);
  not gc12 (wc12, n_209);
  and g546 (n_309, wc13, n_214);
  not gc13 (wc13, n_215);
  and g547 (n_312, wc14, n_220);
  not gc14 (wc14, n_221);
  and g548 (n_319, wc15, n_226);
  not gc15 (wc15, n_227);
  or g549 (n_326, wc16, n_145);
  not gc16 (wc16, n_245);
  or g550 (n_392, wc17, n_157);
  not gc17 (wc17, n_255);
  or g551 (n_341, wc18, n_169);
  not gc18 (wc18, n_265);
  or g552 (n_450, wc19, n_181);
  not gc19 (wc19, n_275);
  or g553 (n_356, wc20, n_193);
  not gc20 (wc20, n_285);
  or g554 (n_418, wc21, n_205);
  not gc21 (wc21, n_295);
  or g555 (n_371, wc22, n_217);
  not gc22 (wc22, n_305);
  or g556 (n_502, wc23, n_229);
  not gc23 (wc23, n_315);
  or g557 (n_514, wc24, n_123);
  not gc24 (wc24, n_126);
  or g558 (n_515, wc25, n_133);
  not gc25 (wc25, n_128);
  or g559 (n_518, wc26, n_129);
  not gc26 (wc26, n_130);
  or g560 (n_519, wc27, n_139);
  not gc27 (wc27, n_134);
  or g561 (n_522, wc28, n_135);
  not gc28 (wc28, n_136);
  or g562 (n_524, wc29, n_145);
  not gc29 (wc29, n_140);
  or g563 (n_527, wc30, n_141);
  not gc30 (wc30, n_142);
  or g564 (n_528, wc31, n_151);
  not gc31 (wc31, n_146);
  or g565 (n_531, wc32, n_147);
  not gc32 (wc32, n_148);
  or g566 (n_533, wc33, n_157);
  not gc33 (wc33, n_152);
  or g567 (n_536, wc34, n_153);
  not gc34 (wc34, n_154);
  or g568 (n_539, wc35, n_163);
  not gc35 (wc35, n_158);
  or g569 (n_542, wc36, n_159);
  not gc36 (wc36, n_160);
  or g570 (n_544, wc37, n_169);
  not gc37 (wc37, n_164);
  or g571 (n_547, wc38, n_165);
  not gc38 (wc38, n_166);
  or g572 (n_548, wc39, n_175);
  not gc39 (wc39, n_170);
  or g573 (n_551, wc40, n_171);
  not gc40 (wc40, n_172);
  or g574 (n_553, wc41, n_181);
  not gc41 (wc41, n_176);
  or g575 (n_556, wc42, n_177);
  not gc42 (wc42, n_178);
  or g576 (n_559, wc43, n_187);
  not gc43 (wc43, n_182);
  or g577 (n_562, wc44, n_183);
  not gc44 (wc44, n_184);
  or g578 (n_564, wc45, n_193);
  not gc45 (wc45, n_188);
  or g579 (n_567, wc46, n_189);
  not gc46 (wc46, n_190);
  or g580 (n_569, wc47, n_199);
  not gc47 (wc47, n_194);
  or g581 (n_572, wc48, n_195);
  not gc48 (wc48, n_196);
  or g582 (n_574, wc49, n_205);
  not gc49 (wc49, n_200);
  or g583 (n_577, wc50, n_201);
  not gc50 (wc50, n_202);
  or g584 (n_580, wc51, n_211);
  not gc51 (wc51, n_206);
  or g585 (n_583, wc52, n_207);
  not gc52 (wc52, n_208);
  or g586 (n_585, wc53, n_217);
  not gc53 (wc53, n_212);
  or g587 (n_588, wc54, n_213);
  not gc54 (wc54, n_214);
  or g588 (n_589, wc55, n_223);
  not gc55 (wc55, n_218);
  or g589 (n_592, wc56, n_219);
  not gc56 (wc56, n_220);
  or g590 (n_594, wc57, n_229);
  not gc57 (wc57, n_224);
  or g591 (n_597, wc58, n_225);
  not gc58 (wc58, n_226);
  or g592 (n_600, wc59, n_235);
  not gc59 (wc59, n_230);
  and g593 (n_250, wc60, n_247);
  not gc60 (wc60, n_242);
  and g594 (n_260, wc61, n_257);
  not gc61 (wc61, n_252);
  and g595 (n_270, wc62, n_267);
  not gc62 (wc62, n_262);
  and g596 (n_280, wc63, n_277);
  not gc63 (wc63, n_272);
  and g597 (n_290, wc64, n_287);
  not gc64 (wc64, n_282);
  and g598 (n_300, wc65, n_297);
  not gc65 (wc65, n_292);
  and g599 (n_310, wc66, n_307);
  not gc66 (wc66, n_302);
  and g600 (n_320, wc67, n_317);
  not gc67 (wc67, n_312);
  and g601 (n_401, wc68, n_265);
  not gc68 (wc68, n_337);
  and g602 (n_459, wc69, n_285);
  not gc69 (wc69, n_352);
  and g603 (n_431, wc70, n_305);
  not gc70 (wc70, n_367);
  xor g604 (Z[1], n_120, n_514);
  or g605 (n_603, wc71, n_231);
  not gc71 (wc71, n_232);
  or g606 (n_238, wc72, n_133);
  not gc72 (wc72, n_236);
  and g607 (n_328, wc73, n_140);
  not gc73 (wc73, n_243);
  and g608 (n_332, wc74, n_249);
  not gc74 (wc74, n_250);
  and g609 (n_394, wc75, n_152);
  not gc75 (wc75, n_253);
  and g610 (n_334, wc76, n_259);
  not gc76 (wc76, n_260);
  and g611 (n_342, wc77, n_164);
  not gc77 (wc77, n_263);
  and g612 (n_346, wc78, n_269);
  not gc78 (wc78, n_270);
  and g613 (n_452, wc79, n_176);
  not gc79 (wc79, n_273);
  and g614 (n_349, wc80, n_279);
  not gc80 (wc80, n_280);
  and g615 (n_357, wc81, n_188);
  not gc81 (wc81, n_283);
  and g616 (n_361, wc82, n_289);
  not gc82 (wc82, n_290);
  and g617 (n_419, wc83, n_200);
  not gc83 (wc83, n_293);
  and g618 (n_364, wc84, n_299);
  not gc84 (wc84, n_300);
  and g619 (n_372, wc85, n_212);
  not gc85 (wc85, n_303);
  and g620 (n_376, wc86, n_309);
  not gc86 (wc86, n_310);
  and g621 (n_504, wc87, n_224);
  not gc87 (wc87, n_313);
  and g622 (n_379, wc88, n_319);
  not gc88 (wc88, n_320);
  or g623 (n_466, wc89, n_199);
  not gc89 (wc89, n_413);
  or g624 (n_474, n_418, wc90);
  not gc90 (wc90, n_413);
  or g625 (n_478, wc91, n_367);
  not gc91 (wc91, n_413);
  and g626 (n_339, wc92, n_265);
  not gc92 (wc92, n_334);
  and g627 (n_354, wc93, n_285);
  not gc93 (wc93, n_349);
  and g628 (n_369, wc94, n_305);
  not gc94 (wc94, n_364);
  or g629 (n_324, wc95, n_139);
  not gc95 (wc95, n_322);
  or g630 (n_329, n_326, wc96);
  not gc96 (wc96, n_322);
  or g631 (n_333, n_330, wc97);
  not gc97 (wc97, n_322);
  and g632 (n_399, wc98, n_158);
  not gc98 (wc98, n_335);
  and g633 (n_402, wc99, n_262);
  not gc99 (wc99, n_339);
  and g634 (n_405, n_342, wc100);
  not gc100 (wc100, n_343);
  and g635 (n_408, n_346, wc101);
  not gc101 (wc101, n_347);
  and g636 (n_457, wc102, n_182);
  not gc102 (wc102, n_350);
  and g637 (n_460, wc103, n_282);
  not gc103 (wc103, n_354);
  and g638 (n_463, n_357, wc104);
  not gc104 (wc104, n_358);
  and g639 (n_410, n_361, wc105);
  not gc105 (wc105, n_362);
  and g640 (n_428, wc106, n_206);
  not gc106 (wc106, n_365);
  and g641 (n_433, wc107, n_302);
  not gc107 (wc107, n_369);
  and g642 (n_438, n_372, wc108);
  not gc108 (wc108, n_373);
  and g643 (n_443, n_376, wc109);
  not gc109 (wc109, n_377);
  and g644 (n_509, wc110, n_230);
  not gc110 (wc110, n_380);
  and g645 (n_416, wc111, n_295);
  not gc111 (wc111, n_410);
  and g646 (n_429, wc112, n_426);
  not gc112 (wc112, n_410);
  and g647 (n_434, wc113, n_431);
  not gc113 (wc113, n_410);
  and g648 (n_439, wc114, n_436);
  not gc114 (wc114, n_410);
  and g649 (n_444, wc115, n_441);
  not gc115 (wc115, n_410);
  or g650 (n_390, wc116, n_151);
  not gc116 (wc116, n_388);
  or g651 (n_395, n_392, wc117);
  not gc117 (wc117, n_388);
  or g652 (n_397, wc118, n_337);
  not gc118 (wc118, n_388);
  and g653 (n_468, wc119, n_194);
  not gc119 (wc119, n_411);
  and g654 (n_472, wc120, n_292);
  not gc120 (wc120, n_416);
  and g655 (n_476, n_419, wc121);
  not gc121 (wc121, n_420);
  and g656 (n_480, n_364, wc122);
  not gc122 (wc122, n_423);
  and g657 (n_484, wc123, n_428);
  not gc123 (wc123, n_429);
  and g658 (n_488, wc124, n_433);
  not gc124 (wc124, n_434);
  and g659 (n_492, wc125, n_438);
  not gc125 (wc125, n_439);
  and g660 (n_496, wc126, n_443);
  not gc126 (wc126, n_444);
  or g661 (n_448, wc127, n_175);
  not gc127 (wc127, n_446);
  or g662 (n_453, n_450, wc128);
  not gc128 (wc128, n_446);
  or g663 (n_455, wc129, n_352);
  not gc129 (wc129, n_446);
  or g664 (n_469, n_466, wc130);
  not gc130 (wc130, n_446);
  or g665 (n_473, n_470, wc131);
  not gc131 (wc131, n_446);
  or g666 (n_477, n_474, wc132);
  not gc132 (wc132, n_446);
  or g667 (n_481, n_478, wc133);
  not gc133 (wc133, n_446);
  or g668 (n_485, n_482, wc134);
  not gc134 (wc134, n_446);
  or g669 (n_489, n_486, wc135);
  not gc135 (wc135, n_446);
  or g670 (n_493, n_490, wc136);
  not gc136 (wc136, n_446);
  or g671 (n_497, n_494, wc137);
  not gc137 (wc137, n_446);
  or g672 (n_500, wc138, n_223);
  not gc138 (wc138, n_498);
  or g673 (n_505, n_502, wc139);
  not gc139 (wc139, n_498);
  or g674 (n_507, wc140, n_382);
  not gc140 (wc140, n_498);
endmodule

module add_signed_533_GENERIC(A, B, Z);
  input [37:0] A, B;
  output [37:0] Z;
  wire [37:0] A, B;
  wire [37:0] Z;
  add_signed_533_GENERIC_REAL g1(.A ({A[36], A[36:0]}), .B ({B[36],
       B[36:0]}), .Z (Z));
endmodule

module add_signed_6294_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [53:0] A, B;
  output [54:0] Z;
  wire [53:0] A, B;
  wire [54:0] Z;
  wire n_167, n_168, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436;
  not g3 (Z[54], n_167);
  nand g4 (n_168, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_173, A[1], B[1]);
  nand g13 (n_177, n_173, n_174, n_175);
  xor g14 (n_176, A[1], B[1]);
  nand g16 (n_178, A[2], B[2]);
  nand g17 (n_179, A[2], n_177);
  nand g18 (n_180, B[2], n_177);
  nand g19 (n_182, n_178, n_179, n_180);
  xor g20 (n_181, A[2], B[2]);
  xor g21 (Z[2], n_177, n_181);
  nand g22 (n_183, A[3], B[3]);
  nand g23 (n_184, A[3], n_182);
  nand g24 (n_185, B[3], n_182);
  nand g25 (n_187, n_183, n_184, n_185);
  xor g26 (n_186, A[3], B[3]);
  xor g27 (Z[3], n_182, n_186);
  nand g28 (n_188, A[4], B[4]);
  nand g29 (n_189, A[4], n_187);
  nand g30 (n_190, B[4], n_187);
  nand g31 (n_192, n_188, n_189, n_190);
  xor g32 (n_191, A[4], B[4]);
  xor g33 (Z[4], n_187, n_191);
  nand g34 (n_193, A[5], B[5]);
  nand g35 (n_194, A[5], n_192);
  nand g36 (n_195, B[5], n_192);
  nand g37 (n_197, n_193, n_194, n_195);
  xor g38 (n_196, A[5], B[5]);
  xor g39 (Z[5], n_192, n_196);
  nand g40 (n_198, A[6], B[6]);
  nand g41 (n_199, A[6], n_197);
  nand g42 (n_200, B[6], n_197);
  nand g43 (n_202, n_198, n_199, n_200);
  xor g44 (n_201, A[6], B[6]);
  xor g45 (Z[6], n_197, n_201);
  nand g46 (n_203, A[7], B[7]);
  nand g47 (n_204, A[7], n_202);
  nand g48 (n_205, B[7], n_202);
  nand g49 (n_207, n_203, n_204, n_205);
  xor g50 (n_206, A[7], B[7]);
  xor g51 (Z[7], n_202, n_206);
  nand g52 (n_208, A[8], B[8]);
  nand g53 (n_209, A[8], n_207);
  nand g54 (n_210, B[8], n_207);
  nand g55 (n_212, n_208, n_209, n_210);
  xor g56 (n_211, A[8], B[8]);
  xor g57 (Z[8], n_207, n_211);
  nand g58 (n_213, A[9], B[9]);
  nand g59 (n_214, A[9], n_212);
  nand g60 (n_215, B[9], n_212);
  nand g61 (n_217, n_213, n_214, n_215);
  xor g62 (n_216, A[9], B[9]);
  xor g63 (Z[9], n_212, n_216);
  nand g64 (n_218, A[10], B[10]);
  nand g65 (n_219, A[10], n_217);
  nand g66 (n_220, B[10], n_217);
  nand g67 (n_222, n_218, n_219, n_220);
  xor g68 (n_221, A[10], B[10]);
  xor g69 (Z[10], n_217, n_221);
  nand g70 (n_223, A[11], B[11]);
  nand g71 (n_224, A[11], n_222);
  nand g72 (n_225, B[11], n_222);
  nand g73 (n_227, n_223, n_224, n_225);
  xor g74 (n_226, A[11], B[11]);
  xor g75 (Z[11], n_222, n_226);
  nand g76 (n_228, A[12], B[12]);
  nand g77 (n_229, A[12], n_227);
  nand g78 (n_230, B[12], n_227);
  nand g79 (n_232, n_228, n_229, n_230);
  xor g80 (n_231, A[12], B[12]);
  xor g81 (Z[12], n_227, n_231);
  nand g82 (n_233, A[13], B[13]);
  nand g83 (n_234, A[13], n_232);
  nand g84 (n_235, B[13], n_232);
  nand g85 (n_237, n_233, n_234, n_235);
  xor g86 (n_236, A[13], B[13]);
  xor g87 (Z[13], n_232, n_236);
  nand g88 (n_238, A[14], B[14]);
  nand g89 (n_239, A[14], n_237);
  nand g90 (n_240, B[14], n_237);
  nand g91 (n_242, n_238, n_239, n_240);
  xor g92 (n_241, A[14], B[14]);
  xor g93 (Z[14], n_237, n_241);
  nand g94 (n_243, A[15], B[15]);
  nand g95 (n_244, A[15], n_242);
  nand g96 (n_245, B[15], n_242);
  nand g97 (n_247, n_243, n_244, n_245);
  xor g98 (n_246, A[15], B[15]);
  xor g99 (Z[15], n_242, n_246);
  nand g100 (n_248, A[16], B[16]);
  nand g101 (n_249, A[16], n_247);
  nand g102 (n_250, B[16], n_247);
  nand g103 (n_252, n_248, n_249, n_250);
  xor g104 (n_251, A[16], B[16]);
  xor g105 (Z[16], n_247, n_251);
  nand g106 (n_253, A[17], B[17]);
  nand g107 (n_254, A[17], n_252);
  nand g108 (n_255, B[17], n_252);
  nand g109 (n_257, n_253, n_254, n_255);
  xor g110 (n_256, A[17], B[17]);
  xor g111 (Z[17], n_252, n_256);
  nand g112 (n_258, A[18], B[18]);
  nand g113 (n_259, A[18], n_257);
  nand g114 (n_260, B[18], n_257);
  nand g115 (n_262, n_258, n_259, n_260);
  xor g116 (n_261, A[18], B[18]);
  xor g117 (Z[18], n_257, n_261);
  nand g118 (n_263, A[19], B[19]);
  nand g119 (n_264, A[19], n_262);
  nand g120 (n_265, B[19], n_262);
  nand g121 (n_267, n_263, n_264, n_265);
  xor g122 (n_266, A[19], B[19]);
  xor g123 (Z[19], n_262, n_266);
  nand g124 (n_268, A[20], B[20]);
  nand g125 (n_269, A[20], n_267);
  nand g126 (n_270, B[20], n_267);
  nand g127 (n_272, n_268, n_269, n_270);
  xor g128 (n_271, A[20], B[20]);
  xor g129 (Z[20], n_267, n_271);
  nand g130 (n_273, A[21], B[21]);
  nand g131 (n_274, A[21], n_272);
  nand g132 (n_275, B[21], n_272);
  nand g133 (n_277, n_273, n_274, n_275);
  xor g134 (n_276, A[21], B[21]);
  xor g135 (Z[21], n_272, n_276);
  nand g136 (n_278, A[22], B[22]);
  nand g137 (n_279, A[22], n_277);
  nand g138 (n_280, B[22], n_277);
  nand g139 (n_282, n_278, n_279, n_280);
  xor g140 (n_281, A[22], B[22]);
  xor g141 (Z[22], n_277, n_281);
  nand g142 (n_283, A[23], B[23]);
  nand g143 (n_284, A[23], n_282);
  nand g144 (n_285, B[23], n_282);
  nand g145 (n_287, n_283, n_284, n_285);
  xor g146 (n_286, A[23], B[23]);
  xor g147 (Z[23], n_282, n_286);
  nand g148 (n_288, A[24], B[24]);
  nand g149 (n_289, A[24], n_287);
  nand g150 (n_290, B[24], n_287);
  nand g151 (n_292, n_288, n_289, n_290);
  xor g152 (n_291, A[24], B[24]);
  xor g153 (Z[24], n_287, n_291);
  nand g154 (n_293, A[25], B[25]);
  nand g155 (n_294, A[25], n_292);
  nand g156 (n_295, B[25], n_292);
  nand g157 (n_297, n_293, n_294, n_295);
  xor g158 (n_296, A[25], B[25]);
  xor g159 (Z[25], n_292, n_296);
  nand g160 (n_298, A[26], B[26]);
  nand g161 (n_299, A[26], n_297);
  nand g162 (n_300, B[26], n_297);
  nand g163 (n_302, n_298, n_299, n_300);
  xor g164 (n_301, A[26], B[26]);
  xor g165 (Z[26], n_297, n_301);
  nand g166 (n_303, A[27], B[27]);
  nand g167 (n_304, A[27], n_302);
  nand g168 (n_305, B[27], n_302);
  nand g169 (n_307, n_303, n_304, n_305);
  xor g170 (n_306, A[27], B[27]);
  xor g171 (Z[27], n_302, n_306);
  nand g172 (n_308, A[28], B[28]);
  nand g173 (n_309, A[28], n_307);
  nand g174 (n_310, B[28], n_307);
  nand g175 (n_312, n_308, n_309, n_310);
  xor g176 (n_311, A[28], B[28]);
  xor g177 (Z[28], n_307, n_311);
  nand g178 (n_313, A[29], B[29]);
  nand g179 (n_314, A[29], n_312);
  nand g180 (n_315, B[29], n_312);
  nand g181 (n_317, n_313, n_314, n_315);
  xor g182 (n_316, A[29], B[29]);
  xor g183 (Z[29], n_312, n_316);
  nand g184 (n_318, A[30], B[30]);
  nand g185 (n_319, A[30], n_317);
  nand g186 (n_320, B[30], n_317);
  nand g187 (n_322, n_318, n_319, n_320);
  xor g188 (n_321, A[30], B[30]);
  xor g189 (Z[30], n_317, n_321);
  nand g190 (n_323, A[31], B[31]);
  nand g191 (n_324, A[31], n_322);
  nand g192 (n_325, B[31], n_322);
  nand g193 (n_327, n_323, n_324, n_325);
  xor g194 (n_326, A[31], B[31]);
  xor g195 (Z[31], n_322, n_326);
  nand g196 (n_328, A[32], B[32]);
  nand g197 (n_329, A[32], n_327);
  nand g198 (n_330, B[32], n_327);
  nand g199 (n_332, n_328, n_329, n_330);
  xor g200 (n_331, A[32], B[32]);
  xor g201 (Z[32], n_327, n_331);
  nand g202 (n_333, A[33], B[33]);
  nand g203 (n_334, A[33], n_332);
  nand g204 (n_335, B[33], n_332);
  nand g205 (n_337, n_333, n_334, n_335);
  xor g206 (n_336, A[33], B[33]);
  xor g207 (Z[33], n_332, n_336);
  nand g208 (n_338, A[34], B[34]);
  nand g209 (n_339, A[34], n_337);
  nand g210 (n_340, B[34], n_337);
  nand g211 (n_342, n_338, n_339, n_340);
  xor g212 (n_341, A[34], B[34]);
  xor g213 (Z[34], n_337, n_341);
  nand g214 (n_343, A[35], B[35]);
  nand g215 (n_344, A[35], n_342);
  nand g216 (n_345, B[35], n_342);
  nand g217 (n_347, n_343, n_344, n_345);
  xor g218 (n_346, A[35], B[35]);
  xor g219 (Z[35], n_342, n_346);
  nand g220 (n_348, A[36], B[36]);
  nand g221 (n_349, A[36], n_347);
  nand g222 (n_350, B[36], n_347);
  nand g223 (n_352, n_348, n_349, n_350);
  xor g224 (n_351, A[36], B[36]);
  xor g225 (Z[36], n_347, n_351);
  nand g226 (n_353, A[37], B[37]);
  nand g227 (n_354, A[37], n_352);
  nand g228 (n_355, B[37], n_352);
  nand g229 (n_357, n_353, n_354, n_355);
  xor g230 (n_356, A[37], B[37]);
  xor g231 (Z[37], n_352, n_356);
  nand g232 (n_358, A[38], B[38]);
  nand g233 (n_359, A[38], n_357);
  nand g234 (n_360, B[38], n_357);
  nand g235 (n_362, n_358, n_359, n_360);
  xor g236 (n_361, A[38], B[38]);
  xor g237 (Z[38], n_357, n_361);
  nand g238 (n_363, A[39], B[39]);
  nand g239 (n_364, A[39], n_362);
  nand g240 (n_365, B[39], n_362);
  nand g241 (n_367, n_363, n_364, n_365);
  xor g242 (n_366, A[39], B[39]);
  xor g243 (Z[39], n_362, n_366);
  nand g244 (n_368, A[40], B[40]);
  nand g245 (n_369, A[40], n_367);
  nand g246 (n_370, B[40], n_367);
  nand g247 (n_372, n_368, n_369, n_370);
  xor g248 (n_371, A[40], B[40]);
  xor g249 (Z[40], n_367, n_371);
  nand g250 (n_373, A[41], B[41]);
  nand g251 (n_374, A[41], n_372);
  nand g252 (n_375, B[41], n_372);
  nand g253 (n_377, n_373, n_374, n_375);
  xor g254 (n_376, A[41], B[41]);
  xor g255 (Z[41], n_372, n_376);
  nand g256 (n_378, A[42], B[42]);
  nand g257 (n_379, A[42], n_377);
  nand g258 (n_380, B[42], n_377);
  nand g259 (n_382, n_378, n_379, n_380);
  xor g260 (n_381, A[42], B[42]);
  xor g261 (Z[42], n_377, n_381);
  nand g262 (n_383, A[43], B[43]);
  nand g263 (n_384, A[43], n_382);
  nand g264 (n_385, B[43], n_382);
  nand g265 (n_387, n_383, n_384, n_385);
  xor g266 (n_386, A[43], B[43]);
  xor g267 (Z[43], n_382, n_386);
  nand g268 (n_388, A[44], B[44]);
  nand g269 (n_389, A[44], n_387);
  nand g270 (n_390, B[44], n_387);
  nand g271 (n_392, n_388, n_389, n_390);
  xor g272 (n_391, A[44], B[44]);
  xor g273 (Z[44], n_387, n_391);
  nand g274 (n_393, A[45], B[45]);
  nand g275 (n_394, A[45], n_392);
  nand g276 (n_395, B[45], n_392);
  nand g277 (n_397, n_393, n_394, n_395);
  xor g278 (n_396, A[45], B[45]);
  xor g279 (Z[45], n_392, n_396);
  nand g280 (n_398, A[46], B[46]);
  nand g281 (n_399, A[46], n_397);
  nand g282 (n_400, B[46], n_397);
  nand g283 (n_402, n_398, n_399, n_400);
  xor g284 (n_401, A[46], B[46]);
  xor g285 (Z[46], n_397, n_401);
  nand g286 (n_403, A[47], B[47]);
  nand g287 (n_404, A[47], n_402);
  nand g288 (n_405, B[47], n_402);
  nand g289 (n_407, n_403, n_404, n_405);
  xor g290 (n_406, A[47], B[47]);
  xor g291 (Z[47], n_402, n_406);
  nand g292 (n_408, A[48], B[48]);
  nand g293 (n_409, A[48], n_407);
  nand g294 (n_410, B[48], n_407);
  nand g295 (n_412, n_408, n_409, n_410);
  xor g296 (n_411, A[48], B[48]);
  xor g297 (Z[48], n_407, n_411);
  nand g298 (n_413, A[49], B[49]);
  nand g299 (n_414, A[49], n_412);
  nand g300 (n_415, B[49], n_412);
  nand g301 (n_417, n_413, n_414, n_415);
  xor g302 (n_416, A[49], B[49]);
  xor g303 (Z[49], n_412, n_416);
  nand g304 (n_418, A[50], B[50]);
  nand g305 (n_419, A[50], n_417);
  nand g306 (n_420, B[50], n_417);
  nand g307 (n_422, n_418, n_419, n_420);
  xor g308 (n_421, A[50], B[50]);
  xor g309 (Z[50], n_417, n_421);
  nand g310 (n_423, A[51], B[51]);
  nand g311 (n_424, A[51], n_422);
  nand g312 (n_425, B[51], n_422);
  nand g313 (n_427, n_423, n_424, n_425);
  xor g314 (n_426, A[51], B[51]);
  xor g315 (Z[51], n_422, n_426);
  nand g316 (n_428, A[52], B[52]);
  nand g317 (n_429, A[52], n_427);
  nand g318 (n_430, B[52], n_427);
  nand g319 (n_432, n_428, n_429, n_430);
  xor g320 (n_431, A[52], B[52]);
  xor g321 (Z[52], n_427, n_431);
  nand g325 (n_167, n_433, n_434, n_435);
  xor g327 (Z[53], n_432, n_436);
  or g329 (n_433, A[53], B[53]);
  xor g330 (n_436, A[53], B[53]);
  or g331 (n_174, wc, n_168);
  not gc (wc, A[1]);
  or g332 (n_175, wc0, n_168);
  not gc0 (wc0, B[1]);
  xnor g333 (Z[1], n_168, n_176);
  or g334 (n_434, A[53], wc1);
  not gc1 (wc1, n_432);
  or g335 (n_435, B[53], wc2);
  not gc2 (wc2, n_432);
endmodule

module add_signed_6294_GENERIC(A, B, Z);
  input [53:0] A, B;
  output [54:0] Z;
  wire [53:0] A, B;
  wire [54:0] Z;
  add_signed_6294_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_6294_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [53:0] A, B;
  output [54:0] Z;
  wire [53:0] A, B;
  wire [54:0] Z;
  wire n_167, n_168, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436;
  not g3 (Z[54], n_167);
  nand g4 (n_168, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_173, A[1], B[1]);
  nand g13 (n_177, n_173, n_174, n_175);
  xor g14 (n_176, A[1], B[1]);
  nand g16 (n_178, A[2], B[2]);
  nand g17 (n_179, A[2], n_177);
  nand g18 (n_180, B[2], n_177);
  nand g19 (n_182, n_178, n_179, n_180);
  xor g20 (n_181, A[2], B[2]);
  xor g21 (Z[2], n_177, n_181);
  nand g22 (n_183, A[3], B[3]);
  nand g23 (n_184, A[3], n_182);
  nand g24 (n_185, B[3], n_182);
  nand g25 (n_187, n_183, n_184, n_185);
  xor g26 (n_186, A[3], B[3]);
  xor g27 (Z[3], n_182, n_186);
  nand g28 (n_188, A[4], B[4]);
  nand g29 (n_189, A[4], n_187);
  nand g30 (n_190, B[4], n_187);
  nand g31 (n_192, n_188, n_189, n_190);
  xor g32 (n_191, A[4], B[4]);
  xor g33 (Z[4], n_187, n_191);
  nand g34 (n_193, A[5], B[5]);
  nand g35 (n_194, A[5], n_192);
  nand g36 (n_195, B[5], n_192);
  nand g37 (n_197, n_193, n_194, n_195);
  xor g38 (n_196, A[5], B[5]);
  xor g39 (Z[5], n_192, n_196);
  nand g40 (n_198, A[6], B[6]);
  nand g41 (n_199, A[6], n_197);
  nand g42 (n_200, B[6], n_197);
  nand g43 (n_202, n_198, n_199, n_200);
  xor g44 (n_201, A[6], B[6]);
  xor g45 (Z[6], n_197, n_201);
  nand g46 (n_203, A[7], B[7]);
  nand g47 (n_204, A[7], n_202);
  nand g48 (n_205, B[7], n_202);
  nand g49 (n_207, n_203, n_204, n_205);
  xor g50 (n_206, A[7], B[7]);
  xor g51 (Z[7], n_202, n_206);
  nand g52 (n_208, A[8], B[8]);
  nand g53 (n_209, A[8], n_207);
  nand g54 (n_210, B[8], n_207);
  nand g55 (n_212, n_208, n_209, n_210);
  xor g56 (n_211, A[8], B[8]);
  xor g57 (Z[8], n_207, n_211);
  nand g58 (n_213, A[9], B[9]);
  nand g59 (n_214, A[9], n_212);
  nand g60 (n_215, B[9], n_212);
  nand g61 (n_217, n_213, n_214, n_215);
  xor g62 (n_216, A[9], B[9]);
  xor g63 (Z[9], n_212, n_216);
  nand g64 (n_218, A[10], B[10]);
  nand g65 (n_219, A[10], n_217);
  nand g66 (n_220, B[10], n_217);
  nand g67 (n_222, n_218, n_219, n_220);
  xor g68 (n_221, A[10], B[10]);
  xor g69 (Z[10], n_217, n_221);
  nand g70 (n_223, A[11], B[11]);
  nand g71 (n_224, A[11], n_222);
  nand g72 (n_225, B[11], n_222);
  nand g73 (n_227, n_223, n_224, n_225);
  xor g74 (n_226, A[11], B[11]);
  xor g75 (Z[11], n_222, n_226);
  nand g76 (n_228, A[12], B[12]);
  nand g77 (n_229, A[12], n_227);
  nand g78 (n_230, B[12], n_227);
  nand g79 (n_232, n_228, n_229, n_230);
  xor g80 (n_231, A[12], B[12]);
  xor g81 (Z[12], n_227, n_231);
  nand g82 (n_233, A[13], B[13]);
  nand g83 (n_234, A[13], n_232);
  nand g84 (n_235, B[13], n_232);
  nand g85 (n_237, n_233, n_234, n_235);
  xor g86 (n_236, A[13], B[13]);
  xor g87 (Z[13], n_232, n_236);
  nand g88 (n_238, A[14], B[14]);
  nand g89 (n_239, A[14], n_237);
  nand g90 (n_240, B[14], n_237);
  nand g91 (n_242, n_238, n_239, n_240);
  xor g92 (n_241, A[14], B[14]);
  xor g93 (Z[14], n_237, n_241);
  nand g94 (n_243, A[15], B[15]);
  nand g95 (n_244, A[15], n_242);
  nand g96 (n_245, B[15], n_242);
  nand g97 (n_247, n_243, n_244, n_245);
  xor g98 (n_246, A[15], B[15]);
  xor g99 (Z[15], n_242, n_246);
  nand g100 (n_248, A[16], B[16]);
  nand g101 (n_249, A[16], n_247);
  nand g102 (n_250, B[16], n_247);
  nand g103 (n_252, n_248, n_249, n_250);
  xor g104 (n_251, A[16], B[16]);
  xor g105 (Z[16], n_247, n_251);
  nand g106 (n_253, A[17], B[17]);
  nand g107 (n_254, A[17], n_252);
  nand g108 (n_255, B[17], n_252);
  nand g109 (n_257, n_253, n_254, n_255);
  xor g110 (n_256, A[17], B[17]);
  xor g111 (Z[17], n_252, n_256);
  nand g112 (n_258, A[18], B[18]);
  nand g113 (n_259, A[18], n_257);
  nand g114 (n_260, B[18], n_257);
  nand g115 (n_262, n_258, n_259, n_260);
  xor g116 (n_261, A[18], B[18]);
  xor g117 (Z[18], n_257, n_261);
  nand g118 (n_263, A[19], B[19]);
  nand g119 (n_264, A[19], n_262);
  nand g120 (n_265, B[19], n_262);
  nand g121 (n_267, n_263, n_264, n_265);
  xor g122 (n_266, A[19], B[19]);
  xor g123 (Z[19], n_262, n_266);
  nand g124 (n_268, A[20], B[20]);
  nand g125 (n_269, A[20], n_267);
  nand g126 (n_270, B[20], n_267);
  nand g127 (n_272, n_268, n_269, n_270);
  xor g128 (n_271, A[20], B[20]);
  xor g129 (Z[20], n_267, n_271);
  nand g130 (n_273, A[21], B[21]);
  nand g131 (n_274, A[21], n_272);
  nand g132 (n_275, B[21], n_272);
  nand g133 (n_277, n_273, n_274, n_275);
  xor g134 (n_276, A[21], B[21]);
  xor g135 (Z[21], n_272, n_276);
  nand g136 (n_278, A[22], B[22]);
  nand g137 (n_279, A[22], n_277);
  nand g138 (n_280, B[22], n_277);
  nand g139 (n_282, n_278, n_279, n_280);
  xor g140 (n_281, A[22], B[22]);
  xor g141 (Z[22], n_277, n_281);
  nand g142 (n_283, A[23], B[23]);
  nand g143 (n_284, A[23], n_282);
  nand g144 (n_285, B[23], n_282);
  nand g145 (n_287, n_283, n_284, n_285);
  xor g146 (n_286, A[23], B[23]);
  xor g147 (Z[23], n_282, n_286);
  nand g148 (n_288, A[24], B[24]);
  nand g149 (n_289, A[24], n_287);
  nand g150 (n_290, B[24], n_287);
  nand g151 (n_292, n_288, n_289, n_290);
  xor g152 (n_291, A[24], B[24]);
  xor g153 (Z[24], n_287, n_291);
  nand g154 (n_293, A[25], B[25]);
  nand g155 (n_294, A[25], n_292);
  nand g156 (n_295, B[25], n_292);
  nand g157 (n_297, n_293, n_294, n_295);
  xor g158 (n_296, A[25], B[25]);
  xor g159 (Z[25], n_292, n_296);
  nand g160 (n_298, A[26], B[26]);
  nand g161 (n_299, A[26], n_297);
  nand g162 (n_300, B[26], n_297);
  nand g163 (n_302, n_298, n_299, n_300);
  xor g164 (n_301, A[26], B[26]);
  xor g165 (Z[26], n_297, n_301);
  nand g166 (n_303, A[27], B[27]);
  nand g167 (n_304, A[27], n_302);
  nand g168 (n_305, B[27], n_302);
  nand g169 (n_307, n_303, n_304, n_305);
  xor g170 (n_306, A[27], B[27]);
  xor g171 (Z[27], n_302, n_306);
  nand g172 (n_308, A[28], B[28]);
  nand g173 (n_309, A[28], n_307);
  nand g174 (n_310, B[28], n_307);
  nand g175 (n_312, n_308, n_309, n_310);
  xor g176 (n_311, A[28], B[28]);
  xor g177 (Z[28], n_307, n_311);
  nand g178 (n_313, A[29], B[29]);
  nand g179 (n_314, A[29], n_312);
  nand g180 (n_315, B[29], n_312);
  nand g181 (n_317, n_313, n_314, n_315);
  xor g182 (n_316, A[29], B[29]);
  xor g183 (Z[29], n_312, n_316);
  nand g184 (n_318, A[30], B[30]);
  nand g185 (n_319, A[30], n_317);
  nand g186 (n_320, B[30], n_317);
  nand g187 (n_322, n_318, n_319, n_320);
  xor g188 (n_321, A[30], B[30]);
  xor g189 (Z[30], n_317, n_321);
  nand g190 (n_323, A[31], B[31]);
  nand g191 (n_324, A[31], n_322);
  nand g192 (n_325, B[31], n_322);
  nand g193 (n_327, n_323, n_324, n_325);
  xor g194 (n_326, A[31], B[31]);
  xor g195 (Z[31], n_322, n_326);
  nand g196 (n_328, A[32], B[32]);
  nand g197 (n_329, A[32], n_327);
  nand g198 (n_330, B[32], n_327);
  nand g199 (n_332, n_328, n_329, n_330);
  xor g200 (n_331, A[32], B[32]);
  xor g201 (Z[32], n_327, n_331);
  nand g202 (n_333, A[33], B[33]);
  nand g203 (n_334, A[33], n_332);
  nand g204 (n_335, B[33], n_332);
  nand g205 (n_337, n_333, n_334, n_335);
  xor g206 (n_336, A[33], B[33]);
  xor g207 (Z[33], n_332, n_336);
  nand g208 (n_338, A[34], B[34]);
  nand g209 (n_339, A[34], n_337);
  nand g210 (n_340, B[34], n_337);
  nand g211 (n_342, n_338, n_339, n_340);
  xor g212 (n_341, A[34], B[34]);
  xor g213 (Z[34], n_337, n_341);
  nand g214 (n_343, A[35], B[35]);
  nand g215 (n_344, A[35], n_342);
  nand g216 (n_345, B[35], n_342);
  nand g217 (n_347, n_343, n_344, n_345);
  xor g218 (n_346, A[35], B[35]);
  xor g219 (Z[35], n_342, n_346);
  nand g220 (n_348, A[36], B[36]);
  nand g221 (n_349, A[36], n_347);
  nand g222 (n_350, B[36], n_347);
  nand g223 (n_352, n_348, n_349, n_350);
  xor g224 (n_351, A[36], B[36]);
  xor g225 (Z[36], n_347, n_351);
  nand g226 (n_353, A[37], B[37]);
  nand g227 (n_354, A[37], n_352);
  nand g228 (n_355, B[37], n_352);
  nand g229 (n_357, n_353, n_354, n_355);
  xor g230 (n_356, A[37], B[37]);
  xor g231 (Z[37], n_352, n_356);
  nand g232 (n_358, A[38], B[38]);
  nand g233 (n_359, A[38], n_357);
  nand g234 (n_360, B[38], n_357);
  nand g235 (n_362, n_358, n_359, n_360);
  xor g236 (n_361, A[38], B[38]);
  xor g237 (Z[38], n_357, n_361);
  nand g238 (n_363, A[39], B[39]);
  nand g239 (n_364, A[39], n_362);
  nand g240 (n_365, B[39], n_362);
  nand g241 (n_367, n_363, n_364, n_365);
  xor g242 (n_366, A[39], B[39]);
  xor g243 (Z[39], n_362, n_366);
  nand g244 (n_368, A[40], B[40]);
  nand g245 (n_369, A[40], n_367);
  nand g246 (n_370, B[40], n_367);
  nand g247 (n_372, n_368, n_369, n_370);
  xor g248 (n_371, A[40], B[40]);
  xor g249 (Z[40], n_367, n_371);
  nand g250 (n_373, A[41], B[41]);
  nand g251 (n_374, A[41], n_372);
  nand g252 (n_375, B[41], n_372);
  nand g253 (n_377, n_373, n_374, n_375);
  xor g254 (n_376, A[41], B[41]);
  xor g255 (Z[41], n_372, n_376);
  nand g256 (n_378, A[42], B[42]);
  nand g257 (n_379, A[42], n_377);
  nand g258 (n_380, B[42], n_377);
  nand g259 (n_382, n_378, n_379, n_380);
  xor g260 (n_381, A[42], B[42]);
  xor g261 (Z[42], n_377, n_381);
  nand g262 (n_383, A[43], B[43]);
  nand g263 (n_384, A[43], n_382);
  nand g264 (n_385, B[43], n_382);
  nand g265 (n_387, n_383, n_384, n_385);
  xor g266 (n_386, A[43], B[43]);
  xor g267 (Z[43], n_382, n_386);
  nand g268 (n_388, A[44], B[44]);
  nand g269 (n_389, A[44], n_387);
  nand g270 (n_390, B[44], n_387);
  nand g271 (n_392, n_388, n_389, n_390);
  xor g272 (n_391, A[44], B[44]);
  xor g273 (Z[44], n_387, n_391);
  nand g274 (n_393, A[45], B[45]);
  nand g275 (n_394, A[45], n_392);
  nand g276 (n_395, B[45], n_392);
  nand g277 (n_397, n_393, n_394, n_395);
  xor g278 (n_396, A[45], B[45]);
  xor g279 (Z[45], n_392, n_396);
  nand g280 (n_398, A[46], B[46]);
  nand g281 (n_399, A[46], n_397);
  nand g282 (n_400, B[46], n_397);
  nand g283 (n_402, n_398, n_399, n_400);
  xor g284 (n_401, A[46], B[46]);
  xor g285 (Z[46], n_397, n_401);
  nand g286 (n_403, A[47], B[47]);
  nand g287 (n_404, A[47], n_402);
  nand g288 (n_405, B[47], n_402);
  nand g289 (n_407, n_403, n_404, n_405);
  xor g290 (n_406, A[47], B[47]);
  xor g291 (Z[47], n_402, n_406);
  nand g292 (n_408, A[48], B[48]);
  nand g293 (n_409, A[48], n_407);
  nand g294 (n_410, B[48], n_407);
  nand g295 (n_412, n_408, n_409, n_410);
  xor g296 (n_411, A[48], B[48]);
  xor g297 (Z[48], n_407, n_411);
  nand g298 (n_413, A[49], B[49]);
  nand g299 (n_414, A[49], n_412);
  nand g300 (n_415, B[49], n_412);
  nand g301 (n_417, n_413, n_414, n_415);
  xor g302 (n_416, A[49], B[49]);
  xor g303 (Z[49], n_412, n_416);
  nand g304 (n_418, A[50], B[50]);
  nand g305 (n_419, A[50], n_417);
  nand g306 (n_420, B[50], n_417);
  nand g307 (n_422, n_418, n_419, n_420);
  xor g308 (n_421, A[50], B[50]);
  xor g309 (Z[50], n_417, n_421);
  nand g310 (n_423, A[51], B[51]);
  nand g311 (n_424, A[51], n_422);
  nand g312 (n_425, B[51], n_422);
  nand g313 (n_427, n_423, n_424, n_425);
  xor g314 (n_426, A[51], B[51]);
  xor g315 (Z[51], n_422, n_426);
  nand g316 (n_428, A[52], B[52]);
  nand g317 (n_429, A[52], n_427);
  nand g318 (n_430, B[52], n_427);
  nand g319 (n_432, n_428, n_429, n_430);
  xor g320 (n_431, A[52], B[52]);
  xor g321 (Z[52], n_427, n_431);
  nand g325 (n_167, n_433, n_434, n_435);
  xor g327 (Z[53], n_432, n_436);
  or g329 (n_433, A[53], B[53]);
  xor g330 (n_436, A[53], B[53]);
  or g331 (n_174, wc, n_168);
  not gc (wc, A[1]);
  or g332 (n_175, wc0, n_168);
  not gc0 (wc0, B[1]);
  xnor g333 (Z[1], n_168, n_176);
  or g334 (n_434, A[53], wc1);
  not gc1 (wc1, n_432);
  or g335 (n_435, B[53], wc2);
  not gc2 (wc2, n_432);
endmodule

module add_signed_6294_1_GENERIC(A, B, Z);
  input [53:0] A, B;
  output [54:0] Z;
  wire [53:0] A, B;
  wire [54:0] Z;
  add_signed_6294_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_6784_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [52:0] A, B;
  output [53:0] Z;
  wire [52:0] A, B;
  wire [53:0] Z;
  wire n_164, n_165, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367;
  wire n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428;
  not g3 (Z[53], n_164);
  nand g4 (n_165, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_170, A[1], B[1]);
  nand g13 (n_174, n_170, n_171, n_172);
  xor g14 (n_173, A[1], B[1]);
  nand g16 (n_175, A[2], B[2]);
  nand g17 (n_176, A[2], n_174);
  nand g18 (n_177, B[2], n_174);
  nand g19 (n_179, n_175, n_176, n_177);
  xor g20 (n_178, A[2], B[2]);
  xor g21 (Z[2], n_174, n_178);
  nand g22 (n_180, A[3], B[3]);
  nand g23 (n_181, A[3], n_179);
  nand g24 (n_182, B[3], n_179);
  nand g25 (n_184, n_180, n_181, n_182);
  xor g26 (n_183, A[3], B[3]);
  xor g27 (Z[3], n_179, n_183);
  nand g28 (n_185, A[4], B[4]);
  nand g29 (n_186, A[4], n_184);
  nand g30 (n_187, B[4], n_184);
  nand g31 (n_189, n_185, n_186, n_187);
  xor g32 (n_188, A[4], B[4]);
  xor g33 (Z[4], n_184, n_188);
  nand g34 (n_190, A[5], B[5]);
  nand g35 (n_191, A[5], n_189);
  nand g36 (n_192, B[5], n_189);
  nand g37 (n_194, n_190, n_191, n_192);
  xor g38 (n_193, A[5], B[5]);
  xor g39 (Z[5], n_189, n_193);
  nand g40 (n_195, A[6], B[6]);
  nand g41 (n_196, A[6], n_194);
  nand g42 (n_197, B[6], n_194);
  nand g43 (n_199, n_195, n_196, n_197);
  xor g44 (n_198, A[6], B[6]);
  xor g45 (Z[6], n_194, n_198);
  nand g46 (n_200, A[7], B[7]);
  nand g47 (n_201, A[7], n_199);
  nand g48 (n_202, B[7], n_199);
  nand g49 (n_204, n_200, n_201, n_202);
  xor g50 (n_203, A[7], B[7]);
  xor g51 (Z[7], n_199, n_203);
  nand g52 (n_205, A[8], B[8]);
  nand g53 (n_206, A[8], n_204);
  nand g54 (n_207, B[8], n_204);
  nand g55 (n_209, n_205, n_206, n_207);
  xor g56 (n_208, A[8], B[8]);
  xor g57 (Z[8], n_204, n_208);
  nand g58 (n_210, A[9], B[9]);
  nand g59 (n_211, A[9], n_209);
  nand g60 (n_212, B[9], n_209);
  nand g61 (n_214, n_210, n_211, n_212);
  xor g62 (n_213, A[9], B[9]);
  xor g63 (Z[9], n_209, n_213);
  nand g64 (n_215, A[10], B[10]);
  nand g65 (n_216, A[10], n_214);
  nand g66 (n_217, B[10], n_214);
  nand g67 (n_219, n_215, n_216, n_217);
  xor g68 (n_218, A[10], B[10]);
  xor g69 (Z[10], n_214, n_218);
  nand g70 (n_220, A[11], B[11]);
  nand g71 (n_221, A[11], n_219);
  nand g72 (n_222, B[11], n_219);
  nand g73 (n_224, n_220, n_221, n_222);
  xor g74 (n_223, A[11], B[11]);
  xor g75 (Z[11], n_219, n_223);
  nand g76 (n_225, A[12], B[12]);
  nand g77 (n_226, A[12], n_224);
  nand g78 (n_227, B[12], n_224);
  nand g79 (n_229, n_225, n_226, n_227);
  xor g80 (n_228, A[12], B[12]);
  xor g81 (Z[12], n_224, n_228);
  nand g82 (n_230, A[13], B[13]);
  nand g83 (n_231, A[13], n_229);
  nand g84 (n_232, B[13], n_229);
  nand g85 (n_234, n_230, n_231, n_232);
  xor g86 (n_233, A[13], B[13]);
  xor g87 (Z[13], n_229, n_233);
  nand g88 (n_235, A[14], B[14]);
  nand g89 (n_236, A[14], n_234);
  nand g90 (n_237, B[14], n_234);
  nand g91 (n_239, n_235, n_236, n_237);
  xor g92 (n_238, A[14], B[14]);
  xor g93 (Z[14], n_234, n_238);
  nand g94 (n_240, A[15], B[15]);
  nand g95 (n_241, A[15], n_239);
  nand g96 (n_242, B[15], n_239);
  nand g97 (n_244, n_240, n_241, n_242);
  xor g98 (n_243, A[15], B[15]);
  xor g99 (Z[15], n_239, n_243);
  nand g100 (n_245, A[16], B[16]);
  nand g101 (n_246, A[16], n_244);
  nand g102 (n_247, B[16], n_244);
  nand g103 (n_249, n_245, n_246, n_247);
  xor g104 (n_248, A[16], B[16]);
  xor g105 (Z[16], n_244, n_248);
  nand g106 (n_250, A[17], B[17]);
  nand g107 (n_251, A[17], n_249);
  nand g108 (n_252, B[17], n_249);
  nand g109 (n_254, n_250, n_251, n_252);
  xor g110 (n_253, A[17], B[17]);
  xor g111 (Z[17], n_249, n_253);
  nand g112 (n_255, A[18], B[18]);
  nand g113 (n_256, A[18], n_254);
  nand g114 (n_257, B[18], n_254);
  nand g115 (n_259, n_255, n_256, n_257);
  xor g116 (n_258, A[18], B[18]);
  xor g117 (Z[18], n_254, n_258);
  nand g118 (n_260, A[19], B[19]);
  nand g119 (n_261, A[19], n_259);
  nand g120 (n_262, B[19], n_259);
  nand g121 (n_264, n_260, n_261, n_262);
  xor g122 (n_263, A[19], B[19]);
  xor g123 (Z[19], n_259, n_263);
  nand g124 (n_265, A[20], B[20]);
  nand g125 (n_266, A[20], n_264);
  nand g126 (n_267, B[20], n_264);
  nand g127 (n_269, n_265, n_266, n_267);
  xor g128 (n_268, A[20], B[20]);
  xor g129 (Z[20], n_264, n_268);
  nand g130 (n_270, A[21], B[21]);
  nand g131 (n_271, A[21], n_269);
  nand g132 (n_272, B[21], n_269);
  nand g133 (n_274, n_270, n_271, n_272);
  xor g134 (n_273, A[21], B[21]);
  xor g135 (Z[21], n_269, n_273);
  nand g136 (n_275, A[22], B[22]);
  nand g137 (n_276, A[22], n_274);
  nand g138 (n_277, B[22], n_274);
  nand g139 (n_279, n_275, n_276, n_277);
  xor g140 (n_278, A[22], B[22]);
  xor g141 (Z[22], n_274, n_278);
  nand g142 (n_280, A[23], B[23]);
  nand g143 (n_281, A[23], n_279);
  nand g144 (n_282, B[23], n_279);
  nand g145 (n_284, n_280, n_281, n_282);
  xor g146 (n_283, A[23], B[23]);
  xor g147 (Z[23], n_279, n_283);
  nand g148 (n_285, A[24], B[24]);
  nand g149 (n_286, A[24], n_284);
  nand g150 (n_287, B[24], n_284);
  nand g151 (n_289, n_285, n_286, n_287);
  xor g152 (n_288, A[24], B[24]);
  xor g153 (Z[24], n_284, n_288);
  nand g154 (n_290, A[25], B[25]);
  nand g155 (n_291, A[25], n_289);
  nand g156 (n_292, B[25], n_289);
  nand g157 (n_294, n_290, n_291, n_292);
  xor g158 (n_293, A[25], B[25]);
  xor g159 (Z[25], n_289, n_293);
  nand g160 (n_295, A[26], B[26]);
  nand g161 (n_296, A[26], n_294);
  nand g162 (n_297, B[26], n_294);
  nand g163 (n_299, n_295, n_296, n_297);
  xor g164 (n_298, A[26], B[26]);
  xor g165 (Z[26], n_294, n_298);
  nand g166 (n_300, A[27], B[27]);
  nand g167 (n_301, A[27], n_299);
  nand g168 (n_302, B[27], n_299);
  nand g169 (n_304, n_300, n_301, n_302);
  xor g170 (n_303, A[27], B[27]);
  xor g171 (Z[27], n_299, n_303);
  nand g172 (n_305, A[28], B[28]);
  nand g173 (n_306, A[28], n_304);
  nand g174 (n_307, B[28], n_304);
  nand g175 (n_309, n_305, n_306, n_307);
  xor g176 (n_308, A[28], B[28]);
  xor g177 (Z[28], n_304, n_308);
  nand g178 (n_310, A[29], B[29]);
  nand g179 (n_311, A[29], n_309);
  nand g180 (n_312, B[29], n_309);
  nand g181 (n_314, n_310, n_311, n_312);
  xor g182 (n_313, A[29], B[29]);
  xor g183 (Z[29], n_309, n_313);
  nand g184 (n_315, A[30], B[30]);
  nand g185 (n_316, A[30], n_314);
  nand g186 (n_317, B[30], n_314);
  nand g187 (n_319, n_315, n_316, n_317);
  xor g188 (n_318, A[30], B[30]);
  xor g189 (Z[30], n_314, n_318);
  nand g190 (n_320, A[31], B[31]);
  nand g191 (n_321, A[31], n_319);
  nand g192 (n_322, B[31], n_319);
  nand g193 (n_324, n_320, n_321, n_322);
  xor g194 (n_323, A[31], B[31]);
  xor g195 (Z[31], n_319, n_323);
  nand g196 (n_325, A[32], B[32]);
  nand g197 (n_326, A[32], n_324);
  nand g198 (n_327, B[32], n_324);
  nand g199 (n_329, n_325, n_326, n_327);
  xor g200 (n_328, A[32], B[32]);
  xor g201 (Z[32], n_324, n_328);
  nand g202 (n_330, A[33], B[33]);
  nand g203 (n_331, A[33], n_329);
  nand g204 (n_332, B[33], n_329);
  nand g205 (n_334, n_330, n_331, n_332);
  xor g206 (n_333, A[33], B[33]);
  xor g207 (Z[33], n_329, n_333);
  nand g208 (n_335, A[34], B[34]);
  nand g209 (n_336, A[34], n_334);
  nand g210 (n_337, B[34], n_334);
  nand g211 (n_339, n_335, n_336, n_337);
  xor g212 (n_338, A[34], B[34]);
  xor g213 (Z[34], n_334, n_338);
  nand g214 (n_340, A[35], B[35]);
  nand g215 (n_341, A[35], n_339);
  nand g216 (n_342, B[35], n_339);
  nand g217 (n_344, n_340, n_341, n_342);
  xor g218 (n_343, A[35], B[35]);
  xor g219 (Z[35], n_339, n_343);
  nand g220 (n_345, A[36], B[36]);
  nand g221 (n_346, A[36], n_344);
  nand g222 (n_347, B[36], n_344);
  nand g223 (n_349, n_345, n_346, n_347);
  xor g224 (n_348, A[36], B[36]);
  xor g225 (Z[36], n_344, n_348);
  nand g226 (n_350, A[37], B[37]);
  nand g227 (n_351, A[37], n_349);
  nand g228 (n_352, B[37], n_349);
  nand g229 (n_354, n_350, n_351, n_352);
  xor g230 (n_353, A[37], B[37]);
  xor g231 (Z[37], n_349, n_353);
  nand g232 (n_355, A[38], B[38]);
  nand g233 (n_356, A[38], n_354);
  nand g234 (n_357, B[38], n_354);
  nand g235 (n_359, n_355, n_356, n_357);
  xor g236 (n_358, A[38], B[38]);
  xor g237 (Z[38], n_354, n_358);
  nand g238 (n_360, A[39], B[39]);
  nand g239 (n_361, A[39], n_359);
  nand g240 (n_362, B[39], n_359);
  nand g241 (n_364, n_360, n_361, n_362);
  xor g242 (n_363, A[39], B[39]);
  xor g243 (Z[39], n_359, n_363);
  nand g244 (n_365, A[40], B[40]);
  nand g245 (n_366, A[40], n_364);
  nand g246 (n_367, B[40], n_364);
  nand g247 (n_369, n_365, n_366, n_367);
  xor g248 (n_368, A[40], B[40]);
  xor g249 (Z[40], n_364, n_368);
  nand g250 (n_370, A[41], B[41]);
  nand g251 (n_371, A[41], n_369);
  nand g252 (n_372, B[41], n_369);
  nand g253 (n_374, n_370, n_371, n_372);
  xor g254 (n_373, A[41], B[41]);
  xor g255 (Z[41], n_369, n_373);
  nand g256 (n_375, A[42], B[42]);
  nand g257 (n_376, A[42], n_374);
  nand g258 (n_377, B[42], n_374);
  nand g259 (n_379, n_375, n_376, n_377);
  xor g260 (n_378, A[42], B[42]);
  xor g261 (Z[42], n_374, n_378);
  nand g262 (n_380, A[43], B[43]);
  nand g263 (n_381, A[43], n_379);
  nand g264 (n_382, B[43], n_379);
  nand g265 (n_384, n_380, n_381, n_382);
  xor g266 (n_383, A[43], B[43]);
  xor g267 (Z[43], n_379, n_383);
  nand g268 (n_385, A[44], B[44]);
  nand g269 (n_386, A[44], n_384);
  nand g270 (n_387, B[44], n_384);
  nand g271 (n_389, n_385, n_386, n_387);
  xor g272 (n_388, A[44], B[44]);
  xor g273 (Z[44], n_384, n_388);
  nand g274 (n_390, A[45], B[45]);
  nand g275 (n_391, A[45], n_389);
  nand g276 (n_392, B[45], n_389);
  nand g277 (n_394, n_390, n_391, n_392);
  xor g278 (n_393, A[45], B[45]);
  xor g279 (Z[45], n_389, n_393);
  nand g280 (n_395, A[46], B[46]);
  nand g281 (n_396, A[46], n_394);
  nand g282 (n_397, B[46], n_394);
  nand g283 (n_399, n_395, n_396, n_397);
  xor g284 (n_398, A[46], B[46]);
  xor g285 (Z[46], n_394, n_398);
  nand g286 (n_400, A[47], B[47]);
  nand g287 (n_401, A[47], n_399);
  nand g288 (n_402, B[47], n_399);
  nand g289 (n_404, n_400, n_401, n_402);
  xor g290 (n_403, A[47], B[47]);
  xor g291 (Z[47], n_399, n_403);
  nand g292 (n_405, A[48], B[48]);
  nand g293 (n_406, A[48], n_404);
  nand g294 (n_407, B[48], n_404);
  nand g295 (n_409, n_405, n_406, n_407);
  xor g296 (n_408, A[48], B[48]);
  xor g297 (Z[48], n_404, n_408);
  nand g298 (n_410, A[49], B[49]);
  nand g299 (n_411, A[49], n_409);
  nand g300 (n_412, B[49], n_409);
  nand g301 (n_414, n_410, n_411, n_412);
  xor g302 (n_413, A[49], B[49]);
  xor g303 (Z[49], n_409, n_413);
  nand g304 (n_415, A[50], B[50]);
  nand g305 (n_416, A[50], n_414);
  nand g306 (n_417, B[50], n_414);
  nand g307 (n_419, n_415, n_416, n_417);
  xor g308 (n_418, A[50], B[50]);
  xor g309 (Z[50], n_414, n_418);
  nand g310 (n_420, A[51], B[51]);
  nand g311 (n_421, A[51], n_419);
  nand g312 (n_422, B[51], n_419);
  nand g313 (n_424, n_420, n_421, n_422);
  xor g314 (n_423, A[51], B[51]);
  xor g315 (Z[51], n_419, n_423);
  nand g319 (n_164, n_425, n_426, n_427);
  xor g321 (Z[52], n_424, n_428);
  or g323 (n_425, A[52], B[52]);
  xor g324 (n_428, A[52], B[52]);
  or g325 (n_171, wc, n_165);
  not gc (wc, A[1]);
  or g326 (n_172, wc0, n_165);
  not gc0 (wc0, B[1]);
  xnor g327 (Z[1], n_165, n_173);
  or g328 (n_426, A[52], wc1);
  not gc1 (wc1, n_424);
  or g329 (n_427, B[52], wc2);
  not gc2 (wc2, n_424);
endmodule

module add_signed_6784_GENERIC(A, B, Z);
  input [52:0] A, B;
  output [53:0] Z;
  wire [52:0] A, B;
  wire [53:0] Z;
  add_signed_6784_GENERIC_REAL g1(.A ({A[52:2], A[0], A[0]}), .B (B),
       .Z (Z));
endmodule

module add_signed_6784_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [52:0] A, B;
  output [53:0] Z;
  wire [52:0] A, B;
  wire [53:0] Z;
  wire n_164, n_165, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367;
  wire n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428;
  not g3 (Z[53], n_164);
  nand g4 (n_165, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_170, A[1], B[1]);
  nand g13 (n_174, n_170, n_171, n_172);
  xor g14 (n_173, A[1], B[1]);
  nand g16 (n_175, A[2], B[2]);
  nand g17 (n_176, A[2], n_174);
  nand g18 (n_177, B[2], n_174);
  nand g19 (n_179, n_175, n_176, n_177);
  xor g20 (n_178, A[2], B[2]);
  xor g21 (Z[2], n_174, n_178);
  nand g22 (n_180, A[3], B[3]);
  nand g23 (n_181, A[3], n_179);
  nand g24 (n_182, B[3], n_179);
  nand g25 (n_184, n_180, n_181, n_182);
  xor g26 (n_183, A[3], B[3]);
  xor g27 (Z[3], n_179, n_183);
  nand g28 (n_185, A[4], B[4]);
  nand g29 (n_186, A[4], n_184);
  nand g30 (n_187, B[4], n_184);
  nand g31 (n_189, n_185, n_186, n_187);
  xor g32 (n_188, A[4], B[4]);
  xor g33 (Z[4], n_184, n_188);
  nand g34 (n_190, A[5], B[5]);
  nand g35 (n_191, A[5], n_189);
  nand g36 (n_192, B[5], n_189);
  nand g37 (n_194, n_190, n_191, n_192);
  xor g38 (n_193, A[5], B[5]);
  xor g39 (Z[5], n_189, n_193);
  nand g40 (n_195, A[6], B[6]);
  nand g41 (n_196, A[6], n_194);
  nand g42 (n_197, B[6], n_194);
  nand g43 (n_199, n_195, n_196, n_197);
  xor g44 (n_198, A[6], B[6]);
  xor g45 (Z[6], n_194, n_198);
  nand g46 (n_200, A[7], B[7]);
  nand g47 (n_201, A[7], n_199);
  nand g48 (n_202, B[7], n_199);
  nand g49 (n_204, n_200, n_201, n_202);
  xor g50 (n_203, A[7], B[7]);
  xor g51 (Z[7], n_199, n_203);
  nand g52 (n_205, A[8], B[8]);
  nand g53 (n_206, A[8], n_204);
  nand g54 (n_207, B[8], n_204);
  nand g55 (n_209, n_205, n_206, n_207);
  xor g56 (n_208, A[8], B[8]);
  xor g57 (Z[8], n_204, n_208);
  nand g58 (n_210, A[9], B[9]);
  nand g59 (n_211, A[9], n_209);
  nand g60 (n_212, B[9], n_209);
  nand g61 (n_214, n_210, n_211, n_212);
  xor g62 (n_213, A[9], B[9]);
  xor g63 (Z[9], n_209, n_213);
  nand g64 (n_215, A[10], B[10]);
  nand g65 (n_216, A[10], n_214);
  nand g66 (n_217, B[10], n_214);
  nand g67 (n_219, n_215, n_216, n_217);
  xor g68 (n_218, A[10], B[10]);
  xor g69 (Z[10], n_214, n_218);
  nand g70 (n_220, A[11], B[11]);
  nand g71 (n_221, A[11], n_219);
  nand g72 (n_222, B[11], n_219);
  nand g73 (n_224, n_220, n_221, n_222);
  xor g74 (n_223, A[11], B[11]);
  xor g75 (Z[11], n_219, n_223);
  nand g76 (n_225, A[12], B[12]);
  nand g77 (n_226, A[12], n_224);
  nand g78 (n_227, B[12], n_224);
  nand g79 (n_229, n_225, n_226, n_227);
  xor g80 (n_228, A[12], B[12]);
  xor g81 (Z[12], n_224, n_228);
  nand g82 (n_230, A[13], B[13]);
  nand g83 (n_231, A[13], n_229);
  nand g84 (n_232, B[13], n_229);
  nand g85 (n_234, n_230, n_231, n_232);
  xor g86 (n_233, A[13], B[13]);
  xor g87 (Z[13], n_229, n_233);
  nand g88 (n_235, A[14], B[14]);
  nand g89 (n_236, A[14], n_234);
  nand g90 (n_237, B[14], n_234);
  nand g91 (n_239, n_235, n_236, n_237);
  xor g92 (n_238, A[14], B[14]);
  xor g93 (Z[14], n_234, n_238);
  nand g94 (n_240, A[15], B[15]);
  nand g95 (n_241, A[15], n_239);
  nand g96 (n_242, B[15], n_239);
  nand g97 (n_244, n_240, n_241, n_242);
  xor g98 (n_243, A[15], B[15]);
  xor g99 (Z[15], n_239, n_243);
  nand g100 (n_245, A[16], B[16]);
  nand g101 (n_246, A[16], n_244);
  nand g102 (n_247, B[16], n_244);
  nand g103 (n_249, n_245, n_246, n_247);
  xor g104 (n_248, A[16], B[16]);
  xor g105 (Z[16], n_244, n_248);
  nand g106 (n_250, A[17], B[17]);
  nand g107 (n_251, A[17], n_249);
  nand g108 (n_252, B[17], n_249);
  nand g109 (n_254, n_250, n_251, n_252);
  xor g110 (n_253, A[17], B[17]);
  xor g111 (Z[17], n_249, n_253);
  nand g112 (n_255, A[18], B[18]);
  nand g113 (n_256, A[18], n_254);
  nand g114 (n_257, B[18], n_254);
  nand g115 (n_259, n_255, n_256, n_257);
  xor g116 (n_258, A[18], B[18]);
  xor g117 (Z[18], n_254, n_258);
  nand g118 (n_260, A[19], B[19]);
  nand g119 (n_261, A[19], n_259);
  nand g120 (n_262, B[19], n_259);
  nand g121 (n_264, n_260, n_261, n_262);
  xor g122 (n_263, A[19], B[19]);
  xor g123 (Z[19], n_259, n_263);
  nand g124 (n_265, A[20], B[20]);
  nand g125 (n_266, A[20], n_264);
  nand g126 (n_267, B[20], n_264);
  nand g127 (n_269, n_265, n_266, n_267);
  xor g128 (n_268, A[20], B[20]);
  xor g129 (Z[20], n_264, n_268);
  nand g130 (n_270, A[21], B[21]);
  nand g131 (n_271, A[21], n_269);
  nand g132 (n_272, B[21], n_269);
  nand g133 (n_274, n_270, n_271, n_272);
  xor g134 (n_273, A[21], B[21]);
  xor g135 (Z[21], n_269, n_273);
  nand g136 (n_275, A[22], B[22]);
  nand g137 (n_276, A[22], n_274);
  nand g138 (n_277, B[22], n_274);
  nand g139 (n_279, n_275, n_276, n_277);
  xor g140 (n_278, A[22], B[22]);
  xor g141 (Z[22], n_274, n_278);
  nand g142 (n_280, A[23], B[23]);
  nand g143 (n_281, A[23], n_279);
  nand g144 (n_282, B[23], n_279);
  nand g145 (n_284, n_280, n_281, n_282);
  xor g146 (n_283, A[23], B[23]);
  xor g147 (Z[23], n_279, n_283);
  nand g148 (n_285, A[24], B[24]);
  nand g149 (n_286, A[24], n_284);
  nand g150 (n_287, B[24], n_284);
  nand g151 (n_289, n_285, n_286, n_287);
  xor g152 (n_288, A[24], B[24]);
  xor g153 (Z[24], n_284, n_288);
  nand g154 (n_290, A[25], B[25]);
  nand g155 (n_291, A[25], n_289);
  nand g156 (n_292, B[25], n_289);
  nand g157 (n_294, n_290, n_291, n_292);
  xor g158 (n_293, A[25], B[25]);
  xor g159 (Z[25], n_289, n_293);
  nand g160 (n_295, A[26], B[26]);
  nand g161 (n_296, A[26], n_294);
  nand g162 (n_297, B[26], n_294);
  nand g163 (n_299, n_295, n_296, n_297);
  xor g164 (n_298, A[26], B[26]);
  xor g165 (Z[26], n_294, n_298);
  nand g166 (n_300, A[27], B[27]);
  nand g167 (n_301, A[27], n_299);
  nand g168 (n_302, B[27], n_299);
  nand g169 (n_304, n_300, n_301, n_302);
  xor g170 (n_303, A[27], B[27]);
  xor g171 (Z[27], n_299, n_303);
  nand g172 (n_305, A[28], B[28]);
  nand g173 (n_306, A[28], n_304);
  nand g174 (n_307, B[28], n_304);
  nand g175 (n_309, n_305, n_306, n_307);
  xor g176 (n_308, A[28], B[28]);
  xor g177 (Z[28], n_304, n_308);
  nand g178 (n_310, A[29], B[29]);
  nand g179 (n_311, A[29], n_309);
  nand g180 (n_312, B[29], n_309);
  nand g181 (n_314, n_310, n_311, n_312);
  xor g182 (n_313, A[29], B[29]);
  xor g183 (Z[29], n_309, n_313);
  nand g184 (n_315, A[30], B[30]);
  nand g185 (n_316, A[30], n_314);
  nand g186 (n_317, B[30], n_314);
  nand g187 (n_319, n_315, n_316, n_317);
  xor g188 (n_318, A[30], B[30]);
  xor g189 (Z[30], n_314, n_318);
  nand g190 (n_320, A[31], B[31]);
  nand g191 (n_321, A[31], n_319);
  nand g192 (n_322, B[31], n_319);
  nand g193 (n_324, n_320, n_321, n_322);
  xor g194 (n_323, A[31], B[31]);
  xor g195 (Z[31], n_319, n_323);
  nand g196 (n_325, A[32], B[32]);
  nand g197 (n_326, A[32], n_324);
  nand g198 (n_327, B[32], n_324);
  nand g199 (n_329, n_325, n_326, n_327);
  xor g200 (n_328, A[32], B[32]);
  xor g201 (Z[32], n_324, n_328);
  nand g202 (n_330, A[33], B[33]);
  nand g203 (n_331, A[33], n_329);
  nand g204 (n_332, B[33], n_329);
  nand g205 (n_334, n_330, n_331, n_332);
  xor g206 (n_333, A[33], B[33]);
  xor g207 (Z[33], n_329, n_333);
  nand g208 (n_335, A[34], B[34]);
  nand g209 (n_336, A[34], n_334);
  nand g210 (n_337, B[34], n_334);
  nand g211 (n_339, n_335, n_336, n_337);
  xor g212 (n_338, A[34], B[34]);
  xor g213 (Z[34], n_334, n_338);
  nand g214 (n_340, A[35], B[35]);
  nand g215 (n_341, A[35], n_339);
  nand g216 (n_342, B[35], n_339);
  nand g217 (n_344, n_340, n_341, n_342);
  xor g218 (n_343, A[35], B[35]);
  xor g219 (Z[35], n_339, n_343);
  nand g220 (n_345, A[36], B[36]);
  nand g221 (n_346, A[36], n_344);
  nand g222 (n_347, B[36], n_344);
  nand g223 (n_349, n_345, n_346, n_347);
  xor g224 (n_348, A[36], B[36]);
  xor g225 (Z[36], n_344, n_348);
  nand g226 (n_350, A[37], B[37]);
  nand g227 (n_351, A[37], n_349);
  nand g228 (n_352, B[37], n_349);
  nand g229 (n_354, n_350, n_351, n_352);
  xor g230 (n_353, A[37], B[37]);
  xor g231 (Z[37], n_349, n_353);
  nand g232 (n_355, A[38], B[38]);
  nand g233 (n_356, A[38], n_354);
  nand g234 (n_357, B[38], n_354);
  nand g235 (n_359, n_355, n_356, n_357);
  xor g236 (n_358, A[38], B[38]);
  xor g237 (Z[38], n_354, n_358);
  nand g238 (n_360, A[39], B[39]);
  nand g239 (n_361, A[39], n_359);
  nand g240 (n_362, B[39], n_359);
  nand g241 (n_364, n_360, n_361, n_362);
  xor g242 (n_363, A[39], B[39]);
  xor g243 (Z[39], n_359, n_363);
  nand g244 (n_365, A[40], B[40]);
  nand g245 (n_366, A[40], n_364);
  nand g246 (n_367, B[40], n_364);
  nand g247 (n_369, n_365, n_366, n_367);
  xor g248 (n_368, A[40], B[40]);
  xor g249 (Z[40], n_364, n_368);
  nand g250 (n_370, A[41], B[41]);
  nand g251 (n_371, A[41], n_369);
  nand g252 (n_372, B[41], n_369);
  nand g253 (n_374, n_370, n_371, n_372);
  xor g254 (n_373, A[41], B[41]);
  xor g255 (Z[41], n_369, n_373);
  nand g256 (n_375, A[42], B[42]);
  nand g257 (n_376, A[42], n_374);
  nand g258 (n_377, B[42], n_374);
  nand g259 (n_379, n_375, n_376, n_377);
  xor g260 (n_378, A[42], B[42]);
  xor g261 (Z[42], n_374, n_378);
  nand g262 (n_380, A[43], B[43]);
  nand g263 (n_381, A[43], n_379);
  nand g264 (n_382, B[43], n_379);
  nand g265 (n_384, n_380, n_381, n_382);
  xor g266 (n_383, A[43], B[43]);
  xor g267 (Z[43], n_379, n_383);
  nand g268 (n_385, A[44], B[44]);
  nand g269 (n_386, A[44], n_384);
  nand g270 (n_387, B[44], n_384);
  nand g271 (n_389, n_385, n_386, n_387);
  xor g272 (n_388, A[44], B[44]);
  xor g273 (Z[44], n_384, n_388);
  nand g274 (n_390, A[45], B[45]);
  nand g275 (n_391, A[45], n_389);
  nand g276 (n_392, B[45], n_389);
  nand g277 (n_394, n_390, n_391, n_392);
  xor g278 (n_393, A[45], B[45]);
  xor g279 (Z[45], n_389, n_393);
  nand g280 (n_395, A[46], B[46]);
  nand g281 (n_396, A[46], n_394);
  nand g282 (n_397, B[46], n_394);
  nand g283 (n_399, n_395, n_396, n_397);
  xor g284 (n_398, A[46], B[46]);
  xor g285 (Z[46], n_394, n_398);
  nand g286 (n_400, A[47], B[47]);
  nand g287 (n_401, A[47], n_399);
  nand g288 (n_402, B[47], n_399);
  nand g289 (n_404, n_400, n_401, n_402);
  xor g290 (n_403, A[47], B[47]);
  xor g291 (Z[47], n_399, n_403);
  nand g292 (n_405, A[48], B[48]);
  nand g293 (n_406, A[48], n_404);
  nand g294 (n_407, B[48], n_404);
  nand g295 (n_409, n_405, n_406, n_407);
  xor g296 (n_408, A[48], B[48]);
  xor g297 (Z[48], n_404, n_408);
  nand g298 (n_410, A[49], B[49]);
  nand g299 (n_411, A[49], n_409);
  nand g300 (n_412, B[49], n_409);
  nand g301 (n_414, n_410, n_411, n_412);
  xor g302 (n_413, A[49], B[49]);
  xor g303 (Z[49], n_409, n_413);
  nand g304 (n_415, A[50], B[50]);
  nand g305 (n_416, A[50], n_414);
  nand g306 (n_417, B[50], n_414);
  nand g307 (n_419, n_415, n_416, n_417);
  xor g308 (n_418, A[50], B[50]);
  xor g309 (Z[50], n_414, n_418);
  nand g310 (n_420, A[51], B[51]);
  nand g311 (n_421, A[51], n_419);
  nand g312 (n_422, B[51], n_419);
  nand g313 (n_424, n_420, n_421, n_422);
  xor g314 (n_423, A[51], B[51]);
  xor g315 (Z[51], n_419, n_423);
  nand g319 (n_164, n_425, n_426, n_427);
  xor g321 (Z[52], n_424, n_428);
  or g323 (n_425, A[52], B[52]);
  xor g324 (n_428, A[52], B[52]);
  or g325 (n_171, wc, n_165);
  not gc (wc, A[1]);
  or g326 (n_172, wc0, n_165);
  not gc0 (wc0, B[1]);
  xnor g327 (Z[1], n_165, n_173);
  or g328 (n_426, A[52], wc1);
  not gc1 (wc1, n_424);
  or g329 (n_427, B[52], wc2);
  not gc2 (wc2, n_424);
endmodule

module add_signed_6784_1_GENERIC(A, B, Z);
  input [52:0] A, B;
  output [53:0] Z;
  wire [52:0] A, B;
  wire [53:0] Z;
  add_signed_6784_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_7256_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [50:0] A, B;
  output [51:0] Z;
  wire [50:0] A, B;
  wire [51:0] Z;
  wire n_158, n_159, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412;
  not g3 (Z[51], n_158);
  nand g4 (n_159, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_164, A[1], B[1]);
  nand g13 (n_168, n_164, n_165, n_166);
  xor g14 (n_167, A[1], B[1]);
  nand g16 (n_169, A[2], B[2]);
  nand g17 (n_170, A[2], n_168);
  nand g18 (n_171, B[2], n_168);
  nand g19 (n_173, n_169, n_170, n_171);
  xor g20 (n_172, A[2], B[2]);
  xor g21 (Z[2], n_168, n_172);
  nand g22 (n_174, A[3], B[3]);
  nand g23 (n_175, A[3], n_173);
  nand g24 (n_176, B[3], n_173);
  nand g25 (n_178, n_174, n_175, n_176);
  xor g26 (n_177, A[3], B[3]);
  xor g27 (Z[3], n_173, n_177);
  nand g28 (n_179, A[4], B[4]);
  nand g29 (n_180, A[4], n_178);
  nand g30 (n_181, B[4], n_178);
  nand g31 (n_183, n_179, n_180, n_181);
  xor g32 (n_182, A[4], B[4]);
  xor g33 (Z[4], n_178, n_182);
  nand g34 (n_184, A[5], B[5]);
  nand g35 (n_185, A[5], n_183);
  nand g36 (n_186, B[5], n_183);
  nand g37 (n_188, n_184, n_185, n_186);
  xor g38 (n_187, A[5], B[5]);
  xor g39 (Z[5], n_183, n_187);
  nand g40 (n_189, A[6], B[6]);
  nand g41 (n_190, A[6], n_188);
  nand g42 (n_191, B[6], n_188);
  nand g43 (n_193, n_189, n_190, n_191);
  xor g44 (n_192, A[6], B[6]);
  xor g45 (Z[6], n_188, n_192);
  nand g46 (n_194, A[7], B[7]);
  nand g47 (n_195, A[7], n_193);
  nand g48 (n_196, B[7], n_193);
  nand g49 (n_198, n_194, n_195, n_196);
  xor g50 (n_197, A[7], B[7]);
  xor g51 (Z[7], n_193, n_197);
  nand g52 (n_199, A[8], B[8]);
  nand g53 (n_200, A[8], n_198);
  nand g54 (n_201, B[8], n_198);
  nand g55 (n_203, n_199, n_200, n_201);
  xor g56 (n_202, A[8], B[8]);
  xor g57 (Z[8], n_198, n_202);
  nand g58 (n_204, A[9], B[9]);
  nand g59 (n_205, A[9], n_203);
  nand g60 (n_206, B[9], n_203);
  nand g61 (n_208, n_204, n_205, n_206);
  xor g62 (n_207, A[9], B[9]);
  xor g63 (Z[9], n_203, n_207);
  nand g64 (n_209, A[10], B[10]);
  nand g65 (n_210, A[10], n_208);
  nand g66 (n_211, B[10], n_208);
  nand g67 (n_213, n_209, n_210, n_211);
  xor g68 (n_212, A[10], B[10]);
  xor g69 (Z[10], n_208, n_212);
  nand g70 (n_214, A[11], B[11]);
  nand g71 (n_215, A[11], n_213);
  nand g72 (n_216, B[11], n_213);
  nand g73 (n_218, n_214, n_215, n_216);
  xor g74 (n_217, A[11], B[11]);
  xor g75 (Z[11], n_213, n_217);
  nand g76 (n_219, A[12], B[12]);
  nand g77 (n_220, A[12], n_218);
  nand g78 (n_221, B[12], n_218);
  nand g79 (n_223, n_219, n_220, n_221);
  xor g80 (n_222, A[12], B[12]);
  xor g81 (Z[12], n_218, n_222);
  nand g82 (n_224, A[13], B[13]);
  nand g83 (n_225, A[13], n_223);
  nand g84 (n_226, B[13], n_223);
  nand g85 (n_228, n_224, n_225, n_226);
  xor g86 (n_227, A[13], B[13]);
  xor g87 (Z[13], n_223, n_227);
  nand g88 (n_229, A[14], B[14]);
  nand g89 (n_230, A[14], n_228);
  nand g90 (n_231, B[14], n_228);
  nand g91 (n_233, n_229, n_230, n_231);
  xor g92 (n_232, A[14], B[14]);
  xor g93 (Z[14], n_228, n_232);
  nand g94 (n_234, A[15], B[15]);
  nand g95 (n_235, A[15], n_233);
  nand g96 (n_236, B[15], n_233);
  nand g97 (n_238, n_234, n_235, n_236);
  xor g98 (n_237, A[15], B[15]);
  xor g99 (Z[15], n_233, n_237);
  nand g100 (n_239, A[16], B[16]);
  nand g101 (n_240, A[16], n_238);
  nand g102 (n_241, B[16], n_238);
  nand g103 (n_243, n_239, n_240, n_241);
  xor g104 (n_242, A[16], B[16]);
  xor g105 (Z[16], n_238, n_242);
  nand g106 (n_244, A[17], B[17]);
  nand g107 (n_245, A[17], n_243);
  nand g108 (n_246, B[17], n_243);
  nand g109 (n_248, n_244, n_245, n_246);
  xor g110 (n_247, A[17], B[17]);
  xor g111 (Z[17], n_243, n_247);
  nand g112 (n_249, A[18], B[18]);
  nand g113 (n_250, A[18], n_248);
  nand g114 (n_251, B[18], n_248);
  nand g115 (n_253, n_249, n_250, n_251);
  xor g116 (n_252, A[18], B[18]);
  xor g117 (Z[18], n_248, n_252);
  nand g118 (n_254, A[19], B[19]);
  nand g119 (n_255, A[19], n_253);
  nand g120 (n_256, B[19], n_253);
  nand g121 (n_258, n_254, n_255, n_256);
  xor g122 (n_257, A[19], B[19]);
  xor g123 (Z[19], n_253, n_257);
  nand g124 (n_259, A[20], B[20]);
  nand g125 (n_260, A[20], n_258);
  nand g126 (n_261, B[20], n_258);
  nand g127 (n_263, n_259, n_260, n_261);
  xor g128 (n_262, A[20], B[20]);
  xor g129 (Z[20], n_258, n_262);
  nand g130 (n_264, A[21], B[21]);
  nand g131 (n_265, A[21], n_263);
  nand g132 (n_266, B[21], n_263);
  nand g133 (n_268, n_264, n_265, n_266);
  xor g134 (n_267, A[21], B[21]);
  xor g135 (Z[21], n_263, n_267);
  nand g136 (n_269, A[22], B[22]);
  nand g137 (n_270, A[22], n_268);
  nand g138 (n_271, B[22], n_268);
  nand g139 (n_273, n_269, n_270, n_271);
  xor g140 (n_272, A[22], B[22]);
  xor g141 (Z[22], n_268, n_272);
  nand g142 (n_274, A[23], B[23]);
  nand g143 (n_275, A[23], n_273);
  nand g144 (n_276, B[23], n_273);
  nand g145 (n_278, n_274, n_275, n_276);
  xor g146 (n_277, A[23], B[23]);
  xor g147 (Z[23], n_273, n_277);
  nand g148 (n_279, A[24], B[24]);
  nand g149 (n_280, A[24], n_278);
  nand g150 (n_281, B[24], n_278);
  nand g151 (n_283, n_279, n_280, n_281);
  xor g152 (n_282, A[24], B[24]);
  xor g153 (Z[24], n_278, n_282);
  nand g154 (n_284, A[25], B[25]);
  nand g155 (n_285, A[25], n_283);
  nand g156 (n_286, B[25], n_283);
  nand g157 (n_288, n_284, n_285, n_286);
  xor g158 (n_287, A[25], B[25]);
  xor g159 (Z[25], n_283, n_287);
  nand g160 (n_289, A[26], B[26]);
  nand g161 (n_290, A[26], n_288);
  nand g162 (n_291, B[26], n_288);
  nand g163 (n_293, n_289, n_290, n_291);
  xor g164 (n_292, A[26], B[26]);
  xor g165 (Z[26], n_288, n_292);
  nand g166 (n_294, A[27], B[27]);
  nand g167 (n_295, A[27], n_293);
  nand g168 (n_296, B[27], n_293);
  nand g169 (n_298, n_294, n_295, n_296);
  xor g170 (n_297, A[27], B[27]);
  xor g171 (Z[27], n_293, n_297);
  nand g172 (n_299, A[28], B[28]);
  nand g173 (n_300, A[28], n_298);
  nand g174 (n_301, B[28], n_298);
  nand g175 (n_303, n_299, n_300, n_301);
  xor g176 (n_302, A[28], B[28]);
  xor g177 (Z[28], n_298, n_302);
  nand g178 (n_304, A[29], B[29]);
  nand g179 (n_305, A[29], n_303);
  nand g180 (n_306, B[29], n_303);
  nand g181 (n_308, n_304, n_305, n_306);
  xor g182 (n_307, A[29], B[29]);
  xor g183 (Z[29], n_303, n_307);
  nand g184 (n_309, A[30], B[30]);
  nand g185 (n_310, A[30], n_308);
  nand g186 (n_311, B[30], n_308);
  nand g187 (n_313, n_309, n_310, n_311);
  xor g188 (n_312, A[30], B[30]);
  xor g189 (Z[30], n_308, n_312);
  nand g190 (n_314, A[31], B[31]);
  nand g191 (n_315, A[31], n_313);
  nand g192 (n_316, B[31], n_313);
  nand g193 (n_318, n_314, n_315, n_316);
  xor g194 (n_317, A[31], B[31]);
  xor g195 (Z[31], n_313, n_317);
  nand g196 (n_319, A[32], B[32]);
  nand g197 (n_320, A[32], n_318);
  nand g198 (n_321, B[32], n_318);
  nand g199 (n_323, n_319, n_320, n_321);
  xor g200 (n_322, A[32], B[32]);
  xor g201 (Z[32], n_318, n_322);
  nand g202 (n_324, A[33], B[33]);
  nand g203 (n_325, A[33], n_323);
  nand g204 (n_326, B[33], n_323);
  nand g205 (n_328, n_324, n_325, n_326);
  xor g206 (n_327, A[33], B[33]);
  xor g207 (Z[33], n_323, n_327);
  nand g208 (n_329, A[34], B[34]);
  nand g209 (n_330, A[34], n_328);
  nand g210 (n_331, B[34], n_328);
  nand g211 (n_333, n_329, n_330, n_331);
  xor g212 (n_332, A[34], B[34]);
  xor g213 (Z[34], n_328, n_332);
  nand g214 (n_334, A[35], B[35]);
  nand g215 (n_335, A[35], n_333);
  nand g216 (n_336, B[35], n_333);
  nand g217 (n_338, n_334, n_335, n_336);
  xor g218 (n_337, A[35], B[35]);
  xor g219 (Z[35], n_333, n_337);
  nand g220 (n_339, A[36], B[36]);
  nand g221 (n_340, A[36], n_338);
  nand g222 (n_341, B[36], n_338);
  nand g223 (n_343, n_339, n_340, n_341);
  xor g224 (n_342, A[36], B[36]);
  xor g225 (Z[36], n_338, n_342);
  nand g226 (n_344, A[37], B[37]);
  nand g227 (n_345, A[37], n_343);
  nand g228 (n_346, B[37], n_343);
  nand g229 (n_348, n_344, n_345, n_346);
  xor g230 (n_347, A[37], B[37]);
  xor g231 (Z[37], n_343, n_347);
  nand g232 (n_349, A[38], B[38]);
  nand g233 (n_350, A[38], n_348);
  nand g234 (n_351, B[38], n_348);
  nand g235 (n_353, n_349, n_350, n_351);
  xor g236 (n_352, A[38], B[38]);
  xor g237 (Z[38], n_348, n_352);
  nand g238 (n_354, A[39], B[39]);
  nand g239 (n_355, A[39], n_353);
  nand g240 (n_356, B[39], n_353);
  nand g241 (n_358, n_354, n_355, n_356);
  xor g242 (n_357, A[39], B[39]);
  xor g243 (Z[39], n_353, n_357);
  nand g244 (n_359, A[40], B[40]);
  nand g245 (n_360, A[40], n_358);
  nand g246 (n_361, B[40], n_358);
  nand g247 (n_363, n_359, n_360, n_361);
  xor g248 (n_362, A[40], B[40]);
  xor g249 (Z[40], n_358, n_362);
  nand g250 (n_364, A[41], B[41]);
  nand g251 (n_365, A[41], n_363);
  nand g252 (n_366, B[41], n_363);
  nand g253 (n_368, n_364, n_365, n_366);
  xor g254 (n_367, A[41], B[41]);
  xor g255 (Z[41], n_363, n_367);
  nand g256 (n_369, A[42], B[42]);
  nand g257 (n_370, A[42], n_368);
  nand g258 (n_371, B[42], n_368);
  nand g259 (n_373, n_369, n_370, n_371);
  xor g260 (n_372, A[42], B[42]);
  xor g261 (Z[42], n_368, n_372);
  nand g262 (n_374, A[43], B[43]);
  nand g263 (n_375, A[43], n_373);
  nand g264 (n_376, B[43], n_373);
  nand g265 (n_378, n_374, n_375, n_376);
  xor g266 (n_377, A[43], B[43]);
  xor g267 (Z[43], n_373, n_377);
  nand g268 (n_379, A[44], B[44]);
  nand g269 (n_380, A[44], n_378);
  nand g270 (n_381, B[44], n_378);
  nand g271 (n_383, n_379, n_380, n_381);
  xor g272 (n_382, A[44], B[44]);
  xor g273 (Z[44], n_378, n_382);
  nand g274 (n_384, A[45], B[45]);
  nand g275 (n_385, A[45], n_383);
  nand g276 (n_386, B[45], n_383);
  nand g277 (n_388, n_384, n_385, n_386);
  xor g278 (n_387, A[45], B[45]);
  xor g279 (Z[45], n_383, n_387);
  nand g280 (n_389, A[46], B[46]);
  nand g281 (n_390, A[46], n_388);
  nand g282 (n_391, B[46], n_388);
  nand g283 (n_393, n_389, n_390, n_391);
  xor g284 (n_392, A[46], B[46]);
  xor g285 (Z[46], n_388, n_392);
  nand g286 (n_394, A[47], B[47]);
  nand g287 (n_395, A[47], n_393);
  nand g288 (n_396, B[47], n_393);
  nand g289 (n_398, n_394, n_395, n_396);
  xor g290 (n_397, A[47], B[47]);
  xor g291 (Z[47], n_393, n_397);
  nand g292 (n_399, A[48], B[48]);
  nand g293 (n_400, A[48], n_398);
  nand g294 (n_401, B[48], n_398);
  nand g295 (n_403, n_399, n_400, n_401);
  xor g296 (n_402, A[48], B[48]);
  xor g297 (Z[48], n_398, n_402);
  nand g298 (n_404, A[49], B[49]);
  nand g299 (n_405, A[49], n_403);
  nand g300 (n_406, B[49], n_403);
  nand g301 (n_408, n_404, n_405, n_406);
  xor g302 (n_407, A[49], B[49]);
  xor g303 (Z[49], n_403, n_407);
  nand g307 (n_158, n_409, n_410, n_411);
  xor g309 (Z[50], n_408, n_412);
  or g311 (n_409, A[50], B[50]);
  xor g312 (n_412, A[50], B[50]);
  or g313 (n_165, wc, n_159);
  not gc (wc, A[1]);
  or g314 (n_166, wc0, n_159);
  not gc0 (wc0, B[1]);
  xnor g315 (Z[1], n_159, n_167);
  or g316 (n_410, A[50], wc1);
  not gc1 (wc1, n_408);
  or g317 (n_411, B[50], wc2);
  not gc2 (wc2, n_408);
endmodule

module add_signed_7256_GENERIC(A, B, Z);
  input [50:0] A, B;
  output [51:0] Z;
  wire [50:0] A, B;
  wire [51:0] Z;
  add_signed_7256_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_7256_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [50:0] A, B;
  output [51:0] Z;
  wire [50:0] A, B;
  wire [51:0] Z;
  wire n_158, n_159, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412;
  not g3 (Z[51], n_158);
  nand g4 (n_159, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_164, A[1], B[1]);
  nand g13 (n_168, n_164, n_165, n_166);
  xor g14 (n_167, A[1], B[1]);
  nand g16 (n_169, A[2], B[2]);
  nand g17 (n_170, A[2], n_168);
  nand g18 (n_171, B[2], n_168);
  nand g19 (n_173, n_169, n_170, n_171);
  xor g20 (n_172, A[2], B[2]);
  xor g21 (Z[2], n_168, n_172);
  nand g22 (n_174, A[3], B[3]);
  nand g23 (n_175, A[3], n_173);
  nand g24 (n_176, B[3], n_173);
  nand g25 (n_178, n_174, n_175, n_176);
  xor g26 (n_177, A[3], B[3]);
  xor g27 (Z[3], n_173, n_177);
  nand g28 (n_179, A[4], B[4]);
  nand g29 (n_180, A[4], n_178);
  nand g30 (n_181, B[4], n_178);
  nand g31 (n_183, n_179, n_180, n_181);
  xor g32 (n_182, A[4], B[4]);
  xor g33 (Z[4], n_178, n_182);
  nand g34 (n_184, A[5], B[5]);
  nand g35 (n_185, A[5], n_183);
  nand g36 (n_186, B[5], n_183);
  nand g37 (n_188, n_184, n_185, n_186);
  xor g38 (n_187, A[5], B[5]);
  xor g39 (Z[5], n_183, n_187);
  nand g40 (n_189, A[6], B[6]);
  nand g41 (n_190, A[6], n_188);
  nand g42 (n_191, B[6], n_188);
  nand g43 (n_193, n_189, n_190, n_191);
  xor g44 (n_192, A[6], B[6]);
  xor g45 (Z[6], n_188, n_192);
  nand g46 (n_194, A[7], B[7]);
  nand g47 (n_195, A[7], n_193);
  nand g48 (n_196, B[7], n_193);
  nand g49 (n_198, n_194, n_195, n_196);
  xor g50 (n_197, A[7], B[7]);
  xor g51 (Z[7], n_193, n_197);
  nand g52 (n_199, A[8], B[8]);
  nand g53 (n_200, A[8], n_198);
  nand g54 (n_201, B[8], n_198);
  nand g55 (n_203, n_199, n_200, n_201);
  xor g56 (n_202, A[8], B[8]);
  xor g57 (Z[8], n_198, n_202);
  nand g58 (n_204, A[9], B[9]);
  nand g59 (n_205, A[9], n_203);
  nand g60 (n_206, B[9], n_203);
  nand g61 (n_208, n_204, n_205, n_206);
  xor g62 (n_207, A[9], B[9]);
  xor g63 (Z[9], n_203, n_207);
  nand g64 (n_209, A[10], B[10]);
  nand g65 (n_210, A[10], n_208);
  nand g66 (n_211, B[10], n_208);
  nand g67 (n_213, n_209, n_210, n_211);
  xor g68 (n_212, A[10], B[10]);
  xor g69 (Z[10], n_208, n_212);
  nand g70 (n_214, A[11], B[11]);
  nand g71 (n_215, A[11], n_213);
  nand g72 (n_216, B[11], n_213);
  nand g73 (n_218, n_214, n_215, n_216);
  xor g74 (n_217, A[11], B[11]);
  xor g75 (Z[11], n_213, n_217);
  nand g76 (n_219, A[12], B[12]);
  nand g77 (n_220, A[12], n_218);
  nand g78 (n_221, B[12], n_218);
  nand g79 (n_223, n_219, n_220, n_221);
  xor g80 (n_222, A[12], B[12]);
  xor g81 (Z[12], n_218, n_222);
  nand g82 (n_224, A[13], B[13]);
  nand g83 (n_225, A[13], n_223);
  nand g84 (n_226, B[13], n_223);
  nand g85 (n_228, n_224, n_225, n_226);
  xor g86 (n_227, A[13], B[13]);
  xor g87 (Z[13], n_223, n_227);
  nand g88 (n_229, A[14], B[14]);
  nand g89 (n_230, A[14], n_228);
  nand g90 (n_231, B[14], n_228);
  nand g91 (n_233, n_229, n_230, n_231);
  xor g92 (n_232, A[14], B[14]);
  xor g93 (Z[14], n_228, n_232);
  nand g94 (n_234, A[15], B[15]);
  nand g95 (n_235, A[15], n_233);
  nand g96 (n_236, B[15], n_233);
  nand g97 (n_238, n_234, n_235, n_236);
  xor g98 (n_237, A[15], B[15]);
  xor g99 (Z[15], n_233, n_237);
  nand g100 (n_239, A[16], B[16]);
  nand g101 (n_240, A[16], n_238);
  nand g102 (n_241, B[16], n_238);
  nand g103 (n_243, n_239, n_240, n_241);
  xor g104 (n_242, A[16], B[16]);
  xor g105 (Z[16], n_238, n_242);
  nand g106 (n_244, A[17], B[17]);
  nand g107 (n_245, A[17], n_243);
  nand g108 (n_246, B[17], n_243);
  nand g109 (n_248, n_244, n_245, n_246);
  xor g110 (n_247, A[17], B[17]);
  xor g111 (Z[17], n_243, n_247);
  nand g112 (n_249, A[18], B[18]);
  nand g113 (n_250, A[18], n_248);
  nand g114 (n_251, B[18], n_248);
  nand g115 (n_253, n_249, n_250, n_251);
  xor g116 (n_252, A[18], B[18]);
  xor g117 (Z[18], n_248, n_252);
  nand g118 (n_254, A[19], B[19]);
  nand g119 (n_255, A[19], n_253);
  nand g120 (n_256, B[19], n_253);
  nand g121 (n_258, n_254, n_255, n_256);
  xor g122 (n_257, A[19], B[19]);
  xor g123 (Z[19], n_253, n_257);
  nand g124 (n_259, A[20], B[20]);
  nand g125 (n_260, A[20], n_258);
  nand g126 (n_261, B[20], n_258);
  nand g127 (n_263, n_259, n_260, n_261);
  xor g128 (n_262, A[20], B[20]);
  xor g129 (Z[20], n_258, n_262);
  nand g130 (n_264, A[21], B[21]);
  nand g131 (n_265, A[21], n_263);
  nand g132 (n_266, B[21], n_263);
  nand g133 (n_268, n_264, n_265, n_266);
  xor g134 (n_267, A[21], B[21]);
  xor g135 (Z[21], n_263, n_267);
  nand g136 (n_269, A[22], B[22]);
  nand g137 (n_270, A[22], n_268);
  nand g138 (n_271, B[22], n_268);
  nand g139 (n_273, n_269, n_270, n_271);
  xor g140 (n_272, A[22], B[22]);
  xor g141 (Z[22], n_268, n_272);
  nand g142 (n_274, A[23], B[23]);
  nand g143 (n_275, A[23], n_273);
  nand g144 (n_276, B[23], n_273);
  nand g145 (n_278, n_274, n_275, n_276);
  xor g146 (n_277, A[23], B[23]);
  xor g147 (Z[23], n_273, n_277);
  nand g148 (n_279, A[24], B[24]);
  nand g149 (n_280, A[24], n_278);
  nand g150 (n_281, B[24], n_278);
  nand g151 (n_283, n_279, n_280, n_281);
  xor g152 (n_282, A[24], B[24]);
  xor g153 (Z[24], n_278, n_282);
  nand g154 (n_284, A[25], B[25]);
  nand g155 (n_285, A[25], n_283);
  nand g156 (n_286, B[25], n_283);
  nand g157 (n_288, n_284, n_285, n_286);
  xor g158 (n_287, A[25], B[25]);
  xor g159 (Z[25], n_283, n_287);
  nand g160 (n_289, A[26], B[26]);
  nand g161 (n_290, A[26], n_288);
  nand g162 (n_291, B[26], n_288);
  nand g163 (n_293, n_289, n_290, n_291);
  xor g164 (n_292, A[26], B[26]);
  xor g165 (Z[26], n_288, n_292);
  nand g166 (n_294, A[27], B[27]);
  nand g167 (n_295, A[27], n_293);
  nand g168 (n_296, B[27], n_293);
  nand g169 (n_298, n_294, n_295, n_296);
  xor g170 (n_297, A[27], B[27]);
  xor g171 (Z[27], n_293, n_297);
  nand g172 (n_299, A[28], B[28]);
  nand g173 (n_300, A[28], n_298);
  nand g174 (n_301, B[28], n_298);
  nand g175 (n_303, n_299, n_300, n_301);
  xor g176 (n_302, A[28], B[28]);
  xor g177 (Z[28], n_298, n_302);
  nand g178 (n_304, A[29], B[29]);
  nand g179 (n_305, A[29], n_303);
  nand g180 (n_306, B[29], n_303);
  nand g181 (n_308, n_304, n_305, n_306);
  xor g182 (n_307, A[29], B[29]);
  xor g183 (Z[29], n_303, n_307);
  nand g184 (n_309, A[30], B[30]);
  nand g185 (n_310, A[30], n_308);
  nand g186 (n_311, B[30], n_308);
  nand g187 (n_313, n_309, n_310, n_311);
  xor g188 (n_312, A[30], B[30]);
  xor g189 (Z[30], n_308, n_312);
  nand g190 (n_314, A[31], B[31]);
  nand g191 (n_315, A[31], n_313);
  nand g192 (n_316, B[31], n_313);
  nand g193 (n_318, n_314, n_315, n_316);
  xor g194 (n_317, A[31], B[31]);
  xor g195 (Z[31], n_313, n_317);
  nand g196 (n_319, A[32], B[32]);
  nand g197 (n_320, A[32], n_318);
  nand g198 (n_321, B[32], n_318);
  nand g199 (n_323, n_319, n_320, n_321);
  xor g200 (n_322, A[32], B[32]);
  xor g201 (Z[32], n_318, n_322);
  nand g202 (n_324, A[33], B[33]);
  nand g203 (n_325, A[33], n_323);
  nand g204 (n_326, B[33], n_323);
  nand g205 (n_328, n_324, n_325, n_326);
  xor g206 (n_327, A[33], B[33]);
  xor g207 (Z[33], n_323, n_327);
  nand g208 (n_329, A[34], B[34]);
  nand g209 (n_330, A[34], n_328);
  nand g210 (n_331, B[34], n_328);
  nand g211 (n_333, n_329, n_330, n_331);
  xor g212 (n_332, A[34], B[34]);
  xor g213 (Z[34], n_328, n_332);
  nand g214 (n_334, A[35], B[35]);
  nand g215 (n_335, A[35], n_333);
  nand g216 (n_336, B[35], n_333);
  nand g217 (n_338, n_334, n_335, n_336);
  xor g218 (n_337, A[35], B[35]);
  xor g219 (Z[35], n_333, n_337);
  nand g220 (n_339, A[36], B[36]);
  nand g221 (n_340, A[36], n_338);
  nand g222 (n_341, B[36], n_338);
  nand g223 (n_343, n_339, n_340, n_341);
  xor g224 (n_342, A[36], B[36]);
  xor g225 (Z[36], n_338, n_342);
  nand g226 (n_344, A[37], B[37]);
  nand g227 (n_345, A[37], n_343);
  nand g228 (n_346, B[37], n_343);
  nand g229 (n_348, n_344, n_345, n_346);
  xor g230 (n_347, A[37], B[37]);
  xor g231 (Z[37], n_343, n_347);
  nand g232 (n_349, A[38], B[38]);
  nand g233 (n_350, A[38], n_348);
  nand g234 (n_351, B[38], n_348);
  nand g235 (n_353, n_349, n_350, n_351);
  xor g236 (n_352, A[38], B[38]);
  xor g237 (Z[38], n_348, n_352);
  nand g238 (n_354, A[39], B[39]);
  nand g239 (n_355, A[39], n_353);
  nand g240 (n_356, B[39], n_353);
  nand g241 (n_358, n_354, n_355, n_356);
  xor g242 (n_357, A[39], B[39]);
  xor g243 (Z[39], n_353, n_357);
  nand g244 (n_359, A[40], B[40]);
  nand g245 (n_360, A[40], n_358);
  nand g246 (n_361, B[40], n_358);
  nand g247 (n_363, n_359, n_360, n_361);
  xor g248 (n_362, A[40], B[40]);
  xor g249 (Z[40], n_358, n_362);
  nand g250 (n_364, A[41], B[41]);
  nand g251 (n_365, A[41], n_363);
  nand g252 (n_366, B[41], n_363);
  nand g253 (n_368, n_364, n_365, n_366);
  xor g254 (n_367, A[41], B[41]);
  xor g255 (Z[41], n_363, n_367);
  nand g256 (n_369, A[42], B[42]);
  nand g257 (n_370, A[42], n_368);
  nand g258 (n_371, B[42], n_368);
  nand g259 (n_373, n_369, n_370, n_371);
  xor g260 (n_372, A[42], B[42]);
  xor g261 (Z[42], n_368, n_372);
  nand g262 (n_374, A[43], B[43]);
  nand g263 (n_375, A[43], n_373);
  nand g264 (n_376, B[43], n_373);
  nand g265 (n_378, n_374, n_375, n_376);
  xor g266 (n_377, A[43], B[43]);
  xor g267 (Z[43], n_373, n_377);
  nand g268 (n_379, A[44], B[44]);
  nand g269 (n_380, A[44], n_378);
  nand g270 (n_381, B[44], n_378);
  nand g271 (n_383, n_379, n_380, n_381);
  xor g272 (n_382, A[44], B[44]);
  xor g273 (Z[44], n_378, n_382);
  nand g274 (n_384, A[45], B[45]);
  nand g275 (n_385, A[45], n_383);
  nand g276 (n_386, B[45], n_383);
  nand g277 (n_388, n_384, n_385, n_386);
  xor g278 (n_387, A[45], B[45]);
  xor g279 (Z[45], n_383, n_387);
  nand g280 (n_389, A[46], B[46]);
  nand g281 (n_390, A[46], n_388);
  nand g282 (n_391, B[46], n_388);
  nand g283 (n_393, n_389, n_390, n_391);
  xor g284 (n_392, A[46], B[46]);
  xor g285 (Z[46], n_388, n_392);
  nand g286 (n_394, A[47], B[47]);
  nand g287 (n_395, A[47], n_393);
  nand g288 (n_396, B[47], n_393);
  nand g289 (n_398, n_394, n_395, n_396);
  xor g290 (n_397, A[47], B[47]);
  xor g291 (Z[47], n_393, n_397);
  nand g292 (n_399, A[48], B[48]);
  nand g293 (n_400, A[48], n_398);
  nand g294 (n_401, B[48], n_398);
  nand g295 (n_403, n_399, n_400, n_401);
  xor g296 (n_402, A[48], B[48]);
  xor g297 (Z[48], n_398, n_402);
  nand g298 (n_404, A[49], B[49]);
  nand g299 (n_405, A[49], n_403);
  nand g300 (n_406, B[49], n_403);
  nand g301 (n_408, n_404, n_405, n_406);
  xor g302 (n_407, A[49], B[49]);
  xor g303 (Z[49], n_403, n_407);
  nand g307 (n_158, n_409, n_410, n_411);
  xor g309 (Z[50], n_408, n_412);
  or g311 (n_409, A[50], B[50]);
  xor g312 (n_412, A[50], B[50]);
  or g313 (n_165, wc, n_159);
  not gc (wc, A[1]);
  or g314 (n_166, wc0, n_159);
  not gc0 (wc0, B[1]);
  xnor g315 (Z[1], n_159, n_167);
  or g316 (n_410, A[50], wc1);
  not gc1 (wc1, n_408);
  or g317 (n_411, B[50], wc2);
  not gc2 (wc2, n_408);
endmodule

module add_signed_7256_1_GENERIC(A, B, Z);
  input [50:0] A, B;
  output [51:0] Z;
  wire [50:0] A, B;
  wire [51:0] Z;
  add_signed_7256_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_7719_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [49:0] A, B;
  output [50:0] Z;
  wire [49:0] A, B;
  wire [50:0] Z;
  wire n_155, n_156, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404;
  not g3 (Z[50], n_155);
  nand g4 (n_156, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_161, A[1], B[1]);
  nand g13 (n_165, n_161, n_162, n_163);
  xor g14 (n_164, A[1], B[1]);
  nand g16 (n_166, A[2], B[2]);
  nand g17 (n_167, A[2], n_165);
  nand g18 (n_168, B[2], n_165);
  nand g19 (n_170, n_166, n_167, n_168);
  xor g20 (n_169, A[2], B[2]);
  xor g21 (Z[2], n_165, n_169);
  nand g22 (n_171, A[3], B[3]);
  nand g23 (n_172, A[3], n_170);
  nand g24 (n_173, B[3], n_170);
  nand g25 (n_175, n_171, n_172, n_173);
  xor g26 (n_174, A[3], B[3]);
  xor g27 (Z[3], n_170, n_174);
  nand g28 (n_176, A[4], B[4]);
  nand g29 (n_177, A[4], n_175);
  nand g30 (n_178, B[4], n_175);
  nand g31 (n_180, n_176, n_177, n_178);
  xor g32 (n_179, A[4], B[4]);
  xor g33 (Z[4], n_175, n_179);
  nand g34 (n_181, A[5], B[5]);
  nand g35 (n_182, A[5], n_180);
  nand g36 (n_183, B[5], n_180);
  nand g37 (n_185, n_181, n_182, n_183);
  xor g38 (n_184, A[5], B[5]);
  xor g39 (Z[5], n_180, n_184);
  nand g40 (n_186, A[6], B[6]);
  nand g41 (n_187, A[6], n_185);
  nand g42 (n_188, B[6], n_185);
  nand g43 (n_190, n_186, n_187, n_188);
  xor g44 (n_189, A[6], B[6]);
  xor g45 (Z[6], n_185, n_189);
  nand g46 (n_191, A[7], B[7]);
  nand g47 (n_192, A[7], n_190);
  nand g48 (n_193, B[7], n_190);
  nand g49 (n_195, n_191, n_192, n_193);
  xor g50 (n_194, A[7], B[7]);
  xor g51 (Z[7], n_190, n_194);
  nand g52 (n_196, A[8], B[8]);
  nand g53 (n_197, A[8], n_195);
  nand g54 (n_198, B[8], n_195);
  nand g55 (n_200, n_196, n_197, n_198);
  xor g56 (n_199, A[8], B[8]);
  xor g57 (Z[8], n_195, n_199);
  nand g58 (n_201, A[9], B[9]);
  nand g59 (n_202, A[9], n_200);
  nand g60 (n_203, B[9], n_200);
  nand g61 (n_205, n_201, n_202, n_203);
  xor g62 (n_204, A[9], B[9]);
  xor g63 (Z[9], n_200, n_204);
  nand g64 (n_206, A[10], B[10]);
  nand g65 (n_207, A[10], n_205);
  nand g66 (n_208, B[10], n_205);
  nand g67 (n_210, n_206, n_207, n_208);
  xor g68 (n_209, A[10], B[10]);
  xor g69 (Z[10], n_205, n_209);
  nand g70 (n_211, A[11], B[11]);
  nand g71 (n_212, A[11], n_210);
  nand g72 (n_213, B[11], n_210);
  nand g73 (n_215, n_211, n_212, n_213);
  xor g74 (n_214, A[11], B[11]);
  xor g75 (Z[11], n_210, n_214);
  nand g76 (n_216, A[12], B[12]);
  nand g77 (n_217, A[12], n_215);
  nand g78 (n_218, B[12], n_215);
  nand g79 (n_220, n_216, n_217, n_218);
  xor g80 (n_219, A[12], B[12]);
  xor g81 (Z[12], n_215, n_219);
  nand g82 (n_221, A[13], B[13]);
  nand g83 (n_222, A[13], n_220);
  nand g84 (n_223, B[13], n_220);
  nand g85 (n_225, n_221, n_222, n_223);
  xor g86 (n_224, A[13], B[13]);
  xor g87 (Z[13], n_220, n_224);
  nand g88 (n_226, A[14], B[14]);
  nand g89 (n_227, A[14], n_225);
  nand g90 (n_228, B[14], n_225);
  nand g91 (n_230, n_226, n_227, n_228);
  xor g92 (n_229, A[14], B[14]);
  xor g93 (Z[14], n_225, n_229);
  nand g94 (n_231, A[15], B[15]);
  nand g95 (n_232, A[15], n_230);
  nand g96 (n_233, B[15], n_230);
  nand g97 (n_235, n_231, n_232, n_233);
  xor g98 (n_234, A[15], B[15]);
  xor g99 (Z[15], n_230, n_234);
  nand g100 (n_236, A[16], B[16]);
  nand g101 (n_237, A[16], n_235);
  nand g102 (n_238, B[16], n_235);
  nand g103 (n_240, n_236, n_237, n_238);
  xor g104 (n_239, A[16], B[16]);
  xor g105 (Z[16], n_235, n_239);
  nand g106 (n_241, A[17], B[17]);
  nand g107 (n_242, A[17], n_240);
  nand g108 (n_243, B[17], n_240);
  nand g109 (n_245, n_241, n_242, n_243);
  xor g110 (n_244, A[17], B[17]);
  xor g111 (Z[17], n_240, n_244);
  nand g112 (n_246, A[18], B[18]);
  nand g113 (n_247, A[18], n_245);
  nand g114 (n_248, B[18], n_245);
  nand g115 (n_250, n_246, n_247, n_248);
  xor g116 (n_249, A[18], B[18]);
  xor g117 (Z[18], n_245, n_249);
  nand g118 (n_251, A[19], B[19]);
  nand g119 (n_252, A[19], n_250);
  nand g120 (n_253, B[19], n_250);
  nand g121 (n_255, n_251, n_252, n_253);
  xor g122 (n_254, A[19], B[19]);
  xor g123 (Z[19], n_250, n_254);
  nand g124 (n_256, A[20], B[20]);
  nand g125 (n_257, A[20], n_255);
  nand g126 (n_258, B[20], n_255);
  nand g127 (n_260, n_256, n_257, n_258);
  xor g128 (n_259, A[20], B[20]);
  xor g129 (Z[20], n_255, n_259);
  nand g130 (n_261, A[21], B[21]);
  nand g131 (n_262, A[21], n_260);
  nand g132 (n_263, B[21], n_260);
  nand g133 (n_265, n_261, n_262, n_263);
  xor g134 (n_264, A[21], B[21]);
  xor g135 (Z[21], n_260, n_264);
  nand g136 (n_266, A[22], B[22]);
  nand g137 (n_267, A[22], n_265);
  nand g138 (n_268, B[22], n_265);
  nand g139 (n_270, n_266, n_267, n_268);
  xor g140 (n_269, A[22], B[22]);
  xor g141 (Z[22], n_265, n_269);
  nand g142 (n_271, A[23], B[23]);
  nand g143 (n_272, A[23], n_270);
  nand g144 (n_273, B[23], n_270);
  nand g145 (n_275, n_271, n_272, n_273);
  xor g146 (n_274, A[23], B[23]);
  xor g147 (Z[23], n_270, n_274);
  nand g148 (n_276, A[24], B[24]);
  nand g149 (n_277, A[24], n_275);
  nand g150 (n_278, B[24], n_275);
  nand g151 (n_280, n_276, n_277, n_278);
  xor g152 (n_279, A[24], B[24]);
  xor g153 (Z[24], n_275, n_279);
  nand g154 (n_281, A[25], B[25]);
  nand g155 (n_282, A[25], n_280);
  nand g156 (n_283, B[25], n_280);
  nand g157 (n_285, n_281, n_282, n_283);
  xor g158 (n_284, A[25], B[25]);
  xor g159 (Z[25], n_280, n_284);
  nand g160 (n_286, A[26], B[26]);
  nand g161 (n_287, A[26], n_285);
  nand g162 (n_288, B[26], n_285);
  nand g163 (n_290, n_286, n_287, n_288);
  xor g164 (n_289, A[26], B[26]);
  xor g165 (Z[26], n_285, n_289);
  nand g166 (n_291, A[27], B[27]);
  nand g167 (n_292, A[27], n_290);
  nand g168 (n_293, B[27], n_290);
  nand g169 (n_295, n_291, n_292, n_293);
  xor g170 (n_294, A[27], B[27]);
  xor g171 (Z[27], n_290, n_294);
  nand g172 (n_296, A[28], B[28]);
  nand g173 (n_297, A[28], n_295);
  nand g174 (n_298, B[28], n_295);
  nand g175 (n_300, n_296, n_297, n_298);
  xor g176 (n_299, A[28], B[28]);
  xor g177 (Z[28], n_295, n_299);
  nand g178 (n_301, A[29], B[29]);
  nand g179 (n_302, A[29], n_300);
  nand g180 (n_303, B[29], n_300);
  nand g181 (n_305, n_301, n_302, n_303);
  xor g182 (n_304, A[29], B[29]);
  xor g183 (Z[29], n_300, n_304);
  nand g184 (n_306, A[30], B[30]);
  nand g185 (n_307, A[30], n_305);
  nand g186 (n_308, B[30], n_305);
  nand g187 (n_310, n_306, n_307, n_308);
  xor g188 (n_309, A[30], B[30]);
  xor g189 (Z[30], n_305, n_309);
  nand g190 (n_311, A[31], B[31]);
  nand g191 (n_312, A[31], n_310);
  nand g192 (n_313, B[31], n_310);
  nand g193 (n_315, n_311, n_312, n_313);
  xor g194 (n_314, A[31], B[31]);
  xor g195 (Z[31], n_310, n_314);
  nand g196 (n_316, A[32], B[32]);
  nand g197 (n_317, A[32], n_315);
  nand g198 (n_318, B[32], n_315);
  nand g199 (n_320, n_316, n_317, n_318);
  xor g200 (n_319, A[32], B[32]);
  xor g201 (Z[32], n_315, n_319);
  nand g202 (n_321, A[33], B[33]);
  nand g203 (n_322, A[33], n_320);
  nand g204 (n_323, B[33], n_320);
  nand g205 (n_325, n_321, n_322, n_323);
  xor g206 (n_324, A[33], B[33]);
  xor g207 (Z[33], n_320, n_324);
  nand g208 (n_326, A[34], B[34]);
  nand g209 (n_327, A[34], n_325);
  nand g210 (n_328, B[34], n_325);
  nand g211 (n_330, n_326, n_327, n_328);
  xor g212 (n_329, A[34], B[34]);
  xor g213 (Z[34], n_325, n_329);
  nand g214 (n_331, A[35], B[35]);
  nand g215 (n_332, A[35], n_330);
  nand g216 (n_333, B[35], n_330);
  nand g217 (n_335, n_331, n_332, n_333);
  xor g218 (n_334, A[35], B[35]);
  xor g219 (Z[35], n_330, n_334);
  nand g220 (n_336, A[36], B[36]);
  nand g221 (n_337, A[36], n_335);
  nand g222 (n_338, B[36], n_335);
  nand g223 (n_340, n_336, n_337, n_338);
  xor g224 (n_339, A[36], B[36]);
  xor g225 (Z[36], n_335, n_339);
  nand g226 (n_341, A[37], B[37]);
  nand g227 (n_342, A[37], n_340);
  nand g228 (n_343, B[37], n_340);
  nand g229 (n_345, n_341, n_342, n_343);
  xor g230 (n_344, A[37], B[37]);
  xor g231 (Z[37], n_340, n_344);
  nand g232 (n_346, A[38], B[38]);
  nand g233 (n_347, A[38], n_345);
  nand g234 (n_348, B[38], n_345);
  nand g235 (n_350, n_346, n_347, n_348);
  xor g236 (n_349, A[38], B[38]);
  xor g237 (Z[38], n_345, n_349);
  nand g238 (n_351, A[39], B[39]);
  nand g239 (n_352, A[39], n_350);
  nand g240 (n_353, B[39], n_350);
  nand g241 (n_355, n_351, n_352, n_353);
  xor g242 (n_354, A[39], B[39]);
  xor g243 (Z[39], n_350, n_354);
  nand g244 (n_356, A[40], B[40]);
  nand g245 (n_357, A[40], n_355);
  nand g246 (n_358, B[40], n_355);
  nand g247 (n_360, n_356, n_357, n_358);
  xor g248 (n_359, A[40], B[40]);
  xor g249 (Z[40], n_355, n_359);
  nand g250 (n_361, A[41], B[41]);
  nand g251 (n_362, A[41], n_360);
  nand g252 (n_363, B[41], n_360);
  nand g253 (n_365, n_361, n_362, n_363);
  xor g254 (n_364, A[41], B[41]);
  xor g255 (Z[41], n_360, n_364);
  nand g256 (n_366, A[42], B[42]);
  nand g257 (n_367, A[42], n_365);
  nand g258 (n_368, B[42], n_365);
  nand g259 (n_370, n_366, n_367, n_368);
  xor g260 (n_369, A[42], B[42]);
  xor g261 (Z[42], n_365, n_369);
  nand g262 (n_371, A[43], B[43]);
  nand g263 (n_372, A[43], n_370);
  nand g264 (n_373, B[43], n_370);
  nand g265 (n_375, n_371, n_372, n_373);
  xor g266 (n_374, A[43], B[43]);
  xor g267 (Z[43], n_370, n_374);
  nand g268 (n_376, A[44], B[44]);
  nand g269 (n_377, A[44], n_375);
  nand g270 (n_378, B[44], n_375);
  nand g271 (n_380, n_376, n_377, n_378);
  xor g272 (n_379, A[44], B[44]);
  xor g273 (Z[44], n_375, n_379);
  nand g274 (n_381, A[45], B[45]);
  nand g275 (n_382, A[45], n_380);
  nand g276 (n_383, B[45], n_380);
  nand g277 (n_385, n_381, n_382, n_383);
  xor g278 (n_384, A[45], B[45]);
  xor g279 (Z[45], n_380, n_384);
  nand g280 (n_386, A[46], B[46]);
  nand g281 (n_387, A[46], n_385);
  nand g282 (n_388, B[46], n_385);
  nand g283 (n_390, n_386, n_387, n_388);
  xor g284 (n_389, A[46], B[46]);
  xor g285 (Z[46], n_385, n_389);
  nand g286 (n_391, A[47], B[47]);
  nand g287 (n_392, A[47], n_390);
  nand g288 (n_393, B[47], n_390);
  nand g289 (n_395, n_391, n_392, n_393);
  xor g290 (n_394, A[47], B[47]);
  xor g291 (Z[47], n_390, n_394);
  nand g292 (n_396, A[48], B[48]);
  nand g293 (n_397, A[48], n_395);
  nand g294 (n_398, B[48], n_395);
  nand g295 (n_400, n_396, n_397, n_398);
  xor g296 (n_399, A[48], B[48]);
  xor g297 (Z[48], n_395, n_399);
  nand g301 (n_155, n_401, n_402, n_403);
  xor g303 (Z[49], n_400, n_404);
  or g305 (n_401, A[49], B[49]);
  xor g306 (n_404, A[49], B[49]);
  or g307 (n_162, wc, n_156);
  not gc (wc, A[1]);
  or g308 (n_163, wc0, n_156);
  not gc0 (wc0, B[1]);
  xnor g309 (Z[1], n_156, n_164);
  or g310 (n_402, A[49], wc1);
  not gc1 (wc1, n_400);
  or g311 (n_403, B[49], wc2);
  not gc2 (wc2, n_400);
endmodule

module add_signed_7719_GENERIC(A, B, Z);
  input [49:0] A, B;
  output [50:0] Z;
  wire [49:0] A, B;
  wire [50:0] Z;
  add_signed_7719_GENERIC_REAL g1(.A ({A[49:2], A[0], A[0]}), .B (B),
       .Z (Z));
endmodule

module add_signed_7719_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [49:0] A, B;
  output [50:0] Z;
  wire [49:0] A, B;
  wire [50:0] Z;
  wire n_155, n_156, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262;
  wire n_263, n_264, n_265, n_266, n_267, n_268, n_269, n_270;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_279, n_280, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_295, n_296, n_297, n_298, n_299, n_300, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404;
  not g3 (Z[50], n_155);
  nand g4 (n_156, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_161, A[1], B[1]);
  nand g13 (n_165, n_161, n_162, n_163);
  xor g14 (n_164, A[1], B[1]);
  nand g16 (n_166, A[2], B[2]);
  nand g17 (n_167, A[2], n_165);
  nand g18 (n_168, B[2], n_165);
  nand g19 (n_170, n_166, n_167, n_168);
  xor g20 (n_169, A[2], B[2]);
  xor g21 (Z[2], n_165, n_169);
  nand g22 (n_171, A[3], B[3]);
  nand g23 (n_172, A[3], n_170);
  nand g24 (n_173, B[3], n_170);
  nand g25 (n_175, n_171, n_172, n_173);
  xor g26 (n_174, A[3], B[3]);
  xor g27 (Z[3], n_170, n_174);
  nand g28 (n_176, A[4], B[4]);
  nand g29 (n_177, A[4], n_175);
  nand g30 (n_178, B[4], n_175);
  nand g31 (n_180, n_176, n_177, n_178);
  xor g32 (n_179, A[4], B[4]);
  xor g33 (Z[4], n_175, n_179);
  nand g34 (n_181, A[5], B[5]);
  nand g35 (n_182, A[5], n_180);
  nand g36 (n_183, B[5], n_180);
  nand g37 (n_185, n_181, n_182, n_183);
  xor g38 (n_184, A[5], B[5]);
  xor g39 (Z[5], n_180, n_184);
  nand g40 (n_186, A[6], B[6]);
  nand g41 (n_187, A[6], n_185);
  nand g42 (n_188, B[6], n_185);
  nand g43 (n_190, n_186, n_187, n_188);
  xor g44 (n_189, A[6], B[6]);
  xor g45 (Z[6], n_185, n_189);
  nand g46 (n_191, A[7], B[7]);
  nand g47 (n_192, A[7], n_190);
  nand g48 (n_193, B[7], n_190);
  nand g49 (n_195, n_191, n_192, n_193);
  xor g50 (n_194, A[7], B[7]);
  xor g51 (Z[7], n_190, n_194);
  nand g52 (n_196, A[8], B[8]);
  nand g53 (n_197, A[8], n_195);
  nand g54 (n_198, B[8], n_195);
  nand g55 (n_200, n_196, n_197, n_198);
  xor g56 (n_199, A[8], B[8]);
  xor g57 (Z[8], n_195, n_199);
  nand g58 (n_201, A[9], B[9]);
  nand g59 (n_202, A[9], n_200);
  nand g60 (n_203, B[9], n_200);
  nand g61 (n_205, n_201, n_202, n_203);
  xor g62 (n_204, A[9], B[9]);
  xor g63 (Z[9], n_200, n_204);
  nand g64 (n_206, A[10], B[10]);
  nand g65 (n_207, A[10], n_205);
  nand g66 (n_208, B[10], n_205);
  nand g67 (n_210, n_206, n_207, n_208);
  xor g68 (n_209, A[10], B[10]);
  xor g69 (Z[10], n_205, n_209);
  nand g70 (n_211, A[11], B[11]);
  nand g71 (n_212, A[11], n_210);
  nand g72 (n_213, B[11], n_210);
  nand g73 (n_215, n_211, n_212, n_213);
  xor g74 (n_214, A[11], B[11]);
  xor g75 (Z[11], n_210, n_214);
  nand g76 (n_216, A[12], B[12]);
  nand g77 (n_217, A[12], n_215);
  nand g78 (n_218, B[12], n_215);
  nand g79 (n_220, n_216, n_217, n_218);
  xor g80 (n_219, A[12], B[12]);
  xor g81 (Z[12], n_215, n_219);
  nand g82 (n_221, A[13], B[13]);
  nand g83 (n_222, A[13], n_220);
  nand g84 (n_223, B[13], n_220);
  nand g85 (n_225, n_221, n_222, n_223);
  xor g86 (n_224, A[13], B[13]);
  xor g87 (Z[13], n_220, n_224);
  nand g88 (n_226, A[14], B[14]);
  nand g89 (n_227, A[14], n_225);
  nand g90 (n_228, B[14], n_225);
  nand g91 (n_230, n_226, n_227, n_228);
  xor g92 (n_229, A[14], B[14]);
  xor g93 (Z[14], n_225, n_229);
  nand g94 (n_231, A[15], B[15]);
  nand g95 (n_232, A[15], n_230);
  nand g96 (n_233, B[15], n_230);
  nand g97 (n_235, n_231, n_232, n_233);
  xor g98 (n_234, A[15], B[15]);
  xor g99 (Z[15], n_230, n_234);
  nand g100 (n_236, A[16], B[16]);
  nand g101 (n_237, A[16], n_235);
  nand g102 (n_238, B[16], n_235);
  nand g103 (n_240, n_236, n_237, n_238);
  xor g104 (n_239, A[16], B[16]);
  xor g105 (Z[16], n_235, n_239);
  nand g106 (n_241, A[17], B[17]);
  nand g107 (n_242, A[17], n_240);
  nand g108 (n_243, B[17], n_240);
  nand g109 (n_245, n_241, n_242, n_243);
  xor g110 (n_244, A[17], B[17]);
  xor g111 (Z[17], n_240, n_244);
  nand g112 (n_246, A[18], B[18]);
  nand g113 (n_247, A[18], n_245);
  nand g114 (n_248, B[18], n_245);
  nand g115 (n_250, n_246, n_247, n_248);
  xor g116 (n_249, A[18], B[18]);
  xor g117 (Z[18], n_245, n_249);
  nand g118 (n_251, A[19], B[19]);
  nand g119 (n_252, A[19], n_250);
  nand g120 (n_253, B[19], n_250);
  nand g121 (n_255, n_251, n_252, n_253);
  xor g122 (n_254, A[19], B[19]);
  xor g123 (Z[19], n_250, n_254);
  nand g124 (n_256, A[20], B[20]);
  nand g125 (n_257, A[20], n_255);
  nand g126 (n_258, B[20], n_255);
  nand g127 (n_260, n_256, n_257, n_258);
  xor g128 (n_259, A[20], B[20]);
  xor g129 (Z[20], n_255, n_259);
  nand g130 (n_261, A[21], B[21]);
  nand g131 (n_262, A[21], n_260);
  nand g132 (n_263, B[21], n_260);
  nand g133 (n_265, n_261, n_262, n_263);
  xor g134 (n_264, A[21], B[21]);
  xor g135 (Z[21], n_260, n_264);
  nand g136 (n_266, A[22], B[22]);
  nand g137 (n_267, A[22], n_265);
  nand g138 (n_268, B[22], n_265);
  nand g139 (n_270, n_266, n_267, n_268);
  xor g140 (n_269, A[22], B[22]);
  xor g141 (Z[22], n_265, n_269);
  nand g142 (n_271, A[23], B[23]);
  nand g143 (n_272, A[23], n_270);
  nand g144 (n_273, B[23], n_270);
  nand g145 (n_275, n_271, n_272, n_273);
  xor g146 (n_274, A[23], B[23]);
  xor g147 (Z[23], n_270, n_274);
  nand g148 (n_276, A[24], B[24]);
  nand g149 (n_277, A[24], n_275);
  nand g150 (n_278, B[24], n_275);
  nand g151 (n_280, n_276, n_277, n_278);
  xor g152 (n_279, A[24], B[24]);
  xor g153 (Z[24], n_275, n_279);
  nand g154 (n_281, A[25], B[25]);
  nand g155 (n_282, A[25], n_280);
  nand g156 (n_283, B[25], n_280);
  nand g157 (n_285, n_281, n_282, n_283);
  xor g158 (n_284, A[25], B[25]);
  xor g159 (Z[25], n_280, n_284);
  nand g160 (n_286, A[26], B[26]);
  nand g161 (n_287, A[26], n_285);
  nand g162 (n_288, B[26], n_285);
  nand g163 (n_290, n_286, n_287, n_288);
  xor g164 (n_289, A[26], B[26]);
  xor g165 (Z[26], n_285, n_289);
  nand g166 (n_291, A[27], B[27]);
  nand g167 (n_292, A[27], n_290);
  nand g168 (n_293, B[27], n_290);
  nand g169 (n_295, n_291, n_292, n_293);
  xor g170 (n_294, A[27], B[27]);
  xor g171 (Z[27], n_290, n_294);
  nand g172 (n_296, A[28], B[28]);
  nand g173 (n_297, A[28], n_295);
  nand g174 (n_298, B[28], n_295);
  nand g175 (n_300, n_296, n_297, n_298);
  xor g176 (n_299, A[28], B[28]);
  xor g177 (Z[28], n_295, n_299);
  nand g178 (n_301, A[29], B[29]);
  nand g179 (n_302, A[29], n_300);
  nand g180 (n_303, B[29], n_300);
  nand g181 (n_305, n_301, n_302, n_303);
  xor g182 (n_304, A[29], B[29]);
  xor g183 (Z[29], n_300, n_304);
  nand g184 (n_306, A[30], B[30]);
  nand g185 (n_307, A[30], n_305);
  nand g186 (n_308, B[30], n_305);
  nand g187 (n_310, n_306, n_307, n_308);
  xor g188 (n_309, A[30], B[30]);
  xor g189 (Z[30], n_305, n_309);
  nand g190 (n_311, A[31], B[31]);
  nand g191 (n_312, A[31], n_310);
  nand g192 (n_313, B[31], n_310);
  nand g193 (n_315, n_311, n_312, n_313);
  xor g194 (n_314, A[31], B[31]);
  xor g195 (Z[31], n_310, n_314);
  nand g196 (n_316, A[32], B[32]);
  nand g197 (n_317, A[32], n_315);
  nand g198 (n_318, B[32], n_315);
  nand g199 (n_320, n_316, n_317, n_318);
  xor g200 (n_319, A[32], B[32]);
  xor g201 (Z[32], n_315, n_319);
  nand g202 (n_321, A[33], B[33]);
  nand g203 (n_322, A[33], n_320);
  nand g204 (n_323, B[33], n_320);
  nand g205 (n_325, n_321, n_322, n_323);
  xor g206 (n_324, A[33], B[33]);
  xor g207 (Z[33], n_320, n_324);
  nand g208 (n_326, A[34], B[34]);
  nand g209 (n_327, A[34], n_325);
  nand g210 (n_328, B[34], n_325);
  nand g211 (n_330, n_326, n_327, n_328);
  xor g212 (n_329, A[34], B[34]);
  xor g213 (Z[34], n_325, n_329);
  nand g214 (n_331, A[35], B[35]);
  nand g215 (n_332, A[35], n_330);
  nand g216 (n_333, B[35], n_330);
  nand g217 (n_335, n_331, n_332, n_333);
  xor g218 (n_334, A[35], B[35]);
  xor g219 (Z[35], n_330, n_334);
  nand g220 (n_336, A[36], B[36]);
  nand g221 (n_337, A[36], n_335);
  nand g222 (n_338, B[36], n_335);
  nand g223 (n_340, n_336, n_337, n_338);
  xor g224 (n_339, A[36], B[36]);
  xor g225 (Z[36], n_335, n_339);
  nand g226 (n_341, A[37], B[37]);
  nand g227 (n_342, A[37], n_340);
  nand g228 (n_343, B[37], n_340);
  nand g229 (n_345, n_341, n_342, n_343);
  xor g230 (n_344, A[37], B[37]);
  xor g231 (Z[37], n_340, n_344);
  nand g232 (n_346, A[38], B[38]);
  nand g233 (n_347, A[38], n_345);
  nand g234 (n_348, B[38], n_345);
  nand g235 (n_350, n_346, n_347, n_348);
  xor g236 (n_349, A[38], B[38]);
  xor g237 (Z[38], n_345, n_349);
  nand g238 (n_351, A[39], B[39]);
  nand g239 (n_352, A[39], n_350);
  nand g240 (n_353, B[39], n_350);
  nand g241 (n_355, n_351, n_352, n_353);
  xor g242 (n_354, A[39], B[39]);
  xor g243 (Z[39], n_350, n_354);
  nand g244 (n_356, A[40], B[40]);
  nand g245 (n_357, A[40], n_355);
  nand g246 (n_358, B[40], n_355);
  nand g247 (n_360, n_356, n_357, n_358);
  xor g248 (n_359, A[40], B[40]);
  xor g249 (Z[40], n_355, n_359);
  nand g250 (n_361, A[41], B[41]);
  nand g251 (n_362, A[41], n_360);
  nand g252 (n_363, B[41], n_360);
  nand g253 (n_365, n_361, n_362, n_363);
  xor g254 (n_364, A[41], B[41]);
  xor g255 (Z[41], n_360, n_364);
  nand g256 (n_366, A[42], B[42]);
  nand g257 (n_367, A[42], n_365);
  nand g258 (n_368, B[42], n_365);
  nand g259 (n_370, n_366, n_367, n_368);
  xor g260 (n_369, A[42], B[42]);
  xor g261 (Z[42], n_365, n_369);
  nand g262 (n_371, A[43], B[43]);
  nand g263 (n_372, A[43], n_370);
  nand g264 (n_373, B[43], n_370);
  nand g265 (n_375, n_371, n_372, n_373);
  xor g266 (n_374, A[43], B[43]);
  xor g267 (Z[43], n_370, n_374);
  nand g268 (n_376, A[44], B[44]);
  nand g269 (n_377, A[44], n_375);
  nand g270 (n_378, B[44], n_375);
  nand g271 (n_380, n_376, n_377, n_378);
  xor g272 (n_379, A[44], B[44]);
  xor g273 (Z[44], n_375, n_379);
  nand g274 (n_381, A[45], B[45]);
  nand g275 (n_382, A[45], n_380);
  nand g276 (n_383, B[45], n_380);
  nand g277 (n_385, n_381, n_382, n_383);
  xor g278 (n_384, A[45], B[45]);
  xor g279 (Z[45], n_380, n_384);
  nand g280 (n_386, A[46], B[46]);
  nand g281 (n_387, A[46], n_385);
  nand g282 (n_388, B[46], n_385);
  nand g283 (n_390, n_386, n_387, n_388);
  xor g284 (n_389, A[46], B[46]);
  xor g285 (Z[46], n_385, n_389);
  nand g286 (n_391, A[47], B[47]);
  nand g287 (n_392, A[47], n_390);
  nand g288 (n_393, B[47], n_390);
  nand g289 (n_395, n_391, n_392, n_393);
  xor g290 (n_394, A[47], B[47]);
  xor g291 (Z[47], n_390, n_394);
  nand g292 (n_396, A[48], B[48]);
  nand g293 (n_397, A[48], n_395);
  nand g294 (n_398, B[48], n_395);
  nand g295 (n_400, n_396, n_397, n_398);
  xor g296 (n_399, A[48], B[48]);
  xor g297 (Z[48], n_395, n_399);
  nand g301 (n_155, n_401, n_402, n_403);
  xor g303 (Z[49], n_400, n_404);
  or g305 (n_401, A[49], B[49]);
  xor g306 (n_404, A[49], B[49]);
  or g307 (n_162, wc, n_156);
  not gc (wc, A[1]);
  or g308 (n_163, wc0, n_156);
  not gc0 (wc0, B[1]);
  xnor g309 (Z[1], n_156, n_164);
  or g310 (n_402, A[49], wc1);
  not gc1 (wc1, n_400);
  or g311 (n_403, B[49], wc2);
  not gc2 (wc2, n_400);
endmodule

module add_signed_7719_1_GENERIC(A, B, Z);
  input [49:0] A, B;
  output [50:0] Z;
  wire [49:0] A, B;
  wire [50:0] Z;
  add_signed_7719_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_80_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [28:0] A, B;
  output [29:0] Z;
  wire [28:0] A, B;
  wire [29:0] Z;
  wire n_92, n_93, n_96, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_106, n_107, n_108, n_109, n_110, n_112, n_113;
  wire n_114, n_115, n_116, n_118, n_119, n_120, n_121, n_122;
  wire n_124, n_125, n_126, n_127, n_128, n_130, n_131, n_132;
  wire n_133, n_134, n_136, n_137, n_138, n_139, n_140, n_142;
  wire n_143, n_144, n_145, n_146, n_148, n_149, n_150, n_151;
  wire n_152, n_154, n_155, n_156, n_157, n_158, n_160, n_161;
  wire n_162, n_163, n_164, n_166, n_167, n_168, n_169, n_170;
  wire n_172, n_173, n_174, n_175, n_176, n_178, n_179, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_188, n_190, n_192;
  wire n_193, n_195, n_196, n_198, n_200, n_202, n_203, n_205;
  wire n_206, n_208, n_210, n_212, n_213, n_215, n_216, n_218;
  wire n_220, n_222, n_223, n_225, n_226, n_228, n_230, n_232;
  wire n_233, n_235, n_236, n_238, n_240, n_242, n_243, n_245;
  wire n_247, n_248, n_249, n_251, n_252, n_253, n_255, n_256;
  wire n_257, n_258, n_260, n_262, n_264, n_265, n_266, n_268;
  wire n_269, n_270, n_272, n_273, n_275, n_277, n_279, n_280;
  wire n_281, n_283, n_284, n_285, n_287, n_288, n_289, n_290;
  wire n_292, n_293, n_295, n_296, n_297, n_299, n_300, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_318, n_321;
  wire n_323, n_324, n_325, n_328, n_331, n_333, n_334, n_336;
  wire n_338, n_339, n_340, n_342, n_343, n_345, n_346, n_347;
  wire n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355;
  wire n_356, n_358, n_359, n_360, n_362, n_363, n_364, n_366;
  wire n_367, n_368, n_370, n_371, n_372, n_374, n_375, n_376;
  wire n_377, n_379, n_380, n_381, n_383, n_384, n_385, n_386;
  wire n_388, n_389, n_390, n_392, n_393, n_394, n_395, n_397;
  wire n_398, n_400, n_401, n_403, n_404, n_405, n_406, n_408;
  wire n_409, n_410, n_412, n_413, n_414, n_415, n_417, n_418;
  wire n_420, n_421, n_423, n_424, n_425, n_426, n_428, n_429;
  wire n_430, n_431, n_433, n_434, n_435, n_436, n_438, n_439;
  wire n_441, n_442;
  not g3 (Z[29], n_92);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_93, A[0], B[0]);
  nor g9 (n_96, A[1], B[1]);
  nand g10 (n_99, A[1], B[1]);
  nor g11 (n_106, A[2], B[2]);
  nand g12 (n_101, A[2], B[2]);
  nor g13 (n_102, A[3], B[3]);
  nand g14 (n_103, A[3], B[3]);
  nor g15 (n_112, A[4], B[4]);
  nand g16 (n_107, A[4], B[4]);
  nor g17 (n_108, A[5], B[5]);
  nand g18 (n_109, A[5], B[5]);
  nor g19 (n_118, A[6], B[6]);
  nand g20 (n_113, A[6], B[6]);
  nor g21 (n_114, A[7], B[7]);
  nand g22 (n_115, A[7], B[7]);
  nor g23 (n_124, A[8], B[8]);
  nand g24 (n_119, A[8], B[8]);
  nor g25 (n_120, A[9], B[9]);
  nand g26 (n_121, A[9], B[9]);
  nor g27 (n_130, A[10], B[10]);
  nand g28 (n_125, A[10], B[10]);
  nor g29 (n_126, A[11], B[11]);
  nand g30 (n_127, A[11], B[11]);
  nor g31 (n_136, A[12], B[12]);
  nand g32 (n_131, A[12], B[12]);
  nor g33 (n_132, A[13], B[13]);
  nand g34 (n_133, A[13], B[13]);
  nor g35 (n_142, A[14], B[14]);
  nand g36 (n_137, A[14], B[14]);
  nor g37 (n_138, A[15], B[15]);
  nand g38 (n_139, A[15], B[15]);
  nor g39 (n_148, A[16], B[16]);
  nand g40 (n_143, A[16], B[16]);
  nor g41 (n_144, A[17], B[17]);
  nand g42 (n_145, A[17], B[17]);
  nor g43 (n_154, A[18], B[18]);
  nand g44 (n_149, A[18], B[18]);
  nor g45 (n_150, A[19], B[19]);
  nand g46 (n_151, A[19], B[19]);
  nor g47 (n_160, A[20], B[20]);
  nand g48 (n_155, A[20], B[20]);
  nor g49 (n_156, A[21], B[21]);
  nand g50 (n_157, A[21], B[21]);
  nor g51 (n_166, A[22], B[22]);
  nand g52 (n_161, A[22], B[22]);
  nor g53 (n_162, A[23], B[23]);
  nand g54 (n_163, A[23], B[23]);
  nor g55 (n_172, A[24], B[24]);
  nand g56 (n_167, A[24], B[24]);
  nor g57 (n_168, A[25], B[25]);
  nand g58 (n_169, A[25], B[25]);
  nor g59 (n_178, A[26], B[26]);
  nand g60 (n_173, A[26], B[26]);
  nor g61 (n_174, A[27], B[27]);
  nand g62 (n_175, A[27], B[27]);
  nand g67 (n_179, n_99, n_100);
  nor g68 (n_104, n_101, n_102);
  nor g71 (n_182, n_106, n_102);
  nor g72 (n_110, n_107, n_108);
  nor g75 (n_188, n_112, n_108);
  nor g76 (n_116, n_113, n_114);
  nor g79 (n_190, n_118, n_114);
  nor g80 (n_122, n_119, n_120);
  nor g83 (n_198, n_124, n_120);
  nor g84 (n_128, n_125, n_126);
  nor g87 (n_200, n_130, n_126);
  nor g88 (n_134, n_131, n_132);
  nor g91 (n_208, n_136, n_132);
  nor g92 (n_140, n_137, n_138);
  nor g95 (n_210, n_142, n_138);
  nor g96 (n_146, n_143, n_144);
  nor g99 (n_218, n_148, n_144);
  nor g100 (n_152, n_149, n_150);
  nor g103 (n_220, n_154, n_150);
  nor g104 (n_158, n_155, n_156);
  nor g107 (n_228, n_160, n_156);
  nor g108 (n_164, n_161, n_162);
  nor g111 (n_230, n_166, n_162);
  nor g112 (n_170, n_167, n_168);
  nor g115 (n_238, n_172, n_168);
  nor g116 (n_176, n_173, n_174);
  nor g119 (n_240, n_178, n_174);
  nand g122 (n_379, n_101, n_181);
  nand g123 (n_184, n_182, n_179);
  nand g124 (n_245, n_183, n_184);
  nor g125 (n_186, n_118, n_185);
  nand g134 (n_253, n_188, n_190);
  nor g135 (n_196, n_130, n_195);
  nand g144 (n_260, n_198, n_200);
  nor g145 (n_206, n_142, n_205);
  nand g154 (n_268, n_208, n_210);
  nor g155 (n_216, n_154, n_215);
  nand g164 (n_275, n_218, n_220);
  nor g165 (n_226, n_166, n_225);
  nand g174 (n_283, n_228, n_230);
  nor g175 (n_236, n_178, n_235);
  nand g184 (n_292, n_238, n_240);
  nand g187 (n_383, n_107, n_247);
  nand g188 (n_248, n_188, n_245);
  nand g189 (n_385, n_185, n_248);
  nand g192 (n_388, n_251, n_252);
  nand g195 (n_293, n_255, n_256);
  nor g196 (n_258, n_136, n_257);
  nor g199 (n_303, n_136, n_260);
  nor g205 (n_266, n_264, n_257);
  nor g208 (n_309, n_260, n_264);
  nor g209 (n_270, n_268, n_257);
  nor g212 (n_312, n_260, n_268);
  nor g213 (n_273, n_160, n_272);
  nor g216 (n_346, n_160, n_275);
  nor g222 (n_281, n_279, n_272);
  nor g225 (n_352, n_275, n_279);
  nor g226 (n_285, n_283, n_272);
  nor g229 (n_318, n_275, n_283);
  nor g230 (n_290, n_287, n_288);
  nor g233 (n_331, n_287, n_292);
  nand g236 (n_392, n_119, n_295);
  nand g237 (n_296, n_198, n_293);
  nand g238 (n_394, n_195, n_296);
  nand g241 (n_397, n_299, n_300);
  nand g244 (n_400, n_257, n_302);
  nand g245 (n_305, n_303, n_293);
  nand g246 (n_403, n_304, n_305);
  nand g247 (n_308, n_306, n_293);
  nand g248 (n_405, n_307, n_308);
  nand g249 (n_311, n_309, n_293);
  nand g250 (n_408, n_310, n_311);
  nand g251 (n_314, n_312, n_293);
  nand g252 (n_336, n_313, n_314);
  nor g253 (n_316, n_172, n_315);
  nand g262 (n_360, n_238, n_318);
  nor g263 (n_325, n_323, n_315);
  nor g268 (n_328, n_292, n_315);
  nand g277 (n_372, n_318, n_331);
  nand g280 (n_412, n_143, n_338);
  nand g281 (n_339, n_218, n_336);
  nand g282 (n_414, n_215, n_339);
  nand g285 (n_417, n_342, n_343);
  nand g288 (n_420, n_272, n_345);
  nand g289 (n_348, n_346, n_336);
  nand g290 (n_423, n_347, n_348);
  nand g291 (n_351, n_349, n_336);
  nand g292 (n_425, n_350, n_351);
  nand g293 (n_354, n_352, n_336);
  nand g294 (n_428, n_353, n_354);
  nand g295 (n_355, n_318, n_336);
  nand g296 (n_430, n_315, n_355);
  nand g299 (n_433, n_358, n_359);
  nand g302 (n_435, n_362, n_363);
  nand g305 (n_438, n_366, n_367);
  nand g308 (n_441, n_370, n_371);
  nand g311 (n_92, n_374, n_375);
  xnor g315 (Z[2], n_179, n_377);
  xnor g318 (Z[3], n_379, n_380);
  xnor g320 (Z[4], n_245, n_381);
  xnor g323 (Z[5], n_383, n_384);
  xnor g325 (Z[6], n_385, n_386);
  xnor g328 (Z[7], n_388, n_389);
  xnor g330 (Z[8], n_293, n_390);
  xnor g333 (Z[9], n_392, n_393);
  xnor g335 (Z[10], n_394, n_395);
  xnor g338 (Z[11], n_397, n_398);
  xnor g341 (Z[12], n_400, n_401);
  xnor g344 (Z[13], n_403, n_404);
  xnor g346 (Z[14], n_405, n_406);
  xnor g349 (Z[15], n_408, n_409);
  xnor g351 (Z[16], n_336, n_410);
  xnor g354 (Z[17], n_412, n_413);
  xnor g356 (Z[18], n_414, n_415);
  xnor g359 (Z[19], n_417, n_418);
  xnor g362 (Z[20], n_420, n_421);
  xnor g365 (Z[21], n_423, n_424);
  xnor g367 (Z[22], n_425, n_426);
  xnor g370 (Z[23], n_428, n_429);
  xnor g372 (Z[24], n_430, n_431);
  xnor g375 (Z[25], n_433, n_434);
  xnor g377 (Z[26], n_435, n_436);
  xnor g380 (Z[27], n_438, n_439);
  xnor g383 (Z[28], n_441, n_442);
  and g386 (n_287, A[28], B[28]);
  or g387 (n_289, A[28], B[28]);
  and g388 (n_215, wc, n_145);
  not gc (wc, n_146);
  and g389 (n_222, wc0, n_151);
  not gc0 (wc0, n_152);
  and g390 (n_225, wc1, n_157);
  not gc1 (wc1, n_158);
  and g391 (n_232, wc2, n_163);
  not gc2 (wc2, n_164);
  and g392 (n_235, wc3, n_169);
  not gc3 (wc3, n_170);
  and g393 (n_242, wc4, n_175);
  not gc4 (wc4, n_176);
  and g394 (n_195, wc5, n_121);
  not gc5 (wc5, n_122);
  and g395 (n_202, wc6, n_127);
  not gc6 (wc6, n_128);
  and g396 (n_205, wc7, n_133);
  not gc7 (wc7, n_134);
  and g397 (n_212, wc8, n_139);
  not gc8 (wc8, n_140);
  and g398 (n_185, wc9, n_109);
  not gc9 (wc9, n_110);
  and g399 (n_192, wc10, n_115);
  not gc10 (wc10, n_116);
  and g400 (n_183, wc11, n_103);
  not gc11 (wc11, n_104);
  or g401 (n_100, n_93, n_96);
  or g402 (n_249, wc12, n_118);
  not gc12 (wc12, n_188);
  or g403 (n_297, wc13, n_130);
  not gc13 (wc13, n_198);
  or g404 (n_264, wc14, n_142);
  not gc14 (wc14, n_208);
  or g405 (n_340, wc15, n_154);
  not gc15 (wc15, n_218);
  or g406 (n_279, wc16, n_166);
  not gc16 (wc16, n_228);
  or g407 (n_323, wc17, n_178);
  not gc17 (wc17, n_238);
  or g408 (n_376, wc18, n_96);
  not gc18 (wc18, n_99);
  or g409 (n_377, wc19, n_106);
  not gc19 (wc19, n_101);
  or g410 (n_380, wc20, n_102);
  not gc20 (wc20, n_103);
  or g411 (n_381, wc21, n_112);
  not gc21 (wc21, n_107);
  or g412 (n_384, wc22, n_108);
  not gc22 (wc22, n_109);
  or g413 (n_386, wc23, n_118);
  not gc23 (wc23, n_113);
  or g414 (n_389, wc24, n_114);
  not gc24 (wc24, n_115);
  or g415 (n_390, wc25, n_124);
  not gc25 (wc25, n_119);
  or g416 (n_393, wc26, n_120);
  not gc26 (wc26, n_121);
  or g417 (n_395, wc27, n_130);
  not gc27 (wc27, n_125);
  or g418 (n_398, wc28, n_126);
  not gc28 (wc28, n_127);
  or g419 (n_401, wc29, n_136);
  not gc29 (wc29, n_131);
  or g420 (n_404, wc30, n_132);
  not gc30 (wc30, n_133);
  or g421 (n_406, wc31, n_142);
  not gc31 (wc31, n_137);
  or g422 (n_409, wc32, n_138);
  not gc32 (wc32, n_139);
  or g423 (n_410, wc33, n_148);
  not gc33 (wc33, n_143);
  or g424 (n_413, wc34, n_144);
  not gc34 (wc34, n_145);
  or g425 (n_415, wc35, n_154);
  not gc35 (wc35, n_149);
  or g426 (n_418, wc36, n_150);
  not gc36 (wc36, n_151);
  or g427 (n_421, wc37, n_160);
  not gc37 (wc37, n_155);
  or g428 (n_424, wc38, n_156);
  not gc38 (wc38, n_157);
  or g429 (n_426, wc39, n_166);
  not gc39 (wc39, n_161);
  or g430 (n_429, wc40, n_162);
  not gc40 (wc40, n_163);
  or g431 (n_431, wc41, n_172);
  not gc41 (wc41, n_167);
  or g432 (n_434, wc42, n_168);
  not gc42 (wc42, n_169);
  or g433 (n_436, wc43, n_178);
  not gc43 (wc43, n_173);
  or g434 (n_439, wc44, n_174);
  not gc44 (wc44, n_175);
  and g435 (n_223, wc45, n_220);
  not gc45 (wc45, n_215);
  and g436 (n_233, wc46, n_230);
  not gc46 (wc46, n_225);
  and g437 (n_243, wc47, n_240);
  not gc47 (wc47, n_235);
  and g438 (n_203, wc48, n_200);
  not gc48 (wc48, n_195);
  and g439 (n_213, wc49, n_210);
  not gc49 (wc49, n_205);
  and g440 (n_193, wc50, n_190);
  not gc50 (wc50, n_185);
  and g441 (n_306, wc51, n_208);
  not gc51 (wc51, n_260);
  and g442 (n_349, wc52, n_228);
  not gc52 (wc52, n_275);
  xor g443 (Z[1], n_93, n_376);
  or g444 (n_442, wc53, n_287);
  not gc53 (wc53, n_289);
  and g445 (n_272, wc54, n_222);
  not gc54 (wc54, n_223);
  and g446 (n_284, wc55, n_232);
  not gc55 (wc55, n_233);
  and g447 (n_288, wc56, n_242);
  not gc56 (wc56, n_243);
  and g448 (n_257, wc57, n_202);
  not gc57 (wc57, n_203);
  and g449 (n_269, wc58, n_212);
  not gc58 (wc58, n_213);
  and g450 (n_255, wc59, n_192);
  not gc59 (wc59, n_193);
  or g451 (n_181, wc60, n_106);
  not gc60 (wc60, n_179);
  and g452 (n_251, wc61, n_113);
  not gc61 (wc61, n_186);
  and g453 (n_299, wc62, n_125);
  not gc62 (wc62, n_196);
  and g454 (n_265, wc63, n_137);
  not gc63 (wc63, n_206);
  and g455 (n_342, wc64, n_149);
  not gc64 (wc64, n_216);
  and g456 (n_280, wc65, n_161);
  not gc65 (wc65, n_226);
  and g457 (n_324, wc66, n_173);
  not gc66 (wc66, n_236);
  or g458 (n_356, wc67, n_172);
  not gc67 (wc67, n_318);
  or g459 (n_364, n_323, wc68);
  not gc68 (wc68, n_318);
  or g460 (n_368, wc69, n_292);
  not gc69 (wc69, n_318);
  and g461 (n_262, wc70, n_208);
  not gc70 (wc70, n_257);
  and g462 (n_277, wc71, n_228);
  not gc71 (wc71, n_272);
  and g463 (n_315, n_284, wc72);
  not gc72 (wc72, n_285);
  and g464 (n_333, n_289, wc73);
  not gc73 (wc73, n_290);
  and g465 (n_313, n_269, wc74);
  not gc74 (wc74, n_270);
  or g466 (n_256, n_253, wc75);
  not gc75 (wc75, n_245);
  or g467 (n_247, wc76, n_112);
  not gc76 (wc76, n_245);
  or g468 (n_252, n_249, wc77);
  not gc77 (wc77, n_245);
  and g469 (n_304, wc78, n_131);
  not gc78 (wc78, n_258);
  and g470 (n_307, wc79, n_205);
  not gc79 (wc79, n_262);
  and g471 (n_310, n_265, wc80);
  not gc80 (wc80, n_266);
  and g472 (n_347, wc81, n_155);
  not gc81 (wc81, n_273);
  and g473 (n_350, wc82, n_225);
  not gc82 (wc82, n_277);
  and g474 (n_353, n_280, wc83);
  not gc83 (wc83, n_281);
  and g475 (n_334, wc84, n_331);
  not gc84 (wc84, n_315);
  and g476 (n_321, wc85, n_238);
  not gc85 (wc85, n_315);
  and g477 (n_374, wc86, n_333);
  not gc86 (wc86, n_334);
  or g478 (n_295, wc87, n_124);
  not gc87 (wc87, n_293);
  or g479 (n_300, n_297, wc88);
  not gc88 (wc88, n_293);
  or g480 (n_302, wc89, n_260);
  not gc89 (wc89, n_293);
  and g481 (n_358, wc90, n_167);
  not gc90 (wc90, n_316);
  and g482 (n_362, wc91, n_235);
  not gc91 (wc91, n_321);
  and g483 (n_366, n_324, wc92);
  not gc92 (wc92, n_325);
  and g484 (n_370, n_288, wc93);
  not gc93 (wc93, n_328);
  or g485 (n_375, n_372, wc94);
  not gc94 (wc94, n_336);
  or g486 (n_338, wc95, n_148);
  not gc95 (wc95, n_336);
  or g487 (n_343, n_340, wc96);
  not gc96 (wc96, n_336);
  or g488 (n_345, wc97, n_275);
  not gc97 (wc97, n_336);
  or g489 (n_359, n_356, wc98);
  not gc98 (wc98, n_336);
  or g490 (n_363, n_360, wc99);
  not gc99 (wc99, n_336);
  or g491 (n_367, n_364, wc100);
  not gc100 (wc100, n_336);
  or g492 (n_371, n_368, wc101);
  not gc101 (wc101, n_336);
endmodule

module add_signed_80_GENERIC(A, B, Z);
  input [28:0] A, B;
  output [29:0] Z;
  wire [28:0] A, B;
  wire [29:0] Z;
  add_signed_80_GENERIC_REAL g1(.A ({A[27], A[27:0]}), .B ({B[27],
       B[27:0]}), .Z (Z));
endmodule

module add_signed_8959_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [20:0] A, B;
  output [18:0] Z;
  wire [20:0] A, B;
  wire [18:0] Z;
  wire n_64, n_66, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_76, n_77, n_78, n_79, n_80, n_82, n_83, n_84;
  wire n_85, n_86, n_88, n_89, n_90, n_91, n_92, n_94;
  wire n_95, n_96, n_97, n_98, n_100, n_101, n_102, n_103;
  wire n_104, n_106, n_107, n_108, n_109, n_110, n_112, n_113;
  wire n_114, n_115, n_116, n_118, n_119, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_128, n_130, n_132, n_133, n_135;
  wire n_136, n_138, n_140, n_142, n_143, n_145, n_146, n_148;
  wire n_150, n_152, n_153, n_155, n_156, n_157, n_160, n_162;
  wire n_164, n_165, n_166, n_168, n_169, n_170, n_172, n_173;
  wire n_174, n_175, n_177, n_179, n_181, n_182, n_183, n_185;
  wire n_186, n_187, n_189, n_191, n_192, n_193, n_195, n_196;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_213, n_214;
  wire n_219, n_220, n_222, n_223, n_224, n_226, n_227, n_228;
  wire n_229, n_231, n_232, n_233, n_235, n_236, n_237, n_238;
  wire n_240, n_241, n_243, n_244, n_246, n_247, n_248, n_249;
  wire n_251, n_252, n_253, n_255, n_256, n_257, n_258;
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_64, A[0], B[0]);
  nor g9 (n_66, A[1], B[1]);
  nand g10 (n_69, A[1], B[1]);
  nor g11 (n_76, A[2], B[2]);
  nand g12 (n_71, A[2], B[2]);
  nor g13 (n_72, A[3], B[3]);
  nand g14 (n_73, A[3], B[3]);
  nor g15 (n_82, A[4], B[4]);
  nand g16 (n_77, A[4], B[4]);
  nor g17 (n_78, A[5], B[5]);
  nand g18 (n_79, A[5], B[5]);
  nor g19 (n_88, A[6], B[6]);
  nand g20 (n_83, A[6], B[6]);
  nor g21 (n_84, A[7], B[7]);
  nand g22 (n_85, A[7], B[7]);
  nor g23 (n_94, A[8], B[8]);
  nand g24 (n_89, A[8], B[8]);
  nor g25 (n_90, A[9], B[9]);
  nand g26 (n_91, A[9], B[9]);
  nor g27 (n_100, A[10], B[10]);
  nand g28 (n_95, A[10], B[10]);
  nor g29 (n_96, A[11], B[11]);
  nand g30 (n_97, A[11], B[11]);
  nor g31 (n_106, A[12], B[12]);
  nand g32 (n_101, A[12], B[12]);
  nor g33 (n_102, A[13], B[13]);
  nand g34 (n_103, A[13], B[13]);
  nor g35 (n_112, A[14], B[14]);
  nand g36 (n_107, A[14], B[14]);
  nor g37 (n_108, A[15], B[15]);
  nand g38 (n_109, A[15], B[15]);
  nor g39 (n_118, A[16], B[16]);
  nand g40 (n_113, A[16], B[16]);
  nor g41 (n_114, A[17], B[17]);
  nand g42 (n_115, A[17], B[17]);
  nand g47 (n_119, n_69, n_70);
  nor g48 (n_74, n_71, n_72);
  nor g51 (n_122, n_76, n_72);
  nor g52 (n_80, n_77, n_78);
  nor g55 (n_128, n_82, n_78);
  nor g56 (n_86, n_83, n_84);
  nor g59 (n_130, n_88, n_84);
  nor g60 (n_92, n_89, n_90);
  nor g63 (n_138, n_94, n_90);
  nor g64 (n_98, n_95, n_96);
  nor g67 (n_140, n_100, n_96);
  nor g68 (n_104, n_101, n_102);
  nor g71 (n_148, n_106, n_102);
  nor g72 (n_110, n_107, n_108);
  nor g75 (n_150, n_112, n_108);
  nor g76 (n_116, n_113, n_114);
  nor g79 (n_160, n_118, n_114);
  nand g82 (n_222, n_71, n_121);
  nand g83 (n_124, n_122, n_119);
  nand g84 (n_162, n_123, n_124);
  nor g85 (n_126, n_88, n_125);
  nand g94 (n_170, n_128, n_130);
  nor g95 (n_136, n_100, n_135);
  nand g104 (n_177, n_138, n_140);
  nor g105 (n_146, n_112, n_145);
  nand g114 (n_185, n_148, n_150);
  nand g122 (n_226, n_77, n_164);
  nand g123 (n_165, n_128, n_162);
  nand g124 (n_228, n_125, n_165);
  nand g127 (n_231, n_168, n_169);
  nand g130 (n_189, n_172, n_173);
  nor g131 (n_175, n_106, n_174);
  nor g134 (n_199, n_106, n_177);
  nor g140 (n_183, n_181, n_174);
  nor g143 (n_205, n_177, n_181);
  nor g144 (n_187, n_185, n_174);
  nor g147 (n_208, n_177, n_185);
  nand g150 (n_235, n_89, n_191);
  nand g151 (n_192, n_138, n_189);
  nand g152 (n_237, n_135, n_192);
  nand g155 (n_240, n_195, n_196);
  nand g158 (n_243, n_174, n_198);
  nand g159 (n_201, n_199, n_189);
  nand g160 (n_246, n_200, n_201);
  nand g161 (n_204, n_202, n_189);
  nand g162 (n_248, n_203, n_204);
  nand g163 (n_207, n_205, n_189);
  nand g164 (n_251, n_206, n_207);
  nand g165 (n_210, n_208, n_189);
  nand g166 (n_211, n_209, n_210);
  nand g169 (n_255, n_113, n_213);
  nand g170 (n_214, n_160, n_211);
  nand g171 (n_257, n_156, n_214);
  xnor g178 (Z[2], n_119, n_220);
  xnor g181 (Z[3], n_222, n_223);
  xnor g183 (Z[4], n_162, n_224);
  xnor g186 (Z[5], n_226, n_227);
  xnor g188 (Z[6], n_228, n_229);
  xnor g191 (Z[7], n_231, n_232);
  xnor g193 (Z[8], n_189, n_233);
  xnor g196 (Z[9], n_235, n_236);
  xnor g198 (Z[10], n_237, n_238);
  xnor g201 (Z[11], n_240, n_241);
  xnor g204 (Z[12], n_243, n_244);
  xnor g207 (Z[13], n_246, n_247);
  xnor g209 (Z[14], n_248, n_249);
  xnor g212 (Z[15], n_251, n_252);
  xnor g214 (Z[16], n_211, n_253);
  xnor g217 (Z[17], n_255, n_256);
  xnor g219 (Z[18], n_257, n_258);
  and g222 (n_155, A[18], B[18]);
  or g223 (n_157, A[18], B[18]);
  or g224 (n_70, n_64, n_66);
  and g225 (n_123, wc, n_73);
  not gc (wc, n_74);
  and g226 (n_125, wc0, n_79);
  not gc0 (wc0, n_80);
  and g227 (n_132, wc1, n_85);
  not gc1 (wc1, n_86);
  and g228 (n_135, wc2, n_91);
  not gc2 (wc2, n_92);
  and g229 (n_142, wc3, n_97);
  not gc3 (wc3, n_98);
  and g230 (n_145, wc4, n_103);
  not gc4 (wc4, n_104);
  and g231 (n_152, wc5, n_109);
  not gc5 (wc5, n_110);
  and g232 (n_156, wc6, n_115);
  not gc6 (wc6, n_116);
  or g233 (n_166, wc7, n_88);
  not gc7 (wc7, n_128);
  or g234 (n_193, wc8, n_100);
  not gc8 (wc8, n_138);
  or g235 (n_181, wc9, n_112);
  not gc9 (wc9, n_148);
  or g236 (n_219, wc10, n_66);
  not gc10 (wc10, n_69);
  or g237 (n_220, wc11, n_76);
  not gc11 (wc11, n_71);
  or g238 (n_223, wc12, n_72);
  not gc12 (wc12, n_73);
  or g239 (n_224, wc13, n_82);
  not gc13 (wc13, n_77);
  or g240 (n_227, wc14, n_78);
  not gc14 (wc14, n_79);
  or g241 (n_229, wc15, n_88);
  not gc15 (wc15, n_83);
  or g242 (n_232, wc16, n_84);
  not gc16 (wc16, n_85);
  or g243 (n_233, wc17, n_94);
  not gc17 (wc17, n_89);
  or g244 (n_236, wc18, n_90);
  not gc18 (wc18, n_91);
  or g245 (n_238, wc19, n_100);
  not gc19 (wc19, n_95);
  or g246 (n_241, wc20, n_96);
  not gc20 (wc20, n_97);
  or g247 (n_244, wc21, n_106);
  not gc21 (wc21, n_101);
  or g248 (n_247, wc22, n_102);
  not gc22 (wc22, n_103);
  or g249 (n_249, wc23, n_112);
  not gc23 (wc23, n_107);
  or g250 (n_252, wc24, n_108);
  not gc24 (wc24, n_109);
  or g251 (n_253, wc25, n_118);
  not gc25 (wc25, n_113);
  or g252 (n_256, wc26, n_114);
  not gc26 (wc26, n_115);
  and g253 (n_133, wc27, n_130);
  not gc27 (wc27, n_125);
  and g254 (n_143, wc28, n_140);
  not gc28 (wc28, n_135);
  and g255 (n_153, wc29, n_150);
  not gc29 (wc29, n_145);
  and g256 (n_202, wc30, n_148);
  not gc30 (wc30, n_177);
  xor g257 (Z[1], n_64, n_219);
  or g258 (n_258, wc31, n_155);
  not gc31 (wc31, n_157);
  or g259 (n_121, wc32, n_76);
  not gc32 (wc32, n_119);
  and g260 (n_168, wc33, n_83);
  not gc33 (wc33, n_126);
  and g261 (n_172, wc34, n_132);
  not gc34 (wc34, n_133);
  and g262 (n_195, wc35, n_95);
  not gc35 (wc35, n_136);
  and g263 (n_174, wc36, n_142);
  not gc36 (wc36, n_143);
  and g264 (n_182, wc37, n_107);
  not gc37 (wc37, n_146);
  and g265 (n_186, wc38, n_152);
  not gc38 (wc38, n_153);
  and g266 (n_179, wc39, n_148);
  not gc39 (wc39, n_174);
  or g267 (n_164, wc40, n_82);
  not gc40 (wc40, n_162);
  or g268 (n_169, n_166, wc41);
  not gc41 (wc41, n_162);
  or g269 (n_173, n_170, wc42);
  not gc42 (wc42, n_162);
  and g270 (n_200, wc43, n_101);
  not gc43 (wc43, n_175);
  and g271 (n_203, wc44, n_145);
  not gc44 (wc44, n_179);
  and g272 (n_206, n_182, wc45);
  not gc45 (wc45, n_183);
  and g273 (n_209, n_186, wc46);
  not gc46 (wc46, n_187);
  or g274 (n_191, wc47, n_94);
  not gc47 (wc47, n_189);
  or g275 (n_196, n_193, wc48);
  not gc48 (wc48, n_189);
  or g276 (n_198, wc49, n_177);
  not gc49 (wc49, n_189);
  or g277 (n_213, wc50, n_118);
  not gc50 (wc50, n_211);
endmodule

module add_signed_8959_GENERIC(A, B, Z);
  input [20:0] A, B;
  output [18:0] Z;
  wire [20:0] A, B;
  wire [18:0] Z;
  add_signed_8959_GENERIC_REAL g1(.A (A), .B ({B[20:19], B[17],
       B[17:0]}), .Z (Z));
endmodule

module add_signed_8959_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [20:0] A, B;
  output [18:0] Z;
  wire [20:0] A, B;
  wire [18:0] Z;
  wire n_64, n_66, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_76, n_77, n_78, n_79, n_80, n_82, n_83, n_84;
  wire n_85, n_86, n_88, n_89, n_90, n_91, n_92, n_94;
  wire n_95, n_96, n_97, n_98, n_100, n_101, n_102, n_103;
  wire n_104, n_106, n_107, n_108, n_109, n_110, n_112, n_113;
  wire n_114, n_115, n_116, n_118, n_119, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_128, n_130, n_132, n_133, n_135;
  wire n_136, n_138, n_140, n_142, n_143, n_145, n_146, n_148;
  wire n_150, n_152, n_153, n_155, n_156, n_157, n_160, n_162;
  wire n_164, n_165, n_166, n_168, n_169, n_170, n_172, n_173;
  wire n_174, n_175, n_177, n_179, n_181, n_182, n_183, n_185;
  wire n_186, n_187, n_189, n_191, n_192, n_193, n_195, n_196;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_213, n_214;
  wire n_219, n_220, n_222, n_223, n_224, n_226, n_227, n_228;
  wire n_229, n_231, n_232, n_233, n_235, n_236, n_237, n_238;
  wire n_240, n_241, n_243, n_244, n_246, n_247, n_248, n_249;
  wire n_251, n_252, n_253, n_255, n_256, n_257, n_258;
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_64, A[0], B[0]);
  nor g9 (n_66, A[1], B[1]);
  nand g10 (n_69, A[1], B[1]);
  nor g11 (n_76, A[2], B[2]);
  nand g12 (n_71, A[2], B[2]);
  nor g13 (n_72, A[3], B[3]);
  nand g14 (n_73, A[3], B[3]);
  nor g15 (n_82, A[4], B[4]);
  nand g16 (n_77, A[4], B[4]);
  nor g17 (n_78, A[5], B[5]);
  nand g18 (n_79, A[5], B[5]);
  nor g19 (n_88, A[6], B[6]);
  nand g20 (n_83, A[6], B[6]);
  nor g21 (n_84, A[7], B[7]);
  nand g22 (n_85, A[7], B[7]);
  nor g23 (n_94, A[8], B[8]);
  nand g24 (n_89, A[8], B[8]);
  nor g25 (n_90, A[9], B[9]);
  nand g26 (n_91, A[9], B[9]);
  nor g27 (n_100, A[10], B[10]);
  nand g28 (n_95, A[10], B[10]);
  nor g29 (n_96, A[11], B[11]);
  nand g30 (n_97, A[11], B[11]);
  nor g31 (n_106, A[12], B[12]);
  nand g32 (n_101, A[12], B[12]);
  nor g33 (n_102, A[13], B[13]);
  nand g34 (n_103, A[13], B[13]);
  nor g35 (n_112, A[14], B[14]);
  nand g36 (n_107, A[14], B[14]);
  nor g37 (n_108, A[15], B[15]);
  nand g38 (n_109, A[15], B[15]);
  nor g39 (n_118, A[16], B[16]);
  nand g40 (n_113, A[16], B[16]);
  nor g41 (n_114, A[17], B[17]);
  nand g42 (n_115, A[17], B[17]);
  nand g47 (n_119, n_69, n_70);
  nor g48 (n_74, n_71, n_72);
  nor g51 (n_122, n_76, n_72);
  nor g52 (n_80, n_77, n_78);
  nor g55 (n_128, n_82, n_78);
  nor g56 (n_86, n_83, n_84);
  nor g59 (n_130, n_88, n_84);
  nor g60 (n_92, n_89, n_90);
  nor g63 (n_138, n_94, n_90);
  nor g64 (n_98, n_95, n_96);
  nor g67 (n_140, n_100, n_96);
  nor g68 (n_104, n_101, n_102);
  nor g71 (n_148, n_106, n_102);
  nor g72 (n_110, n_107, n_108);
  nor g75 (n_150, n_112, n_108);
  nor g76 (n_116, n_113, n_114);
  nor g79 (n_160, n_118, n_114);
  nand g82 (n_222, n_71, n_121);
  nand g83 (n_124, n_122, n_119);
  nand g84 (n_162, n_123, n_124);
  nor g85 (n_126, n_88, n_125);
  nand g94 (n_170, n_128, n_130);
  nor g95 (n_136, n_100, n_135);
  nand g104 (n_177, n_138, n_140);
  nor g105 (n_146, n_112, n_145);
  nand g114 (n_185, n_148, n_150);
  nand g122 (n_226, n_77, n_164);
  nand g123 (n_165, n_128, n_162);
  nand g124 (n_228, n_125, n_165);
  nand g127 (n_231, n_168, n_169);
  nand g130 (n_189, n_172, n_173);
  nor g131 (n_175, n_106, n_174);
  nor g134 (n_199, n_106, n_177);
  nor g140 (n_183, n_181, n_174);
  nor g143 (n_205, n_177, n_181);
  nor g144 (n_187, n_185, n_174);
  nor g147 (n_208, n_177, n_185);
  nand g150 (n_235, n_89, n_191);
  nand g151 (n_192, n_138, n_189);
  nand g152 (n_237, n_135, n_192);
  nand g155 (n_240, n_195, n_196);
  nand g158 (n_243, n_174, n_198);
  nand g159 (n_201, n_199, n_189);
  nand g160 (n_246, n_200, n_201);
  nand g161 (n_204, n_202, n_189);
  nand g162 (n_248, n_203, n_204);
  nand g163 (n_207, n_205, n_189);
  nand g164 (n_251, n_206, n_207);
  nand g165 (n_210, n_208, n_189);
  nand g166 (n_211, n_209, n_210);
  nand g169 (n_255, n_113, n_213);
  nand g170 (n_214, n_160, n_211);
  nand g171 (n_257, n_156, n_214);
  xnor g178 (Z[2], n_119, n_220);
  xnor g181 (Z[3], n_222, n_223);
  xnor g183 (Z[4], n_162, n_224);
  xnor g186 (Z[5], n_226, n_227);
  xnor g188 (Z[6], n_228, n_229);
  xnor g191 (Z[7], n_231, n_232);
  xnor g193 (Z[8], n_189, n_233);
  xnor g196 (Z[9], n_235, n_236);
  xnor g198 (Z[10], n_237, n_238);
  xnor g201 (Z[11], n_240, n_241);
  xnor g204 (Z[12], n_243, n_244);
  xnor g207 (Z[13], n_246, n_247);
  xnor g209 (Z[14], n_248, n_249);
  xnor g212 (Z[15], n_251, n_252);
  xnor g214 (Z[16], n_211, n_253);
  xnor g217 (Z[17], n_255, n_256);
  xnor g219 (Z[18], n_257, n_258);
  and g222 (n_155, A[18], B[18]);
  or g223 (n_157, A[18], B[18]);
  or g224 (n_70, n_64, n_66);
  and g225 (n_123, wc, n_73);
  not gc (wc, n_74);
  and g226 (n_125, wc0, n_79);
  not gc0 (wc0, n_80);
  and g227 (n_132, wc1, n_85);
  not gc1 (wc1, n_86);
  and g228 (n_135, wc2, n_91);
  not gc2 (wc2, n_92);
  and g229 (n_142, wc3, n_97);
  not gc3 (wc3, n_98);
  and g230 (n_145, wc4, n_103);
  not gc4 (wc4, n_104);
  and g231 (n_152, wc5, n_109);
  not gc5 (wc5, n_110);
  and g232 (n_156, wc6, n_115);
  not gc6 (wc6, n_116);
  or g233 (n_166, wc7, n_88);
  not gc7 (wc7, n_128);
  or g234 (n_193, wc8, n_100);
  not gc8 (wc8, n_138);
  or g235 (n_181, wc9, n_112);
  not gc9 (wc9, n_148);
  or g236 (n_219, wc10, n_66);
  not gc10 (wc10, n_69);
  or g237 (n_220, wc11, n_76);
  not gc11 (wc11, n_71);
  or g238 (n_223, wc12, n_72);
  not gc12 (wc12, n_73);
  or g239 (n_224, wc13, n_82);
  not gc13 (wc13, n_77);
  or g240 (n_227, wc14, n_78);
  not gc14 (wc14, n_79);
  or g241 (n_229, wc15, n_88);
  not gc15 (wc15, n_83);
  or g242 (n_232, wc16, n_84);
  not gc16 (wc16, n_85);
  or g243 (n_233, wc17, n_94);
  not gc17 (wc17, n_89);
  or g244 (n_236, wc18, n_90);
  not gc18 (wc18, n_91);
  or g245 (n_238, wc19, n_100);
  not gc19 (wc19, n_95);
  or g246 (n_241, wc20, n_96);
  not gc20 (wc20, n_97);
  or g247 (n_244, wc21, n_106);
  not gc21 (wc21, n_101);
  or g248 (n_247, wc22, n_102);
  not gc22 (wc22, n_103);
  or g249 (n_249, wc23, n_112);
  not gc23 (wc23, n_107);
  or g250 (n_252, wc24, n_108);
  not gc24 (wc24, n_109);
  or g251 (n_253, wc25, n_118);
  not gc25 (wc25, n_113);
  or g252 (n_256, wc26, n_114);
  not gc26 (wc26, n_115);
  and g253 (n_133, wc27, n_130);
  not gc27 (wc27, n_125);
  and g254 (n_143, wc28, n_140);
  not gc28 (wc28, n_135);
  and g255 (n_153, wc29, n_150);
  not gc29 (wc29, n_145);
  and g256 (n_202, wc30, n_148);
  not gc30 (wc30, n_177);
  xor g257 (Z[1], n_64, n_219);
  or g258 (n_258, wc31, n_155);
  not gc31 (wc31, n_157);
  or g259 (n_121, wc32, n_76);
  not gc32 (wc32, n_119);
  and g260 (n_168, wc33, n_83);
  not gc33 (wc33, n_126);
  and g261 (n_172, wc34, n_132);
  not gc34 (wc34, n_133);
  and g262 (n_195, wc35, n_95);
  not gc35 (wc35, n_136);
  and g263 (n_174, wc36, n_142);
  not gc36 (wc36, n_143);
  and g264 (n_182, wc37, n_107);
  not gc37 (wc37, n_146);
  and g265 (n_186, wc38, n_152);
  not gc38 (wc38, n_153);
  and g266 (n_179, wc39, n_148);
  not gc39 (wc39, n_174);
  or g267 (n_164, wc40, n_82);
  not gc40 (wc40, n_162);
  or g268 (n_169, n_166, wc41);
  not gc41 (wc41, n_162);
  or g269 (n_173, n_170, wc42);
  not gc42 (wc42, n_162);
  and g270 (n_200, wc43, n_101);
  not gc43 (wc43, n_175);
  and g271 (n_203, wc44, n_145);
  not gc44 (wc44, n_179);
  and g272 (n_206, n_182, wc45);
  not gc45 (wc45, n_183);
  and g273 (n_209, n_186, wc46);
  not gc46 (wc46, n_187);
  or g274 (n_191, wc47, n_94);
  not gc47 (wc47, n_189);
  or g275 (n_196, n_193, wc48);
  not gc48 (wc48, n_189);
  or g276 (n_198, wc49, n_177);
  not gc49 (wc49, n_189);
  or g277 (n_213, wc50, n_118);
  not gc50 (wc50, n_211);
endmodule

module add_signed_8959_1_GENERIC(A, B, Z);
  input [20:0] A, B;
  output [18:0] Z;
  wire [20:0] A, B;
  wire [18:0] Z;
  add_signed_8959_1_GENERIC_REAL g1(.A (A), .B ({B[20:19], B[17],
       B[17:0]}), .Z (Z));
endmodule

module add_signed_8959_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [20:0] A, B;
  output [18:0] Z;
  wire [20:0] A, B;
  wire [18:0] Z;
  wire n_64, n_66, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_76, n_77, n_78, n_79, n_80, n_82, n_83, n_84;
  wire n_85, n_86, n_88, n_89, n_90, n_91, n_92, n_94;
  wire n_95, n_96, n_97, n_98, n_100, n_101, n_102, n_103;
  wire n_104, n_106, n_107, n_108, n_109, n_110, n_112, n_113;
  wire n_114, n_115, n_116, n_118, n_119, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_128, n_130, n_132, n_133, n_135;
  wire n_136, n_138, n_140, n_142, n_143, n_145, n_146, n_148;
  wire n_150, n_152, n_153, n_155, n_156, n_157, n_160, n_162;
  wire n_164, n_165, n_166, n_168, n_169, n_170, n_172, n_173;
  wire n_174, n_175, n_177, n_179, n_181, n_182, n_183, n_185;
  wire n_186, n_187, n_189, n_191, n_192, n_193, n_195, n_196;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_213, n_214;
  wire n_219, n_220, n_222, n_223, n_224, n_226, n_227, n_228;
  wire n_229, n_231, n_232, n_233, n_235, n_236, n_237, n_238;
  wire n_240, n_241, n_243, n_244, n_246, n_247, n_248, n_249;
  wire n_251, n_252, n_253, n_255, n_256, n_257, n_258;
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_64, A[0], B[0]);
  nor g9 (n_66, A[1], B[1]);
  nand g10 (n_69, A[1], B[1]);
  nor g11 (n_76, A[2], B[2]);
  nand g12 (n_71, A[2], B[2]);
  nor g13 (n_72, A[3], B[3]);
  nand g14 (n_73, A[3], B[3]);
  nor g15 (n_82, A[4], B[4]);
  nand g16 (n_77, A[4], B[4]);
  nor g17 (n_78, A[5], B[5]);
  nand g18 (n_79, A[5], B[5]);
  nor g19 (n_88, A[6], B[6]);
  nand g20 (n_83, A[6], B[6]);
  nor g21 (n_84, A[7], B[7]);
  nand g22 (n_85, A[7], B[7]);
  nor g23 (n_94, A[8], B[8]);
  nand g24 (n_89, A[8], B[8]);
  nor g25 (n_90, A[9], B[9]);
  nand g26 (n_91, A[9], B[9]);
  nor g27 (n_100, A[10], B[10]);
  nand g28 (n_95, A[10], B[10]);
  nor g29 (n_96, A[11], B[11]);
  nand g30 (n_97, A[11], B[11]);
  nor g31 (n_106, A[12], B[12]);
  nand g32 (n_101, A[12], B[12]);
  nor g33 (n_102, A[13], B[13]);
  nand g34 (n_103, A[13], B[13]);
  nor g35 (n_112, A[14], B[14]);
  nand g36 (n_107, A[14], B[14]);
  nor g37 (n_108, A[15], B[15]);
  nand g38 (n_109, A[15], B[15]);
  nor g39 (n_118, A[16], B[16]);
  nand g40 (n_113, A[16], B[16]);
  nor g41 (n_114, A[17], B[17]);
  nand g42 (n_115, A[17], B[17]);
  nand g47 (n_119, n_69, n_70);
  nor g48 (n_74, n_71, n_72);
  nor g51 (n_122, n_76, n_72);
  nor g52 (n_80, n_77, n_78);
  nor g55 (n_128, n_82, n_78);
  nor g56 (n_86, n_83, n_84);
  nor g59 (n_130, n_88, n_84);
  nor g60 (n_92, n_89, n_90);
  nor g63 (n_138, n_94, n_90);
  nor g64 (n_98, n_95, n_96);
  nor g67 (n_140, n_100, n_96);
  nor g68 (n_104, n_101, n_102);
  nor g71 (n_148, n_106, n_102);
  nor g72 (n_110, n_107, n_108);
  nor g75 (n_150, n_112, n_108);
  nor g76 (n_116, n_113, n_114);
  nor g79 (n_160, n_118, n_114);
  nand g82 (n_222, n_71, n_121);
  nand g83 (n_124, n_122, n_119);
  nand g84 (n_162, n_123, n_124);
  nor g85 (n_126, n_88, n_125);
  nand g94 (n_170, n_128, n_130);
  nor g95 (n_136, n_100, n_135);
  nand g104 (n_177, n_138, n_140);
  nor g105 (n_146, n_112, n_145);
  nand g114 (n_185, n_148, n_150);
  nand g122 (n_226, n_77, n_164);
  nand g123 (n_165, n_128, n_162);
  nand g124 (n_228, n_125, n_165);
  nand g127 (n_231, n_168, n_169);
  nand g130 (n_189, n_172, n_173);
  nor g131 (n_175, n_106, n_174);
  nor g134 (n_199, n_106, n_177);
  nor g140 (n_183, n_181, n_174);
  nor g143 (n_205, n_177, n_181);
  nor g144 (n_187, n_185, n_174);
  nor g147 (n_208, n_177, n_185);
  nand g150 (n_235, n_89, n_191);
  nand g151 (n_192, n_138, n_189);
  nand g152 (n_237, n_135, n_192);
  nand g155 (n_240, n_195, n_196);
  nand g158 (n_243, n_174, n_198);
  nand g159 (n_201, n_199, n_189);
  nand g160 (n_246, n_200, n_201);
  nand g161 (n_204, n_202, n_189);
  nand g162 (n_248, n_203, n_204);
  nand g163 (n_207, n_205, n_189);
  nand g164 (n_251, n_206, n_207);
  nand g165 (n_210, n_208, n_189);
  nand g166 (n_211, n_209, n_210);
  nand g169 (n_255, n_113, n_213);
  nand g170 (n_214, n_160, n_211);
  nand g171 (n_257, n_156, n_214);
  xnor g178 (Z[2], n_119, n_220);
  xnor g181 (Z[3], n_222, n_223);
  xnor g183 (Z[4], n_162, n_224);
  xnor g186 (Z[5], n_226, n_227);
  xnor g188 (Z[6], n_228, n_229);
  xnor g191 (Z[7], n_231, n_232);
  xnor g193 (Z[8], n_189, n_233);
  xnor g196 (Z[9], n_235, n_236);
  xnor g198 (Z[10], n_237, n_238);
  xnor g201 (Z[11], n_240, n_241);
  xnor g204 (Z[12], n_243, n_244);
  xnor g207 (Z[13], n_246, n_247);
  xnor g209 (Z[14], n_248, n_249);
  xnor g212 (Z[15], n_251, n_252);
  xnor g214 (Z[16], n_211, n_253);
  xnor g217 (Z[17], n_255, n_256);
  xnor g219 (Z[18], n_257, n_258);
  and g222 (n_155, A[18], B[18]);
  or g223 (n_157, A[18], B[18]);
  or g224 (n_70, n_64, n_66);
  and g225 (n_123, wc, n_73);
  not gc (wc, n_74);
  and g226 (n_125, wc0, n_79);
  not gc0 (wc0, n_80);
  and g227 (n_132, wc1, n_85);
  not gc1 (wc1, n_86);
  and g228 (n_135, wc2, n_91);
  not gc2 (wc2, n_92);
  and g229 (n_142, wc3, n_97);
  not gc3 (wc3, n_98);
  and g230 (n_145, wc4, n_103);
  not gc4 (wc4, n_104);
  and g231 (n_152, wc5, n_109);
  not gc5 (wc5, n_110);
  and g232 (n_156, wc6, n_115);
  not gc6 (wc6, n_116);
  or g233 (n_166, wc7, n_88);
  not gc7 (wc7, n_128);
  or g234 (n_193, wc8, n_100);
  not gc8 (wc8, n_138);
  or g235 (n_181, wc9, n_112);
  not gc9 (wc9, n_148);
  or g236 (n_219, wc10, n_66);
  not gc10 (wc10, n_69);
  or g237 (n_220, wc11, n_76);
  not gc11 (wc11, n_71);
  or g238 (n_223, wc12, n_72);
  not gc12 (wc12, n_73);
  or g239 (n_224, wc13, n_82);
  not gc13 (wc13, n_77);
  or g240 (n_227, wc14, n_78);
  not gc14 (wc14, n_79);
  or g241 (n_229, wc15, n_88);
  not gc15 (wc15, n_83);
  or g242 (n_232, wc16, n_84);
  not gc16 (wc16, n_85);
  or g243 (n_233, wc17, n_94);
  not gc17 (wc17, n_89);
  or g244 (n_236, wc18, n_90);
  not gc18 (wc18, n_91);
  or g245 (n_238, wc19, n_100);
  not gc19 (wc19, n_95);
  or g246 (n_241, wc20, n_96);
  not gc20 (wc20, n_97);
  or g247 (n_244, wc21, n_106);
  not gc21 (wc21, n_101);
  or g248 (n_247, wc22, n_102);
  not gc22 (wc22, n_103);
  or g249 (n_249, wc23, n_112);
  not gc23 (wc23, n_107);
  or g250 (n_252, wc24, n_108);
  not gc24 (wc24, n_109);
  or g251 (n_253, wc25, n_118);
  not gc25 (wc25, n_113);
  or g252 (n_256, wc26, n_114);
  not gc26 (wc26, n_115);
  and g253 (n_133, wc27, n_130);
  not gc27 (wc27, n_125);
  and g254 (n_143, wc28, n_140);
  not gc28 (wc28, n_135);
  and g255 (n_153, wc29, n_150);
  not gc29 (wc29, n_145);
  and g256 (n_202, wc30, n_148);
  not gc30 (wc30, n_177);
  xor g257 (Z[1], n_64, n_219);
  or g258 (n_258, wc31, n_155);
  not gc31 (wc31, n_157);
  or g259 (n_121, wc32, n_76);
  not gc32 (wc32, n_119);
  and g260 (n_168, wc33, n_83);
  not gc33 (wc33, n_126);
  and g261 (n_172, wc34, n_132);
  not gc34 (wc34, n_133);
  and g262 (n_195, wc35, n_95);
  not gc35 (wc35, n_136);
  and g263 (n_174, wc36, n_142);
  not gc36 (wc36, n_143);
  and g264 (n_182, wc37, n_107);
  not gc37 (wc37, n_146);
  and g265 (n_186, wc38, n_152);
  not gc38 (wc38, n_153);
  and g266 (n_179, wc39, n_148);
  not gc39 (wc39, n_174);
  or g267 (n_164, wc40, n_82);
  not gc40 (wc40, n_162);
  or g268 (n_169, n_166, wc41);
  not gc41 (wc41, n_162);
  or g269 (n_173, n_170, wc42);
  not gc42 (wc42, n_162);
  and g270 (n_200, wc43, n_101);
  not gc43 (wc43, n_175);
  and g271 (n_203, wc44, n_145);
  not gc44 (wc44, n_179);
  and g272 (n_206, n_182, wc45);
  not gc45 (wc45, n_183);
  and g273 (n_209, n_186, wc46);
  not gc46 (wc46, n_187);
  or g274 (n_191, wc47, n_94);
  not gc47 (wc47, n_189);
  or g275 (n_196, n_193, wc48);
  not gc48 (wc48, n_189);
  or g276 (n_198, wc49, n_177);
  not gc49 (wc49, n_189);
  or g277 (n_213, wc50, n_118);
  not gc50 (wc50, n_211);
endmodule

module add_signed_8959_2_GENERIC(A, B, Z);
  input [20:0] A, B;
  output [18:0] Z;
  wire [20:0] A, B;
  wire [18:0] Z;
  add_signed_8959_2_GENERIC_REAL g1(.A (A), .B ({B[20:19], B[17],
       B[17:0]}), .Z (Z));
endmodule

module add_signed_9024_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [31:0] A, B;
  output [30:0] Z;
  wire [31:0] A, B;
  wire [30:0] Z;
  wire n_99, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214;
  wire n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230;
  wire n_231, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246;
  wire n_247, n_248, n_252;
  nand g4 (n_99, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_104, A[1], B[1]);
  nand g13 (n_108, n_104, n_105, n_106);
  xor g14 (n_107, A[1], B[1]);
  nand g16 (n_109, A[2], B[2]);
  nand g17 (n_110, A[2], n_108);
  nand g18 (n_111, B[2], n_108);
  nand g19 (n_113, n_109, n_110, n_111);
  xor g20 (n_112, A[2], B[2]);
  xor g21 (Z[2], n_108, n_112);
  nand g22 (n_114, A[3], B[3]);
  nand g23 (n_115, A[3], n_113);
  nand g24 (n_116, B[3], n_113);
  nand g25 (n_118, n_114, n_115, n_116);
  xor g26 (n_117, A[3], B[3]);
  xor g27 (Z[3], n_113, n_117);
  nand g28 (n_119, A[4], B[4]);
  nand g29 (n_120, A[4], n_118);
  nand g30 (n_121, B[4], n_118);
  nand g31 (n_123, n_119, n_120, n_121);
  xor g32 (n_122, A[4], B[4]);
  xor g33 (Z[4], n_118, n_122);
  nand g34 (n_124, A[5], B[5]);
  nand g35 (n_125, A[5], n_123);
  nand g36 (n_126, B[5], n_123);
  nand g37 (n_128, n_124, n_125, n_126);
  xor g38 (n_127, A[5], B[5]);
  xor g39 (Z[5], n_123, n_127);
  nand g40 (n_129, A[6], B[6]);
  nand g41 (n_130, A[6], n_128);
  nand g42 (n_131, B[6], n_128);
  nand g43 (n_133, n_129, n_130, n_131);
  xor g44 (n_132, A[6], B[6]);
  xor g45 (Z[6], n_128, n_132);
  nand g46 (n_134, A[7], B[7]);
  nand g47 (n_135, A[7], n_133);
  nand g48 (n_136, B[7], n_133);
  nand g49 (n_138, n_134, n_135, n_136);
  xor g50 (n_137, A[7], B[7]);
  xor g51 (Z[7], n_133, n_137);
  nand g52 (n_139, A[8], B[8]);
  nand g53 (n_140, A[8], n_138);
  nand g54 (n_141, B[8], n_138);
  nand g55 (n_143, n_139, n_140, n_141);
  xor g56 (n_142, A[8], B[8]);
  xor g57 (Z[8], n_138, n_142);
  nand g58 (n_144, A[9], B[9]);
  nand g59 (n_145, A[9], n_143);
  nand g60 (n_146, B[9], n_143);
  nand g61 (n_148, n_144, n_145, n_146);
  xor g62 (n_147, A[9], B[9]);
  xor g63 (Z[9], n_143, n_147);
  nand g64 (n_149, A[10], B[10]);
  nand g65 (n_150, A[10], n_148);
  nand g66 (n_151, B[10], n_148);
  nand g67 (n_153, n_149, n_150, n_151);
  xor g68 (n_152, A[10], B[10]);
  xor g69 (Z[10], n_148, n_152);
  nand g70 (n_154, A[11], B[11]);
  nand g71 (n_155, A[11], n_153);
  nand g72 (n_156, B[11], n_153);
  nand g73 (n_158, n_154, n_155, n_156);
  xor g74 (n_157, A[11], B[11]);
  xor g75 (Z[11], n_153, n_157);
  nand g76 (n_159, A[12], B[12]);
  nand g77 (n_160, A[12], n_158);
  nand g78 (n_161, B[12], n_158);
  nand g79 (n_163, n_159, n_160, n_161);
  xor g80 (n_162, A[12], B[12]);
  xor g81 (Z[12], n_158, n_162);
  nand g82 (n_164, A[13], B[13]);
  nand g83 (n_165, A[13], n_163);
  nand g84 (n_166, B[13], n_163);
  nand g85 (n_168, n_164, n_165, n_166);
  xor g86 (n_167, A[13], B[13]);
  xor g87 (Z[13], n_163, n_167);
  nand g88 (n_169, A[14], B[14]);
  nand g89 (n_170, A[14], n_168);
  nand g90 (n_171, B[14], n_168);
  nand g91 (n_173, n_169, n_170, n_171);
  xor g92 (n_172, A[14], B[14]);
  xor g93 (Z[14], n_168, n_172);
  nand g94 (n_174, A[15], B[15]);
  nand g95 (n_175, A[15], n_173);
  nand g96 (n_176, B[15], n_173);
  nand g97 (n_178, n_174, n_175, n_176);
  xor g98 (n_177, A[15], B[15]);
  xor g99 (Z[15], n_173, n_177);
  nand g100 (n_179, A[16], B[16]);
  nand g101 (n_180, A[16], n_178);
  nand g102 (n_181, B[16], n_178);
  nand g103 (n_183, n_179, n_180, n_181);
  xor g104 (n_182, A[16], B[16]);
  xor g105 (Z[16], n_178, n_182);
  nand g106 (n_184, A[17], B[17]);
  nand g107 (n_185, A[17], n_183);
  nand g108 (n_186, B[17], n_183);
  nand g109 (n_188, n_184, n_185, n_186);
  xor g110 (n_187, A[17], B[17]);
  xor g111 (Z[17], n_183, n_187);
  nand g112 (n_189, A[18], B[18]);
  nand g113 (n_190, A[18], n_188);
  nand g114 (n_191, B[18], n_188);
  nand g115 (n_193, n_189, n_190, n_191);
  xor g116 (n_192, A[18], B[18]);
  xor g117 (Z[18], n_188, n_192);
  nand g118 (n_194, A[19], B[19]);
  nand g119 (n_195, A[19], n_193);
  nand g120 (n_196, B[19], n_193);
  nand g121 (n_198, n_194, n_195, n_196);
  xor g122 (n_197, A[19], B[19]);
  xor g123 (Z[19], n_193, n_197);
  nand g124 (n_199, A[20], B[20]);
  nand g125 (n_200, A[20], n_198);
  nand g126 (n_201, B[20], n_198);
  nand g127 (n_203, n_199, n_200, n_201);
  xor g128 (n_202, A[20], B[20]);
  xor g129 (Z[20], n_198, n_202);
  nand g130 (n_204, A[21], B[21]);
  nand g131 (n_205, A[21], n_203);
  nand g132 (n_206, B[21], n_203);
  nand g133 (n_208, n_204, n_205, n_206);
  xor g134 (n_207, A[21], B[21]);
  xor g135 (Z[21], n_203, n_207);
  nand g136 (n_209, A[22], B[22]);
  nand g137 (n_210, A[22], n_208);
  nand g138 (n_211, B[22], n_208);
  nand g139 (n_213, n_209, n_210, n_211);
  xor g140 (n_212, A[22], B[22]);
  xor g141 (Z[22], n_208, n_212);
  nand g142 (n_214, A[23], B[23]);
  nand g143 (n_215, A[23], n_213);
  nand g144 (n_216, B[23], n_213);
  nand g145 (n_218, n_214, n_215, n_216);
  xor g146 (n_217, A[23], B[23]);
  xor g147 (Z[23], n_213, n_217);
  nand g148 (n_219, A[24], B[24]);
  nand g149 (n_220, A[24], n_218);
  nand g150 (n_221, B[24], n_218);
  nand g151 (n_223, n_219, n_220, n_221);
  xor g152 (n_222, A[24], B[24]);
  xor g153 (Z[24], n_218, n_222);
  nand g154 (n_224, A[25], B[25]);
  nand g155 (n_225, A[25], n_223);
  nand g156 (n_226, B[25], n_223);
  nand g157 (n_228, n_224, n_225, n_226);
  xor g158 (n_227, A[25], B[25]);
  xor g159 (Z[25], n_223, n_227);
  nand g160 (n_229, A[26], B[26]);
  nand g161 (n_230, A[26], n_228);
  nand g162 (n_231, B[26], n_228);
  nand g163 (n_233, n_229, n_230, n_231);
  xor g164 (n_232, A[26], B[26]);
  xor g165 (Z[26], n_228, n_232);
  nand g166 (n_234, A[27], B[27]);
  nand g167 (n_235, A[27], n_233);
  nand g168 (n_236, B[27], n_233);
  nand g169 (n_238, n_234, n_235, n_236);
  xor g170 (n_237, A[27], B[27]);
  xor g171 (Z[27], n_233, n_237);
  nand g172 (n_239, A[28], B[28]);
  nand g173 (n_240, A[28], n_238);
  nand g174 (n_241, B[28], n_238);
  nand g175 (n_243, n_239, n_240, n_241);
  xor g176 (n_242, A[28], B[28]);
  xor g177 (Z[28], n_238, n_242);
  nand g178 (n_244, A[29], B[29]);
  nand g179 (n_245, A[29], n_243);
  nand g180 (n_246, B[29], n_243);
  nand g181 (n_248, n_244, n_245, n_246);
  xor g182 (n_247, A[29], B[29]);
  xor g183 (Z[29], n_243, n_247);
  xor g189 (Z[30], n_248, n_252);
  xor g191 (n_252, A[30], B[30]);
  or g192 (n_105, wc, n_99);
  not gc (wc, A[1]);
  or g193 (n_106, wc0, n_99);
  not gc0 (wc0, B[1]);
  xnor g194 (Z[1], n_99, n_107);
endmodule

module add_signed_9024_GENERIC(A, B, Z);
  input [31:0] A, B;
  output [30:0] Z;
  wire [31:0] A, B;
  wire [30:0] Z;
  add_signed_9024_GENERIC_REAL g1(.A ({A[31], A[28], A[28], A[28:0]}),
       .B ({B[31], B[28], B[28], B[28:0]}), .Z (Z));
endmodule

module add_signed_9027_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [27:0] A, B;
  output [26:0] Z;
  wire [27:0] A, B;
  wire [26:0] Z;
  wire n_87, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_220;
  nand g4 (n_87, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_92, A[1], B[1]);
  nand g13 (n_96, n_92, n_93, n_94);
  xor g14 (n_95, A[1], B[1]);
  nand g16 (n_97, A[2], B[2]);
  nand g17 (n_98, A[2], n_96);
  nand g18 (n_99, B[2], n_96);
  nand g19 (n_101, n_97, n_98, n_99);
  xor g20 (n_100, A[2], B[2]);
  xor g21 (Z[2], n_96, n_100);
  nand g22 (n_102, A[3], B[3]);
  nand g23 (n_103, A[3], n_101);
  nand g24 (n_104, B[3], n_101);
  nand g25 (n_106, n_102, n_103, n_104);
  xor g26 (n_105, A[3], B[3]);
  xor g27 (Z[3], n_101, n_105);
  nand g28 (n_107, A[4], B[4]);
  nand g29 (n_108, A[4], n_106);
  nand g30 (n_109, B[4], n_106);
  nand g31 (n_111, n_107, n_108, n_109);
  xor g32 (n_110, A[4], B[4]);
  xor g33 (Z[4], n_106, n_110);
  nand g34 (n_112, A[5], B[5]);
  nand g35 (n_113, A[5], n_111);
  nand g36 (n_114, B[5], n_111);
  nand g37 (n_116, n_112, n_113, n_114);
  xor g38 (n_115, A[5], B[5]);
  xor g39 (Z[5], n_111, n_115);
  nand g40 (n_117, A[6], B[6]);
  nand g41 (n_118, A[6], n_116);
  nand g42 (n_119, B[6], n_116);
  nand g43 (n_121, n_117, n_118, n_119);
  xor g44 (n_120, A[6], B[6]);
  xor g45 (Z[6], n_116, n_120);
  nand g46 (n_122, A[7], B[7]);
  nand g47 (n_123, A[7], n_121);
  nand g48 (n_124, B[7], n_121);
  nand g49 (n_126, n_122, n_123, n_124);
  xor g50 (n_125, A[7], B[7]);
  xor g51 (Z[7], n_121, n_125);
  nand g52 (n_127, A[8], B[8]);
  nand g53 (n_128, A[8], n_126);
  nand g54 (n_129, B[8], n_126);
  nand g55 (n_131, n_127, n_128, n_129);
  xor g56 (n_130, A[8], B[8]);
  xor g57 (Z[8], n_126, n_130);
  nand g58 (n_132, A[9], B[9]);
  nand g59 (n_133, A[9], n_131);
  nand g60 (n_134, B[9], n_131);
  nand g61 (n_136, n_132, n_133, n_134);
  xor g62 (n_135, A[9], B[9]);
  xor g63 (Z[9], n_131, n_135);
  nand g64 (n_137, A[10], B[10]);
  nand g65 (n_138, A[10], n_136);
  nand g66 (n_139, B[10], n_136);
  nand g67 (n_141, n_137, n_138, n_139);
  xor g68 (n_140, A[10], B[10]);
  xor g69 (Z[10], n_136, n_140);
  nand g70 (n_142, A[11], B[11]);
  nand g71 (n_143, A[11], n_141);
  nand g72 (n_144, B[11], n_141);
  nand g73 (n_146, n_142, n_143, n_144);
  xor g74 (n_145, A[11], B[11]);
  xor g75 (Z[11], n_141, n_145);
  nand g76 (n_147, A[12], B[12]);
  nand g77 (n_148, A[12], n_146);
  nand g78 (n_149, B[12], n_146);
  nand g79 (n_151, n_147, n_148, n_149);
  xor g80 (n_150, A[12], B[12]);
  xor g81 (Z[12], n_146, n_150);
  nand g82 (n_152, A[13], B[13]);
  nand g83 (n_153, A[13], n_151);
  nand g84 (n_154, B[13], n_151);
  nand g85 (n_156, n_152, n_153, n_154);
  xor g86 (n_155, A[13], B[13]);
  xor g87 (Z[13], n_151, n_155);
  nand g88 (n_157, A[14], B[14]);
  nand g89 (n_158, A[14], n_156);
  nand g90 (n_159, B[14], n_156);
  nand g91 (n_161, n_157, n_158, n_159);
  xor g92 (n_160, A[14], B[14]);
  xor g93 (Z[14], n_156, n_160);
  nand g94 (n_162, A[15], B[15]);
  nand g95 (n_163, A[15], n_161);
  nand g96 (n_164, B[15], n_161);
  nand g97 (n_166, n_162, n_163, n_164);
  xor g98 (n_165, A[15], B[15]);
  xor g99 (Z[15], n_161, n_165);
  nand g100 (n_167, A[16], B[16]);
  nand g101 (n_168, A[16], n_166);
  nand g102 (n_169, B[16], n_166);
  nand g103 (n_171, n_167, n_168, n_169);
  xor g104 (n_170, A[16], B[16]);
  xor g105 (Z[16], n_166, n_170);
  nand g106 (n_172, A[17], B[17]);
  nand g107 (n_173, A[17], n_171);
  nand g108 (n_174, B[17], n_171);
  nand g109 (n_176, n_172, n_173, n_174);
  xor g110 (n_175, A[17], B[17]);
  xor g111 (Z[17], n_171, n_175);
  nand g112 (n_177, A[18], B[18]);
  nand g113 (n_178, A[18], n_176);
  nand g114 (n_179, B[18], n_176);
  nand g115 (n_181, n_177, n_178, n_179);
  xor g116 (n_180, A[18], B[18]);
  xor g117 (Z[18], n_176, n_180);
  nand g118 (n_182, A[19], B[19]);
  nand g119 (n_183, A[19], n_181);
  nand g120 (n_184, B[19], n_181);
  nand g121 (n_186, n_182, n_183, n_184);
  xor g122 (n_185, A[19], B[19]);
  xor g123 (Z[19], n_181, n_185);
  nand g124 (n_187, A[20], B[20]);
  nand g125 (n_188, A[20], n_186);
  nand g126 (n_189, B[20], n_186);
  nand g127 (n_191, n_187, n_188, n_189);
  xor g128 (n_190, A[20], B[20]);
  xor g129 (Z[20], n_186, n_190);
  nand g130 (n_192, A[21], B[21]);
  nand g131 (n_193, A[21], n_191);
  nand g132 (n_194, B[21], n_191);
  nand g133 (n_196, n_192, n_193, n_194);
  xor g134 (n_195, A[21], B[21]);
  xor g135 (Z[21], n_191, n_195);
  nand g136 (n_197, A[22], B[22]);
  nand g137 (n_198, A[22], n_196);
  nand g138 (n_199, B[22], n_196);
  nand g139 (n_201, n_197, n_198, n_199);
  xor g140 (n_200, A[22], B[22]);
  xor g141 (Z[22], n_196, n_200);
  nand g142 (n_202, A[23], B[23]);
  nand g143 (n_203, A[23], n_201);
  nand g144 (n_204, B[23], n_201);
  nand g145 (n_206, n_202, n_203, n_204);
  xor g146 (n_205, A[23], B[23]);
  xor g147 (Z[23], n_201, n_205);
  nand g148 (n_207, A[24], B[24]);
  nand g149 (n_208, A[24], n_206);
  nand g150 (n_209, B[24], n_206);
  nand g151 (n_211, n_207, n_208, n_209);
  xor g152 (n_210, A[24], B[24]);
  xor g153 (Z[24], n_206, n_210);
  nand g154 (n_212, A[25], B[25]);
  nand g155 (n_213, A[25], n_211);
  nand g156 (n_214, B[25], n_211);
  nand g157 (n_216, n_212, n_213, n_214);
  xor g158 (n_215, A[25], B[25]);
  xor g159 (Z[25], n_211, n_215);
  xor g165 (Z[26], n_216, n_220);
  xor g167 (n_220, A[26], B[26]);
  or g168 (n_93, wc, n_87);
  not gc (wc, A[1]);
  or g169 (n_94, wc0, n_87);
  not gc0 (wc0, B[1]);
  xnor g170 (Z[1], n_87, n_95);
endmodule

module add_signed_9027_GENERIC(A, B, Z);
  input [27:0] A, B;
  output [26:0] Z;
  wire [27:0] A, B;
  wire [26:0] Z;
  add_signed_9027_GENERIC_REAL g1(.A ({A[27], A[23], A[23], A[23],
       A[23:0]}), .B ({B[27], B[23], B[23], B[23], B[23:0]}), .Z (Z));
endmodule

module add_signed_9030_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [21:0] A, B;
  output [20:0] Z;
  wire [21:0] A, B;
  wire [20:0] Z;
  wire n_69, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_172;
  nand g4 (n_69, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_74, A[1], B[1]);
  nand g13 (n_78, n_74, n_75, n_76);
  xor g14 (n_77, A[1], B[1]);
  nand g16 (n_79, A[2], B[2]);
  nand g17 (n_80, A[2], n_78);
  nand g18 (n_81, B[2], n_78);
  nand g19 (n_83, n_79, n_80, n_81);
  xor g20 (n_82, A[2], B[2]);
  xor g21 (Z[2], n_78, n_82);
  nand g22 (n_84, A[3], B[3]);
  nand g23 (n_85, A[3], n_83);
  nand g24 (n_86, B[3], n_83);
  nand g25 (n_88, n_84, n_85, n_86);
  xor g26 (n_87, A[3], B[3]);
  xor g27 (Z[3], n_83, n_87);
  nand g28 (n_89, A[4], B[4]);
  nand g29 (n_90, A[4], n_88);
  nand g30 (n_91, B[4], n_88);
  nand g31 (n_93, n_89, n_90, n_91);
  xor g32 (n_92, A[4], B[4]);
  xor g33 (Z[4], n_88, n_92);
  nand g34 (n_94, A[5], B[5]);
  nand g35 (n_95, A[5], n_93);
  nand g36 (n_96, B[5], n_93);
  nand g37 (n_98, n_94, n_95, n_96);
  xor g38 (n_97, A[5], B[5]);
  xor g39 (Z[5], n_93, n_97);
  nand g40 (n_99, A[6], B[6]);
  nand g41 (n_100, A[6], n_98);
  nand g42 (n_101, B[6], n_98);
  nand g43 (n_103, n_99, n_100, n_101);
  xor g44 (n_102, A[6], B[6]);
  xor g45 (Z[6], n_98, n_102);
  nand g46 (n_104, A[7], B[7]);
  nand g47 (n_105, A[7], n_103);
  nand g48 (n_106, B[7], n_103);
  nand g49 (n_108, n_104, n_105, n_106);
  xor g50 (n_107, A[7], B[7]);
  xor g51 (Z[7], n_103, n_107);
  nand g52 (n_109, A[8], B[8]);
  nand g53 (n_110, A[8], n_108);
  nand g54 (n_111, B[8], n_108);
  nand g55 (n_113, n_109, n_110, n_111);
  xor g56 (n_112, A[8], B[8]);
  xor g57 (Z[8], n_108, n_112);
  nand g58 (n_114, A[9], B[9]);
  nand g59 (n_115, A[9], n_113);
  nand g60 (n_116, B[9], n_113);
  nand g61 (n_118, n_114, n_115, n_116);
  xor g62 (n_117, A[9], B[9]);
  xor g63 (Z[9], n_113, n_117);
  nand g64 (n_119, A[10], B[10]);
  nand g65 (n_120, A[10], n_118);
  nand g66 (n_121, B[10], n_118);
  nand g67 (n_123, n_119, n_120, n_121);
  xor g68 (n_122, A[10], B[10]);
  xor g69 (Z[10], n_118, n_122);
  nand g70 (n_124, A[11], B[11]);
  nand g71 (n_125, A[11], n_123);
  nand g72 (n_126, B[11], n_123);
  nand g73 (n_128, n_124, n_125, n_126);
  xor g74 (n_127, A[11], B[11]);
  xor g75 (Z[11], n_123, n_127);
  nand g76 (n_129, A[12], B[12]);
  nand g77 (n_130, A[12], n_128);
  nand g78 (n_131, B[12], n_128);
  nand g79 (n_133, n_129, n_130, n_131);
  xor g80 (n_132, A[12], B[12]);
  xor g81 (Z[12], n_128, n_132);
  nand g82 (n_134, A[13], B[13]);
  nand g83 (n_135, A[13], n_133);
  nand g84 (n_136, B[13], n_133);
  nand g85 (n_138, n_134, n_135, n_136);
  xor g86 (n_137, A[13], B[13]);
  xor g87 (Z[13], n_133, n_137);
  nand g88 (n_139, A[14], B[14]);
  nand g89 (n_140, A[14], n_138);
  nand g90 (n_141, B[14], n_138);
  nand g91 (n_143, n_139, n_140, n_141);
  xor g92 (n_142, A[14], B[14]);
  xor g93 (Z[14], n_138, n_142);
  nand g94 (n_144, A[15], B[15]);
  nand g95 (n_145, A[15], n_143);
  nand g96 (n_146, B[15], n_143);
  nand g97 (n_148, n_144, n_145, n_146);
  xor g98 (n_147, A[15], B[15]);
  xor g99 (Z[15], n_143, n_147);
  nand g100 (n_149, A[16], B[16]);
  nand g101 (n_150, A[16], n_148);
  nand g102 (n_151, B[16], n_148);
  nand g103 (n_153, n_149, n_150, n_151);
  xor g104 (n_152, A[16], B[16]);
  xor g105 (Z[16], n_148, n_152);
  nand g106 (n_154, A[17], B[17]);
  nand g107 (n_155, A[17], n_153);
  nand g108 (n_156, B[17], n_153);
  nand g109 (n_158, n_154, n_155, n_156);
  xor g110 (n_157, A[17], B[17]);
  xor g111 (Z[17], n_153, n_157);
  nand g112 (n_159, A[18], B[18]);
  nand g113 (n_160, A[18], n_158);
  nand g114 (n_161, B[18], n_158);
  nand g115 (n_163, n_159, n_160, n_161);
  xor g116 (n_162, A[18], B[18]);
  xor g117 (Z[18], n_158, n_162);
  nand g118 (n_164, A[19], B[19]);
  nand g119 (n_165, A[19], n_163);
  nand g120 (n_166, B[19], n_163);
  nand g121 (n_168, n_164, n_165, n_166);
  xor g122 (n_167, A[19], B[19]);
  xor g123 (Z[19], n_163, n_167);
  xor g129 (Z[20], n_168, n_172);
  xor g131 (n_172, A[20], B[20]);
  or g132 (n_75, wc, n_69);
  not gc (wc, A[1]);
  or g133 (n_76, wc0, n_69);
  not gc0 (wc0, B[1]);
  xnor g134 (Z[1], n_69, n_77);
endmodule

module add_signed_9030_GENERIC(A, B, Z);
  input [21:0] A, B;
  output [20:0] Z;
  wire [21:0] A, B;
  wire [20:0] Z;
  add_signed_9030_GENERIC_REAL g1(.A ({A[21], A[18], A[18], A[18:0]}),
       .B ({B[21], B[18], B[18], B[18:0]}), .Z (Z));
endmodule

module add_signed_9092_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [32:0] A, B;
  output [31:0] Z;
  wire [32:0] A, B;
  wire [31:0] Z;
  wire n_102, n_105, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_115, n_116, n_117, n_118, n_119, n_121, n_122, n_123;
  wire n_124, n_125, n_127, n_128, n_129, n_130, n_131, n_133;
  wire n_134, n_135, n_136, n_137, n_139, n_140, n_141, n_142;
  wire n_143, n_145, n_146, n_147, n_148, n_149, n_151, n_152;
  wire n_153, n_154, n_155, n_157, n_158, n_159, n_160, n_161;
  wire n_163, n_164, n_165, n_166, n_167, n_169, n_170, n_171;
  wire n_172, n_173, n_175, n_176, n_177, n_178, n_179, n_181;
  wire n_182, n_183, n_184, n_185, n_187, n_188, n_189, n_190;
  wire n_191, n_193, n_194, n_195, n_196, n_199, n_200, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_209, n_211, n_213;
  wire n_214, n_216, n_217, n_219, n_221, n_223, n_224, n_226;
  wire n_227, n_229, n_231, n_233, n_234, n_236, n_237, n_239;
  wire n_241, n_243, n_244, n_246, n_247, n_249, n_251, n_253;
  wire n_254, n_256, n_257, n_259, n_261, n_263, n_264, n_266;
  wire n_267, n_269, n_276, n_278, n_279, n_280, n_282, n_283;
  wire n_284, n_286, n_287, n_288, n_289, n_291, n_293, n_295;
  wire n_296, n_297, n_299, n_300, n_301, n_303, n_304, n_306;
  wire n_308, n_310, n_311, n_312, n_314, n_315, n_316, n_318;
  wire n_319, n_321, n_323, n_325, n_326, n_327, n_333, n_335;
  wire n_336, n_337, n_339, n_340, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_358, n_361, n_363, n_364, n_365;
  wire n_368, n_371, n_373, n_374, n_376, n_378, n_379, n_381;
  wire n_383, n_384, n_391, n_393, n_394, n_395, n_397, n_398;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_413, n_414, n_415, n_417;
  wire n_418, n_419, n_421, n_422, n_423, n_425, n_426, n_427;
  wire n_429, n_430, n_431, n_433, n_434, n_435, n_437, n_438;
  wire n_443, n_444, n_446, n_447, n_448, n_450, n_451, n_452;
  wire n_453, n_455, n_456, n_457, n_459, n_460, n_461, n_462;
  wire n_464, n_465, n_467, n_468, n_470, n_471, n_472, n_473;
  wire n_475, n_476, n_477, n_479, n_480, n_481, n_482, n_484;
  wire n_485, n_487, n_488, n_490, n_491, n_492, n_493, n_495;
  wire n_496, n_497, n_498, n_500, n_501, n_502, n_503, n_505;
  wire n_506, n_508, n_509, n_511, n_512, n_513, n_514, n_516;
  wire n_517;
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_102, A[0], B[0]);
  nor g9 (n_105, A[1], B[1]);
  nand g10 (n_108, A[1], B[1]);
  nor g11 (n_115, A[2], B[2]);
  nand g12 (n_110, A[2], B[2]);
  nor g13 (n_111, A[3], B[3]);
  nand g14 (n_112, A[3], B[3]);
  nor g15 (n_121, A[4], B[4]);
  nand g16 (n_116, A[4], B[4]);
  nor g17 (n_117, A[5], B[5]);
  nand g18 (n_118, A[5], B[5]);
  nor g19 (n_127, A[6], B[6]);
  nand g20 (n_122, A[6], B[6]);
  nor g21 (n_123, A[7], B[7]);
  nand g22 (n_124, A[7], B[7]);
  nor g23 (n_133, A[8], B[8]);
  nand g24 (n_128, A[8], B[8]);
  nor g25 (n_129, A[9], B[9]);
  nand g26 (n_130, A[9], B[9]);
  nor g27 (n_139, A[10], B[10]);
  nand g28 (n_134, A[10], B[10]);
  nor g29 (n_135, A[11], B[11]);
  nand g30 (n_136, A[11], B[11]);
  nor g31 (n_145, A[12], B[12]);
  nand g32 (n_140, A[12], B[12]);
  nor g33 (n_141, A[13], B[13]);
  nand g34 (n_142, A[13], B[13]);
  nor g35 (n_151, A[14], B[14]);
  nand g36 (n_146, A[14], B[14]);
  nor g37 (n_147, A[15], B[15]);
  nand g38 (n_148, A[15], B[15]);
  nor g39 (n_157, A[16], B[16]);
  nand g40 (n_152, A[16], B[16]);
  nor g41 (n_153, A[17], B[17]);
  nand g42 (n_154, A[17], B[17]);
  nor g43 (n_163, A[18], B[18]);
  nand g44 (n_158, A[18], B[18]);
  nor g45 (n_159, A[19], B[19]);
  nand g46 (n_160, A[19], B[19]);
  nor g47 (n_169, A[20], B[20]);
  nand g48 (n_164, A[20], B[20]);
  nor g49 (n_165, A[21], B[21]);
  nand g50 (n_166, A[21], B[21]);
  nor g51 (n_175, A[22], B[22]);
  nand g52 (n_170, A[22], B[22]);
  nor g53 (n_171, A[23], B[23]);
  nand g54 (n_172, A[23], B[23]);
  nor g55 (n_181, A[24], B[24]);
  nand g56 (n_176, A[24], B[24]);
  nor g57 (n_177, A[25], B[25]);
  nand g58 (n_178, A[25], B[25]);
  nor g59 (n_187, A[26], B[26]);
  nand g60 (n_182, A[26], B[26]);
  nor g61 (n_183, A[27], B[27]);
  nand g62 (n_184, A[27], B[27]);
  nor g63 (n_193, A[28], B[28]);
  nand g64 (n_188, A[28], B[28]);
  nor g65 (n_189, A[29], B[29]);
  nand g66 (n_190, A[29], B[29]);
  nor g67 (n_199, A[30], B[30]);
  nand g68 (n_194, A[30], B[30]);
  nand g73 (n_200, n_108, n_109);
  nor g74 (n_113, n_110, n_111);
  nor g77 (n_203, n_115, n_111);
  nor g78 (n_119, n_116, n_117);
  nor g81 (n_209, n_121, n_117);
  nor g82 (n_125, n_122, n_123);
  nor g85 (n_211, n_127, n_123);
  nor g86 (n_131, n_128, n_129);
  nor g89 (n_219, n_133, n_129);
  nor g90 (n_137, n_134, n_135);
  nor g93 (n_221, n_139, n_135);
  nor g94 (n_143, n_140, n_141);
  nor g97 (n_229, n_145, n_141);
  nor g98 (n_149, n_146, n_147);
  nor g101 (n_231, n_151, n_147);
  nor g102 (n_155, n_152, n_153);
  nor g105 (n_239, n_157, n_153);
  nor g106 (n_161, n_158, n_159);
  nor g109 (n_241, n_163, n_159);
  nor g110 (n_167, n_164, n_165);
  nor g113 (n_249, n_169, n_165);
  nor g114 (n_173, n_170, n_171);
  nor g117 (n_251, n_175, n_171);
  nor g118 (n_179, n_176, n_177);
  nor g121 (n_259, n_181, n_177);
  nor g122 (n_185, n_182, n_183);
  nor g125 (n_261, n_187, n_183);
  nor g126 (n_191, n_188, n_189);
  nor g129 (n_269, n_193, n_189);
  nand g136 (n_446, n_110, n_202);
  nand g137 (n_205, n_203, n_200);
  nand g138 (n_276, n_204, n_205);
  nor g139 (n_207, n_127, n_206);
  nand g148 (n_284, n_209, n_211);
  nor g149 (n_217, n_139, n_216);
  nand g158 (n_291, n_219, n_221);
  nor g159 (n_227, n_151, n_226);
  nand g168 (n_299, n_229, n_231);
  nor g169 (n_237, n_163, n_236);
  nand g178 (n_306, n_239, n_241);
  nor g179 (n_247, n_175, n_246);
  nand g188 (n_314, n_249, n_251);
  nor g189 (n_257, n_187, n_256);
  nand g198 (n_321, n_259, n_261);
  nor g199 (n_267, n_199, n_266);
  nand g211 (n_450, n_116, n_278);
  nand g212 (n_279, n_209, n_276);
  nand g213 (n_452, n_206, n_279);
  nand g216 (n_455, n_282, n_283);
  nand g219 (n_333, n_286, n_287);
  nor g220 (n_289, n_145, n_288);
  nor g223 (n_343, n_145, n_291);
  nor g229 (n_297, n_295, n_288);
  nor g232 (n_349, n_291, n_295);
  nor g233 (n_301, n_299, n_288);
  nor g236 (n_352, n_291, n_299);
  nor g237 (n_304, n_169, n_303);
  nor g240 (n_401, n_169, n_306);
  nor g246 (n_312, n_310, n_303);
  nor g249 (n_407, n_306, n_310);
  nor g250 (n_316, n_314, n_303);
  nor g253 (n_358, n_306, n_314);
  nor g254 (n_319, n_193, n_318);
  nor g257 (n_371, n_193, n_321);
  nor g263 (n_327, n_325, n_318);
  nor g266 (n_381, n_321, n_325);
  nand g273 (n_459, n_128, n_335);
  nand g274 (n_336, n_219, n_333);
  nand g275 (n_461, n_216, n_336);
  nand g278 (n_464, n_339, n_340);
  nand g281 (n_467, n_288, n_342);
  nand g282 (n_345, n_343, n_333);
  nand g283 (n_470, n_344, n_345);
  nand g284 (n_348, n_346, n_333);
  nand g285 (n_472, n_347, n_348);
  nand g286 (n_351, n_349, n_333);
  nand g287 (n_475, n_350, n_351);
  nand g288 (n_354, n_352, n_333);
  nand g289 (n_391, n_353, n_354);
  nor g290 (n_356, n_181, n_355);
  nand g299 (n_415, n_259, n_358);
  nor g300 (n_365, n_363, n_355);
  nor g305 (n_368, n_321, n_355);
  nand g314 (n_427, n_358, n_371);
  nand g319 (n_431, n_358, n_376);
  nand g324 (n_435, n_358, n_381);
  nand g332 (n_479, n_152, n_393);
  nand g333 (n_394, n_239, n_391);
  nand g334 (n_481, n_236, n_394);
  nand g337 (n_484, n_397, n_398);
  nand g340 (n_487, n_303, n_400);
  nand g341 (n_403, n_401, n_391);
  nand g342 (n_490, n_402, n_403);
  nand g343 (n_406, n_404, n_391);
  nand g344 (n_492, n_405, n_406);
  nand g345 (n_409, n_407, n_391);
  nand g346 (n_495, n_408, n_409);
  nand g347 (n_410, n_358, n_391);
  nand g348 (n_497, n_355, n_410);
  nand g351 (n_500, n_413, n_414);
  nand g354 (n_502, n_417, n_418);
  nand g357 (n_505, n_421, n_422);
  nand g360 (n_508, n_425, n_426);
  nand g363 (n_511, n_429, n_430);
  nand g366 (n_513, n_433, n_434);
  nand g369 (n_516, n_437, n_438);
  xnor g376 (Z[2], n_200, n_444);
  xnor g379 (Z[3], n_446, n_447);
  xnor g381 (Z[4], n_276, n_448);
  xnor g384 (Z[5], n_450, n_451);
  xnor g386 (Z[6], n_452, n_453);
  xnor g389 (Z[7], n_455, n_456);
  xnor g391 (Z[8], n_333, n_457);
  xnor g394 (Z[9], n_459, n_460);
  xnor g396 (Z[10], n_461, n_462);
  xnor g399 (Z[11], n_464, n_465);
  xnor g402 (Z[12], n_467, n_468);
  xnor g405 (Z[13], n_470, n_471);
  xnor g407 (Z[14], n_472, n_473);
  xnor g410 (Z[15], n_475, n_476);
  xnor g412 (Z[16], n_391, n_477);
  xnor g415 (Z[17], n_479, n_480);
  xnor g417 (Z[18], n_481, n_482);
  xnor g420 (Z[19], n_484, n_485);
  xnor g423 (Z[20], n_487, n_488);
  xnor g426 (Z[21], n_490, n_491);
  xnor g428 (Z[22], n_492, n_493);
  xnor g431 (Z[23], n_495, n_496);
  xnor g433 (Z[24], n_497, n_498);
  xnor g436 (Z[25], n_500, n_501);
  xnor g438 (Z[26], n_502, n_503);
  xnor g441 (Z[27], n_505, n_506);
  xnor g444 (Z[28], n_508, n_509);
  xnor g447 (Z[29], n_511, n_512);
  xnor g449 (Z[30], n_513, n_514);
  xnor g452 (Z[31], n_516, n_517);
  and g455 (n_195, A[31], B[31]);
  or g456 (n_196, A[31], B[31]);
  or g457 (n_109, n_102, n_105);
  and g458 (n_204, wc, n_112);
  not gc (wc, n_113);
  and g459 (n_206, wc0, n_118);
  not gc0 (wc0, n_119);
  and g460 (n_213, wc1, n_124);
  not gc1 (wc1, n_125);
  and g461 (n_216, wc2, n_130);
  not gc2 (wc2, n_131);
  and g462 (n_223, wc3, n_136);
  not gc3 (wc3, n_137);
  and g463 (n_226, wc4, n_142);
  not gc4 (wc4, n_143);
  and g464 (n_233, wc5, n_148);
  not gc5 (wc5, n_149);
  and g465 (n_236, wc6, n_154);
  not gc6 (wc6, n_155);
  and g466 (n_243, wc7, n_160);
  not gc7 (wc7, n_161);
  and g467 (n_246, wc8, n_166);
  not gc8 (wc8, n_167);
  and g468 (n_253, wc9, n_172);
  not gc9 (wc9, n_173);
  and g469 (n_256, wc10, n_178);
  not gc10 (wc10, n_179);
  and g470 (n_263, wc11, n_184);
  not gc11 (wc11, n_185);
  and g471 (n_266, wc12, n_190);
  not gc12 (wc12, n_191);
  or g472 (n_280, wc13, n_127);
  not gc13 (wc13, n_209);
  or g473 (n_337, wc14, n_139);
  not gc14 (wc14, n_219);
  or g474 (n_295, wc15, n_151);
  not gc15 (wc15, n_229);
  or g475 (n_395, wc16, n_163);
  not gc16 (wc16, n_239);
  or g476 (n_310, wc17, n_175);
  not gc17 (wc17, n_249);
  or g477 (n_363, wc18, n_187);
  not gc18 (wc18, n_259);
  or g478 (n_325, wc19, n_199);
  not gc19 (wc19, n_269);
  or g479 (n_443, wc20, n_105);
  not gc20 (wc20, n_108);
  or g480 (n_444, wc21, n_115);
  not gc21 (wc21, n_110);
  or g481 (n_447, wc22, n_111);
  not gc22 (wc22, n_112);
  or g482 (n_448, wc23, n_121);
  not gc23 (wc23, n_116);
  or g483 (n_451, wc24, n_117);
  not gc24 (wc24, n_118);
  or g484 (n_453, wc25, n_127);
  not gc25 (wc25, n_122);
  or g485 (n_456, wc26, n_123);
  not gc26 (wc26, n_124);
  or g486 (n_457, wc27, n_133);
  not gc27 (wc27, n_128);
  or g487 (n_460, wc28, n_129);
  not gc28 (wc28, n_130);
  or g488 (n_462, wc29, n_139);
  not gc29 (wc29, n_134);
  or g489 (n_465, wc30, n_135);
  not gc30 (wc30, n_136);
  or g490 (n_468, wc31, n_145);
  not gc31 (wc31, n_140);
  or g491 (n_471, wc32, n_141);
  not gc32 (wc32, n_142);
  or g492 (n_473, wc33, n_151);
  not gc33 (wc33, n_146);
  or g493 (n_476, wc34, n_147);
  not gc34 (wc34, n_148);
  or g494 (n_477, wc35, n_157);
  not gc35 (wc35, n_152);
  or g495 (n_480, wc36, n_153);
  not gc36 (wc36, n_154);
  or g496 (n_482, wc37, n_163);
  not gc37 (wc37, n_158);
  or g497 (n_485, wc38, n_159);
  not gc38 (wc38, n_160);
  or g498 (n_488, wc39, n_169);
  not gc39 (wc39, n_164);
  or g499 (n_491, wc40, n_165);
  not gc40 (wc40, n_166);
  or g500 (n_493, wc41, n_175);
  not gc41 (wc41, n_170);
  or g501 (n_496, wc42, n_171);
  not gc42 (wc42, n_172);
  or g502 (n_498, wc43, n_181);
  not gc43 (wc43, n_176);
  or g503 (n_501, wc44, n_177);
  not gc44 (wc44, n_178);
  or g504 (n_503, wc45, n_187);
  not gc45 (wc45, n_182);
  or g505 (n_506, wc46, n_183);
  not gc46 (wc46, n_184);
  or g506 (n_509, wc47, n_193);
  not gc47 (wc47, n_188);
  or g507 (n_512, wc48, n_189);
  not gc48 (wc48, n_190);
  or g508 (n_514, wc49, n_199);
  not gc49 (wc49, n_194);
  and g509 (n_214, wc50, n_211);
  not gc50 (wc50, n_206);
  and g510 (n_224, wc51, n_221);
  not gc51 (wc51, n_216);
  and g511 (n_234, wc52, n_231);
  not gc52 (wc52, n_226);
  and g512 (n_244, wc53, n_241);
  not gc53 (wc53, n_236);
  and g513 (n_254, wc54, n_251);
  not gc54 (wc54, n_246);
  and g514 (n_264, wc55, n_261);
  not gc55 (wc55, n_256);
  and g515 (n_346, wc56, n_229);
  not gc56 (wc56, n_291);
  and g516 (n_404, wc57, n_249);
  not gc57 (wc57, n_306);
  and g517 (n_376, wc58, n_269);
  not gc58 (wc58, n_321);
  xor g518 (Z[1], n_102, n_443);
  or g519 (n_517, wc59, n_195);
  not gc59 (wc59, n_196);
  or g520 (n_202, wc60, n_115);
  not gc60 (wc60, n_200);
  and g521 (n_282, wc61, n_122);
  not gc61 (wc61, n_207);
  and g522 (n_286, wc62, n_213);
  not gc62 (wc62, n_214);
  and g523 (n_339, wc63, n_134);
  not gc63 (wc63, n_217);
  and g524 (n_288, wc64, n_223);
  not gc64 (wc64, n_224);
  and g525 (n_296, wc65, n_146);
  not gc65 (wc65, n_227);
  and g526 (n_300, wc66, n_233);
  not gc66 (wc66, n_234);
  and g527 (n_397, wc67, n_158);
  not gc67 (wc67, n_237);
  and g528 (n_303, wc68, n_243);
  not gc68 (wc68, n_244);
  and g529 (n_311, wc69, n_170);
  not gc69 (wc69, n_247);
  and g530 (n_315, wc70, n_253);
  not gc70 (wc70, n_254);
  and g531 (n_364, wc71, n_182);
  not gc71 (wc71, n_257);
  and g532 (n_318, wc72, n_263);
  not gc72 (wc72, n_264);
  and g533 (n_326, wc73, n_194);
  not gc73 (wc73, n_267);
  or g534 (n_411, wc74, n_181);
  not gc74 (wc74, n_358);
  or g535 (n_419, n_363, wc75);
  not gc75 (wc75, n_358);
  or g536 (n_423, wc76, n_321);
  not gc76 (wc76, n_358);
  and g537 (n_293, wc77, n_229);
  not gc77 (wc77, n_288);
  and g538 (n_308, wc78, n_249);
  not gc78 (wc78, n_303);
  and g539 (n_323, wc79, n_269);
  not gc79 (wc79, n_318);
  or g540 (n_278, wc80, n_121);
  not gc80 (wc80, n_276);
  or g541 (n_283, n_280, wc81);
  not gc81 (wc81, n_276);
  or g542 (n_287, n_284, wc82);
  not gc82 (wc82, n_276);
  and g543 (n_344, wc83, n_140);
  not gc83 (wc83, n_289);
  and g544 (n_347, wc84, n_226);
  not gc84 (wc84, n_293);
  and g545 (n_350, n_296, wc85);
  not gc85 (wc85, n_297);
  and g546 (n_353, n_300, wc86);
  not gc86 (wc86, n_301);
  and g547 (n_402, wc87, n_164);
  not gc87 (wc87, n_304);
  and g548 (n_405, wc88, n_246);
  not gc88 (wc88, n_308);
  and g549 (n_408, n_311, wc89);
  not gc89 (wc89, n_312);
  and g550 (n_355, n_315, wc90);
  not gc90 (wc90, n_316);
  and g551 (n_373, wc91, n_188);
  not gc91 (wc91, n_319);
  and g552 (n_378, wc92, n_266);
  not gc92 (wc92, n_323);
  and g553 (n_383, n_326, wc93);
  not gc93 (wc93, n_327);
  and g554 (n_361, wc94, n_259);
  not gc94 (wc94, n_355);
  and g555 (n_374, wc95, n_371);
  not gc95 (wc95, n_355);
  and g556 (n_379, wc96, n_376);
  not gc96 (wc96, n_355);
  and g557 (n_384, wc97, n_381);
  not gc97 (wc97, n_355);
  or g558 (n_335, wc98, n_133);
  not gc98 (wc98, n_333);
  or g559 (n_340, n_337, wc99);
  not gc99 (wc99, n_333);
  or g560 (n_342, wc100, n_291);
  not gc100 (wc100, n_333);
  and g561 (n_413, wc101, n_176);
  not gc101 (wc101, n_356);
  and g562 (n_417, wc102, n_256);
  not gc102 (wc102, n_361);
  and g563 (n_421, n_364, wc103);
  not gc103 (wc103, n_365);
  and g564 (n_425, n_318, wc104);
  not gc104 (wc104, n_368);
  and g565 (n_429, wc105, n_373);
  not gc105 (wc105, n_374);
  and g566 (n_433, wc106, n_378);
  not gc106 (wc106, n_379);
  and g567 (n_437, wc107, n_383);
  not gc107 (wc107, n_384);
  or g568 (n_393, wc108, n_157);
  not gc108 (wc108, n_391);
  or g569 (n_398, n_395, wc109);
  not gc109 (wc109, n_391);
  or g570 (n_400, wc110, n_306);
  not gc110 (wc110, n_391);
  or g571 (n_414, n_411, wc111);
  not gc111 (wc111, n_391);
  or g572 (n_418, n_415, wc112);
  not gc112 (wc112, n_391);
  or g573 (n_422, n_419, wc113);
  not gc113 (wc113, n_391);
  or g574 (n_426, n_423, wc114);
  not gc114 (wc114, n_391);
  or g575 (n_430, n_427, wc115);
  not gc115 (wc115, n_391);
  or g576 (n_434, n_431, wc116);
  not gc116 (wc116, n_391);
  or g577 (n_438, n_435, wc117);
  not gc117 (wc117, n_391);
endmodule

module add_signed_9092_GENERIC(A, B, Z);
  input [32:0] A, B;
  output [31:0] Z;
  wire [32:0] A, B;
  wire [31:0] Z;
  add_signed_9092_GENERIC_REAL g1(.A ({A[32], A[30], A[30:0]}), .B
       ({B[32], B[30], B[30:0]}), .Z (Z));
endmodule

module add_signed_9095_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [23:0] A, B;
  output [22:0] Z;
  wire [23:0] A, B;
  wire [22:0] Z;
  wire n_75, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_188;
  nand g4 (n_75, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_120, A[9], B[9]);
  nand g59 (n_121, A[9], n_119);
  nand g60 (n_122, B[9], n_119);
  nand g61 (n_124, n_120, n_121, n_122);
  xor g62 (n_123, A[9], B[9]);
  xor g63 (Z[9], n_119, n_123);
  nand g64 (n_125, A[10], B[10]);
  nand g65 (n_126, A[10], n_124);
  nand g66 (n_127, B[10], n_124);
  nand g67 (n_129, n_125, n_126, n_127);
  xor g68 (n_128, A[10], B[10]);
  xor g69 (Z[10], n_124, n_128);
  nand g70 (n_130, A[11], B[11]);
  nand g71 (n_131, A[11], n_129);
  nand g72 (n_132, B[11], n_129);
  nand g73 (n_134, n_130, n_131, n_132);
  xor g74 (n_133, A[11], B[11]);
  xor g75 (Z[11], n_129, n_133);
  nand g76 (n_135, A[12], B[12]);
  nand g77 (n_136, A[12], n_134);
  nand g78 (n_137, B[12], n_134);
  nand g79 (n_139, n_135, n_136, n_137);
  xor g80 (n_138, A[12], B[12]);
  xor g81 (Z[12], n_134, n_138);
  nand g82 (n_140, A[13], B[13]);
  nand g83 (n_141, A[13], n_139);
  nand g84 (n_142, B[13], n_139);
  nand g85 (n_144, n_140, n_141, n_142);
  xor g86 (n_143, A[13], B[13]);
  xor g87 (Z[13], n_139, n_143);
  nand g88 (n_145, A[14], B[14]);
  nand g89 (n_146, A[14], n_144);
  nand g90 (n_147, B[14], n_144);
  nand g91 (n_149, n_145, n_146, n_147);
  xor g92 (n_148, A[14], B[14]);
  xor g93 (Z[14], n_144, n_148);
  nand g94 (n_150, A[15], B[15]);
  nand g95 (n_151, A[15], n_149);
  nand g96 (n_152, B[15], n_149);
  nand g97 (n_154, n_150, n_151, n_152);
  xor g98 (n_153, A[15], B[15]);
  xor g99 (Z[15], n_149, n_153);
  nand g100 (n_155, A[16], B[16]);
  nand g101 (n_156, A[16], n_154);
  nand g102 (n_157, B[16], n_154);
  nand g103 (n_159, n_155, n_156, n_157);
  xor g104 (n_158, A[16], B[16]);
  xor g105 (Z[16], n_154, n_158);
  nand g106 (n_160, A[17], B[17]);
  nand g107 (n_161, A[17], n_159);
  nand g108 (n_162, B[17], n_159);
  nand g109 (n_164, n_160, n_161, n_162);
  xor g110 (n_163, A[17], B[17]);
  xor g111 (Z[17], n_159, n_163);
  nand g112 (n_165, A[18], B[18]);
  nand g113 (n_166, A[18], n_164);
  nand g114 (n_167, B[18], n_164);
  nand g115 (n_169, n_165, n_166, n_167);
  xor g116 (n_168, A[18], B[18]);
  xor g117 (Z[18], n_164, n_168);
  nand g118 (n_170, A[19], B[19]);
  nand g119 (n_171, A[19], n_169);
  nand g120 (n_172, B[19], n_169);
  nand g121 (n_174, n_170, n_171, n_172);
  xor g122 (n_173, A[19], B[19]);
  xor g123 (Z[19], n_169, n_173);
  nand g124 (n_175, A[20], B[20]);
  nand g125 (n_176, A[20], n_174);
  nand g126 (n_177, B[20], n_174);
  nand g127 (n_179, n_175, n_176, n_177);
  xor g128 (n_178, A[20], B[20]);
  xor g129 (Z[20], n_174, n_178);
  nand g130 (n_180, A[21], B[21]);
  nand g131 (n_181, A[21], n_179);
  nand g132 (n_182, B[21], n_179);
  nand g133 (n_184, n_180, n_181, n_182);
  xor g134 (n_183, A[21], B[21]);
  xor g135 (Z[21], n_179, n_183);
  xor g141 (Z[22], n_184, n_188);
  xor g143 (n_188, A[22], B[22]);
  or g144 (n_81, wc, n_75);
  not gc (wc, A[1]);
  or g145 (n_82, wc0, n_75);
  not gc0 (wc0, B[1]);
  xnor g146 (Z[1], n_75, n_83);
endmodule

module add_signed_9095_GENERIC(A, B, Z);
  input [23:0] A, B;
  output [22:0] Z;
  wire [23:0] A, B;
  wire [22:0] Z;
  add_signed_9095_GENERIC_REAL g1(.A ({A[23], A[20], A[20], A[20:0]}),
       .B ({B[23], B[20], B[20], B[20:0]}), .Z (Z));
endmodule

module add_signed_9162_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [24:0] A, B;
  output [23:0] Z;
  wire [24:0] A, B;
  wire [23:0] Z;
  wire n_78, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_196;
  nand g4 (n_78, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_83, A[1], B[1]);
  nand g13 (n_87, n_83, n_84, n_85);
  xor g14 (n_86, A[1], B[1]);
  nand g16 (n_88, A[2], B[2]);
  nand g17 (n_89, A[2], n_87);
  nand g18 (n_90, B[2], n_87);
  nand g19 (n_92, n_88, n_89, n_90);
  xor g20 (n_91, A[2], B[2]);
  xor g21 (Z[2], n_87, n_91);
  nand g22 (n_93, A[3], B[3]);
  nand g23 (n_94, A[3], n_92);
  nand g24 (n_95, B[3], n_92);
  nand g25 (n_97, n_93, n_94, n_95);
  xor g26 (n_96, A[3], B[3]);
  xor g27 (Z[3], n_92, n_96);
  nand g28 (n_98, A[4], B[4]);
  nand g29 (n_99, A[4], n_97);
  nand g30 (n_100, B[4], n_97);
  nand g31 (n_102, n_98, n_99, n_100);
  xor g32 (n_101, A[4], B[4]);
  xor g33 (Z[4], n_97, n_101);
  nand g34 (n_103, A[5], B[5]);
  nand g35 (n_104, A[5], n_102);
  nand g36 (n_105, B[5], n_102);
  nand g37 (n_107, n_103, n_104, n_105);
  xor g38 (n_106, A[5], B[5]);
  xor g39 (Z[5], n_102, n_106);
  nand g40 (n_108, A[6], B[6]);
  nand g41 (n_109, A[6], n_107);
  nand g42 (n_110, B[6], n_107);
  nand g43 (n_112, n_108, n_109, n_110);
  xor g44 (n_111, A[6], B[6]);
  xor g45 (Z[6], n_107, n_111);
  nand g46 (n_113, A[7], B[7]);
  nand g47 (n_114, A[7], n_112);
  nand g48 (n_115, B[7], n_112);
  nand g49 (n_117, n_113, n_114, n_115);
  xor g50 (n_116, A[7], B[7]);
  xor g51 (Z[7], n_112, n_116);
  nand g52 (n_118, A[8], B[8]);
  nand g53 (n_119, A[8], n_117);
  nand g54 (n_120, B[8], n_117);
  nand g55 (n_122, n_118, n_119, n_120);
  xor g56 (n_121, A[8], B[8]);
  xor g57 (Z[8], n_117, n_121);
  nand g58 (n_123, A[9], B[9]);
  nand g59 (n_124, A[9], n_122);
  nand g60 (n_125, B[9], n_122);
  nand g61 (n_127, n_123, n_124, n_125);
  xor g62 (n_126, A[9], B[9]);
  xor g63 (Z[9], n_122, n_126);
  nand g64 (n_128, A[10], B[10]);
  nand g65 (n_129, A[10], n_127);
  nand g66 (n_130, B[10], n_127);
  nand g67 (n_132, n_128, n_129, n_130);
  xor g68 (n_131, A[10], B[10]);
  xor g69 (Z[10], n_127, n_131);
  nand g70 (n_133, A[11], B[11]);
  nand g71 (n_134, A[11], n_132);
  nand g72 (n_135, B[11], n_132);
  nand g73 (n_137, n_133, n_134, n_135);
  xor g74 (n_136, A[11], B[11]);
  xor g75 (Z[11], n_132, n_136);
  nand g76 (n_138, A[12], B[12]);
  nand g77 (n_139, A[12], n_137);
  nand g78 (n_140, B[12], n_137);
  nand g79 (n_142, n_138, n_139, n_140);
  xor g80 (n_141, A[12], B[12]);
  xor g81 (Z[12], n_137, n_141);
  nand g82 (n_143, A[13], B[13]);
  nand g83 (n_144, A[13], n_142);
  nand g84 (n_145, B[13], n_142);
  nand g85 (n_147, n_143, n_144, n_145);
  xor g86 (n_146, A[13], B[13]);
  xor g87 (Z[13], n_142, n_146);
  nand g88 (n_148, A[14], B[14]);
  nand g89 (n_149, A[14], n_147);
  nand g90 (n_150, B[14], n_147);
  nand g91 (n_152, n_148, n_149, n_150);
  xor g92 (n_151, A[14], B[14]);
  xor g93 (Z[14], n_147, n_151);
  nand g94 (n_153, A[15], B[15]);
  nand g95 (n_154, A[15], n_152);
  nand g96 (n_155, B[15], n_152);
  nand g97 (n_157, n_153, n_154, n_155);
  xor g98 (n_156, A[15], B[15]);
  xor g99 (Z[15], n_152, n_156);
  nand g100 (n_158, A[16], B[16]);
  nand g101 (n_159, A[16], n_157);
  nand g102 (n_160, B[16], n_157);
  nand g103 (n_162, n_158, n_159, n_160);
  xor g104 (n_161, A[16], B[16]);
  xor g105 (Z[16], n_157, n_161);
  nand g106 (n_163, A[17], B[17]);
  nand g107 (n_164, A[17], n_162);
  nand g108 (n_165, B[17], n_162);
  nand g109 (n_167, n_163, n_164, n_165);
  xor g110 (n_166, A[17], B[17]);
  xor g111 (Z[17], n_162, n_166);
  nand g112 (n_168, A[18], B[18]);
  nand g113 (n_169, A[18], n_167);
  nand g114 (n_170, B[18], n_167);
  nand g115 (n_172, n_168, n_169, n_170);
  xor g116 (n_171, A[18], B[18]);
  xor g117 (Z[18], n_167, n_171);
  nand g118 (n_173, A[19], B[19]);
  nand g119 (n_174, A[19], n_172);
  nand g120 (n_175, B[19], n_172);
  nand g121 (n_177, n_173, n_174, n_175);
  xor g122 (n_176, A[19], B[19]);
  xor g123 (Z[19], n_172, n_176);
  nand g124 (n_178, A[20], B[20]);
  nand g125 (n_179, A[20], n_177);
  nand g126 (n_180, B[20], n_177);
  nand g127 (n_182, n_178, n_179, n_180);
  xor g128 (n_181, A[20], B[20]);
  xor g129 (Z[20], n_177, n_181);
  nand g130 (n_183, A[21], B[21]);
  nand g131 (n_184, A[21], n_182);
  nand g132 (n_185, B[21], n_182);
  nand g133 (n_187, n_183, n_184, n_185);
  xor g134 (n_186, A[21], B[21]);
  xor g135 (Z[21], n_182, n_186);
  nand g136 (n_188, A[22], B[22]);
  nand g137 (n_189, A[22], n_187);
  nand g138 (n_190, B[22], n_187);
  nand g139 (n_192, n_188, n_189, n_190);
  xor g140 (n_191, A[22], B[22]);
  xor g141 (Z[22], n_187, n_191);
  xor g147 (Z[23], n_192, n_196);
  xor g149 (n_196, A[23], B[23]);
  or g150 (n_84, wc, n_78);
  not gc (wc, A[1]);
  or g151 (n_85, wc0, n_78);
  not gc0 (wc0, B[1]);
  xnor g152 (Z[1], n_78, n_86);
endmodule

module add_signed_9162_GENERIC(A, B, Z);
  input [24:0] A, B;
  output [23:0] Z;
  wire [24:0] A, B;
  wire [23:0] Z;
  add_signed_9162_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_9196_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [35:0] A, B;
  output [34:0] Z;
  wire [35:0] A, B;
  wire [34:0] Z;
  wire n_111, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_284;
  nand g4 (n_111, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_116, A[1], B[1]);
  nand g13 (n_120, n_116, n_117, n_118);
  xor g14 (n_119, A[1], B[1]);
  nand g16 (n_121, A[2], B[2]);
  nand g17 (n_122, A[2], n_120);
  nand g18 (n_123, B[2], n_120);
  nand g19 (n_125, n_121, n_122, n_123);
  xor g20 (n_124, A[2], B[2]);
  xor g21 (Z[2], n_120, n_124);
  nand g22 (n_126, A[3], B[3]);
  nand g23 (n_127, A[3], n_125);
  nand g24 (n_128, B[3], n_125);
  nand g25 (n_130, n_126, n_127, n_128);
  xor g26 (n_129, A[3], B[3]);
  xor g27 (Z[3], n_125, n_129);
  nand g28 (n_131, A[4], B[4]);
  nand g29 (n_132, A[4], n_130);
  nand g30 (n_133, B[4], n_130);
  nand g31 (n_135, n_131, n_132, n_133);
  xor g32 (n_134, A[4], B[4]);
  xor g33 (Z[4], n_130, n_134);
  nand g34 (n_136, A[5], B[5]);
  nand g35 (n_137, A[5], n_135);
  nand g36 (n_138, B[5], n_135);
  nand g37 (n_140, n_136, n_137, n_138);
  xor g38 (n_139, A[5], B[5]);
  xor g39 (Z[5], n_135, n_139);
  nand g40 (n_141, A[6], B[6]);
  nand g41 (n_142, A[6], n_140);
  nand g42 (n_143, B[6], n_140);
  nand g43 (n_145, n_141, n_142, n_143);
  xor g44 (n_144, A[6], B[6]);
  xor g45 (Z[6], n_140, n_144);
  nand g46 (n_146, A[7], B[7]);
  nand g47 (n_147, A[7], n_145);
  nand g48 (n_148, B[7], n_145);
  nand g49 (n_150, n_146, n_147, n_148);
  xor g50 (n_149, A[7], B[7]);
  xor g51 (Z[7], n_145, n_149);
  nand g52 (n_151, A[8], B[8]);
  nand g53 (n_152, A[8], n_150);
  nand g54 (n_153, B[8], n_150);
  nand g55 (n_155, n_151, n_152, n_153);
  xor g56 (n_154, A[8], B[8]);
  xor g57 (Z[8], n_150, n_154);
  nand g58 (n_156, A[9], B[9]);
  nand g59 (n_157, A[9], n_155);
  nand g60 (n_158, B[9], n_155);
  nand g61 (n_160, n_156, n_157, n_158);
  xor g62 (n_159, A[9], B[9]);
  xor g63 (Z[9], n_155, n_159);
  nand g64 (n_161, A[10], B[10]);
  nand g65 (n_162, A[10], n_160);
  nand g66 (n_163, B[10], n_160);
  nand g67 (n_165, n_161, n_162, n_163);
  xor g68 (n_164, A[10], B[10]);
  xor g69 (Z[10], n_160, n_164);
  nand g70 (n_166, A[11], B[11]);
  nand g71 (n_167, A[11], n_165);
  nand g72 (n_168, B[11], n_165);
  nand g73 (n_170, n_166, n_167, n_168);
  xor g74 (n_169, A[11], B[11]);
  xor g75 (Z[11], n_165, n_169);
  nand g76 (n_171, A[12], B[12]);
  nand g77 (n_172, A[12], n_170);
  nand g78 (n_173, B[12], n_170);
  nand g79 (n_175, n_171, n_172, n_173);
  xor g80 (n_174, A[12], B[12]);
  xor g81 (Z[12], n_170, n_174);
  nand g82 (n_176, A[13], B[13]);
  nand g83 (n_177, A[13], n_175);
  nand g84 (n_178, B[13], n_175);
  nand g85 (n_180, n_176, n_177, n_178);
  xor g86 (n_179, A[13], B[13]);
  xor g87 (Z[13], n_175, n_179);
  nand g88 (n_181, A[14], B[14]);
  nand g89 (n_182, A[14], n_180);
  nand g90 (n_183, B[14], n_180);
  nand g91 (n_185, n_181, n_182, n_183);
  xor g92 (n_184, A[14], B[14]);
  xor g93 (Z[14], n_180, n_184);
  nand g94 (n_186, A[15], B[15]);
  nand g95 (n_187, A[15], n_185);
  nand g96 (n_188, B[15], n_185);
  nand g97 (n_190, n_186, n_187, n_188);
  xor g98 (n_189, A[15], B[15]);
  xor g99 (Z[15], n_185, n_189);
  nand g100 (n_191, A[16], B[16]);
  nand g101 (n_192, A[16], n_190);
  nand g102 (n_193, B[16], n_190);
  nand g103 (n_195, n_191, n_192, n_193);
  xor g104 (n_194, A[16], B[16]);
  xor g105 (Z[16], n_190, n_194);
  nand g106 (n_196, A[17], B[17]);
  nand g107 (n_197, A[17], n_195);
  nand g108 (n_198, B[17], n_195);
  nand g109 (n_200, n_196, n_197, n_198);
  xor g110 (n_199, A[17], B[17]);
  xor g111 (Z[17], n_195, n_199);
  nand g112 (n_201, A[18], B[18]);
  nand g113 (n_202, A[18], n_200);
  nand g114 (n_203, B[18], n_200);
  nand g115 (n_205, n_201, n_202, n_203);
  xor g116 (n_204, A[18], B[18]);
  xor g117 (Z[18], n_200, n_204);
  nand g118 (n_206, A[19], B[19]);
  nand g119 (n_207, A[19], n_205);
  nand g120 (n_208, B[19], n_205);
  nand g121 (n_210, n_206, n_207, n_208);
  xor g122 (n_209, A[19], B[19]);
  xor g123 (Z[19], n_205, n_209);
  nand g124 (n_211, A[20], B[20]);
  nand g125 (n_212, A[20], n_210);
  nand g126 (n_213, B[20], n_210);
  nand g127 (n_215, n_211, n_212, n_213);
  xor g128 (n_214, A[20], B[20]);
  xor g129 (Z[20], n_210, n_214);
  nand g130 (n_216, A[21], B[21]);
  nand g131 (n_217, A[21], n_215);
  nand g132 (n_218, B[21], n_215);
  nand g133 (n_220, n_216, n_217, n_218);
  xor g134 (n_219, A[21], B[21]);
  xor g135 (Z[21], n_215, n_219);
  nand g136 (n_221, A[22], B[22]);
  nand g137 (n_222, A[22], n_220);
  nand g138 (n_223, B[22], n_220);
  nand g139 (n_225, n_221, n_222, n_223);
  xor g140 (n_224, A[22], B[22]);
  xor g141 (Z[22], n_220, n_224);
  nand g142 (n_226, A[23], B[23]);
  nand g143 (n_227, A[23], n_225);
  nand g144 (n_228, B[23], n_225);
  nand g145 (n_230, n_226, n_227, n_228);
  xor g146 (n_229, A[23], B[23]);
  xor g147 (Z[23], n_225, n_229);
  nand g148 (n_231, A[24], B[24]);
  nand g149 (n_232, A[24], n_230);
  nand g150 (n_233, B[24], n_230);
  nand g151 (n_235, n_231, n_232, n_233);
  xor g152 (n_234, A[24], B[24]);
  xor g153 (Z[24], n_230, n_234);
  nand g154 (n_236, A[25], B[25]);
  nand g155 (n_237, A[25], n_235);
  nand g156 (n_238, B[25], n_235);
  nand g157 (n_240, n_236, n_237, n_238);
  xor g158 (n_239, A[25], B[25]);
  xor g159 (Z[25], n_235, n_239);
  nand g160 (n_241, A[26], B[26]);
  nand g161 (n_242, A[26], n_240);
  nand g162 (n_243, B[26], n_240);
  nand g163 (n_245, n_241, n_242, n_243);
  xor g164 (n_244, A[26], B[26]);
  xor g165 (Z[26], n_240, n_244);
  nand g166 (n_246, A[27], B[27]);
  nand g167 (n_247, A[27], n_245);
  nand g168 (n_248, B[27], n_245);
  nand g169 (n_250, n_246, n_247, n_248);
  xor g170 (n_249, A[27], B[27]);
  xor g171 (Z[27], n_245, n_249);
  nand g172 (n_251, A[28], B[28]);
  nand g173 (n_252, A[28], n_250);
  nand g174 (n_253, B[28], n_250);
  nand g175 (n_255, n_251, n_252, n_253);
  xor g176 (n_254, A[28], B[28]);
  xor g177 (Z[28], n_250, n_254);
  nand g178 (n_256, A[29], B[29]);
  nand g179 (n_257, A[29], n_255);
  nand g180 (n_258, B[29], n_255);
  nand g181 (n_260, n_256, n_257, n_258);
  xor g182 (n_259, A[29], B[29]);
  xor g183 (Z[29], n_255, n_259);
  nand g184 (n_261, A[30], B[30]);
  nand g185 (n_262, A[30], n_260);
  nand g186 (n_263, B[30], n_260);
  nand g187 (n_265, n_261, n_262, n_263);
  xor g188 (n_264, A[30], B[30]);
  xor g189 (Z[30], n_260, n_264);
  nand g190 (n_266, A[31], B[31]);
  nand g191 (n_267, A[31], n_265);
  nand g192 (n_268, B[31], n_265);
  nand g193 (n_270, n_266, n_267, n_268);
  xor g194 (n_269, A[31], B[31]);
  xor g195 (Z[31], n_265, n_269);
  nand g196 (n_271, A[32], B[32]);
  nand g197 (n_272, A[32], n_270);
  nand g198 (n_273, B[32], n_270);
  nand g199 (n_275, n_271, n_272, n_273);
  xor g200 (n_274, A[32], B[32]);
  xor g201 (Z[32], n_270, n_274);
  nand g202 (n_276, A[33], B[33]);
  nand g203 (n_277, A[33], n_275);
  nand g204 (n_278, B[33], n_275);
  nand g205 (n_280, n_276, n_277, n_278);
  xor g206 (n_279, A[33], B[33]);
  xor g207 (Z[33], n_275, n_279);
  xor g213 (Z[34], n_280, n_284);
  xor g215 (n_284, A[34], B[34]);
  or g216 (n_117, wc, n_111);
  not gc (wc, A[1]);
  or g217 (n_118, wc0, n_111);
  not gc0 (wc0, B[1]);
  xnor g218 (Z[1], n_111, n_119);
endmodule

module add_signed_9196_GENERIC(A, B, Z);
  input [35:0] A, B;
  output [34:0] Z;
  wire [35:0] A, B;
  wire [34:0] Z;
  add_signed_9196_GENERIC_REAL g1(.A ({A[35], A[32], A[32], A[32:0]}),
       .B ({B[35], B[32], B[32], B[32:0]}), .Z (Z));
endmodule

module add_signed_9238_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [33:0] A, B;
  output [32:0] Z;
  wire [33:0] A, B;
  wire [32:0] Z;
  wire n_105, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_268;
  nand g4 (n_105, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_110, A[1], B[1]);
  nand g13 (n_114, n_110, n_111, n_112);
  xor g14 (n_113, A[1], B[1]);
  nand g16 (n_115, A[2], B[2]);
  nand g17 (n_116, A[2], n_114);
  nand g18 (n_117, B[2], n_114);
  nand g19 (n_119, n_115, n_116, n_117);
  xor g20 (n_118, A[2], B[2]);
  xor g21 (Z[2], n_114, n_118);
  nand g22 (n_120, A[3], B[3]);
  nand g23 (n_121, A[3], n_119);
  nand g24 (n_122, B[3], n_119);
  nand g25 (n_124, n_120, n_121, n_122);
  xor g26 (n_123, A[3], B[3]);
  xor g27 (Z[3], n_119, n_123);
  nand g28 (n_125, A[4], B[4]);
  nand g29 (n_126, A[4], n_124);
  nand g30 (n_127, B[4], n_124);
  nand g31 (n_129, n_125, n_126, n_127);
  xor g32 (n_128, A[4], B[4]);
  xor g33 (Z[4], n_124, n_128);
  nand g34 (n_130, A[5], B[5]);
  nand g35 (n_131, A[5], n_129);
  nand g36 (n_132, B[5], n_129);
  nand g37 (n_134, n_130, n_131, n_132);
  xor g38 (n_133, A[5], B[5]);
  xor g39 (Z[5], n_129, n_133);
  nand g40 (n_135, A[6], B[6]);
  nand g41 (n_136, A[6], n_134);
  nand g42 (n_137, B[6], n_134);
  nand g43 (n_139, n_135, n_136, n_137);
  xor g44 (n_138, A[6], B[6]);
  xor g45 (Z[6], n_134, n_138);
  nand g46 (n_140, A[7], B[7]);
  nand g47 (n_141, A[7], n_139);
  nand g48 (n_142, B[7], n_139);
  nand g49 (n_144, n_140, n_141, n_142);
  xor g50 (n_143, A[7], B[7]);
  xor g51 (Z[7], n_139, n_143);
  nand g52 (n_145, A[8], B[8]);
  nand g53 (n_146, A[8], n_144);
  nand g54 (n_147, B[8], n_144);
  nand g55 (n_149, n_145, n_146, n_147);
  xor g56 (n_148, A[8], B[8]);
  xor g57 (Z[8], n_144, n_148);
  nand g58 (n_150, A[9], B[9]);
  nand g59 (n_151, A[9], n_149);
  nand g60 (n_152, B[9], n_149);
  nand g61 (n_154, n_150, n_151, n_152);
  xor g62 (n_153, A[9], B[9]);
  xor g63 (Z[9], n_149, n_153);
  nand g64 (n_155, A[10], B[10]);
  nand g65 (n_156, A[10], n_154);
  nand g66 (n_157, B[10], n_154);
  nand g67 (n_159, n_155, n_156, n_157);
  xor g68 (n_158, A[10], B[10]);
  xor g69 (Z[10], n_154, n_158);
  nand g70 (n_160, A[11], B[11]);
  nand g71 (n_161, A[11], n_159);
  nand g72 (n_162, B[11], n_159);
  nand g73 (n_164, n_160, n_161, n_162);
  xor g74 (n_163, A[11], B[11]);
  xor g75 (Z[11], n_159, n_163);
  nand g76 (n_165, A[12], B[12]);
  nand g77 (n_166, A[12], n_164);
  nand g78 (n_167, B[12], n_164);
  nand g79 (n_169, n_165, n_166, n_167);
  xor g80 (n_168, A[12], B[12]);
  xor g81 (Z[12], n_164, n_168);
  nand g82 (n_170, A[13], B[13]);
  nand g83 (n_171, A[13], n_169);
  nand g84 (n_172, B[13], n_169);
  nand g85 (n_174, n_170, n_171, n_172);
  xor g86 (n_173, A[13], B[13]);
  xor g87 (Z[13], n_169, n_173);
  nand g88 (n_175, A[14], B[14]);
  nand g89 (n_176, A[14], n_174);
  nand g90 (n_177, B[14], n_174);
  nand g91 (n_179, n_175, n_176, n_177);
  xor g92 (n_178, A[14], B[14]);
  xor g93 (Z[14], n_174, n_178);
  nand g94 (n_180, A[15], B[15]);
  nand g95 (n_181, A[15], n_179);
  nand g96 (n_182, B[15], n_179);
  nand g97 (n_184, n_180, n_181, n_182);
  xor g98 (n_183, A[15], B[15]);
  xor g99 (Z[15], n_179, n_183);
  nand g100 (n_185, A[16], B[16]);
  nand g101 (n_186, A[16], n_184);
  nand g102 (n_187, B[16], n_184);
  nand g103 (n_189, n_185, n_186, n_187);
  xor g104 (n_188, A[16], B[16]);
  xor g105 (Z[16], n_184, n_188);
  nand g106 (n_190, A[17], B[17]);
  nand g107 (n_191, A[17], n_189);
  nand g108 (n_192, B[17], n_189);
  nand g109 (n_194, n_190, n_191, n_192);
  xor g110 (n_193, A[17], B[17]);
  xor g111 (Z[17], n_189, n_193);
  nand g112 (n_195, A[18], B[18]);
  nand g113 (n_196, A[18], n_194);
  nand g114 (n_197, B[18], n_194);
  nand g115 (n_199, n_195, n_196, n_197);
  xor g116 (n_198, A[18], B[18]);
  xor g117 (Z[18], n_194, n_198);
  nand g118 (n_200, A[19], B[19]);
  nand g119 (n_201, A[19], n_199);
  nand g120 (n_202, B[19], n_199);
  nand g121 (n_204, n_200, n_201, n_202);
  xor g122 (n_203, A[19], B[19]);
  xor g123 (Z[19], n_199, n_203);
  nand g124 (n_205, A[20], B[20]);
  nand g125 (n_206, A[20], n_204);
  nand g126 (n_207, B[20], n_204);
  nand g127 (n_209, n_205, n_206, n_207);
  xor g128 (n_208, A[20], B[20]);
  xor g129 (Z[20], n_204, n_208);
  nand g130 (n_210, A[21], B[21]);
  nand g131 (n_211, A[21], n_209);
  nand g132 (n_212, B[21], n_209);
  nand g133 (n_214, n_210, n_211, n_212);
  xor g134 (n_213, A[21], B[21]);
  xor g135 (Z[21], n_209, n_213);
  nand g136 (n_215, A[22], B[22]);
  nand g137 (n_216, A[22], n_214);
  nand g138 (n_217, B[22], n_214);
  nand g139 (n_219, n_215, n_216, n_217);
  xor g140 (n_218, A[22], B[22]);
  xor g141 (Z[22], n_214, n_218);
  nand g142 (n_220, A[23], B[23]);
  nand g143 (n_221, A[23], n_219);
  nand g144 (n_222, B[23], n_219);
  nand g145 (n_224, n_220, n_221, n_222);
  xor g146 (n_223, A[23], B[23]);
  xor g147 (Z[23], n_219, n_223);
  nand g148 (n_225, A[24], B[24]);
  nand g149 (n_226, A[24], n_224);
  nand g150 (n_227, B[24], n_224);
  nand g151 (n_229, n_225, n_226, n_227);
  xor g152 (n_228, A[24], B[24]);
  xor g153 (Z[24], n_224, n_228);
  nand g154 (n_230, A[25], B[25]);
  nand g155 (n_231, A[25], n_229);
  nand g156 (n_232, B[25], n_229);
  nand g157 (n_234, n_230, n_231, n_232);
  xor g158 (n_233, A[25], B[25]);
  xor g159 (Z[25], n_229, n_233);
  nand g160 (n_235, A[26], B[26]);
  nand g161 (n_236, A[26], n_234);
  nand g162 (n_237, B[26], n_234);
  nand g163 (n_239, n_235, n_236, n_237);
  xor g164 (n_238, A[26], B[26]);
  xor g165 (Z[26], n_234, n_238);
  nand g166 (n_240, A[27], B[27]);
  nand g167 (n_241, A[27], n_239);
  nand g168 (n_242, B[27], n_239);
  nand g169 (n_244, n_240, n_241, n_242);
  xor g170 (n_243, A[27], B[27]);
  xor g171 (Z[27], n_239, n_243);
  nand g172 (n_245, A[28], B[28]);
  nand g173 (n_246, A[28], n_244);
  nand g174 (n_247, B[28], n_244);
  nand g175 (n_249, n_245, n_246, n_247);
  xor g176 (n_248, A[28], B[28]);
  xor g177 (Z[28], n_244, n_248);
  nand g178 (n_250, A[29], B[29]);
  nand g179 (n_251, A[29], n_249);
  nand g180 (n_252, B[29], n_249);
  nand g181 (n_254, n_250, n_251, n_252);
  xor g182 (n_253, A[29], B[29]);
  xor g183 (Z[29], n_249, n_253);
  nand g184 (n_255, A[30], B[30]);
  nand g185 (n_256, A[30], n_254);
  nand g186 (n_257, B[30], n_254);
  nand g187 (n_259, n_255, n_256, n_257);
  xor g188 (n_258, A[30], B[30]);
  xor g189 (Z[30], n_254, n_258);
  nand g190 (n_260, A[31], B[31]);
  nand g191 (n_261, A[31], n_259);
  nand g192 (n_262, B[31], n_259);
  nand g193 (n_264, n_260, n_261, n_262);
  xor g194 (n_263, A[31], B[31]);
  xor g195 (Z[31], n_259, n_263);
  xor g201 (Z[32], n_264, n_268);
  xor g203 (n_268, A[32], B[32]);
  or g204 (n_111, wc, n_105);
  not gc (wc, A[1]);
  or g205 (n_112, wc0, n_105);
  not gc0 (wc0, B[1]);
  xnor g206 (Z[1], n_105, n_113);
endmodule

module add_signed_9238_GENERIC(A, B, Z);
  input [33:0] A, B;
  output [32:0] Z;
  wire [33:0] A, B;
  wire [32:0] Z;
  add_signed_9238_GENERIC_REAL g1(.A ({A[33], A[31], A[31:0]}), .B
       ({B[33], B[31], B[31:0]}), .Z (Z));
endmodule

module add_signed_9277_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [35:0] A, B;
  output [33:0] Z;
  wire [35:0] A, B;
  wire [33:0] Z;
  wire n_109, n_111, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_121, n_122, n_123, n_124, n_125, n_127, n_128, n_129;
  wire n_130, n_131, n_133, n_134, n_135, n_136, n_137, n_139;
  wire n_140, n_141, n_142, n_143, n_145, n_146, n_147, n_148;
  wire n_149, n_151, n_152, n_153, n_154, n_155, n_157, n_158;
  wire n_159, n_160, n_161, n_163, n_164, n_165, n_166, n_167;
  wire n_169, n_170, n_171, n_172, n_173, n_175, n_176, n_177;
  wire n_178, n_179, n_181, n_182, n_183, n_184, n_185, n_187;
  wire n_188, n_189, n_190, n_191, n_193, n_194, n_195, n_196;
  wire n_197, n_199, n_200, n_201, n_202, n_203, n_205, n_206;
  wire n_207, n_208, n_211, n_212, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_221, n_223, n_225, n_226, n_228, n_229;
  wire n_231, n_233, n_235, n_236, n_238, n_239, n_241, n_243;
  wire n_245, n_246, n_248, n_249, n_251, n_253, n_255, n_256;
  wire n_258, n_259, n_261, n_263, n_265, n_266, n_268, n_269;
  wire n_271, n_273, n_275, n_276, n_278, n_279, n_281, n_283;
  wire n_285, n_286, n_288, n_290, n_291, n_292, n_294, n_295;
  wire n_296, n_298, n_299, n_300, n_301, n_303, n_305, n_307;
  wire n_308, n_309, n_311, n_312, n_313, n_315, n_316, n_318;
  wire n_320, n_322, n_323, n_324, n_326, n_327, n_328, n_330;
  wire n_331, n_333, n_335, n_337, n_338, n_339, n_341, n_342;
  wire n_343, n_345, n_347, n_348, n_349, n_351, n_352, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_370, n_373;
  wire n_375, n_376, n_377, n_380, n_383, n_385, n_386, n_388;
  wire n_390, n_391, n_393, n_395, n_396, n_398, n_400, n_401;
  wire n_403, n_405, n_406, n_407, n_409, n_410, n_412, n_413;
  wire n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421;
  wire n_422, n_423, n_425, n_426, n_427, n_429, n_430, n_431;
  wire n_433, n_434, n_435, n_437, n_438, n_439, n_441, n_442;
  wire n_443, n_445, n_446, n_447, n_449, n_450, n_451, n_453;
  wire n_454, n_455, n_457, n_461, n_462, n_464, n_465, n_466;
  wire n_468, n_469, n_470, n_471, n_473, n_474, n_475, n_477;
  wire n_478, n_479, n_480, n_482, n_483, n_485, n_486, n_488;
  wire n_489, n_490, n_491, n_493, n_494, n_495, n_497, n_498;
  wire n_499, n_500, n_502, n_503, n_505, n_506, n_508, n_509;
  wire n_510, n_511, n_513, n_514, n_515, n_516, n_518, n_519;
  wire n_520, n_521, n_523, n_524, n_526, n_527, n_529, n_530;
  wire n_531, n_532, n_534, n_535, n_536, n_538, n_539;
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_109, A[0], B[0]);
  nor g9 (n_111, A[1], B[1]);
  nand g10 (n_114, A[1], B[1]);
  nor g11 (n_121, A[2], B[2]);
  nand g12 (n_116, A[2], B[2]);
  nor g13 (n_117, A[3], B[3]);
  nand g14 (n_118, A[3], B[3]);
  nor g15 (n_127, A[4], B[4]);
  nand g16 (n_122, A[4], B[4]);
  nor g17 (n_123, A[5], B[5]);
  nand g18 (n_124, A[5], B[5]);
  nor g19 (n_133, A[6], B[6]);
  nand g20 (n_128, A[6], B[6]);
  nor g21 (n_129, A[7], B[7]);
  nand g22 (n_130, A[7], B[7]);
  nor g23 (n_139, A[8], B[8]);
  nand g24 (n_134, A[8], B[8]);
  nor g25 (n_135, A[9], B[9]);
  nand g26 (n_136, A[9], B[9]);
  nor g27 (n_145, A[10], B[10]);
  nand g28 (n_140, A[10], B[10]);
  nor g29 (n_141, A[11], B[11]);
  nand g30 (n_142, A[11], B[11]);
  nor g31 (n_151, A[12], B[12]);
  nand g32 (n_146, A[12], B[12]);
  nor g33 (n_147, A[13], B[13]);
  nand g34 (n_148, A[13], B[13]);
  nor g35 (n_157, A[14], B[14]);
  nand g36 (n_152, A[14], B[14]);
  nor g37 (n_153, A[15], B[15]);
  nand g38 (n_154, A[15], B[15]);
  nor g39 (n_163, A[16], B[16]);
  nand g40 (n_158, A[16], B[16]);
  nor g41 (n_159, A[17], B[17]);
  nand g42 (n_160, A[17], B[17]);
  nor g43 (n_169, A[18], B[18]);
  nand g44 (n_164, A[18], B[18]);
  nor g45 (n_165, A[19], B[19]);
  nand g46 (n_166, A[19], B[19]);
  nor g47 (n_175, A[20], B[20]);
  nand g48 (n_170, A[20], B[20]);
  nor g49 (n_171, A[21], B[21]);
  nand g50 (n_172, A[21], B[21]);
  nor g51 (n_181, A[22], B[22]);
  nand g52 (n_176, A[22], B[22]);
  nor g53 (n_177, A[23], B[23]);
  nand g54 (n_178, A[23], B[23]);
  nor g55 (n_187, A[24], B[24]);
  nand g56 (n_182, A[24], B[24]);
  nor g57 (n_183, A[25], B[25]);
  nand g58 (n_184, A[25], B[25]);
  nor g59 (n_193, A[26], B[26]);
  nand g60 (n_188, A[26], B[26]);
  nor g61 (n_189, A[27], B[27]);
  nand g62 (n_190, A[27], B[27]);
  nor g63 (n_199, A[28], B[28]);
  nand g64 (n_194, A[28], B[28]);
  nor g65 (n_195, A[29], B[29]);
  nand g66 (n_196, A[29], B[29]);
  nor g67 (n_205, A[30], B[30]);
  nand g68 (n_200, A[30], B[30]);
  nor g69 (n_201, A[31], B[31]);
  nand g70 (n_202, A[31], B[31]);
  nor g71 (n_211, A[32], B[32]);
  nand g72 (n_206, A[32], B[32]);
  nand g77 (n_212, n_114, n_115);
  nor g78 (n_119, n_116, n_117);
  nor g81 (n_215, n_121, n_117);
  nor g82 (n_125, n_122, n_123);
  nor g85 (n_221, n_127, n_123);
  nor g86 (n_131, n_128, n_129);
  nor g89 (n_223, n_133, n_129);
  nor g90 (n_137, n_134, n_135);
  nor g93 (n_231, n_139, n_135);
  nor g94 (n_143, n_140, n_141);
  nor g97 (n_233, n_145, n_141);
  nor g98 (n_149, n_146, n_147);
  nor g101 (n_241, n_151, n_147);
  nor g102 (n_155, n_152, n_153);
  nor g105 (n_243, n_157, n_153);
  nor g106 (n_161, n_158, n_159);
  nor g109 (n_251, n_163, n_159);
  nor g110 (n_167, n_164, n_165);
  nor g113 (n_253, n_169, n_165);
  nor g114 (n_173, n_170, n_171);
  nor g117 (n_261, n_175, n_171);
  nor g118 (n_179, n_176, n_177);
  nor g121 (n_263, n_181, n_177);
  nor g122 (n_185, n_182, n_183);
  nor g125 (n_271, n_187, n_183);
  nor g126 (n_191, n_188, n_189);
  nor g129 (n_273, n_193, n_189);
  nor g130 (n_197, n_194, n_195);
  nor g133 (n_281, n_199, n_195);
  nor g134 (n_203, n_200, n_201);
  nor g137 (n_283, n_205, n_201);
  nand g144 (n_464, n_116, n_214);
  nand g145 (n_217, n_215, n_212);
  nand g146 (n_288, n_216, n_217);
  nor g147 (n_219, n_133, n_218);
  nand g156 (n_296, n_221, n_223);
  nor g157 (n_229, n_145, n_228);
  nand g166 (n_303, n_231, n_233);
  nor g167 (n_239, n_157, n_238);
  nand g176 (n_311, n_241, n_243);
  nor g177 (n_249, n_169, n_248);
  nand g186 (n_318, n_251, n_253);
  nor g187 (n_259, n_181, n_258);
  nand g196 (n_326, n_261, n_263);
  nor g197 (n_269, n_193, n_268);
  nand g206 (n_333, n_271, n_273);
  nor g207 (n_279, n_205, n_278);
  nand g216 (n_341, n_281, n_283);
  nand g219 (n_468, n_122, n_290);
  nand g220 (n_291, n_221, n_288);
  nand g221 (n_470, n_218, n_291);
  nand g224 (n_473, n_294, n_295);
  nand g227 (n_345, n_298, n_299);
  nor g228 (n_301, n_151, n_300);
  nor g231 (n_355, n_151, n_303);
  nor g237 (n_309, n_307, n_300);
  nor g240 (n_361, n_303, n_307);
  nor g241 (n_313, n_311, n_300);
  nor g244 (n_364, n_303, n_311);
  nor g245 (n_316, n_175, n_315);
  nor g248 (n_413, n_175, n_318);
  nor g254 (n_324, n_322, n_315);
  nor g257 (n_419, n_318, n_322);
  nor g258 (n_328, n_326, n_315);
  nor g261 (n_370, n_318, n_326);
  nor g262 (n_331, n_199, n_330);
  nor g265 (n_383, n_199, n_333);
  nor g271 (n_339, n_337, n_330);
  nor g274 (n_393, n_333, n_337);
  nor g275 (n_343, n_341, n_330);
  nor g278 (n_398, n_333, n_341);
  nand g281 (n_477, n_134, n_347);
  nand g282 (n_348, n_231, n_345);
  nand g283 (n_479, n_228, n_348);
  nand g286 (n_482, n_351, n_352);
  nand g289 (n_485, n_300, n_354);
  nand g290 (n_357, n_355, n_345);
  nand g291 (n_488, n_356, n_357);
  nand g292 (n_360, n_358, n_345);
  nand g293 (n_490, n_359, n_360);
  nand g294 (n_363, n_361, n_345);
  nand g295 (n_493, n_362, n_363);
  nand g296 (n_366, n_364, n_345);
  nand g297 (n_403, n_365, n_366);
  nor g298 (n_368, n_187, n_367);
  nand g307 (n_427, n_271, n_370);
  nor g308 (n_377, n_375, n_367);
  nor g313 (n_380, n_333, n_367);
  nand g322 (n_439, n_370, n_383);
  nand g327 (n_443, n_370, n_388);
  nand g332 (n_447, n_370, n_393);
  nand g337 (n_451, n_370, n_398);
  nand g340 (n_497, n_158, n_405);
  nand g341 (n_406, n_251, n_403);
  nand g342 (n_499, n_248, n_406);
  nand g345 (n_502, n_409, n_410);
  nand g348 (n_505, n_315, n_412);
  nand g349 (n_415, n_413, n_403);
  nand g350 (n_508, n_414, n_415);
  nand g351 (n_418, n_416, n_403);
  nand g352 (n_510, n_417, n_418);
  nand g353 (n_421, n_419, n_403);
  nand g354 (n_513, n_420, n_421);
  nand g355 (n_422, n_370, n_403);
  nand g356 (n_515, n_367, n_422);
  nand g359 (n_518, n_425, n_426);
  nand g362 (n_520, n_429, n_430);
  nand g365 (n_523, n_433, n_434);
  nand g368 (n_526, n_437, n_438);
  nand g371 (n_529, n_441, n_442);
  nand g374 (n_531, n_445, n_446);
  nand g377 (n_534, n_449, n_450);
  nand g380 (n_455, n_453, n_454);
  nand g383 (n_538, n_206, n_457);
  xnor g389 (Z[2], n_212, n_462);
  xnor g392 (Z[3], n_464, n_465);
  xnor g394 (Z[4], n_288, n_466);
  xnor g397 (Z[5], n_468, n_469);
  xnor g399 (Z[6], n_470, n_471);
  xnor g402 (Z[7], n_473, n_474);
  xnor g404 (Z[8], n_345, n_475);
  xnor g407 (Z[9], n_477, n_478);
  xnor g409 (Z[10], n_479, n_480);
  xnor g412 (Z[11], n_482, n_483);
  xnor g415 (Z[12], n_485, n_486);
  xnor g418 (Z[13], n_488, n_489);
  xnor g420 (Z[14], n_490, n_491);
  xnor g423 (Z[15], n_493, n_494);
  xnor g425 (Z[16], n_403, n_495);
  xnor g428 (Z[17], n_497, n_498);
  xnor g430 (Z[18], n_499, n_500);
  xnor g433 (Z[19], n_502, n_503);
  xnor g436 (Z[20], n_505, n_506);
  xnor g439 (Z[21], n_508, n_509);
  xnor g441 (Z[22], n_510, n_511);
  xnor g444 (Z[23], n_513, n_514);
  xnor g446 (Z[24], n_515, n_516);
  xnor g449 (Z[25], n_518, n_519);
  xnor g451 (Z[26], n_520, n_521);
  xnor g454 (Z[27], n_523, n_524);
  xnor g457 (Z[28], n_526, n_527);
  xnor g460 (Z[29], n_529, n_530);
  xnor g462 (Z[30], n_531, n_532);
  xnor g465 (Z[31], n_534, n_535);
  xnor g467 (Z[32], n_455, n_536);
  xnor g470 (Z[33], n_538, n_539);
  and g473 (n_207, A[33], B[33]);
  or g474 (n_208, A[33], B[33]);
  or g475 (n_115, n_109, n_111);
  and g476 (n_216, wc, n_118);
  not gc (wc, n_119);
  and g477 (n_218, wc0, n_124);
  not gc0 (wc0, n_125);
  and g478 (n_225, wc1, n_130);
  not gc1 (wc1, n_131);
  and g479 (n_228, wc2, n_136);
  not gc2 (wc2, n_137);
  and g480 (n_235, wc3, n_142);
  not gc3 (wc3, n_143);
  and g481 (n_238, wc4, n_148);
  not gc4 (wc4, n_149);
  and g482 (n_245, wc5, n_154);
  not gc5 (wc5, n_155);
  and g483 (n_248, wc6, n_160);
  not gc6 (wc6, n_161);
  and g484 (n_255, wc7, n_166);
  not gc7 (wc7, n_167);
  and g485 (n_258, wc8, n_172);
  not gc8 (wc8, n_173);
  and g486 (n_265, wc9, n_178);
  not gc9 (wc9, n_179);
  and g487 (n_268, wc10, n_184);
  not gc10 (wc10, n_185);
  and g488 (n_275, wc11, n_190);
  not gc11 (wc11, n_191);
  and g489 (n_278, wc12, n_196);
  not gc12 (wc12, n_197);
  and g490 (n_285, wc13, n_202);
  not gc13 (wc13, n_203);
  or g491 (n_292, wc14, n_133);
  not gc14 (wc14, n_221);
  or g492 (n_349, wc15, n_145);
  not gc15 (wc15, n_231);
  or g493 (n_307, wc16, n_157);
  not gc16 (wc16, n_241);
  or g494 (n_407, wc17, n_169);
  not gc17 (wc17, n_251);
  or g495 (n_322, wc18, n_181);
  not gc18 (wc18, n_261);
  or g496 (n_375, wc19, n_193);
  not gc19 (wc19, n_271);
  or g497 (n_337, wc20, n_205);
  not gc20 (wc20, n_281);
  or g498 (n_461, wc21, n_111);
  not gc21 (wc21, n_114);
  or g499 (n_462, wc22, n_121);
  not gc22 (wc22, n_116);
  or g500 (n_465, wc23, n_117);
  not gc23 (wc23, n_118);
  or g501 (n_466, wc24, n_127);
  not gc24 (wc24, n_122);
  or g502 (n_469, wc25, n_123);
  not gc25 (wc25, n_124);
  or g503 (n_471, wc26, n_133);
  not gc26 (wc26, n_128);
  or g504 (n_474, wc27, n_129);
  not gc27 (wc27, n_130);
  or g505 (n_475, wc28, n_139);
  not gc28 (wc28, n_134);
  or g506 (n_478, wc29, n_135);
  not gc29 (wc29, n_136);
  or g507 (n_480, wc30, n_145);
  not gc30 (wc30, n_140);
  or g508 (n_483, wc31, n_141);
  not gc31 (wc31, n_142);
  or g509 (n_486, wc32, n_151);
  not gc32 (wc32, n_146);
  or g510 (n_489, wc33, n_147);
  not gc33 (wc33, n_148);
  or g511 (n_491, wc34, n_157);
  not gc34 (wc34, n_152);
  or g512 (n_494, wc35, n_153);
  not gc35 (wc35, n_154);
  or g513 (n_495, wc36, n_163);
  not gc36 (wc36, n_158);
  or g514 (n_498, wc37, n_159);
  not gc37 (wc37, n_160);
  or g515 (n_500, wc38, n_169);
  not gc38 (wc38, n_164);
  or g516 (n_503, wc39, n_165);
  not gc39 (wc39, n_166);
  or g517 (n_506, wc40, n_175);
  not gc40 (wc40, n_170);
  or g518 (n_509, wc41, n_171);
  not gc41 (wc41, n_172);
  or g519 (n_511, wc42, n_181);
  not gc42 (wc42, n_176);
  or g520 (n_514, wc43, n_177);
  not gc43 (wc43, n_178);
  or g521 (n_516, wc44, n_187);
  not gc44 (wc44, n_182);
  or g522 (n_519, wc45, n_183);
  not gc45 (wc45, n_184);
  or g523 (n_521, wc46, n_193);
  not gc46 (wc46, n_188);
  or g524 (n_524, wc47, n_189);
  not gc47 (wc47, n_190);
  or g525 (n_527, wc48, n_199);
  not gc48 (wc48, n_194);
  or g526 (n_530, wc49, n_195);
  not gc49 (wc49, n_196);
  or g527 (n_532, wc50, n_205);
  not gc50 (wc50, n_200);
  or g528 (n_535, wc51, n_201);
  not gc51 (wc51, n_202);
  or g529 (n_536, wc52, n_211);
  not gc52 (wc52, n_206);
  and g530 (n_226, wc53, n_223);
  not gc53 (wc53, n_218);
  and g531 (n_236, wc54, n_233);
  not gc54 (wc54, n_228);
  and g532 (n_246, wc55, n_243);
  not gc55 (wc55, n_238);
  and g533 (n_256, wc56, n_253);
  not gc56 (wc56, n_248);
  and g534 (n_266, wc57, n_263);
  not gc57 (wc57, n_258);
  and g535 (n_276, wc58, n_273);
  not gc58 (wc58, n_268);
  and g536 (n_286, wc59, n_283);
  not gc59 (wc59, n_278);
  and g537 (n_358, wc60, n_241);
  not gc60 (wc60, n_303);
  and g538 (n_416, wc61, n_261);
  not gc61 (wc61, n_318);
  and g539 (n_388, wc62, n_281);
  not gc62 (wc62, n_333);
  xor g540 (Z[1], n_109, n_461);
  or g541 (n_539, wc63, n_207);
  not gc63 (wc63, n_208);
  or g542 (n_214, wc64, n_121);
  not gc64 (wc64, n_212);
  and g543 (n_294, wc65, n_128);
  not gc65 (wc65, n_219);
  and g544 (n_298, wc66, n_225);
  not gc66 (wc66, n_226);
  and g545 (n_351, wc67, n_140);
  not gc67 (wc67, n_229);
  and g546 (n_300, wc68, n_235);
  not gc68 (wc68, n_236);
  and g547 (n_308, wc69, n_152);
  not gc69 (wc69, n_239);
  and g548 (n_312, wc70, n_245);
  not gc70 (wc70, n_246);
  and g549 (n_409, wc71, n_164);
  not gc71 (wc71, n_249);
  and g550 (n_315, wc72, n_255);
  not gc72 (wc72, n_256);
  and g551 (n_323, wc73, n_176);
  not gc73 (wc73, n_259);
  and g552 (n_327, wc74, n_265);
  not gc74 (wc74, n_266);
  and g553 (n_376, wc75, n_188);
  not gc75 (wc75, n_269);
  and g554 (n_330, wc76, n_275);
  not gc76 (wc76, n_276);
  and g555 (n_338, wc77, n_200);
  not gc77 (wc77, n_279);
  and g556 (n_342, wc78, n_285);
  not gc78 (wc78, n_286);
  or g557 (n_423, wc79, n_187);
  not gc79 (wc79, n_370);
  or g558 (n_431, n_375, wc80);
  not gc80 (wc80, n_370);
  or g559 (n_435, wc81, n_333);
  not gc81 (wc81, n_370);
  and g560 (n_305, wc82, n_241);
  not gc82 (wc82, n_300);
  and g561 (n_320, wc83, n_261);
  not gc83 (wc83, n_315);
  and g562 (n_335, wc84, n_281);
  not gc84 (wc84, n_330);
  or g563 (n_290, wc85, n_127);
  not gc85 (wc85, n_288);
  or g564 (n_295, n_292, wc86);
  not gc86 (wc86, n_288);
  or g565 (n_299, n_296, wc87);
  not gc87 (wc87, n_288);
  and g566 (n_356, wc88, n_146);
  not gc88 (wc88, n_301);
  and g567 (n_359, wc89, n_238);
  not gc89 (wc89, n_305);
  and g568 (n_362, n_308, wc90);
  not gc90 (wc90, n_309);
  and g569 (n_365, n_312, wc91);
  not gc91 (wc91, n_313);
  and g570 (n_414, wc92, n_170);
  not gc92 (wc92, n_316);
  and g571 (n_417, wc93, n_258);
  not gc93 (wc93, n_320);
  and g572 (n_420, n_323, wc94);
  not gc94 (wc94, n_324);
  and g573 (n_367, n_327, wc95);
  not gc95 (wc95, n_328);
  and g574 (n_385, wc96, n_194);
  not gc96 (wc96, n_331);
  and g575 (n_390, wc97, n_278);
  not gc97 (wc97, n_335);
  and g576 (n_395, n_338, wc98);
  not gc98 (wc98, n_339);
  and g577 (n_400, n_342, wc99);
  not gc99 (wc99, n_343);
  and g578 (n_373, wc100, n_271);
  not gc100 (wc100, n_367);
  and g579 (n_386, wc101, n_383);
  not gc101 (wc101, n_367);
  and g580 (n_391, wc102, n_388);
  not gc102 (wc102, n_367);
  and g581 (n_396, wc103, n_393);
  not gc103 (wc103, n_367);
  and g582 (n_401, wc104, n_398);
  not gc104 (wc104, n_367);
  or g583 (n_347, wc105, n_139);
  not gc105 (wc105, n_345);
  or g584 (n_352, n_349, wc106);
  not gc106 (wc106, n_345);
  or g585 (n_354, wc107, n_303);
  not gc107 (wc107, n_345);
  and g586 (n_425, wc108, n_182);
  not gc108 (wc108, n_368);
  and g587 (n_429, wc109, n_268);
  not gc109 (wc109, n_373);
  and g588 (n_433, n_376, wc110);
  not gc110 (wc110, n_377);
  and g589 (n_437, n_330, wc111);
  not gc111 (wc111, n_380);
  and g590 (n_441, wc112, n_385);
  not gc112 (wc112, n_386);
  and g591 (n_445, wc113, n_390);
  not gc113 (wc113, n_391);
  and g592 (n_449, wc114, n_395);
  not gc114 (wc114, n_396);
  and g593 (n_453, wc115, n_400);
  not gc115 (wc115, n_401);
  or g594 (n_405, wc116, n_163);
  not gc116 (wc116, n_403);
  or g595 (n_410, n_407, wc117);
  not gc117 (wc117, n_403);
  or g596 (n_412, wc118, n_318);
  not gc118 (wc118, n_403);
  or g597 (n_426, n_423, wc119);
  not gc119 (wc119, n_403);
  or g598 (n_430, n_427, wc120);
  not gc120 (wc120, n_403);
  or g599 (n_434, n_431, wc121);
  not gc121 (wc121, n_403);
  or g600 (n_438, n_435, wc122);
  not gc122 (wc122, n_403);
  or g601 (n_442, n_439, wc123);
  not gc123 (wc123, n_403);
  or g602 (n_446, n_443, wc124);
  not gc124 (wc124, n_403);
  or g603 (n_450, n_447, wc125);
  not gc125 (wc125, n_403);
  or g604 (n_454, n_451, wc126);
  not gc126 (wc126, n_403);
  or g605 (n_457, wc127, n_211);
  not gc127 (wc127, n_455);
endmodule

module add_signed_9277_GENERIC(A, B, Z);
  input [35:0] A, B;
  output [33:0] Z;
  wire [35:0] A, B;
  wire [33:0] Z;
  add_signed_9277_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module bmux_9159_GENERIC_REAL(ctl, in_0, in_1, z);
// synthesis_equation "reg [24:0] temp;always @(*) case(ctl) 1'b0: temp = in_0;1'b1: temp = in_1;endcase assign z = temp;"
  input ctl;
  input [24:0] in_0, in_1;
  output [24:0] z;
  wire ctl;
  wire [24:0] in_0, in_1;
  wire [24:0] z;
  or g26 (z[24], wc, wc1);
  and gc1 (wc1, in_1[24], ctl);
  and gc0 (wc, in_0[24], wc0);
  not gc (wc0, ctl);
  or g27 (z[23], wc2, wc4);
  and gc4 (wc4, in_1[23], ctl);
  and gc3 (wc2, in_0[23], wc3);
  not gc2 (wc3, ctl);
  or g28 (z[22], wc5, wc7);
  and gc7 (wc7, in_1[22], ctl);
  and gc6 (wc5, in_0[22], wc6);
  not gc5 (wc6, ctl);
  or g29 (z[21], wc8, wc10);
  and gc10 (wc10, in_1[21], ctl);
  and gc9 (wc8, in_0[21], wc9);
  not gc8 (wc9, ctl);
  or g30 (z[20], wc11, wc13);
  and gc13 (wc13, in_1[20], ctl);
  and gc12 (wc11, in_0[20], wc12);
  not gc11 (wc12, ctl);
  or g31 (z[19], wc14, wc16);
  and gc16 (wc16, in_1[19], ctl);
  and gc15 (wc14, in_0[19], wc15);
  not gc14 (wc15, ctl);
  or g32 (z[18], wc17, wc19);
  and gc19 (wc19, in_1[18], ctl);
  and gc18 (wc17, in_0[18], wc18);
  not gc17 (wc18, ctl);
  or g33 (z[17], wc20, wc22);
  and gc22 (wc22, in_1[17], ctl);
  and gc21 (wc20, in_0[17], wc21);
  not gc20 (wc21, ctl);
  or g34 (z[16], wc23, wc25);
  and gc25 (wc25, in_1[16], ctl);
  and gc24 (wc23, in_0[16], wc24);
  not gc23 (wc24, ctl);
  or g35 (z[15], wc26, wc28);
  and gc28 (wc28, in_1[15], ctl);
  and gc27 (wc26, in_0[15], wc27);
  not gc26 (wc27, ctl);
  or g36 (z[14], wc29, wc31);
  and gc31 (wc31, in_1[14], ctl);
  and gc30 (wc29, in_0[14], wc30);
  not gc29 (wc30, ctl);
  or g37 (z[13], wc32, wc34);
  and gc34 (wc34, in_1[13], ctl);
  and gc33 (wc32, in_0[13], wc33);
  not gc32 (wc33, ctl);
  or g38 (z[12], wc35, wc37);
  and gc37 (wc37, in_1[12], ctl);
  and gc36 (wc35, in_0[12], wc36);
  not gc35 (wc36, ctl);
  or g39 (z[11], wc38, wc40);
  and gc40 (wc40, in_1[11], ctl);
  and gc39 (wc38, in_0[11], wc39);
  not gc38 (wc39, ctl);
  or g40 (z[10], wc41, wc43);
  and gc43 (wc43, in_1[10], ctl);
  and gc42 (wc41, in_0[10], wc42);
  not gc41 (wc42, ctl);
  or g41 (z[9], wc44, wc46);
  and gc46 (wc46, in_1[9], ctl);
  and gc45 (wc44, in_0[9], wc45);
  not gc44 (wc45, ctl);
  or g42 (z[8], wc47, wc49);
  and gc49 (wc49, in_1[8], ctl);
  and gc48 (wc47, in_0[8], wc48);
  not gc47 (wc48, ctl);
  or g43 (z[7], wc50, wc52);
  and gc52 (wc52, in_1[7], ctl);
  and gc51 (wc50, in_0[7], wc51);
  not gc50 (wc51, ctl);
  or g44 (z[6], wc53, wc55);
  and gc55 (wc55, in_1[6], ctl);
  and gc54 (wc53, in_0[6], wc54);
  not gc53 (wc54, ctl);
  or g45 (z[5], wc56, wc58);
  and gc58 (wc58, in_1[5], ctl);
  and gc57 (wc56, in_0[5], wc57);
  not gc56 (wc57, ctl);
  or g46 (z[4], wc59, wc61);
  and gc61 (wc61, in_1[4], ctl);
  and gc60 (wc59, in_0[4], wc60);
  not gc59 (wc60, ctl);
  or g47 (z[3], wc62, wc64);
  and gc64 (wc64, in_1[3], ctl);
  and gc63 (wc62, in_0[3], wc63);
  not gc62 (wc63, ctl);
  or g48 (z[2], wc65, wc67);
  and gc67 (wc67, in_1[2], ctl);
  and gc66 (wc65, in_0[2], wc66);
  not gc65 (wc66, ctl);
  or g49 (z[1], wc68, wc70);
  and gc70 (wc70, in_1[1], ctl);
  and gc69 (wc68, in_0[1], wc69);
  not gc68 (wc69, ctl);
  or g50 (z[0], wc71, wc73);
  and gc73 (wc73, in_1[0], ctl);
  and gc72 (wc71, in_0[0], wc72);
  not gc71 (wc72, ctl);
endmodule

module bmux_9159_GENERIC(ctl, in_0, in_1, z);
  input ctl;
  input [24:0] in_0, in_1;
  output [24:0] z;
  wire ctl;
  wire [24:0] in_0, in_1;
  wire [24:0] z;
  bmux_9159_GENERIC_REAL g1(.ctl (ctl), .in_0 (in_0), .in_1 (in_1), .z
       (z));
endmodule

module bmux_9159_1_GENERIC_REAL(ctl, in_0, in_1, z);
// synthesis_equation "reg [24:0] temp;always @(*) case(ctl) 1'b0: temp = in_0;1'b1: temp = in_1;endcase assign z = temp;"
  input ctl;
  input [24:0] in_0, in_1;
  output [24:0] z;
  wire ctl;
  wire [24:0] in_0, in_1;
  wire [24:0] z;
  or g26 (z[24], wc, wc1);
  and gc1 (wc1, in_1[24], ctl);
  and gc0 (wc, in_0[24], wc0);
  not gc (wc0, ctl);
  or g27 (z[23], wc2, wc4);
  and gc4 (wc4, in_1[23], ctl);
  and gc3 (wc2, in_0[23], wc3);
  not gc2 (wc3, ctl);
  or g28 (z[22], wc5, wc7);
  and gc7 (wc7, in_1[22], ctl);
  and gc6 (wc5, in_0[22], wc6);
  not gc5 (wc6, ctl);
  or g29 (z[21], wc8, wc10);
  and gc10 (wc10, in_1[21], ctl);
  and gc9 (wc8, in_0[21], wc9);
  not gc8 (wc9, ctl);
  or g30 (z[20], wc11, wc13);
  and gc13 (wc13, in_1[20], ctl);
  and gc12 (wc11, in_0[20], wc12);
  not gc11 (wc12, ctl);
  or g31 (z[19], wc14, wc16);
  and gc16 (wc16, in_1[19], ctl);
  and gc15 (wc14, in_0[19], wc15);
  not gc14 (wc15, ctl);
  or g32 (z[18], wc17, wc19);
  and gc19 (wc19, in_1[18], ctl);
  and gc18 (wc17, in_0[18], wc18);
  not gc17 (wc18, ctl);
  or g33 (z[17], wc20, wc22);
  and gc22 (wc22, in_1[17], ctl);
  and gc21 (wc20, in_0[17], wc21);
  not gc20 (wc21, ctl);
  or g34 (z[16], wc23, wc25);
  and gc25 (wc25, in_1[16], ctl);
  and gc24 (wc23, in_0[16], wc24);
  not gc23 (wc24, ctl);
  or g35 (z[15], wc26, wc28);
  and gc28 (wc28, in_1[15], ctl);
  and gc27 (wc26, in_0[15], wc27);
  not gc26 (wc27, ctl);
  or g36 (z[14], wc29, wc31);
  and gc31 (wc31, in_1[14], ctl);
  and gc30 (wc29, in_0[14], wc30);
  not gc29 (wc30, ctl);
  or g37 (z[13], wc32, wc34);
  and gc34 (wc34, in_1[13], ctl);
  and gc33 (wc32, in_0[13], wc33);
  not gc32 (wc33, ctl);
  or g38 (z[12], wc35, wc37);
  and gc37 (wc37, in_1[12], ctl);
  and gc36 (wc35, in_0[12], wc36);
  not gc35 (wc36, ctl);
  or g39 (z[11], wc38, wc40);
  and gc40 (wc40, in_1[11], ctl);
  and gc39 (wc38, in_0[11], wc39);
  not gc38 (wc39, ctl);
  or g40 (z[10], wc41, wc43);
  and gc43 (wc43, in_1[10], ctl);
  and gc42 (wc41, in_0[10], wc42);
  not gc41 (wc42, ctl);
  or g41 (z[9], wc44, wc46);
  and gc46 (wc46, in_1[9], ctl);
  and gc45 (wc44, in_0[9], wc45);
  not gc44 (wc45, ctl);
  or g42 (z[8], wc47, wc49);
  and gc49 (wc49, in_1[8], ctl);
  and gc48 (wc47, in_0[8], wc48);
  not gc47 (wc48, ctl);
  or g43 (z[7], wc50, wc52);
  and gc52 (wc52, in_1[7], ctl);
  and gc51 (wc50, in_0[7], wc51);
  not gc50 (wc51, ctl);
  or g44 (z[6], wc53, wc55);
  and gc55 (wc55, in_1[6], ctl);
  and gc54 (wc53, in_0[6], wc54);
  not gc53 (wc54, ctl);
  or g45 (z[5], wc56, wc58);
  and gc58 (wc58, in_1[5], ctl);
  and gc57 (wc56, in_0[5], wc57);
  not gc56 (wc57, ctl);
  or g46 (z[4], wc59, wc61);
  and gc61 (wc61, in_1[4], ctl);
  and gc60 (wc59, in_0[4], wc60);
  not gc59 (wc60, ctl);
  or g47 (z[3], wc62, wc64);
  and gc64 (wc64, in_1[3], ctl);
  and gc63 (wc62, in_0[3], wc63);
  not gc62 (wc63, ctl);
  or g48 (z[2], wc65, wc67);
  and gc67 (wc67, in_1[2], ctl);
  and gc66 (wc65, in_0[2], wc66);
  not gc65 (wc66, ctl);
  or g49 (z[1], wc68, wc70);
  and gc70 (wc70, in_1[1], ctl);
  and gc69 (wc68, in_0[1], wc69);
  not gc68 (wc69, ctl);
  or g50 (z[0], wc71, wc73);
  and gc73 (wc73, in_1[0], ctl);
  and gc72 (wc71, in_0[0], wc72);
  not gc71 (wc72, ctl);
endmodule

module bmux_9159_1_GENERIC(ctl, in_0, in_1, z);
  input ctl;
  input [24:0] in_0, in_1;
  output [24:0] z;
  wire ctl;
  wire [24:0] in_0, in_1;
  wire [24:0] z;
  bmux_9159_1_GENERIC_REAL g1(.ctl (ctl), .in_0 (in_0), .in_1 (in_1),
       .z (z));
endmodule

module bmux_9159_2_GENERIC_REAL(ctl, in_0, in_1, z);
// synthesis_equation "reg [24:0] temp;always @(*) case(ctl) 1'b0: temp = in_0;1'b1: temp = in_1;endcase assign z = temp;"
  input ctl;
  input [24:0] in_0, in_1;
  output [24:0] z;
  wire ctl;
  wire [24:0] in_0, in_1;
  wire [24:0] z;
  or g26 (z[24], wc, wc1);
  and gc1 (wc1, in_1[24], ctl);
  and gc0 (wc, in_0[24], wc0);
  not gc (wc0, ctl);
  or g27 (z[23], wc2, wc4);
  and gc4 (wc4, in_1[23], ctl);
  and gc3 (wc2, in_0[23], wc3);
  not gc2 (wc3, ctl);
  or g28 (z[22], wc5, wc7);
  and gc7 (wc7, in_1[22], ctl);
  and gc6 (wc5, in_0[22], wc6);
  not gc5 (wc6, ctl);
  or g29 (z[21], wc8, wc10);
  and gc10 (wc10, in_1[21], ctl);
  and gc9 (wc8, in_0[21], wc9);
  not gc8 (wc9, ctl);
  or g30 (z[20], wc11, wc13);
  and gc13 (wc13, in_1[20], ctl);
  and gc12 (wc11, in_0[20], wc12);
  not gc11 (wc12, ctl);
  or g31 (z[19], wc14, wc16);
  and gc16 (wc16, in_1[19], ctl);
  and gc15 (wc14, in_0[19], wc15);
  not gc14 (wc15, ctl);
  or g32 (z[18], wc17, wc19);
  and gc19 (wc19, in_1[18], ctl);
  and gc18 (wc17, in_0[18], wc18);
  not gc17 (wc18, ctl);
  or g33 (z[17], wc20, wc22);
  and gc22 (wc22, in_1[17], ctl);
  and gc21 (wc20, in_0[17], wc21);
  not gc20 (wc21, ctl);
  or g34 (z[16], wc23, wc25);
  and gc25 (wc25, in_1[16], ctl);
  and gc24 (wc23, in_0[16], wc24);
  not gc23 (wc24, ctl);
  or g35 (z[15], wc26, wc28);
  and gc28 (wc28, in_1[15], ctl);
  and gc27 (wc26, in_0[15], wc27);
  not gc26 (wc27, ctl);
  or g36 (z[14], wc29, wc31);
  and gc31 (wc31, in_1[14], ctl);
  and gc30 (wc29, in_0[14], wc30);
  not gc29 (wc30, ctl);
  or g37 (z[13], wc32, wc34);
  and gc34 (wc34, in_1[13], ctl);
  and gc33 (wc32, in_0[13], wc33);
  not gc32 (wc33, ctl);
  or g38 (z[12], wc35, wc37);
  and gc37 (wc37, in_1[12], ctl);
  and gc36 (wc35, in_0[12], wc36);
  not gc35 (wc36, ctl);
  or g39 (z[11], wc38, wc40);
  and gc40 (wc40, in_1[11], ctl);
  and gc39 (wc38, in_0[11], wc39);
  not gc38 (wc39, ctl);
  or g40 (z[10], wc41, wc43);
  and gc43 (wc43, in_1[10], ctl);
  and gc42 (wc41, in_0[10], wc42);
  not gc41 (wc42, ctl);
  or g41 (z[9], wc44, wc46);
  and gc46 (wc46, in_1[9], ctl);
  and gc45 (wc44, in_0[9], wc45);
  not gc44 (wc45, ctl);
  or g42 (z[8], wc47, wc49);
  and gc49 (wc49, in_1[8], ctl);
  and gc48 (wc47, in_0[8], wc48);
  not gc47 (wc48, ctl);
  or g43 (z[7], wc50, wc52);
  and gc52 (wc52, in_1[7], ctl);
  and gc51 (wc50, in_0[7], wc51);
  not gc50 (wc51, ctl);
  or g44 (z[6], wc53, wc55);
  and gc55 (wc55, in_1[6], ctl);
  and gc54 (wc53, in_0[6], wc54);
  not gc53 (wc54, ctl);
  or g45 (z[5], wc56, wc58);
  and gc58 (wc58, in_1[5], ctl);
  and gc57 (wc56, in_0[5], wc57);
  not gc56 (wc57, ctl);
  or g46 (z[4], wc59, wc61);
  and gc61 (wc61, in_1[4], ctl);
  and gc60 (wc59, in_0[4], wc60);
  not gc59 (wc60, ctl);
  or g47 (z[3], wc62, wc64);
  and gc64 (wc64, in_1[3], ctl);
  and gc63 (wc62, in_0[3], wc63);
  not gc62 (wc63, ctl);
  or g48 (z[2], wc65, wc67);
  and gc67 (wc67, in_1[2], ctl);
  and gc66 (wc65, in_0[2], wc66);
  not gc65 (wc66, ctl);
  or g49 (z[1], wc68, wc70);
  and gc70 (wc70, in_1[1], ctl);
  and gc69 (wc68, in_0[1], wc69);
  not gc68 (wc69, ctl);
  or g50 (z[0], wc71, wc73);
  and gc73 (wc73, in_1[0], ctl);
  and gc72 (wc71, in_0[0], wc72);
  not gc71 (wc72, ctl);
endmodule

module bmux_9159_2_GENERIC(ctl, in_0, in_1, z);
  input ctl;
  input [24:0] in_0, in_1;
  output [24:0] z;
  wire ctl;
  wire [24:0] in_0, in_1;
  wire [24:0] z;
  bmux_9159_2_GENERIC_REAL g1(.ctl (ctl), .in_0 (in_0), .in_1 (in_1),
       .z (z));
endmodule

module bmux_9159_3_GENERIC_REAL(ctl, in_0, in_1, z);
// synthesis_equation "reg [24:0] temp;always @(*) case(ctl) 1'b0: temp = in_0;1'b1: temp = in_1;endcase assign z = temp;"
  input ctl;
  input [24:0] in_0, in_1;
  output [24:0] z;
  wire ctl;
  wire [24:0] in_0, in_1;
  wire [24:0] z;
  or g26 (z[24], wc, wc1);
  and gc1 (wc1, in_1[24], ctl);
  and gc0 (wc, in_0[24], wc0);
  not gc (wc0, ctl);
  or g27 (z[23], wc2, wc4);
  and gc4 (wc4, in_1[23], ctl);
  and gc3 (wc2, in_0[23], wc3);
  not gc2 (wc3, ctl);
  or g28 (z[22], wc5, wc7);
  and gc7 (wc7, in_1[22], ctl);
  and gc6 (wc5, in_0[22], wc6);
  not gc5 (wc6, ctl);
  or g29 (z[21], wc8, wc10);
  and gc10 (wc10, in_1[21], ctl);
  and gc9 (wc8, in_0[21], wc9);
  not gc8 (wc9, ctl);
  or g30 (z[20], wc11, wc13);
  and gc13 (wc13, in_1[20], ctl);
  and gc12 (wc11, in_0[20], wc12);
  not gc11 (wc12, ctl);
  or g31 (z[19], wc14, wc16);
  and gc16 (wc16, in_1[19], ctl);
  and gc15 (wc14, in_0[19], wc15);
  not gc14 (wc15, ctl);
  or g32 (z[18], wc17, wc19);
  and gc19 (wc19, in_1[18], ctl);
  and gc18 (wc17, in_0[18], wc18);
  not gc17 (wc18, ctl);
  or g33 (z[17], wc20, wc22);
  and gc22 (wc22, in_1[17], ctl);
  and gc21 (wc20, in_0[17], wc21);
  not gc20 (wc21, ctl);
  or g34 (z[16], wc23, wc25);
  and gc25 (wc25, in_1[16], ctl);
  and gc24 (wc23, in_0[16], wc24);
  not gc23 (wc24, ctl);
  or g35 (z[15], wc26, wc28);
  and gc28 (wc28, in_1[15], ctl);
  and gc27 (wc26, in_0[15], wc27);
  not gc26 (wc27, ctl);
  or g36 (z[14], wc29, wc31);
  and gc31 (wc31, in_1[14], ctl);
  and gc30 (wc29, in_0[14], wc30);
  not gc29 (wc30, ctl);
  or g37 (z[13], wc32, wc34);
  and gc34 (wc34, in_1[13], ctl);
  and gc33 (wc32, in_0[13], wc33);
  not gc32 (wc33, ctl);
  or g38 (z[12], wc35, wc37);
  and gc37 (wc37, in_1[12], ctl);
  and gc36 (wc35, in_0[12], wc36);
  not gc35 (wc36, ctl);
  or g39 (z[11], wc38, wc40);
  and gc40 (wc40, in_1[11], ctl);
  and gc39 (wc38, in_0[11], wc39);
  not gc38 (wc39, ctl);
  or g40 (z[10], wc41, wc43);
  and gc43 (wc43, in_1[10], ctl);
  and gc42 (wc41, in_0[10], wc42);
  not gc41 (wc42, ctl);
  or g41 (z[9], wc44, wc46);
  and gc46 (wc46, in_1[9], ctl);
  and gc45 (wc44, in_0[9], wc45);
  not gc44 (wc45, ctl);
  or g42 (z[8], wc47, wc49);
  and gc49 (wc49, in_1[8], ctl);
  and gc48 (wc47, in_0[8], wc48);
  not gc47 (wc48, ctl);
  or g43 (z[7], wc50, wc52);
  and gc52 (wc52, in_1[7], ctl);
  and gc51 (wc50, in_0[7], wc51);
  not gc50 (wc51, ctl);
  or g44 (z[6], wc53, wc55);
  and gc55 (wc55, in_1[6], ctl);
  and gc54 (wc53, in_0[6], wc54);
  not gc53 (wc54, ctl);
  or g45 (z[5], wc56, wc58);
  and gc58 (wc58, in_1[5], ctl);
  and gc57 (wc56, in_0[5], wc57);
  not gc56 (wc57, ctl);
  or g46 (z[4], wc59, wc61);
  and gc61 (wc61, in_1[4], ctl);
  and gc60 (wc59, in_0[4], wc60);
  not gc59 (wc60, ctl);
  or g47 (z[3], wc62, wc64);
  and gc64 (wc64, in_1[3], ctl);
  and gc63 (wc62, in_0[3], wc63);
  not gc62 (wc63, ctl);
  or g48 (z[2], wc65, wc67);
  and gc67 (wc67, in_1[2], ctl);
  and gc66 (wc65, in_0[2], wc66);
  not gc65 (wc66, ctl);
  or g49 (z[1], wc68, wc70);
  and gc70 (wc70, in_1[1], ctl);
  and gc69 (wc68, in_0[1], wc69);
  not gc68 (wc69, ctl);
  or g50 (z[0], wc71, wc73);
  and gc73 (wc73, in_1[0], ctl);
  and gc72 (wc71, in_0[0], wc72);
  not gc71 (wc72, ctl);
endmodule

module bmux_9159_3_GENERIC(ctl, in_0, in_1, z);
  input ctl;
  input [24:0] in_0, in_1;
  output [24:0] z;
  wire ctl;
  wire [24:0] in_0, in_1;
  wire [24:0] z;
  bmux_9159_3_GENERIC_REAL g1(.ctl (ctl), .in_0 (in_0), .in_1 (in_1),
       .z (z));
endmodule

module csa_tree_9126_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 26'b0;"
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  wire n_73, n_77, n_78, n_82, n_83, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_222, n_226, n_230;
  assign out_0[0] = in_1[0];
  xor g32 (out_1[0], in_0[0], in_2[0]);
  and g33 (out_0[1], in_0[0], in_2[0]);
  xor g34 (n_136, in_0[1], in_1[1]);
  xor g35 (out_1[1], n_136, in_2[1]);
  nand g36 (n_137, in_0[1], in_1[1]);
  nand g4 (n_138, in_2[1], in_1[1]);
  nand g5 (n_139, in_0[1], in_2[1]);
  nand g37 (out_0[2], n_137, n_138, n_139);
  xor g38 (n_140, in_0[2], in_1[2]);
  xor g39 (out_1[2], n_140, in_2[2]);
  nand g40 (n_141, in_0[2], in_1[2]);
  nand g41 (n_142, in_2[2], in_1[2]);
  nand g42 (n_143, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_141, n_142, n_143);
  xor g43 (n_144, in_0[3], in_1[3]);
  xor g44 (out_1[3], n_144, in_2[3]);
  nand g45 (n_145, in_0[3], in_1[3]);
  nand g46 (n_146, in_2[3], in_1[3]);
  nand g47 (n_147, in_0[3], in_2[3]);
  nand g48 (out_0[4], n_145, n_146, n_147);
  xor g49 (n_148, in_0[4], in_1[4]);
  xor g50 (out_1[4], n_148, in_2[4]);
  nand g51 (n_149, in_0[4], in_1[4]);
  nand g52 (n_150, in_2[4], in_1[4]);
  nand g53 (n_151, in_0[4], in_2[4]);
  nand g54 (out_0[5], n_149, n_150, n_151);
  xor g55 (n_152, in_0[5], in_1[5]);
  xor g56 (out_1[5], n_152, in_2[5]);
  nand g57 (n_153, in_0[5], in_1[5]);
  nand g58 (n_154, in_2[5], in_1[5]);
  nand g59 (n_155, in_0[5], in_2[5]);
  nand g60 (out_0[6], n_153, n_154, n_155);
  xor g61 (n_156, in_0[6], in_1[6]);
  xor g62 (out_1[6], n_156, in_2[6]);
  nand g63 (n_157, in_0[6], in_1[6]);
  nand g64 (n_158, in_2[6], in_1[6]);
  nand g65 (n_159, in_0[6], in_2[6]);
  nand g66 (out_0[7], n_157, n_158, n_159);
  xor g67 (n_160, in_0[7], in_1[7]);
  xor g68 (out_1[7], n_160, in_2[7]);
  nand g69 (n_161, in_0[7], in_1[7]);
  nand g70 (n_162, in_2[7], in_1[7]);
  nand g71 (n_163, in_0[7], in_2[7]);
  nand g72 (out_0[8], n_161, n_162, n_163);
  xor g73 (n_164, in_0[8], in_1[8]);
  xor g74 (out_1[8], n_164, in_2[8]);
  nand g75 (n_165, in_0[8], in_1[8]);
  nand g76 (n_166, in_2[8], in_1[8]);
  nand g77 (n_167, in_0[8], in_2[8]);
  nand g78 (out_0[9], n_165, n_166, n_167);
  xor g79 (n_168, in_0[9], in_1[9]);
  xor g80 (out_1[9], n_168, in_2[9]);
  nand g81 (n_169, in_0[9], in_1[9]);
  nand g82 (n_170, in_2[9], in_1[9]);
  nand g83 (n_171, in_0[9], in_2[9]);
  nand g84 (out_0[10], n_169, n_170, n_171);
  xor g85 (n_172, in_0[10], in_1[10]);
  xor g86 (out_1[10], n_172, in_2[10]);
  nand g87 (n_173, in_0[10], in_1[10]);
  nand g88 (n_174, in_2[10], in_1[10]);
  nand g89 (n_175, in_0[10], in_2[10]);
  nand g90 (out_0[11], n_173, n_174, n_175);
  xor g91 (n_176, in_0[11], in_1[11]);
  xor g92 (out_1[11], n_176, in_2[11]);
  nand g93 (n_177, in_0[11], in_1[11]);
  nand g94 (n_178, in_2[11], in_1[11]);
  nand g95 (n_179, in_0[11], in_2[11]);
  nand g96 (out_0[12], n_177, n_178, n_179);
  xor g97 (n_180, in_0[12], in_1[12]);
  xor g98 (out_1[12], n_180, in_2[12]);
  nand g99 (n_181, in_0[12], in_1[12]);
  nand g100 (n_182, in_2[12], in_1[12]);
  nand g101 (n_183, in_0[12], in_2[12]);
  nand g102 (out_0[13], n_181, n_182, n_183);
  xor g103 (n_184, in_0[13], in_1[13]);
  xor g104 (out_1[13], n_184, in_2[13]);
  nand g105 (n_185, in_0[13], in_1[13]);
  nand g106 (n_186, in_2[13], in_1[13]);
  nand g107 (n_187, in_0[13], in_2[13]);
  nand g108 (out_0[14], n_185, n_186, n_187);
  xor g109 (n_188, in_0[14], in_1[14]);
  xor g110 (out_1[14], n_188, in_2[14]);
  nand g111 (n_189, in_0[14], in_1[14]);
  nand g112 (n_190, in_2[14], in_1[14]);
  nand g113 (n_191, in_0[14], in_2[14]);
  nand g114 (out_0[15], n_189, n_190, n_191);
  xor g115 (n_192, in_0[15], in_1[15]);
  xor g116 (out_1[15], n_192, in_2[15]);
  nand g117 (n_193, in_0[15], in_1[15]);
  nand g118 (n_194, in_2[15], in_1[15]);
  nand g119 (n_195, in_0[15], in_2[15]);
  nand g120 (out_0[16], n_193, n_194, n_195);
  xor g121 (n_196, in_0[16], in_1[16]);
  xor g122 (out_1[16], n_196, in_2[16]);
  nand g123 (n_197, in_0[16], in_1[16]);
  nand g124 (n_198, in_2[16], in_1[16]);
  nand g125 (n_199, in_0[16], in_2[16]);
  nand g126 (out_0[17], n_197, n_198, n_199);
  xor g127 (n_200, in_0[17], in_1[17]);
  xor g128 (out_1[17], n_200, in_2[17]);
  nand g129 (n_201, in_0[17], in_1[17]);
  nand g130 (n_202, in_2[17], in_1[17]);
  nand g131 (n_203, in_0[17], in_2[17]);
  nand g132 (out_0[18], n_201, n_202, n_203);
  xor g133 (n_204, in_0[18], in_1[18]);
  xor g134 (out_1[18], n_204, in_2[18]);
  nand g135 (n_205, in_0[18], in_1[18]);
  nand g136 (n_206, in_2[18], in_1[18]);
  nand g137 (n_207, in_0[18], in_2[18]);
  nand g138 (out_0[19], n_205, n_206, n_207);
  xor g139 (n_208, in_0[19], in_1[19]);
  xor g140 (out_1[19], n_208, in_2[19]);
  nand g141 (n_209, in_0[19], in_1[19]);
  nand g142 (n_210, in_2[19], in_1[19]);
  nand g143 (n_211, in_0[19], in_2[19]);
  nand g144 (out_0[20], n_209, n_210, n_211);
  xor g145 (n_212, in_0[20], in_1[20]);
  xor g146 (out_1[20], n_212, in_2[20]);
  nand g147 (n_213, in_0[20], in_1[20]);
  nand g148 (n_214, in_2[20], in_1[20]);
  nand g149 (n_215, in_0[20], in_2[20]);
  nand g150 (out_0[21], n_213, n_214, n_215);
  xor g151 (n_216, in_0[21], in_1[21]);
  xor g152 (out_1[21], n_216, in_2[21]);
  nand g153 (n_217, in_0[21], in_1[21]);
  nand g154 (n_218, in_2[21], in_1[21]);
  nand g155 (n_219, in_0[21], in_2[21]);
  nand g156 (out_0[22], n_217, n_218, n_219);
  xor g157 (n_73, in_0[22], in_1[22]);
  and g158 (n_78, in_0[22], in_1[22]);
  xor g160 (out_1[22], in_2[22], n_73);
  xor g165 (n_77, in_0[23], in_1[23]);
  and g166 (n_83, in_0[23], in_1[23]);
  nand g170 (n_226, n_78, n_77);
  nand g178 (n_230, n_83, n_82);
  or g181 (n_222, in_2[22], wc);
  not gc (wc, n_73);
  xor g185 (n_82, in_0[24], in_1[24]);
  nor g186 (out_0[25], in_0[24], in_1[24]);
  or g188 (out_0[23], wc0, wc1, n_73);
  not gc1 (wc1, n_222);
  not gc0 (wc0, in_2[22]);
  xnor g189 (out_1[23], n_78, n_77);
  or g190 (out_0[24], wc2, n_77, n_78);
  not gc2 (wc2, n_226);
  xnor g192 (out_1[24], n_83, n_82);
  or g193 (out_1[25], n_82, wc3, n_83);
  not gc3 (wc3, n_230);
endmodule

module csa_tree_9126_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  csa_tree_9126_GENERIC_REAL g1(.in_0 ({in_0[20], in_0[20], in_0[20],
       in_0[20], in_0[20:0]}), .in_1 ({in_1[20], in_1[20], in_1[20],
       in_1[20], in_1[20:0]}), .in_2 (in_2), .out_0 (out_0), .out_1
       (out_1));
endmodule

module csa_tree_9239_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 36'b0;"
  input [34:0] in_0, in_1;
  input [32:0] in_2;
  output [35:0] out_0, out_1;
  wire [34:0] in_0, in_1;
  wire [32:0] in_2;
  wire [35:0] out_0, out_1;
  wire n_103, n_107, n_108, n_112, n_113, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_223, n_224, n_225, n_226, n_227, n_228;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268;
  wire n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276;
  wire n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284;
  wire n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_295, n_296, n_297, n_298, n_299, n_300;
  wire n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308;
  wire n_309, n_312, n_316, n_320;
  assign out_0[0] = in_1[0];
  xor g42 (out_1[0], in_0[0], in_2[0]);
  and g43 (out_0[1], in_0[0], in_2[0]);
  xor g44 (n_186, in_0[1], in_1[1]);
  xor g45 (out_1[1], n_186, in_2[1]);
  nand g46 (n_187, in_0[1], in_1[1]);
  nand g4 (n_188, in_2[1], in_1[1]);
  nand g5 (n_189, in_0[1], in_2[1]);
  nand g47 (out_0[2], n_187, n_188, n_189);
  xor g48 (n_190, in_0[2], in_1[2]);
  xor g49 (out_1[2], n_190, in_2[2]);
  nand g50 (n_191, in_0[2], in_1[2]);
  nand g51 (n_192, in_2[2], in_1[2]);
  nand g52 (n_193, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_191, n_192, n_193);
  xor g53 (n_194, in_0[3], in_1[3]);
  xor g54 (out_1[3], n_194, in_2[3]);
  nand g55 (n_195, in_0[3], in_1[3]);
  nand g56 (n_196, in_2[3], in_1[3]);
  nand g57 (n_197, in_0[3], in_2[3]);
  nand g58 (out_0[4], n_195, n_196, n_197);
  xor g59 (n_198, in_0[4], in_1[4]);
  xor g60 (out_1[4], n_198, in_2[4]);
  nand g61 (n_199, in_0[4], in_1[4]);
  nand g62 (n_200, in_2[4], in_1[4]);
  nand g63 (n_201, in_0[4], in_2[4]);
  nand g64 (out_0[5], n_199, n_200, n_201);
  xor g65 (n_202, in_0[5], in_1[5]);
  xor g66 (out_1[5], n_202, in_2[5]);
  nand g67 (n_203, in_0[5], in_1[5]);
  nand g68 (n_204, in_2[5], in_1[5]);
  nand g69 (n_205, in_0[5], in_2[5]);
  nand g70 (out_0[6], n_203, n_204, n_205);
  xor g71 (n_206, in_0[6], in_1[6]);
  xor g72 (out_1[6], n_206, in_2[6]);
  nand g73 (n_207, in_0[6], in_1[6]);
  nand g74 (n_208, in_2[6], in_1[6]);
  nand g75 (n_209, in_0[6], in_2[6]);
  nand g76 (out_0[7], n_207, n_208, n_209);
  xor g77 (n_210, in_0[7], in_1[7]);
  xor g78 (out_1[7], n_210, in_2[7]);
  nand g79 (n_211, in_0[7], in_1[7]);
  nand g80 (n_212, in_2[7], in_1[7]);
  nand g81 (n_213, in_0[7], in_2[7]);
  nand g82 (out_0[8], n_211, n_212, n_213);
  xor g83 (n_214, in_0[8], in_1[8]);
  xor g84 (out_1[8], n_214, in_2[8]);
  nand g85 (n_215, in_0[8], in_1[8]);
  nand g86 (n_216, in_2[8], in_1[8]);
  nand g87 (n_217, in_0[8], in_2[8]);
  nand g88 (out_0[9], n_215, n_216, n_217);
  xor g89 (n_218, in_0[9], in_1[9]);
  xor g90 (out_1[9], n_218, in_2[9]);
  nand g91 (n_219, in_0[9], in_1[9]);
  nand g92 (n_220, in_2[9], in_1[9]);
  nand g93 (n_221, in_0[9], in_2[9]);
  nand g94 (out_0[10], n_219, n_220, n_221);
  xor g95 (n_222, in_0[10], in_1[10]);
  xor g96 (out_1[10], n_222, in_2[10]);
  nand g97 (n_223, in_0[10], in_1[10]);
  nand g98 (n_224, in_2[10], in_1[10]);
  nand g99 (n_225, in_0[10], in_2[10]);
  nand g100 (out_0[11], n_223, n_224, n_225);
  xor g101 (n_226, in_0[11], in_1[11]);
  xor g102 (out_1[11], n_226, in_2[11]);
  nand g103 (n_227, in_0[11], in_1[11]);
  nand g104 (n_228, in_2[11], in_1[11]);
  nand g105 (n_229, in_0[11], in_2[11]);
  nand g106 (out_0[12], n_227, n_228, n_229);
  xor g107 (n_230, in_0[12], in_1[12]);
  xor g108 (out_1[12], n_230, in_2[12]);
  nand g109 (n_231, in_0[12], in_1[12]);
  nand g110 (n_232, in_2[12], in_1[12]);
  nand g111 (n_233, in_0[12], in_2[12]);
  nand g112 (out_0[13], n_231, n_232, n_233);
  xor g113 (n_234, in_0[13], in_1[13]);
  xor g114 (out_1[13], n_234, in_2[13]);
  nand g115 (n_235, in_0[13], in_1[13]);
  nand g116 (n_236, in_2[13], in_1[13]);
  nand g117 (n_237, in_0[13], in_2[13]);
  nand g118 (out_0[14], n_235, n_236, n_237);
  xor g119 (n_238, in_0[14], in_1[14]);
  xor g120 (out_1[14], n_238, in_2[14]);
  nand g121 (n_239, in_0[14], in_1[14]);
  nand g122 (n_240, in_2[14], in_1[14]);
  nand g123 (n_241, in_0[14], in_2[14]);
  nand g124 (out_0[15], n_239, n_240, n_241);
  xor g125 (n_242, in_0[15], in_1[15]);
  xor g126 (out_1[15], n_242, in_2[15]);
  nand g127 (n_243, in_0[15], in_1[15]);
  nand g128 (n_244, in_2[15], in_1[15]);
  nand g129 (n_245, in_0[15], in_2[15]);
  nand g130 (out_0[16], n_243, n_244, n_245);
  xor g131 (n_246, in_0[16], in_1[16]);
  xor g132 (out_1[16], n_246, in_2[16]);
  nand g133 (n_247, in_0[16], in_1[16]);
  nand g134 (n_248, in_2[16], in_1[16]);
  nand g135 (n_249, in_0[16], in_2[16]);
  nand g136 (out_0[17], n_247, n_248, n_249);
  xor g137 (n_250, in_0[17], in_1[17]);
  xor g138 (out_1[17], n_250, in_2[17]);
  nand g139 (n_251, in_0[17], in_1[17]);
  nand g140 (n_252, in_2[17], in_1[17]);
  nand g141 (n_253, in_0[17], in_2[17]);
  nand g142 (out_0[18], n_251, n_252, n_253);
  xor g143 (n_254, in_0[18], in_1[18]);
  xor g144 (out_1[18], n_254, in_2[18]);
  nand g145 (n_255, in_0[18], in_1[18]);
  nand g146 (n_256, in_2[18], in_1[18]);
  nand g147 (n_257, in_0[18], in_2[18]);
  nand g148 (out_0[19], n_255, n_256, n_257);
  xor g149 (n_258, in_0[19], in_1[19]);
  xor g150 (out_1[19], n_258, in_2[19]);
  nand g151 (n_259, in_0[19], in_1[19]);
  nand g152 (n_260, in_2[19], in_1[19]);
  nand g153 (n_261, in_0[19], in_2[19]);
  nand g154 (out_0[20], n_259, n_260, n_261);
  xor g155 (n_262, in_0[20], in_1[20]);
  xor g156 (out_1[20], n_262, in_2[20]);
  nand g157 (n_263, in_0[20], in_1[20]);
  nand g158 (n_264, in_2[20], in_1[20]);
  nand g159 (n_265, in_0[20], in_2[20]);
  nand g160 (out_0[21], n_263, n_264, n_265);
  xor g161 (n_266, in_0[21], in_1[21]);
  xor g162 (out_1[21], n_266, in_2[21]);
  nand g163 (n_267, in_0[21], in_1[21]);
  nand g164 (n_268, in_2[21], in_1[21]);
  nand g165 (n_269, in_0[21], in_2[21]);
  nand g166 (out_0[22], n_267, n_268, n_269);
  xor g167 (n_270, in_0[22], in_1[22]);
  xor g168 (out_1[22], n_270, in_2[22]);
  nand g169 (n_271, in_0[22], in_1[22]);
  nand g170 (n_272, in_2[22], in_1[22]);
  nand g171 (n_273, in_0[22], in_2[22]);
  nand g172 (out_0[23], n_271, n_272, n_273);
  xor g173 (n_274, in_0[23], in_1[23]);
  xor g174 (out_1[23], n_274, in_2[23]);
  nand g175 (n_275, in_0[23], in_1[23]);
  nand g176 (n_276, in_2[23], in_1[23]);
  nand g177 (n_277, in_0[23], in_2[23]);
  nand g178 (out_0[24], n_275, n_276, n_277);
  xor g179 (n_278, in_0[24], in_1[24]);
  xor g180 (out_1[24], n_278, in_2[24]);
  nand g181 (n_279, in_0[24], in_1[24]);
  nand g182 (n_280, in_2[24], in_1[24]);
  nand g183 (n_281, in_0[24], in_2[24]);
  nand g184 (out_0[25], n_279, n_280, n_281);
  xor g185 (n_282, in_0[25], in_1[25]);
  xor g186 (out_1[25], n_282, in_2[25]);
  nand g187 (n_283, in_0[25], in_1[25]);
  nand g188 (n_284, in_2[25], in_1[25]);
  nand g189 (n_285, in_0[25], in_2[25]);
  nand g190 (out_0[26], n_283, n_284, n_285);
  xor g191 (n_286, in_0[26], in_1[26]);
  xor g192 (out_1[26], n_286, in_2[26]);
  nand g193 (n_287, in_0[26], in_1[26]);
  nand g194 (n_288, in_2[26], in_1[26]);
  nand g195 (n_289, in_0[26], in_2[26]);
  nand g196 (out_0[27], n_287, n_288, n_289);
  xor g197 (n_290, in_0[27], in_1[27]);
  xor g198 (out_1[27], n_290, in_2[27]);
  nand g199 (n_291, in_0[27], in_1[27]);
  nand g200 (n_292, in_2[27], in_1[27]);
  nand g201 (n_293, in_0[27], in_2[27]);
  nand g202 (out_0[28], n_291, n_292, n_293);
  xor g203 (n_294, in_0[28], in_1[28]);
  xor g204 (out_1[28], n_294, in_2[28]);
  nand g205 (n_295, in_0[28], in_1[28]);
  nand g206 (n_296, in_2[28], in_1[28]);
  nand g207 (n_297, in_0[28], in_2[28]);
  nand g208 (out_0[29], n_295, n_296, n_297);
  xor g209 (n_298, in_0[29], in_1[29]);
  xor g210 (out_1[29], n_298, in_2[29]);
  nand g211 (n_299, in_0[29], in_1[29]);
  nand g212 (n_300, in_2[29], in_1[29]);
  nand g213 (n_301, in_0[29], in_2[29]);
  nand g214 (out_0[30], n_299, n_300, n_301);
  xor g215 (n_302, in_0[30], in_1[30]);
  xor g216 (out_1[30], n_302, in_2[30]);
  nand g217 (n_303, in_0[30], in_1[30]);
  nand g218 (n_304, in_2[30], in_1[30]);
  nand g219 (n_305, in_0[30], in_2[30]);
  nand g220 (out_0[31], n_303, n_304, n_305);
  xor g221 (n_306, in_0[31], in_1[31]);
  xor g222 (out_1[31], n_306, in_2[31]);
  nand g223 (n_307, in_0[31], in_1[31]);
  nand g224 (n_308, in_2[31], in_1[31]);
  nand g225 (n_309, in_0[31], in_2[31]);
  nand g226 (out_0[32], n_307, n_308, n_309);
  xor g227 (n_103, in_0[32], in_1[32]);
  and g228 (n_108, in_0[32], in_1[32]);
  xor g230 (out_1[32], in_2[32], n_103);
  xor g235 (n_107, in_0[33], in_1[33]);
  and g236 (n_113, in_0[33], in_1[33]);
  nand g240 (n_316, n_108, n_107);
  nand g248 (n_320, n_113, n_112);
  or g251 (n_312, in_2[32], wc);
  not gc (wc, n_103);
  xor g255 (n_112, in_0[34], in_1[34]);
  nor g256 (out_0[35], in_0[34], in_1[34]);
  or g258 (out_0[33], wc0, wc1, n_103);
  not gc1 (wc1, n_312);
  not gc0 (wc0, in_2[32]);
  xnor g259 (out_1[33], n_108, n_107);
  or g260 (out_0[34], wc2, n_107, n_108);
  not gc2 (wc2, n_316);
  xnor g262 (out_1[34], n_113, n_112);
  or g263 (out_1[35], n_112, wc3, n_113);
  not gc3 (wc3, n_320);
endmodule

module csa_tree_9239_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [34:0] in_0, in_1;
  input [32:0] in_2;
  output [35:0] out_0, out_1;
  wire [34:0] in_0, in_1;
  wire [32:0] in_2;
  wire [35:0] out_0, out_1;
  csa_tree_9239_GENERIC_REAL g1(.in_0 ({in_0[34], in_0[31], in_0[31],
       in_0[31:0]}), .in_1 ({in_1[34], in_1[31], in_1[31],
       in_1[31:0]}), .in_2 (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_add_252_40_group_16906_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [36:0] in_0, in_1;
  input [34:0] in_2;
  output [35:0] out_0;
  wire [36:0] in_0, in_1;
  wire [34:0] in_2;
  wire [35:0] out_0;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_280;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_356, n_363, n_364, n_365, n_366, n_367;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_376, n_377;
  wire n_378, n_379, n_380, n_382, n_383, n_384, n_385, n_386;
  wire n_388, n_389, n_390, n_391, n_392, n_394, n_395, n_396;
  wire n_397, n_398, n_400, n_401, n_402, n_403, n_404, n_406;
  wire n_407, n_408, n_409, n_410, n_412, n_413, n_414, n_415;
  wire n_416, n_418, n_419, n_420, n_421, n_422, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_434;
  wire n_435, n_436, n_437, n_438, n_440, n_441, n_442, n_443;
  wire n_444, n_446, n_447, n_448, n_449, n_450, n_452, n_453;
  wire n_454, n_455, n_456, n_458, n_459, n_460, n_461, n_462;
  wire n_464, n_465, n_466, n_467, n_468, n_469, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_478, n_480, n_482, n_483;
  wire n_485, n_486, n_488, n_490, n_492, n_493, n_495, n_496;
  wire n_498, n_500, n_502, n_503, n_505, n_506, n_508, n_510;
  wire n_512, n_513, n_515, n_516, n_518, n_520, n_522, n_523;
  wire n_525, n_526, n_528, n_530, n_532, n_533, n_535, n_536;
  wire n_538, n_540, n_542, n_543, n_545, n_546, n_548, n_550;
  wire n_552, n_553, n_554, n_556, n_557, n_558, n_560, n_561;
  wire n_562, n_563, n_565, n_567, n_569, n_570, n_571, n_573;
  wire n_574, n_575, n_577, n_578, n_580, n_582, n_584, n_585;
  wire n_586, n_588, n_589, n_590, n_592, n_593, n_595, n_597;
  wire n_599, n_600, n_601, n_603, n_604, n_605, n_607, n_609;
  wire n_610, n_611, n_613, n_614, n_616, n_617, n_618, n_619;
  wire n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627;
  wire n_628, n_629, n_630, n_632, n_635, n_637, n_638, n_639;
  wire n_642, n_645, n_647, n_648, n_650, n_652, n_653, n_655;
  wire n_657, n_658, n_660, n_662, n_663, n_665, n_667, n_668;
  wire n_669, n_671, n_672, n_674, n_675, n_676, n_677, n_678;
  wire n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_687;
  wire n_688, n_689, n_691, n_692, n_693, n_695, n_696, n_697;
  wire n_699, n_700, n_701, n_703, n_704, n_705, n_707, n_708;
  wire n_709, n_711, n_712, n_713, n_715, n_716, n_717, n_719;
  wire n_720, n_721, n_723, n_724, n_725, n_726, n_728, n_729;
  wire n_730, n_732, n_733, n_734, n_735, n_737, n_738, n_739;
  wire n_741, n_742, n_743, n_744, n_746, n_747, n_749, n_750;
  wire n_752, n_753, n_754, n_755, n_757, n_758, n_759, n_761;
  wire n_762, n_763, n_764, n_766, n_767, n_769, n_770, n_772;
  wire n_773, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_785, n_787, n_788, n_790, n_791, n_793;
  wire n_794, n_795, n_796, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_805, n_807, n_808, n_809;
  xor g39 (n_216, in_0[1], in_2[1]);
  and g2 (n_179, in_0[1], in_2[1]);
  xor g40 (n_225, in_0[2], in_2[2]);
  xor g41 (n_215, n_225, in_1[2]);
  nand g3 (n_226, in_0[2], in_2[2]);
  nand g42 (n_227, in_1[2], in_2[2]);
  nand g43 (n_228, in_0[2], in_1[2]);
  nand g44 (n_178, n_226, n_227, n_228);
  xor g45 (n_229, in_0[3], in_2[3]);
  xor g46 (n_214, n_229, in_1[3]);
  nand g47 (n_230, in_0[3], in_2[3]);
  nand g4 (n_231, in_1[3], in_2[3]);
  nand g48 (n_232, in_0[3], in_1[3]);
  nand g49 (n_177, n_230, n_231, n_232);
  xor g50 (n_233, in_0[4], in_2[4]);
  xor g51 (n_213, n_233, in_1[4]);
  nand g52 (n_234, in_0[4], in_2[4]);
  nand g53 (n_235, in_1[4], in_2[4]);
  nand g5 (n_236, in_0[4], in_1[4]);
  nand g54 (n_176, n_234, n_235, n_236);
  xor g55 (n_237, in_0[5], in_2[5]);
  xor g56 (n_212, n_237, in_1[5]);
  nand g57 (n_238, in_0[5], in_2[5]);
  nand g58 (n_239, in_1[5], in_2[5]);
  nand g59 (n_240, in_0[5], in_1[5]);
  nand g6 (n_175, n_238, n_239, n_240);
  xor g60 (n_241, in_0[6], in_2[6]);
  xor g61 (n_211, n_241, in_1[6]);
  nand g62 (n_242, in_0[6], in_2[6]);
  nand g63 (n_243, in_1[6], in_2[6]);
  nand g64 (n_244, in_0[6], in_1[6]);
  nand g65 (n_174, n_242, n_243, n_244);
  xor g66 (n_245, in_0[7], in_2[7]);
  xor g67 (n_210, n_245, in_1[7]);
  nand g68 (n_246, in_0[7], in_2[7]);
  nand g69 (n_247, in_1[7], in_2[7]);
  nand g70 (n_248, in_0[7], in_1[7]);
  nand g71 (n_173, n_246, n_247, n_248);
  xor g72 (n_249, in_0[8], in_2[8]);
  xor g73 (n_209, n_249, in_1[8]);
  nand g74 (n_250, in_0[8], in_2[8]);
  nand g75 (n_251, in_1[8], in_2[8]);
  nand g76 (n_252, in_0[8], in_1[8]);
  nand g77 (n_172, n_250, n_251, n_252);
  xor g78 (n_253, in_0[9], in_2[9]);
  xor g79 (n_208, n_253, in_1[9]);
  nand g80 (n_254, in_0[9], in_2[9]);
  nand g81 (n_255, in_1[9], in_2[9]);
  nand g82 (n_256, in_0[9], in_1[9]);
  nand g83 (n_171, n_254, n_255, n_256);
  xor g84 (n_257, in_0[10], in_2[10]);
  xor g85 (n_207, n_257, in_1[10]);
  nand g86 (n_258, in_0[10], in_2[10]);
  nand g87 (n_217, in_1[10], in_2[10]);
  nand g88 (n_218, in_0[10], in_1[10]);
  nand g89 (n_170, n_258, n_217, n_218);
  xor g90 (n_259, in_0[11], in_2[11]);
  xor g91 (n_206, n_259, in_1[11]);
  nand g92 (n_260, in_0[11], in_2[11]);
  nand g93 (n_261, in_1[11], in_2[11]);
  nand g94 (n_262, in_0[11], in_1[11]);
  nand g95 (n_169, n_260, n_261, n_262);
  xor g96 (n_263, in_0[12], in_2[12]);
  xor g97 (n_205, n_263, in_1[12]);
  nand g98 (n_264, in_0[12], in_2[12]);
  nand g99 (n_265, in_1[12], in_2[12]);
  nand g100 (n_266, in_0[12], in_1[12]);
  nand g101 (n_168, n_264, n_265, n_266);
  xor g102 (n_267, in_0[13], in_2[13]);
  xor g103 (n_204, n_267, in_1[13]);
  nand g104 (n_268, in_0[13], in_2[13]);
  nand g105 (n_269, in_1[13], in_2[13]);
  nand g106 (n_270, in_0[13], in_1[13]);
  nand g107 (n_167, n_268, n_269, n_270);
  xor g108 (n_271, in_0[14], in_2[14]);
  xor g109 (n_203, n_271, in_1[14]);
  nand g110 (n_272, in_0[14], in_2[14]);
  nand g111 (n_273, in_1[14], in_2[14]);
  nand g112 (n_274, in_0[14], in_1[14]);
  nand g113 (n_166, n_272, n_273, n_274);
  xor g114 (n_275, in_0[15], in_2[15]);
  xor g115 (n_202, n_275, in_1[15]);
  nand g116 (n_276, in_0[15], in_2[15]);
  nand g117 (n_277, in_1[15], in_2[15]);
  nand g118 (n_278, in_0[15], in_1[15]);
  nand g119 (n_165, n_276, n_277, n_278);
  xor g120 (n_279, in_0[16], in_2[16]);
  xor g121 (n_201, n_279, in_1[16]);
  nand g122 (n_280, in_0[16], in_2[16]);
  nand g123 (n_281, in_1[16], in_2[16]);
  nand g124 (n_282, in_0[16], in_1[16]);
  nand g125 (n_164, n_280, n_281, n_282);
  xor g126 (n_283, in_0[17], in_2[17]);
  xor g127 (n_200, n_283, in_1[17]);
  nand g128 (n_284, in_0[17], in_2[17]);
  nand g129 (n_285, in_1[17], in_2[17]);
  nand g130 (n_286, in_0[17], in_1[17]);
  nand g131 (n_163, n_284, n_285, n_286);
  xor g132 (n_287, in_0[18], in_2[18]);
  xor g133 (n_199, n_287, in_1[18]);
  nand g134 (n_288, in_0[18], in_2[18]);
  nand g135 (n_289, in_1[18], in_2[18]);
  nand g136 (n_290, in_0[18], in_1[18]);
  nand g137 (n_162, n_288, n_289, n_290);
  xor g138 (n_291, in_0[19], in_2[19]);
  xor g139 (n_198, n_291, in_1[19]);
  nand g140 (n_292, in_0[19], in_2[19]);
  nand g141 (n_293, in_1[19], in_2[19]);
  nand g142 (n_294, in_0[19], in_1[19]);
  nand g143 (n_161, n_292, n_293, n_294);
  xor g144 (n_295, in_0[20], in_2[20]);
  xor g145 (n_197, n_295, in_1[20]);
  nand g146 (n_296, in_0[20], in_2[20]);
  nand g147 (n_297, in_1[20], in_2[20]);
  nand g148 (n_298, in_0[20], in_1[20]);
  nand g149 (n_160, n_296, n_297, n_298);
  xor g150 (n_299, in_0[21], in_2[21]);
  xor g151 (n_196, n_299, in_1[21]);
  nand g152 (n_300, in_0[21], in_2[21]);
  nand g153 (n_301, in_1[21], in_2[21]);
  nand g154 (n_302, in_0[21], in_1[21]);
  nand g155 (n_159, n_300, n_301, n_302);
  xor g156 (n_303, in_0[22], in_2[22]);
  xor g157 (n_195, n_303, in_1[22]);
  nand g158 (n_304, in_0[22], in_2[22]);
  nand g159 (n_305, in_1[22], in_2[22]);
  nand g160 (n_306, in_0[22], in_1[22]);
  nand g161 (n_158, n_304, n_305, n_306);
  xor g162 (n_307, in_0[23], in_2[23]);
  xor g163 (n_194, n_307, in_1[23]);
  nand g164 (n_308, in_0[23], in_2[23]);
  nand g165 (n_309, in_1[23], in_2[23]);
  nand g166 (n_310, in_0[23], in_1[23]);
  nand g167 (n_157, n_308, n_309, n_310);
  xor g168 (n_311, in_0[24], in_2[24]);
  xor g169 (n_193, n_311, in_1[24]);
  nand g170 (n_312, in_0[24], in_2[24]);
  nand g171 (n_313, in_1[24], in_2[24]);
  nand g172 (n_314, in_0[24], in_1[24]);
  nand g173 (n_156, n_312, n_313, n_314);
  xor g174 (n_315, in_0[25], in_2[25]);
  xor g175 (n_192, n_315, in_1[25]);
  nand g176 (n_316, in_0[25], in_2[25]);
  nand g177 (n_317, in_1[25], in_2[25]);
  nand g178 (n_318, in_0[25], in_1[25]);
  nand g179 (n_155, n_316, n_317, n_318);
  xor g180 (n_319, in_0[26], in_2[26]);
  xor g181 (n_191, n_319, in_1[26]);
  nand g182 (n_320, in_0[26], in_2[26]);
  nand g183 (n_321, in_1[26], in_2[26]);
  nand g184 (n_322, in_0[26], in_1[26]);
  nand g185 (n_154, n_320, n_321, n_322);
  xor g186 (n_323, in_0[27], in_2[27]);
  xor g187 (n_190, n_323, in_1[27]);
  nand g188 (n_324, in_0[27], in_2[27]);
  nand g189 (n_325, in_1[27], in_2[27]);
  nand g190 (n_326, in_0[27], in_1[27]);
  nand g191 (n_153, n_324, n_325, n_326);
  xor g192 (n_327, in_0[28], in_2[28]);
  xor g193 (n_189, n_327, in_1[28]);
  nand g194 (n_328, in_0[28], in_2[28]);
  nand g195 (n_329, in_1[28], in_2[28]);
  nand g196 (n_330, in_0[28], in_1[28]);
  nand g197 (n_152, n_328, n_329, n_330);
  xor g198 (n_331, in_0[29], in_2[29]);
  xor g199 (n_188, n_331, in_1[29]);
  nand g200 (n_332, in_0[29], in_2[29]);
  nand g201 (n_333, in_1[29], in_2[29]);
  nand g202 (n_334, in_0[29], in_1[29]);
  nand g203 (n_151, n_332, n_333, n_334);
  xor g204 (n_335, in_0[30], in_2[30]);
  xor g205 (n_187, n_335, in_1[30]);
  nand g206 (n_336, in_0[30], in_2[30]);
  nand g207 (n_337, in_1[30], in_2[30]);
  nand g208 (n_338, in_0[30], in_1[30]);
  nand g209 (n_150, n_336, n_337, n_338);
  xor g210 (n_339, in_0[31], in_2[31]);
  xor g211 (n_186, n_339, in_1[31]);
  nand g212 (n_340, in_0[31], in_2[31]);
  nand g213 (n_341, in_1[31], in_2[31]);
  nand g214 (n_342, in_0[31], in_1[31]);
  nand g215 (n_149, n_340, n_341, n_342);
  xor g216 (n_343, in_0[32], in_2[32]);
  xor g217 (n_185, n_343, in_1[32]);
  nand g218 (n_344, in_0[32], in_2[32]);
  nand g219 (n_345, in_1[32], in_2[32]);
  nand g220 (n_346, in_0[32], in_1[32]);
  nand g221 (n_148, n_344, n_345, n_346);
  xor g222 (n_347, in_0[33], in_2[33]);
  xor g223 (n_184, n_347, in_1[33]);
  nand g224 (n_348, in_0[33], in_2[33]);
  nand g225 (n_349, in_1[33], in_2[33]);
  nand g226 (n_350, in_0[33], in_1[33]);
  nand g227 (n_147, n_348, n_349, n_350);
  nand g235 (n_146, n_352, n_353, n_354);
  xor g239 (n_182, n_356, in_0[34]);
  xor g246 (n_809, in_2[0], in_1[0]);
  nand g247 (n_363, in_2[0], in_1[0]);
  nand g248 (n_364, in_2[0], in_0[0]);
  nand g7 (n_365, in_1[0], in_0[0]);
  nand g8 (n_367, n_363, n_364, n_365);
  nor g9 (n_366, in_1[1], n_216);
  nand g10 (n_369, in_1[1], n_216);
  nor g11 (n_376, n_179, n_215);
  nand g12 (n_371, n_179, n_215);
  nor g13 (n_372, n_178, n_214);
  nand g14 (n_373, n_178, n_214);
  nor g15 (n_382, n_177, n_213);
  nand g16 (n_377, n_177, n_213);
  nor g17 (n_378, n_176, n_212);
  nand g18 (n_379, n_176, n_212);
  nor g19 (n_388, n_175, n_211);
  nand g20 (n_383, n_175, n_211);
  nor g21 (n_384, n_174, n_210);
  nand g22 (n_385, n_174, n_210);
  nor g23 (n_394, n_173, n_209);
  nand g24 (n_389, n_173, n_209);
  nor g25 (n_390, n_172, n_208);
  nand g26 (n_391, n_172, n_208);
  nor g27 (n_400, n_171, n_207);
  nand g28 (n_395, n_171, n_207);
  nor g29 (n_396, n_170, n_206);
  nand g30 (n_397, n_170, n_206);
  nor g31 (n_406, n_169, n_205);
  nand g32 (n_401, n_169, n_205);
  nor g33 (n_402, n_168, n_204);
  nand g34 (n_403, n_168, n_204);
  nor g35 (n_412, n_167, n_203);
  nand g36 (n_407, n_167, n_203);
  nor g37 (n_408, n_166, n_202);
  nand g38 (n_409, n_166, n_202);
  nor g249 (n_418, n_165, n_201);
  nand g250 (n_413, n_165, n_201);
  nor g251 (n_414, n_164, n_200);
  nand g252 (n_415, n_164, n_200);
  nor g253 (n_424, n_163, n_199);
  nand g254 (n_419, n_163, n_199);
  nor g255 (n_420, n_162, n_198);
  nand g256 (n_421, n_162, n_198);
  nor g257 (n_181, n_161, n_197);
  nand g258 (n_425, n_161, n_197);
  nor g259 (n_426, n_160, n_196);
  nand g260 (n_427, n_160, n_196);
  nor g261 (n_434, n_159, n_195);
  nand g262 (n_429, n_159, n_195);
  nor g263 (n_430, n_158, n_194);
  nand g264 (n_431, n_158, n_194);
  nor g265 (n_440, n_157, n_193);
  nand g266 (n_435, n_157, n_193);
  nor g267 (n_436, n_156, n_192);
  nand g268 (n_437, n_156, n_192);
  nor g269 (n_446, n_155, n_191);
  nand g270 (n_441, n_155, n_191);
  nor g271 (n_442, n_154, n_190);
  nand g272 (n_443, n_154, n_190);
  nor g273 (n_452, n_153, n_189);
  nand g274 (n_447, n_153, n_189);
  nor g275 (n_448, n_152, n_188);
  nand g276 (n_449, n_152, n_188);
  nor g277 (n_458, n_151, n_187);
  nand g278 (n_453, n_151, n_187);
  nor g279 (n_454, n_150, n_186);
  nand g280 (n_455, n_150, n_186);
  nor g281 (n_464, n_149, n_185);
  nand g282 (n_459, n_149, n_185);
  nor g283 (n_460, n_148, n_184);
  nand g284 (n_461, n_148, n_184);
  nor g285 (n_468, n_147, n_183);
  nand g286 (n_465, n_147, n_183);
  nand g291 (n_469, n_369, n_370);
  nor g292 (n_374, n_371, n_372);
  nor g295 (n_472, n_376, n_372);
  nor g296 (n_380, n_377, n_378);
  nor g299 (n_478, n_382, n_378);
  nor g300 (n_386, n_383, n_384);
  nor g303 (n_480, n_388, n_384);
  nor g304 (n_392, n_389, n_390);
  nor g307 (n_488, n_394, n_390);
  nor g308 (n_398, n_395, n_396);
  nor g311 (n_490, n_400, n_396);
  nor g312 (n_404, n_401, n_402);
  nor g315 (n_498, n_406, n_402);
  nor g316 (n_410, n_407, n_408);
  nor g319 (n_500, n_412, n_408);
  nor g320 (n_416, n_413, n_414);
  nor g323 (n_508, n_418, n_414);
  nor g324 (n_422, n_419, n_420);
  nor g327 (n_510, n_424, n_420);
  nor g328 (n_428, n_425, n_426);
  nor g331 (n_518, n_181, n_426);
  nor g332 (n_432, n_429, n_430);
  nor g335 (n_520, n_434, n_430);
  nor g336 (n_438, n_435, n_436);
  nor g339 (n_528, n_440, n_436);
  nor g340 (n_444, n_441, n_442);
  nor g343 (n_530, n_446, n_442);
  nor g344 (n_450, n_447, n_448);
  nor g347 (n_538, n_452, n_448);
  nor g348 (n_456, n_453, n_454);
  nor g351 (n_540, n_458, n_454);
  nor g352 (n_462, n_459, n_460);
  nor g355 (n_548, n_464, n_460);
  nand g358 (n_728, n_371, n_471);
  nand g359 (n_474, n_472, n_469);
  nand g360 (n_550, n_473, n_474);
  nor g361 (n_476, n_388, n_475);
  nand g370 (n_558, n_478, n_480);
  nor g371 (n_486, n_400, n_485);
  nand g380 (n_565, n_488, n_490);
  nor g381 (n_496, n_412, n_495);
  nand g390 (n_573, n_498, n_500);
  nor g391 (n_506, n_424, n_505);
  nand g400 (n_580, n_508, n_510);
  nor g401 (n_516, n_434, n_515);
  nand g410 (n_588, n_518, n_520);
  nor g411 (n_526, n_446, n_525);
  nand g420 (n_595, n_528, n_530);
  nor g421 (n_536, n_458, n_535);
  nand g430 (n_603, n_538, n_540);
  nor g431 (n_546, n_468, n_545);
  nand g438 (n_732, n_377, n_552);
  nand g439 (n_553, n_478, n_550);
  nand g440 (n_734, n_475, n_553);
  nand g443 (n_737, n_556, n_557);
  nand g446 (n_607, n_560, n_561);
  nor g447 (n_563, n_406, n_562);
  nor g450 (n_617, n_406, n_565);
  nor g456 (n_571, n_569, n_562);
  nor g459 (n_623, n_565, n_569);
  nor g460 (n_575, n_573, n_562);
  nor g463 (n_626, n_565, n_573);
  nor g464 (n_578, n_181, n_577);
  nor g467 (n_675, n_181, n_580);
  nor g473 (n_586, n_584, n_577);
  nor g476 (n_681, n_580, n_584);
  nor g477 (n_590, n_588, n_577);
  nor g480 (n_632, n_580, n_588);
  nor g481 (n_593, n_452, n_592);
  nor g484 (n_645, n_452, n_595);
  nor g490 (n_601, n_599, n_592);
  nor g493 (n_655, n_595, n_599);
  nor g494 (n_605, n_603, n_592);
  nor g497 (n_660, n_595, n_603);
  nand g500 (n_741, n_389, n_609);
  nand g501 (n_610, n_488, n_607);
  nand g502 (n_743, n_485, n_610);
  nand g505 (n_746, n_613, n_614);
  nand g508 (n_749, n_562, n_616);
  nand g509 (n_619, n_617, n_607);
  nand g510 (n_752, n_618, n_619);
  nand g511 (n_622, n_620, n_607);
  nand g512 (n_754, n_621, n_622);
  nand g513 (n_625, n_623, n_607);
  nand g514 (n_757, n_624, n_625);
  nand g515 (n_628, n_626, n_607);
  nand g516 (n_665, n_627, n_628);
  nor g517 (n_630, n_440, n_629);
  nand g526 (n_689, n_528, n_632);
  nor g527 (n_639, n_637, n_629);
  nor g532 (n_642, n_595, n_629);
  nand g541 (n_701, n_632, n_645);
  nand g546 (n_705, n_632, n_650);
  nand g551 (n_709, n_632, n_655);
  nand g556 (n_713, n_632, n_660);
  nand g559 (n_761, n_413, n_667);
  nand g560 (n_668, n_508, n_665);
  nand g561 (n_763, n_505, n_668);
  nand g564 (n_766, n_671, n_672);
  nand g567 (n_769, n_577, n_674);
  nand g568 (n_677, n_675, n_665);
  nand g569 (n_772, n_676, n_677);
  nand g570 (n_680, n_678, n_665);
  nand g571 (n_774, n_679, n_680);
  nand g572 (n_683, n_681, n_665);
  nand g573 (n_777, n_682, n_683);
  nand g574 (n_684, n_632, n_665);
  nand g575 (n_779, n_629, n_684);
  nand g578 (n_782, n_687, n_688);
  nand g581 (n_784, n_691, n_692);
  nand g584 (n_787, n_695, n_696);
  nand g587 (n_790, n_699, n_700);
  nand g590 (n_793, n_703, n_704);
  nand g593 (n_795, n_707, n_708);
  nand g596 (n_798, n_711, n_712);
  nand g599 (n_717, n_715, n_716);
  nand g602 (n_802, n_459, n_719);
  nand g603 (n_720, n_548, n_717);
  nand g604 (n_804, n_545, n_720);
  nand g607 (n_807, n_723, n_724);
  xnor g609 (out_0[1], n_367, n_725);
  xnor g611 (out_0[2], n_469, n_726);
  xnor g614 (out_0[3], n_728, n_729);
  xnor g616 (out_0[4], n_550, n_730);
  xnor g619 (out_0[5], n_732, n_733);
  xnor g621 (out_0[6], n_734, n_735);
  xnor g624 (out_0[7], n_737, n_738);
  xnor g626 (out_0[8], n_607, n_739);
  xnor g629 (out_0[9], n_741, n_742);
  xnor g631 (out_0[10], n_743, n_744);
  xnor g634 (out_0[11], n_746, n_747);
  xnor g637 (out_0[12], n_749, n_750);
  xnor g640 (out_0[13], n_752, n_753);
  xnor g642 (out_0[14], n_754, n_755);
  xnor g645 (out_0[15], n_757, n_758);
  xnor g647 (out_0[16], n_665, n_759);
  xnor g650 (out_0[17], n_761, n_762);
  xnor g652 (out_0[18], n_763, n_764);
  xnor g655 (out_0[19], n_766, n_767);
  xnor g658 (out_0[20], n_769, n_770);
  xnor g661 (out_0[21], n_772, n_773);
  xnor g663 (out_0[22], n_774, n_775);
  xnor g666 (out_0[23], n_777, n_778);
  xnor g668 (out_0[24], n_779, n_780);
  xnor g671 (out_0[25], n_782, n_783);
  xnor g673 (out_0[26], n_784, n_785);
  xnor g676 (out_0[27], n_787, n_788);
  xnor g679 (out_0[28], n_790, n_791);
  xnor g682 (out_0[29], n_793, n_794);
  xnor g684 (out_0[30], n_795, n_796);
  xnor g687 (out_0[31], n_798, n_799);
  xnor g689 (out_0[32], n_717, n_800);
  xnor g692 (out_0[33], n_802, n_803);
  xnor g694 (out_0[34], n_804, n_805);
  xnor g697 (out_0[35], n_807, n_808);
  xor g698 (out_0[0], in_0[0], n_809);
  xnor g701 (n_351, in_1[34], in_2[34]);
  or g702 (n_352, in_2[34], wc);
  not gc (wc, in_1[34]);
  or g703 (n_353, in_0[34], in_2[34]);
  or g704 (n_354, wc0, in_0[34]);
  not gc0 (wc0, in_1[34]);
  xnor g705 (n_356, in_0[35], in_1[35]);
  xnor g706 (n_183, n_351, in_0[34]);
  or g707 (n_370, n_366, wc1);
  not gc1 (wc1, n_367);
  or g708 (n_725, wc2, n_366);
  not gc2 (wc2, n_369);
  and g709 (n_466, n_146, n_182);
  or g710 (n_467, n_146, n_182);
  and g711 (n_473, wc3, n_373);
  not gc3 (wc3, n_374);
  and g712 (n_475, wc4, n_379);
  not gc4 (wc4, n_380);
  and g713 (n_482, wc5, n_385);
  not gc5 (wc5, n_386);
  and g714 (n_485, wc6, n_391);
  not gc6 (wc6, n_392);
  and g715 (n_492, wc7, n_397);
  not gc7 (wc7, n_398);
  and g716 (n_495, wc8, n_403);
  not gc8 (wc8, n_404);
  and g717 (n_502, wc9, n_409);
  not gc9 (wc9, n_410);
  and g718 (n_505, wc10, n_415);
  not gc10 (wc10, n_416);
  and g719 (n_512, wc11, n_421);
  not gc11 (wc11, n_422);
  and g720 (n_515, wc12, n_427);
  not gc12 (wc12, n_428);
  and g721 (n_522, wc13, n_431);
  not gc13 (wc13, n_432);
  and g722 (n_525, wc14, n_437);
  not gc14 (wc14, n_438);
  and g723 (n_532, wc15, n_443);
  not gc15 (wc15, n_444);
  and g724 (n_535, wc16, n_449);
  not gc16 (wc16, n_450);
  and g725 (n_542, wc17, n_455);
  not gc17 (wc17, n_456);
  and g726 (n_545, wc18, n_461);
  not gc18 (wc18, n_462);
  or g727 (n_554, wc19, n_388);
  not gc19 (wc19, n_478);
  or g728 (n_611, wc20, n_400);
  not gc20 (wc20, n_488);
  or g729 (n_569, wc21, n_412);
  not gc21 (wc21, n_498);
  or g730 (n_669, wc22, n_424);
  not gc22 (wc22, n_508);
  or g731 (n_584, wc23, n_434);
  not gc23 (wc23, n_518);
  or g732 (n_637, wc24, n_446);
  not gc24 (wc24, n_528);
  or g733 (n_599, wc25, n_458);
  not gc25 (wc25, n_538);
  or g734 (n_726, wc26, n_376);
  not gc26 (wc26, n_371);
  or g735 (n_729, wc27, n_372);
  not gc27 (wc27, n_373);
  or g736 (n_730, wc28, n_382);
  not gc28 (wc28, n_377);
  or g737 (n_733, wc29, n_378);
  not gc29 (wc29, n_379);
  or g738 (n_735, wc30, n_388);
  not gc30 (wc30, n_383);
  or g739 (n_738, wc31, n_384);
  not gc31 (wc31, n_385);
  or g740 (n_739, wc32, n_394);
  not gc32 (wc32, n_389);
  or g741 (n_742, wc33, n_390);
  not gc33 (wc33, n_391);
  or g742 (n_744, wc34, n_400);
  not gc34 (wc34, n_395);
  or g743 (n_747, wc35, n_396);
  not gc35 (wc35, n_397);
  or g744 (n_750, wc36, n_406);
  not gc36 (wc36, n_401);
  or g745 (n_753, wc37, n_402);
  not gc37 (wc37, n_403);
  or g746 (n_755, wc38, n_412);
  not gc38 (wc38, n_407);
  or g747 (n_758, wc39, n_408);
  not gc39 (wc39, n_409);
  or g748 (n_759, wc40, n_418);
  not gc40 (wc40, n_413);
  or g749 (n_762, wc41, n_414);
  not gc41 (wc41, n_415);
  or g750 (n_764, wc42, n_424);
  not gc42 (wc42, n_419);
  or g751 (n_767, wc43, n_420);
  not gc43 (wc43, n_421);
  or g752 (n_770, wc44, n_181);
  not gc44 (wc44, n_425);
  or g753 (n_773, wc45, n_426);
  not gc45 (wc45, n_427);
  or g754 (n_775, wc46, n_434);
  not gc46 (wc46, n_429);
  or g755 (n_778, wc47, n_430);
  not gc47 (wc47, n_431);
  or g756 (n_780, wc48, n_440);
  not gc48 (wc48, n_435);
  or g757 (n_783, wc49, n_436);
  not gc49 (wc49, n_437);
  or g758 (n_785, wc50, n_446);
  not gc50 (wc50, n_441);
  or g759 (n_788, wc51, n_442);
  not gc51 (wc51, n_443);
  or g760 (n_791, wc52, n_452);
  not gc52 (wc52, n_447);
  or g761 (n_794, wc53, n_448);
  not gc53 (wc53, n_449);
  or g762 (n_796, wc54, n_458);
  not gc54 (wc54, n_453);
  or g763 (n_799, wc55, n_454);
  not gc55 (wc55, n_455);
  or g764 (n_800, wc56, n_464);
  not gc56 (wc56, n_459);
  or g765 (n_803, wc57, n_460);
  not gc57 (wc57, n_461);
  or g766 (n_471, wc58, n_376);
  not gc58 (wc58, n_469);
  and g767 (n_483, wc59, n_480);
  not gc59 (wc59, n_475);
  and g768 (n_493, wc60, n_490);
  not gc60 (wc60, n_485);
  and g769 (n_503, wc61, n_500);
  not gc61 (wc61, n_495);
  and g770 (n_513, wc62, n_510);
  not gc62 (wc62, n_505);
  and g771 (n_523, wc63, n_520);
  not gc63 (wc63, n_515);
  and g772 (n_533, wc64, n_530);
  not gc64 (wc64, n_525);
  and g773 (n_543, wc65, n_540);
  not gc65 (wc65, n_535);
  or g774 (n_721, wc66, n_468);
  not gc66 (wc66, n_548);
  and g775 (n_620, wc67, n_498);
  not gc67 (wc67, n_565);
  and g776 (n_678, wc68, n_518);
  not gc68 (wc68, n_580);
  and g777 (n_650, wc69, n_538);
  not gc69 (wc69, n_595);
  or g778 (n_805, wc70, n_468);
  not gc70 (wc70, n_465);
  and g779 (n_556, wc71, n_383);
  not gc71 (wc71, n_476);
  and g780 (n_560, wc72, n_482);
  not gc72 (wc72, n_483);
  and g781 (n_613, wc73, n_395);
  not gc73 (wc73, n_486);
  and g782 (n_562, wc74, n_492);
  not gc74 (wc74, n_493);
  and g783 (n_570, wc75, n_407);
  not gc75 (wc75, n_496);
  and g784 (n_574, wc76, n_502);
  not gc76 (wc76, n_503);
  and g785 (n_671, wc77, n_419);
  not gc77 (wc77, n_506);
  and g786 (n_577, wc78, n_512);
  not gc78 (wc78, n_513);
  and g787 (n_585, wc79, n_429);
  not gc79 (wc79, n_516);
  and g788 (n_589, wc80, n_522);
  not gc80 (wc80, n_523);
  and g789 (n_638, wc81, n_441);
  not gc81 (wc81, n_526);
  and g790 (n_592, wc82, n_532);
  not gc82 (wc82, n_533);
  and g791 (n_600, wc83, n_453);
  not gc83 (wc83, n_536);
  and g792 (n_604, wc84, n_542);
  not gc84 (wc84, n_543);
  and g793 (n_723, wc85, n_465);
  not gc85 (wc85, n_546);
  or g794 (n_685, wc86, n_440);
  not gc86 (wc86, n_632);
  or g795 (n_693, n_637, wc87);
  not gc87 (wc87, n_632);
  or g796 (n_697, wc88, n_595);
  not gc88 (wc88, n_632);
  or g797 (n_808, wc89, n_466);
  not gc89 (wc89, n_467);
  or g798 (n_552, wc90, n_382);
  not gc90 (wc90, n_550);
  or g799 (n_557, n_554, wc91);
  not gc91 (wc91, n_550);
  or g800 (n_561, n_558, wc92);
  not gc92 (wc92, n_550);
  and g801 (n_567, wc93, n_498);
  not gc93 (wc93, n_562);
  and g802 (n_582, wc94, n_518);
  not gc94 (wc94, n_577);
  and g803 (n_597, wc95, n_538);
  not gc95 (wc95, n_592);
  and g804 (n_618, wc96, n_401);
  not gc96 (wc96, n_563);
  and g805 (n_621, wc97, n_495);
  not gc97 (wc97, n_567);
  and g806 (n_624, n_570, wc98);
  not gc98 (wc98, n_571);
  and g807 (n_627, n_574, wc99);
  not gc99 (wc99, n_575);
  and g808 (n_676, wc100, n_425);
  not gc100 (wc100, n_578);
  and g809 (n_679, wc101, n_515);
  not gc101 (wc101, n_582);
  and g810 (n_682, n_585, wc102);
  not gc102 (wc102, n_586);
  and g811 (n_629, n_589, wc103);
  not gc103 (wc103, n_590);
  and g812 (n_647, wc104, n_447);
  not gc104 (wc104, n_593);
  and g813 (n_652, wc105, n_535);
  not gc105 (wc105, n_597);
  and g814 (n_657, n_600, wc106);
  not gc106 (wc106, n_601);
  and g815 (n_662, n_604, wc107);
  not gc107 (wc107, n_605);
  or g816 (n_609, wc108, n_394);
  not gc108 (wc108, n_607);
  or g817 (n_614, n_611, wc109);
  not gc109 (wc109, n_607);
  or g818 (n_616, wc110, n_565);
  not gc110 (wc110, n_607);
  and g819 (n_635, wc111, n_528);
  not gc111 (wc111, n_629);
  and g820 (n_648, wc112, n_645);
  not gc112 (wc112, n_629);
  and g821 (n_653, wc113, n_650);
  not gc113 (wc113, n_629);
  and g822 (n_658, wc114, n_655);
  not gc114 (wc114, n_629);
  and g823 (n_663, wc115, n_660);
  not gc115 (wc115, n_629);
  and g824 (n_687, wc116, n_435);
  not gc116 (wc116, n_630);
  and g825 (n_691, wc117, n_525);
  not gc117 (wc117, n_635);
  and g826 (n_695, n_638, wc118);
  not gc118 (wc118, n_639);
  and g827 (n_699, n_592, wc119);
  not gc119 (wc119, n_642);
  and g828 (n_703, wc120, n_647);
  not gc120 (wc120, n_648);
  and g829 (n_707, wc121, n_652);
  not gc121 (wc121, n_653);
  and g830 (n_711, wc122, n_657);
  not gc122 (wc122, n_658);
  and g831 (n_715, wc123, n_662);
  not gc123 (wc123, n_663);
  or g832 (n_667, wc124, n_418);
  not gc124 (wc124, n_665);
  or g833 (n_672, n_669, wc125);
  not gc125 (wc125, n_665);
  or g834 (n_674, wc126, n_580);
  not gc126 (wc126, n_665);
  or g835 (n_688, n_685, wc127);
  not gc127 (wc127, n_665);
  or g836 (n_692, n_689, wc128);
  not gc128 (wc128, n_665);
  or g837 (n_696, n_693, wc129);
  not gc129 (wc129, n_665);
  or g838 (n_700, n_697, wc130);
  not gc130 (wc130, n_665);
  or g839 (n_704, n_701, wc131);
  not gc131 (wc131, n_665);
  or g840 (n_708, n_705, wc132);
  not gc132 (wc132, n_665);
  or g841 (n_712, n_709, wc133);
  not gc133 (wc133, n_665);
  or g842 (n_716, n_713, wc134);
  not gc134 (wc134, n_665);
  or g843 (n_719, wc135, n_464);
  not gc135 (wc135, n_717);
  or g844 (n_724, n_721, wc136);
  not gc136 (wc136, n_717);
endmodule

module csa_tree_add_252_40_group_16906_GENERIC(in_0, in_1, in_2, out_0);
  input [36:0] in_0, in_1;
  input [34:0] in_2;
  output [35:0] out_0;
  wire [36:0] in_0, in_1;
  wire [34:0] in_2;
  wire [35:0] out_0;
  csa_tree_add_252_40_group_16906_GENERIC_REAL g1(.in_0 ({in_0[36],
       in_0[32], in_0[32], in_0[32], in_0[32:0]}), .in_1 ({in_1[36],
       in_1[32], in_1[32], in_1[32], in_1[32:0]}), .in_2 ({in_2[33],
       in_2[33:0]}), .out_0 (out_0));
endmodule

module csa_tree_add_324_40_group_16916_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [22:0] in_0, in_1;
  input [20:0] in_2;
  output [21:0] out_0;
  wire [22:0] in_0, in_1;
  wire [20:0] in_2;
  wire [21:0] out_0;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_216;
  wire n_223, n_224, n_225, n_226, n_227, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_236, n_237, n_238, n_239, n_240;
  wire n_242, n_243, n_244, n_245, n_246, n_248, n_249, n_250;
  wire n_251, n_252, n_254, n_255, n_256, n_257, n_258, n_260;
  wire n_261, n_262, n_264, n_265, n_266, n_267, n_268, n_270;
  wire n_271, n_272, n_273, n_274, n_276, n_277, n_278, n_279;
  wire n_280, n_282, n_283, n_284, n_285, n_286, n_287, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_296, n_298, n_300;
  wire n_301, n_303, n_304, n_306, n_308, n_310, n_311, n_313;
  wire n_314, n_316, n_318, n_320, n_321, n_323, n_324, n_326;
  wire n_328, n_330, n_331, n_333, n_335, n_336, n_337, n_339;
  wire n_340, n_341, n_343, n_344, n_345, n_346, n_348, n_350;
  wire n_352, n_353, n_354, n_356, n_357, n_358, n_360, n_361;
  wire n_363, n_364, n_366, n_367, n_368, n_370, n_371, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381;
  wire n_382, n_383, n_384, n_385, n_386, n_388, n_389, n_390;
  wire n_392, n_393, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_402, n_403, n_404, n_406, n_407, n_408, n_409, n_411;
  wire n_412, n_413, n_415, n_416, n_417, n_418, n_420, n_421;
  wire n_423, n_424, n_426, n_427, n_428, n_429, n_431, n_432;
  wire n_433, n_435, n_436, n_437, n_438, n_440, n_441, n_443;
  wire n_444, n_446, n_447, n_448;
  xor g25 (n_132, in_0[1], in_2[1]);
  and g2 (n_109, in_0[1], in_2[1]);
  xor g26 (n_141, in_0[2], in_2[2]);
  xor g27 (n_131, n_141, in_1[2]);
  nand g3 (n_142, in_0[2], in_2[2]);
  nand g28 (n_143, in_1[2], in_2[2]);
  nand g29 (n_144, in_0[2], in_1[2]);
  nand g30 (n_108, n_142, n_143, n_144);
  xor g31 (n_145, in_0[3], in_2[3]);
  xor g32 (n_130, n_145, in_1[3]);
  nand g33 (n_146, in_0[3], in_2[3]);
  nand g4 (n_147, in_1[3], in_2[3]);
  nand g34 (n_148, in_0[3], in_1[3]);
  nand g35 (n_107, n_146, n_147, n_148);
  xor g36 (n_149, in_0[4], in_2[4]);
  xor g37 (n_129, n_149, in_1[4]);
  nand g38 (n_150, in_0[4], in_2[4]);
  nand g39 (n_151, in_1[4], in_2[4]);
  nand g5 (n_152, in_0[4], in_1[4]);
  nand g40 (n_106, n_150, n_151, n_152);
  xor g41 (n_153, in_0[5], in_2[5]);
  xor g42 (n_128, n_153, in_1[5]);
  nand g43 (n_154, in_0[5], in_2[5]);
  nand g44 (n_155, in_1[5], in_2[5]);
  nand g45 (n_156, in_0[5], in_1[5]);
  nand g6 (n_105, n_154, n_155, n_156);
  xor g46 (n_157, in_0[6], in_2[6]);
  xor g47 (n_127, n_157, in_1[6]);
  nand g48 (n_158, in_0[6], in_2[6]);
  nand g49 (n_159, in_1[6], in_2[6]);
  nand g50 (n_160, in_0[6], in_1[6]);
  nand g51 (n_104, n_158, n_159, n_160);
  xor g52 (n_133, in_0[7], in_2[7]);
  xor g53 (n_126, n_133, in_1[7]);
  nand g54 (n_134, in_0[7], in_2[7]);
  nand g55 (n_161, in_1[7], in_2[7]);
  nand g56 (n_162, in_0[7], in_1[7]);
  nand g57 (n_103, n_134, n_161, n_162);
  xor g58 (n_163, in_0[8], in_2[8]);
  xor g59 (n_125, n_163, in_1[8]);
  nand g60 (n_164, in_0[8], in_2[8]);
  nand g61 (n_165, in_1[8], in_2[8]);
  nand g62 (n_166, in_0[8], in_1[8]);
  nand g63 (n_102, n_164, n_165, n_166);
  xor g64 (n_167, in_0[9], in_2[9]);
  xor g65 (n_124, n_167, in_1[9]);
  nand g66 (n_168, in_0[9], in_2[9]);
  nand g67 (n_169, in_1[9], in_2[9]);
  nand g68 (n_170, in_0[9], in_1[9]);
  nand g69 (n_101, n_168, n_169, n_170);
  xor g70 (n_171, in_0[10], in_2[10]);
  xor g71 (n_123, n_171, in_1[10]);
  nand g72 (n_172, in_0[10], in_2[10]);
  nand g73 (n_173, in_1[10], in_2[10]);
  nand g74 (n_174, in_0[10], in_1[10]);
  nand g75 (n_100, n_172, n_173, n_174);
  xor g76 (n_175, in_0[11], in_2[11]);
  xor g77 (n_122, n_175, in_1[11]);
  nand g78 (n_176, in_0[11], in_2[11]);
  nand g79 (n_177, in_1[11], in_2[11]);
  nand g80 (n_178, in_0[11], in_1[11]);
  nand g81 (n_99, n_176, n_177, n_178);
  xor g82 (n_179, in_0[12], in_2[12]);
  xor g83 (n_121, n_179, in_1[12]);
  nand g84 (n_180, in_0[12], in_2[12]);
  nand g85 (n_181, in_1[12], in_2[12]);
  nand g86 (n_182, in_0[12], in_1[12]);
  nand g87 (n_98, n_180, n_181, n_182);
  xor g88 (n_183, in_0[13], in_2[13]);
  xor g89 (n_120, n_183, in_1[13]);
  nand g90 (n_184, in_0[13], in_2[13]);
  nand g91 (n_185, in_1[13], in_2[13]);
  nand g92 (n_186, in_0[13], in_1[13]);
  nand g93 (n_97, n_184, n_185, n_186);
  xor g94 (n_187, in_0[14], in_2[14]);
  xor g95 (n_119, n_187, in_1[14]);
  nand g96 (n_188, in_0[14], in_2[14]);
  nand g97 (n_189, in_1[14], in_2[14]);
  nand g98 (n_190, in_0[14], in_1[14]);
  nand g99 (n_96, n_188, n_189, n_190);
  xor g100 (n_191, in_0[15], in_2[15]);
  xor g101 (n_118, n_191, in_1[15]);
  nand g102 (n_192, in_0[15], in_2[15]);
  nand g103 (n_193, in_1[15], in_2[15]);
  nand g104 (n_194, in_0[15], in_1[15]);
  nand g105 (n_95, n_192, n_193, n_194);
  xor g106 (n_195, in_0[16], in_2[16]);
  xor g107 (n_117, n_195, in_1[16]);
  nand g108 (n_196, in_0[16], in_2[16]);
  nand g109 (n_197, in_1[16], in_2[16]);
  nand g110 (n_198, in_0[16], in_1[16]);
  nand g111 (n_94, n_196, n_197, n_198);
  xor g112 (n_199, in_0[17], in_2[17]);
  xor g113 (n_116, n_199, in_1[17]);
  nand g114 (n_200, in_0[17], in_2[17]);
  nand g115 (n_201, in_1[17], in_2[17]);
  nand g116 (n_202, in_0[17], in_1[17]);
  nand g117 (n_93, n_200, n_201, n_202);
  xor g118 (n_203, in_0[18], in_2[18]);
  xor g119 (n_115, n_203, in_1[18]);
  nand g120 (n_204, in_0[18], in_2[18]);
  nand g121 (n_205, in_1[18], in_2[18]);
  nand g122 (n_206, in_0[18], in_1[18]);
  nand g123 (n_92, n_204, n_205, n_206);
  xor g124 (n_207, in_0[19], in_2[19]);
  xor g125 (n_114, n_207, in_1[19]);
  nand g126 (n_208, in_0[19], in_2[19]);
  nand g127 (n_209, in_1[19], in_2[19]);
  nand g128 (n_210, in_0[19], in_1[19]);
  nand g129 (n_91, n_208, n_209, n_210);
  nand g137 (n_90, n_212, n_213, n_214);
  xor g141 (n_112, n_216, in_0[20]);
  xor g148 (n_448, in_2[0], in_1[0]);
  nand g149 (n_223, in_2[0], in_1[0]);
  nand g150 (n_224, in_2[0], in_0[0]);
  nand g7 (n_225, in_1[0], in_0[0]);
  nand g8 (n_227, n_223, n_224, n_225);
  nor g9 (n_226, in_1[1], n_132);
  nand g10 (n_229, in_1[1], n_132);
  nor g11 (n_236, n_109, n_131);
  nand g12 (n_231, n_109, n_131);
  nor g13 (n_232, n_108, n_130);
  nand g14 (n_233, n_108, n_130);
  nor g15 (n_242, n_107, n_129);
  nand g16 (n_237, n_107, n_129);
  nor g17 (n_238, n_106, n_128);
  nand g18 (n_239, n_106, n_128);
  nor g19 (n_248, n_105, n_127);
  nand g20 (n_243, n_105, n_127);
  nor g21 (n_244, n_104, n_126);
  nand g22 (n_245, n_104, n_126);
  nor g23 (n_254, n_103, n_125);
  nand g24 (n_249, n_103, n_125);
  nor g151 (n_250, n_102, n_124);
  nand g152 (n_251, n_102, n_124);
  nor g153 (n_260, n_101, n_123);
  nand g154 (n_255, n_101, n_123);
  nor g155 (n_256, n_100, n_122);
  nand g156 (n_257, n_100, n_122);
  nor g157 (n_264, n_99, n_121);
  nand g158 (n_110, n_99, n_121);
  nor g159 (n_111, n_98, n_120);
  nand g160 (n_261, n_98, n_120);
  nor g161 (n_270, n_97, n_119);
  nand g162 (n_265, n_97, n_119);
  nor g163 (n_266, n_96, n_118);
  nand g164 (n_267, n_96, n_118);
  nor g165 (n_276, n_95, n_117);
  nand g166 (n_271, n_95, n_117);
  nor g167 (n_272, n_94, n_116);
  nand g168 (n_273, n_94, n_116);
  nor g169 (n_282, n_93, n_115);
  nand g170 (n_277, n_93, n_115);
  nor g171 (n_278, n_92, n_114);
  nand g172 (n_279, n_92, n_114);
  nor g173 (n_286, n_91, n_113);
  nand g174 (n_283, n_91, n_113);
  nand g179 (n_287, n_229, n_230);
  nor g180 (n_234, n_231, n_232);
  nor g183 (n_290, n_236, n_232);
  nor g184 (n_240, n_237, n_238);
  nor g187 (n_296, n_242, n_238);
  nor g188 (n_246, n_243, n_244);
  nor g191 (n_298, n_248, n_244);
  nor g192 (n_252, n_249, n_250);
  nor g195 (n_306, n_254, n_250);
  nor g196 (n_258, n_255, n_256);
  nor g199 (n_308, n_260, n_256);
  nor g200 (n_262, n_110, n_111);
  nor g203 (n_316, n_264, n_111);
  nor g204 (n_268, n_265, n_266);
  nor g207 (n_318, n_270, n_266);
  nor g208 (n_274, n_271, n_272);
  nor g211 (n_326, n_276, n_272);
  nor g212 (n_280, n_277, n_278);
  nor g215 (n_328, n_282, n_278);
  nand g218 (n_402, n_231, n_289);
  nand g219 (n_292, n_290, n_287);
  nand g220 (n_333, n_291, n_292);
  nor g221 (n_294, n_248, n_293);
  nand g230 (n_341, n_296, n_298);
  nor g231 (n_304, n_260, n_303);
  nand g240 (n_348, n_306, n_308);
  nor g241 (n_314, n_270, n_313);
  nand g250 (n_356, n_316, n_318);
  nor g251 (n_324, n_282, n_323);
  nand g260 (n_363, n_326, n_328);
  nand g263 (n_406, n_237, n_335);
  nand g264 (n_336, n_296, n_333);
  nand g265 (n_408, n_293, n_336);
  nand g268 (n_411, n_339, n_340);
  nand g271 (n_364, n_343, n_344);
  nor g272 (n_346, n_264, n_345);
  nor g275 (n_374, n_264, n_348);
  nor g281 (n_354, n_352, n_345);
  nor g284 (n_380, n_348, n_352);
  nor g285 (n_358, n_356, n_345);
  nor g288 (n_383, n_348, n_356);
  nor g289 (n_361, n_286, n_360);
  nor g292 (n_396, n_286, n_363);
  nand g295 (n_415, n_249, n_366);
  nand g296 (n_367, n_306, n_364);
  nand g297 (n_417, n_303, n_367);
  nand g300 (n_420, n_370, n_371);
  nand g303 (n_423, n_345, n_373);
  nand g304 (n_376, n_374, n_364);
  nand g305 (n_426, n_375, n_376);
  nand g306 (n_379, n_377, n_364);
  nand g307 (n_428, n_378, n_379);
  nand g308 (n_382, n_380, n_364);
  nand g309 (n_431, n_381, n_382);
  nand g310 (n_385, n_383, n_364);
  nand g311 (n_386, n_384, n_385);
  nand g314 (n_435, n_271, n_388);
  nand g315 (n_389, n_326, n_386);
  nand g316 (n_437, n_323, n_389);
  nand g319 (n_440, n_392, n_393);
  nand g322 (n_443, n_360, n_395);
  nand g323 (n_398, n_396, n_386);
  nand g324 (n_446, n_397, n_398);
  xnor g326 (out_0[1], n_227, n_399);
  xnor g328 (out_0[2], n_287, n_400);
  xnor g331 (out_0[3], n_402, n_403);
  xnor g333 (out_0[4], n_333, n_404);
  xnor g336 (out_0[5], n_406, n_407);
  xnor g338 (out_0[6], n_408, n_409);
  xnor g341 (out_0[7], n_411, n_412);
  xnor g343 (out_0[8], n_364, n_413);
  xnor g346 (out_0[9], n_415, n_416);
  xnor g348 (out_0[10], n_417, n_418);
  xnor g351 (out_0[11], n_420, n_421);
  xnor g354 (out_0[12], n_423, n_424);
  xnor g357 (out_0[13], n_426, n_427);
  xnor g359 (out_0[14], n_428, n_429);
  xnor g362 (out_0[15], n_431, n_432);
  xnor g364 (out_0[16], n_386, n_433);
  xnor g367 (out_0[17], n_435, n_436);
  xnor g369 (out_0[18], n_437, n_438);
  xnor g372 (out_0[19], n_440, n_441);
  xnor g375 (out_0[20], n_443, n_444);
  xnor g378 (out_0[21], n_446, n_447);
  xor g379 (out_0[0], in_0[0], n_448);
  xnor g382 (n_211, in_1[20], in_2[20]);
  or g383 (n_212, in_2[20], wc);
  not gc (wc, in_1[20]);
  or g384 (n_213, in_0[20], in_2[20]);
  or g385 (n_214, wc0, in_0[20]);
  not gc0 (wc0, in_1[20]);
  xnor g386 (n_216, in_0[21], in_1[21]);
  xnor g387 (n_113, n_211, in_0[20]);
  or g388 (n_230, n_226, wc1);
  not gc1 (wc1, n_227);
  or g389 (n_399, wc2, n_226);
  not gc2 (wc2, n_229);
  and g390 (n_284, n_90, n_112);
  or g391 (n_285, n_90, n_112);
  and g392 (n_291, wc3, n_233);
  not gc3 (wc3, n_234);
  and g393 (n_293, wc4, n_239);
  not gc4 (wc4, n_240);
  and g394 (n_300, wc5, n_245);
  not gc5 (wc5, n_246);
  and g395 (n_303, wc6, n_251);
  not gc6 (wc6, n_252);
  and g396 (n_310, wc7, n_257);
  not gc7 (wc7, n_258);
  and g397 (n_313, wc8, n_261);
  not gc8 (wc8, n_262);
  and g398 (n_320, wc9, n_267);
  not gc9 (wc9, n_268);
  and g399 (n_323, wc10, n_273);
  not gc10 (wc10, n_274);
  and g400 (n_330, wc11, n_279);
  not gc11 (wc11, n_280);
  or g401 (n_337, wc12, n_248);
  not gc12 (wc12, n_296);
  or g402 (n_368, wc13, n_260);
  not gc13 (wc13, n_306);
  or g403 (n_352, wc14, n_270);
  not gc14 (wc14, n_316);
  or g404 (n_390, wc15, n_282);
  not gc15 (wc15, n_326);
  or g405 (n_400, wc16, n_236);
  not gc16 (wc16, n_231);
  or g406 (n_403, wc17, n_232);
  not gc17 (wc17, n_233);
  or g407 (n_404, wc18, n_242);
  not gc18 (wc18, n_237);
  or g408 (n_407, wc19, n_238);
  not gc19 (wc19, n_239);
  or g409 (n_409, wc20, n_248);
  not gc20 (wc20, n_243);
  or g410 (n_412, wc21, n_244);
  not gc21 (wc21, n_245);
  or g411 (n_413, wc22, n_254);
  not gc22 (wc22, n_249);
  or g412 (n_416, wc23, n_250);
  not gc23 (wc23, n_251);
  or g413 (n_418, wc24, n_260);
  not gc24 (wc24, n_255);
  or g414 (n_421, wc25, n_256);
  not gc25 (wc25, n_257);
  or g415 (n_424, wc26, n_264);
  not gc26 (wc26, n_110);
  or g416 (n_427, wc27, n_111);
  not gc27 (wc27, n_261);
  or g417 (n_429, wc28, n_270);
  not gc28 (wc28, n_265);
  or g418 (n_432, wc29, n_266);
  not gc29 (wc29, n_267);
  or g419 (n_433, wc30, n_276);
  not gc30 (wc30, n_271);
  or g420 (n_436, wc31, n_272);
  not gc31 (wc31, n_273);
  or g421 (n_438, wc32, n_282);
  not gc32 (wc32, n_277);
  or g422 (n_441, wc33, n_278);
  not gc33 (wc33, n_279);
  or g423 (n_289, wc34, n_236);
  not gc34 (wc34, n_287);
  and g424 (n_301, wc35, n_298);
  not gc35 (wc35, n_293);
  and g425 (n_311, wc36, n_308);
  not gc36 (wc36, n_303);
  and g426 (n_321, wc37, n_318);
  not gc37 (wc37, n_313);
  and g427 (n_331, wc38, n_328);
  not gc38 (wc38, n_323);
  and g428 (n_377, wc39, n_316);
  not gc39 (wc39, n_348);
  or g429 (n_444, wc40, n_286);
  not gc40 (wc40, n_283);
  and g430 (n_339, wc41, n_243);
  not gc41 (wc41, n_294);
  and g431 (n_343, wc42, n_300);
  not gc42 (wc42, n_301);
  and g432 (n_370, wc43, n_255);
  not gc43 (wc43, n_304);
  and g433 (n_345, wc44, n_310);
  not gc44 (wc44, n_311);
  and g434 (n_353, wc45, n_265);
  not gc45 (wc45, n_314);
  and g435 (n_357, wc46, n_320);
  not gc46 (wc46, n_321);
  and g436 (n_392, wc47, n_277);
  not gc47 (wc47, n_324);
  and g437 (n_360, wc48, n_330);
  not gc48 (wc48, n_331);
  or g438 (n_447, wc49, n_284);
  not gc49 (wc49, n_285);
  or g439 (n_335, wc50, n_242);
  not gc50 (wc50, n_333);
  or g440 (n_340, n_337, wc51);
  not gc51 (wc51, n_333);
  or g441 (n_344, n_341, wc52);
  not gc52 (wc52, n_333);
  and g442 (n_350, wc53, n_316);
  not gc53 (wc53, n_345);
  and g443 (n_375, wc54, n_110);
  not gc54 (wc54, n_346);
  and g444 (n_378, wc55, n_313);
  not gc55 (wc55, n_350);
  and g445 (n_381, n_353, wc56);
  not gc56 (wc56, n_354);
  and g446 (n_384, n_357, wc57);
  not gc57 (wc57, n_358);
  and g447 (n_397, wc58, n_283);
  not gc58 (wc58, n_361);
  or g448 (n_366, wc59, n_254);
  not gc59 (wc59, n_364);
  or g449 (n_371, n_368, wc60);
  not gc60 (wc60, n_364);
  or g450 (n_373, wc61, n_348);
  not gc61 (wc61, n_364);
  or g451 (n_388, wc62, n_276);
  not gc62 (wc62, n_386);
  or g452 (n_393, n_390, wc63);
  not gc63 (wc63, n_386);
  or g453 (n_395, wc64, n_363);
  not gc64 (wc64, n_386);
endmodule

module csa_tree_add_324_40_group_16916_GENERIC(in_0, in_1, in_2, out_0);
  input [22:0] in_0, in_1;
  input [20:0] in_2;
  output [21:0] out_0;
  wire [22:0] in_0, in_1;
  wire [20:0] in_2;
  wire [21:0] out_0;
  csa_tree_add_324_40_group_16916_GENERIC_REAL g1(.in_0 ({in_0[22],
       in_0[18], in_0[18], in_0[18], in_0[18:0]}), .in_1 ({in_1[22],
       in_1[18], in_1[18], in_1[18], in_1[18:0]}), .in_2 ({in_2[19],
       in_2[19:0]}), .out_0 (out_0));
endmodule

module csa_tree_add_399_40_group_16908_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  wire n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109;
  wire n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117;
  wire n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125;
  wire n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133;
  wire n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150, n_151, n_152, n_159, n_160, n_161, n_162, n_163;
  wire n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171;
  wire n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179;
  wire n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187;
  wire n_188, n_189, n_190, n_191, n_192, n_193, n_194, n_195;
  wire n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203;
  wire n_204, n_205, n_206, n_207, n_208, n_209, n_210, n_211;
  wire n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219;
  wire n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_227;
  wire n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_246, n_253, n_254, n_255, n_256, n_257, n_259;
  wire n_260, n_261, n_262, n_263, n_264, n_266, n_267, n_268;
  wire n_269, n_270, n_272, n_273, n_274, n_275, n_276, n_278;
  wire n_279, n_280, n_281, n_282, n_284, n_285, n_286, n_287;
  wire n_288, n_290, n_291, n_292, n_293, n_294, n_296, n_297;
  wire n_298, n_300, n_301, n_302, n_303, n_304, n_306, n_307;
  wire n_308, n_309, n_310, n_312, n_313, n_314, n_315, n_316;
  wire n_318, n_319, n_320, n_321, n_322, n_324, n_325, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_334, n_336, n_338;
  wire n_339, n_341, n_342, n_344, n_346, n_348, n_349, n_351;
  wire n_352, n_354, n_356, n_358, n_359, n_361, n_362, n_364;
  wire n_366, n_368, n_369, n_371, n_372, n_374, n_376, n_378;
  wire n_379, n_381, n_383, n_384, n_385, n_387, n_388, n_389;
  wire n_391, n_392, n_393, n_394, n_396, n_398, n_400, n_401;
  wire n_402, n_404, n_405, n_406, n_408, n_409, n_411, n_413;
  wire n_415, n_416, n_417, n_419, n_420, n_421, n_423, n_425;
  wire n_426, n_427, n_429, n_430, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_450, n_452, n_453;
  wire n_454, n_456, n_457, n_459, n_460, n_461, n_462, n_463;
  wire n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471;
  wire n_473, n_474, n_475, n_477, n_478, n_479, n_480, n_482;
  wire n_483, n_484, n_486, n_487, n_488, n_489, n_491, n_492;
  wire n_494, n_495, n_497, n_498, n_499, n_500, n_502, n_503;
  wire n_504, n_506, n_507, n_508, n_509, n_511, n_512, n_514;
  wire n_515, n_517, n_518, n_519, n_520, n_522, n_523, n_524;
  wire n_525, n_526;
  xor g28 (n_150, in_2[1], in_0[1]);
  and g2 (n_124, in_2[1], in_0[1]);
  xor g29 (n_159, in_2[2], in_0[2]);
  xor g30 (n_149, n_159, in_1[2]);
  nand g3 (n_160, in_2[2], in_0[2]);
  nand g31 (n_161, in_1[2], in_0[2]);
  nand g32 (n_162, in_2[2], in_1[2]);
  nand g33 (n_123, n_160, n_161, n_162);
  xor g34 (n_163, in_2[3], in_0[3]);
  xor g35 (n_148, n_163, in_1[3]);
  nand g36 (n_164, in_2[3], in_0[3]);
  nand g4 (n_165, in_1[3], in_0[3]);
  nand g37 (n_166, in_2[3], in_1[3]);
  nand g38 (n_122, n_164, n_165, n_166);
  xor g39 (n_167, in_2[4], in_0[4]);
  xor g40 (n_147, n_167, in_1[4]);
  nand g41 (n_168, in_2[4], in_0[4]);
  nand g42 (n_169, in_1[4], in_0[4]);
  nand g5 (n_170, in_2[4], in_1[4]);
  nand g43 (n_121, n_168, n_169, n_170);
  xor g44 (n_171, in_2[5], in_0[5]);
  xor g45 (n_146, n_171, in_1[5]);
  nand g46 (n_172, in_2[5], in_0[5]);
  nand g47 (n_173, in_1[5], in_0[5]);
  nand g48 (n_174, in_2[5], in_1[5]);
  nand g6 (n_120, n_172, n_173, n_174);
  xor g49 (n_175, in_2[6], in_0[6]);
  xor g50 (n_145, n_175, in_1[6]);
  nand g51 (n_176, in_2[6], in_0[6]);
  nand g52 (n_177, in_1[6], in_0[6]);
  nand g53 (n_178, in_2[6], in_1[6]);
  nand g54 (n_119, n_176, n_177, n_178);
  xor g55 (n_179, in_2[7], in_0[7]);
  xor g56 (n_144, n_179, in_1[7]);
  nand g57 (n_180, in_2[7], in_0[7]);
  nand g58 (n_181, in_1[7], in_0[7]);
  nand g59 (n_151, in_2[7], in_1[7]);
  nand g60 (n_118, n_180, n_181, n_151);
  xor g61 (n_152, in_2[8], in_0[8]);
  xor g62 (n_143, n_152, in_1[8]);
  nand g63 (n_182, in_2[8], in_0[8]);
  nand g64 (n_183, in_1[8], in_0[8]);
  nand g65 (n_184, in_2[8], in_1[8]);
  nand g66 (n_117, n_182, n_183, n_184);
  xor g67 (n_185, in_2[9], in_0[9]);
  xor g68 (n_142, n_185, in_1[9]);
  nand g69 (n_186, in_2[9], in_0[9]);
  nand g70 (n_187, in_1[9], in_0[9]);
  nand g71 (n_188, in_2[9], in_1[9]);
  nand g72 (n_116, n_186, n_187, n_188);
  xor g73 (n_189, in_2[10], in_0[10]);
  xor g74 (n_141, n_189, in_1[10]);
  nand g75 (n_190, in_2[10], in_0[10]);
  nand g76 (n_191, in_1[10], in_0[10]);
  nand g77 (n_192, in_2[10], in_1[10]);
  nand g78 (n_115, n_190, n_191, n_192);
  xor g79 (n_193, in_2[11], in_0[11]);
  xor g80 (n_140, n_193, in_1[11]);
  nand g81 (n_194, in_2[11], in_0[11]);
  nand g82 (n_195, in_1[11], in_0[11]);
  nand g83 (n_196, in_2[11], in_1[11]);
  nand g84 (n_114, n_194, n_195, n_196);
  xor g85 (n_197, in_2[12], in_0[12]);
  xor g86 (n_139, n_197, in_1[12]);
  nand g87 (n_198, in_2[12], in_0[12]);
  nand g88 (n_199, in_1[12], in_0[12]);
  nand g89 (n_200, in_2[12], in_1[12]);
  nand g90 (n_113, n_198, n_199, n_200);
  xor g91 (n_201, in_2[13], in_0[13]);
  xor g92 (n_138, n_201, in_1[13]);
  nand g93 (n_202, in_2[13], in_0[13]);
  nand g94 (n_203, in_1[13], in_0[13]);
  nand g95 (n_204, in_2[13], in_1[13]);
  nand g96 (n_112, n_202, n_203, n_204);
  xor g97 (n_205, in_2[14], in_0[14]);
  xor g98 (n_137, n_205, in_1[14]);
  nand g99 (n_206, in_2[14], in_0[14]);
  nand g100 (n_207, in_1[14], in_0[14]);
  nand g101 (n_208, in_2[14], in_1[14]);
  nand g102 (n_111, n_206, n_207, n_208);
  xor g103 (n_209, in_2[15], in_0[15]);
  xor g104 (n_136, n_209, in_1[15]);
  nand g105 (n_210, in_2[15], in_0[15]);
  nand g106 (n_211, in_1[15], in_0[15]);
  nand g107 (n_212, in_2[15], in_1[15]);
  nand g108 (n_110, n_210, n_211, n_212);
  xor g109 (n_213, in_2[16], in_0[16]);
  xor g110 (n_135, n_213, in_1[16]);
  nand g111 (n_214, in_2[16], in_0[16]);
  nand g112 (n_215, in_1[16], in_0[16]);
  nand g113 (n_216, in_2[16], in_1[16]);
  nand g114 (n_109, n_214, n_215, n_216);
  xor g115 (n_217, in_2[17], in_0[17]);
  xor g116 (n_134, n_217, in_1[17]);
  nand g117 (n_218, in_2[17], in_0[17]);
  nand g118 (n_219, in_1[17], in_0[17]);
  nand g119 (n_220, in_2[17], in_1[17]);
  nand g120 (n_108, n_218, n_219, n_220);
  xor g121 (n_221, in_2[18], in_0[18]);
  xor g122 (n_133, n_221, in_1[18]);
  nand g123 (n_222, in_2[18], in_0[18]);
  nand g124 (n_223, in_1[18], in_0[18]);
  nand g125 (n_224, in_2[18], in_1[18]);
  nand g126 (n_107, n_222, n_223, n_224);
  xor g127 (n_225, in_2[19], in_0[19]);
  xor g128 (n_132, n_225, in_1[19]);
  nand g129 (n_226, in_2[19], in_0[19]);
  nand g130 (n_227, in_1[19], in_0[19]);
  nand g131 (n_228, in_2[19], in_1[19]);
  nand g132 (n_131, n_226, n_227, n_228);
  xor g133 (n_229, in_2[20], in_1[20]);
  xor g134 (n_106, n_229, in_0[20]);
  nand g135 (n_230, in_2[20], in_1[20]);
  nand g136 (n_231, in_0[20], in_1[20]);
  nand g137 (n_232, in_2[20], in_0[20]);
  nand g138 (n_130, n_230, n_231, n_232);
  xor g139 (n_233, in_2[21], in_0[21]);
  xor g140 (n_105, n_233, in_1[21]);
  nand g141 (n_234, in_2[21], in_0[21]);
  nand g142 (n_235, in_1[21], in_0[21]);
  nand g143 (n_236, in_2[21], in_1[21]);
  nand g144 (n_104, n_234, n_235, n_236);
  xor g145 (n_237, in_2[22], in_0[22]);
  xor g146 (n_129, n_237, in_1[22]);
  nand g147 (n_238, in_2[22], in_0[22]);
  nand g148 (n_239, in_1[22], in_0[22]);
  nand g149 (n_240, in_2[22], in_1[22]);
  nand g150 (n_128, n_238, n_239, n_240);
  xor g153 (n_241, in_2[23], in_1[23]);
  xor g154 (n_103, n_241, in_0[23]);
  nand g155 (n_242, in_2[23], in_1[23]);
  nand g156 (n_243, in_0[23], in_1[23]);
  nand g157 (n_244, in_2[23], in_0[23]);
  nand g158 (n_127, n_242, n_243, n_244);
  xor g161 (n_246, in_2[23], in_0[24]);
  xor g162 (n_102, n_246, in_1[24]);
  xor g169 (n_526, in_0[0], in_1[0]);
  nand g170 (n_253, in_0[0], in_1[0]);
  nand g171 (n_254, in_0[0], in_2[0]);
  nand g7 (n_255, in_1[0], in_2[0]);
  nand g8 (n_257, n_253, n_254, n_255);
  nor g9 (n_256, in_1[1], n_150);
  nand g10 (n_259, in_1[1], n_150);
  nor g11 (n_266, n_124, n_149);
  nand g12 (n_261, n_124, n_149);
  nor g13 (n_262, n_123, n_148);
  nand g14 (n_263, n_123, n_148);
  nor g15 (n_272, n_122, n_147);
  nand g16 (n_267, n_122, n_147);
  nor g17 (n_268, n_121, n_146);
  nand g18 (n_269, n_121, n_146);
  nor g19 (n_278, n_120, n_145);
  nand g20 (n_273, n_120, n_145);
  nor g21 (n_274, n_119, n_144);
  nand g22 (n_275, n_119, n_144);
  nor g23 (n_284, n_118, n_143);
  nand g24 (n_279, n_118, n_143);
  nor g25 (n_280, n_117, n_142);
  nand g26 (n_281, n_117, n_142);
  nor g27 (n_290, n_116, n_141);
  nand g172 (n_285, n_116, n_141);
  nor g173 (n_286, n_115, n_140);
  nand g174 (n_287, n_115, n_140);
  nor g175 (n_296, n_114, n_139);
  nand g176 (n_291, n_114, n_139);
  nor g177 (n_292, n_113, n_138);
  nand g178 (n_293, n_113, n_138);
  nor g179 (n_300, n_112, n_137);
  nand g180 (n_125, n_112, n_137);
  nor g181 (n_126, n_111, n_136);
  nand g182 (n_297, n_111, n_136);
  nor g183 (n_306, n_110, n_135);
  nand g184 (n_301, n_110, n_135);
  nor g185 (n_302, n_109, n_134);
  nand g186 (n_303, n_109, n_134);
  nor g187 (n_312, n_108, n_133);
  nand g188 (n_307, n_108, n_133);
  nor g189 (n_308, n_107, n_132);
  nand g190 (n_309, n_107, n_132);
  nor g191 (n_318, n_106, n_131);
  nand g192 (n_313, n_106, n_131);
  nor g193 (n_314, n_105, n_130);
  nand g194 (n_315, n_105, n_130);
  nor g195 (n_324, n_104, n_129);
  nand g196 (n_319, n_104, n_129);
  nor g197 (n_320, n_103, n_128);
  nand g198 (n_321, n_103, n_128);
  nand g203 (n_325, n_259, n_260);
  nor g204 (n_264, n_261, n_262);
  nor g207 (n_328, n_266, n_262);
  nor g208 (n_270, n_267, n_268);
  nor g211 (n_334, n_272, n_268);
  nor g212 (n_276, n_273, n_274);
  nor g215 (n_336, n_278, n_274);
  nor g216 (n_282, n_279, n_280);
  nor g219 (n_344, n_284, n_280);
  nor g220 (n_288, n_285, n_286);
  nor g223 (n_346, n_290, n_286);
  nor g224 (n_294, n_291, n_292);
  nor g227 (n_354, n_296, n_292);
  nor g228 (n_298, n_125, n_126);
  nor g231 (n_356, n_300, n_126);
  nor g232 (n_304, n_301, n_302);
  nor g235 (n_364, n_306, n_302);
  nor g236 (n_310, n_307, n_308);
  nor g239 (n_366, n_312, n_308);
  nor g240 (n_316, n_313, n_314);
  nor g243 (n_374, n_318, n_314);
  nor g244 (n_322, n_319, n_320);
  nor g247 (n_376, n_324, n_320);
  nand g250 (n_473, n_261, n_327);
  nand g251 (n_330, n_328, n_325);
  nand g252 (n_381, n_329, n_330);
  nor g253 (n_332, n_278, n_331);
  nand g262 (n_389, n_334, n_336);
  nor g263 (n_342, n_290, n_341);
  nand g272 (n_396, n_344, n_346);
  nor g273 (n_352, n_300, n_351);
  nand g282 (n_404, n_354, n_356);
  nor g283 (n_362, n_312, n_361);
  nand g292 (n_411, n_364, n_366);
  nor g293 (n_372, n_324, n_371);
  nand g302 (n_419, n_374, n_376);
  nand g305 (n_477, n_267, n_383);
  nand g306 (n_384, n_334, n_381);
  nand g307 (n_479, n_331, n_384);
  nand g310 (n_482, n_387, n_388);
  nand g313 (n_423, n_391, n_392);
  nor g314 (n_394, n_296, n_393);
  nor g317 (n_433, n_296, n_396);
  nor g323 (n_402, n_400, n_393);
  nor g326 (n_439, n_396, n_400);
  nor g327 (n_406, n_404, n_393);
  nor g330 (n_442, n_396, n_404);
  nor g331 (n_409, n_318, n_408);
  nor g334 (n_460, n_318, n_411);
  nor g340 (n_417, n_415, n_408);
  nor g343 (n_466, n_411, n_415);
  nor g344 (n_421, n_419, n_408);
  nor g347 (n_448, n_411, n_419);
  nand g350 (n_486, n_279, n_425);
  nand g351 (n_426, n_344, n_423);
  nand g352 (n_488, n_341, n_426);
  nand g355 (n_491, n_429, n_430);
  nand g358 (n_494, n_393, n_432);
  nand g359 (n_435, n_433, n_423);
  nand g360 (n_497, n_434, n_435);
  nand g361 (n_438, n_436, n_423);
  nand g362 (n_499, n_437, n_438);
  nand g363 (n_441, n_439, n_423);
  nand g364 (n_502, n_440, n_441);
  nand g365 (n_444, n_442, n_423);
  nand g366 (n_450, n_443, n_444);
  nand g370 (n_506, n_301, n_452);
  nand g371 (n_453, n_364, n_450);
  nand g372 (n_508, n_361, n_453);
  nand g375 (n_511, n_456, n_457);
  nand g378 (n_514, n_408, n_459);
  nand g379 (n_462, n_460, n_450);
  nand g380 (n_517, n_461, n_462);
  nand g381 (n_465, n_463, n_450);
  nand g382 (n_519, n_464, n_465);
  nand g383 (n_468, n_466, n_450);
  nand g384 (n_522, n_467, n_468);
  nand g385 (n_469, n_448, n_450);
  nand g386 (n_524, n_446, n_469);
  xnor g388 (out_0[1], n_257, n_470);
  xnor g390 (out_0[2], n_325, n_471);
  xnor g393 (out_0[3], n_473, n_474);
  xnor g395 (out_0[4], n_381, n_475);
  xnor g398 (out_0[5], n_477, n_478);
  xnor g400 (out_0[6], n_479, n_480);
  xnor g403 (out_0[7], n_482, n_483);
  xnor g405 (out_0[8], n_423, n_484);
  xnor g408 (out_0[9], n_486, n_487);
  xnor g410 (out_0[10], n_488, n_489);
  xnor g413 (out_0[11], n_491, n_492);
  xnor g416 (out_0[12], n_494, n_495);
  xnor g419 (out_0[13], n_497, n_498);
  xnor g421 (out_0[14], n_499, n_500);
  xnor g424 (out_0[15], n_502, n_503);
  xnor g426 (out_0[16], n_450, n_504);
  xnor g429 (out_0[17], n_506, n_507);
  xnor g431 (out_0[18], n_508, n_509);
  xnor g434 (out_0[19], n_511, n_512);
  xnor g437 (out_0[20], n_514, n_515);
  xnor g440 (out_0[21], n_517, n_518);
  xnor g442 (out_0[22], n_519, n_520);
  xnor g445 (out_0[23], n_522, n_523);
  xnor g447 (out_0[24], n_524, n_525);
  xor g448 (out_0[0], in_2[0], n_526);
  or g449 (n_260, n_256, wc);
  not gc (wc, n_257);
  or g450 (n_470, wc0, n_256);
  not gc0 (wc0, n_259);
  and g451 (n_329, wc1, n_263);
  not gc1 (wc1, n_264);
  and g452 (n_331, wc2, n_269);
  not gc2 (wc2, n_270);
  and g453 (n_338, wc3, n_275);
  not gc3 (wc3, n_276);
  and g454 (n_341, wc4, n_281);
  not gc4 (wc4, n_282);
  and g455 (n_348, wc5, n_287);
  not gc5 (wc5, n_288);
  and g456 (n_351, wc6, n_293);
  not gc6 (wc6, n_294);
  and g457 (n_358, wc7, n_297);
  not gc7 (wc7, n_298);
  and g458 (n_361, wc8, n_303);
  not gc8 (wc8, n_304);
  and g459 (n_368, wc9, n_309);
  not gc9 (wc9, n_310);
  and g460 (n_371, wc10, n_315);
  not gc10 (wc10, n_316);
  or g461 (n_385, wc11, n_278);
  not gc11 (wc11, n_334);
  or g462 (n_427, wc12, n_290);
  not gc12 (wc12, n_344);
  or g463 (n_400, wc13, n_300);
  not gc13 (wc13, n_354);
  or g464 (n_454, wc14, n_312);
  not gc14 (wc14, n_364);
  or g465 (n_415, wc15, n_324);
  not gc15 (wc15, n_374);
  or g466 (n_471, wc16, n_266);
  not gc16 (wc16, n_261);
  or g467 (n_474, wc17, n_262);
  not gc17 (wc17, n_263);
  or g468 (n_475, wc18, n_272);
  not gc18 (wc18, n_267);
  or g469 (n_478, wc19, n_268);
  not gc19 (wc19, n_269);
  or g470 (n_480, wc20, n_278);
  not gc20 (wc20, n_273);
  or g471 (n_483, wc21, n_274);
  not gc21 (wc21, n_275);
  or g472 (n_484, wc22, n_284);
  not gc22 (wc22, n_279);
  or g473 (n_487, wc23, n_280);
  not gc23 (wc23, n_281);
  or g474 (n_489, wc24, n_290);
  not gc24 (wc24, n_285);
  or g475 (n_492, wc25, n_286);
  not gc25 (wc25, n_287);
  or g476 (n_495, wc26, n_296);
  not gc26 (wc26, n_291);
  or g477 (n_498, wc27, n_292);
  not gc27 (wc27, n_293);
  or g478 (n_500, wc28, n_300);
  not gc28 (wc28, n_125);
  or g479 (n_503, wc29, n_126);
  not gc29 (wc29, n_297);
  or g480 (n_504, wc30, n_306);
  not gc30 (wc30, n_301);
  or g481 (n_507, wc31, n_302);
  not gc31 (wc31, n_303);
  or g482 (n_509, wc32, n_312);
  not gc32 (wc32, n_307);
  or g483 (n_512, wc33, n_308);
  not gc33 (wc33, n_309);
  or g484 (n_515, wc34, n_318);
  not gc34 (wc34, n_313);
  or g485 (n_518, wc35, n_314);
  not gc35 (wc35, n_315);
  or g486 (n_520, wc36, n_324);
  not gc36 (wc36, n_319);
  or g487 (n_327, wc37, n_266);
  not gc37 (wc37, n_325);
  and g488 (n_339, wc38, n_336);
  not gc38 (wc38, n_331);
  and g489 (n_349, wc39, n_346);
  not gc39 (wc39, n_341);
  and g490 (n_359, wc40, n_356);
  not gc40 (wc40, n_351);
  and g491 (n_369, wc41, n_366);
  not gc41 (wc41, n_361);
  and g492 (n_436, wc42, n_354);
  not gc42 (wc42, n_396);
  and g493 (n_463, wc43, n_374);
  not gc43 (wc43, n_411);
  and g494 (n_445, n_127, n_102);
  or g495 (n_447, n_127, n_102);
  and g496 (n_378, wc44, n_321);
  not gc44 (wc44, n_322);
  and g497 (n_387, wc45, n_273);
  not gc45 (wc45, n_332);
  and g498 (n_391, wc46, n_338);
  not gc46 (wc46, n_339);
  and g499 (n_429, wc47, n_285);
  not gc47 (wc47, n_342);
  and g500 (n_393, wc48, n_348);
  not gc48 (wc48, n_349);
  and g501 (n_401, wc49, n_125);
  not gc49 (wc49, n_352);
  and g502 (n_405, wc50, n_358);
  not gc50 (wc50, n_359);
  and g503 (n_456, wc51, n_307);
  not gc51 (wc51, n_362);
  and g504 (n_408, wc52, n_368);
  not gc52 (wc52, n_369);
  and g505 (n_416, wc53, n_319);
  not gc53 (wc53, n_372);
  or g506 (n_523, wc54, n_320);
  not gc54 (wc54, n_321);
  and g507 (n_379, wc55, n_376);
  not gc55 (wc55, n_371);
  or g508 (n_383, wc56, n_272);
  not gc56 (wc56, n_381);
  or g509 (n_388, n_385, wc57);
  not gc57 (wc57, n_381);
  or g510 (n_392, n_389, wc58);
  not gc58 (wc58, n_381);
  and g511 (n_398, wc59, n_354);
  not gc59 (wc59, n_393);
  and g512 (n_413, wc60, n_374);
  not gc60 (wc60, n_408);
  and g513 (n_420, wc61, n_378);
  not gc61 (wc61, n_379);
  and g514 (n_434, wc62, n_291);
  not gc62 (wc62, n_394);
  and g515 (n_437, wc63, n_351);
  not gc63 (wc63, n_398);
  and g516 (n_440, n_401, wc64);
  not gc64 (wc64, n_402);
  and g517 (n_443, n_405, wc65);
  not gc65 (wc65, n_406);
  and g518 (n_461, wc66, n_313);
  not gc66 (wc66, n_409);
  and g519 (n_464, wc67, n_371);
  not gc67 (wc67, n_413);
  and g520 (n_467, n_416, wc68);
  not gc68 (wc68, n_417);
  or g521 (n_525, wc69, n_445);
  not gc69 (wc69, n_447);
  or g522 (n_425, wc70, n_284);
  not gc70 (wc70, n_423);
  or g523 (n_430, n_427, wc71);
  not gc71 (wc71, n_423);
  or g524 (n_432, wc72, n_396);
  not gc72 (wc72, n_423);
  and g525 (n_446, n_420, wc73);
  not gc73 (wc73, n_421);
  or g526 (n_452, wc74, n_306);
  not gc74 (wc74, n_450);
  or g527 (n_457, n_454, wc75);
  not gc75 (wc75, n_450);
  or g528 (n_459, wc76, n_411);
  not gc76 (wc76, n_450);
endmodule

module csa_tree_add_399_40_group_16908_GENERIC(in_0, in_1, in_2, out_0);
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  csa_tree_add_399_40_group_16908_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_449_42_group_16912_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [28:0] in_0, in_1;
  input [26:0] in_2;
  output [27:0] out_0;
  wire [28:0] in_0, in_1;
  wire [26:0] in_2;
  wire [27:0] out_0;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_276, n_283, n_284, n_285, n_286;
  wire n_287, n_289, n_290, n_291, n_292, n_293, n_294, n_296;
  wire n_297, n_298, n_299, n_300, n_302, n_303, n_304, n_305;
  wire n_306, n_308, n_309, n_310, n_311, n_312, n_314, n_315;
  wire n_316, n_317, n_318, n_320, n_321, n_322, n_323, n_324;
  wire n_326, n_327, n_328, n_329, n_330, n_332, n_333, n_334;
  wire n_336, n_337, n_338, n_339, n_340, n_342, n_343, n_344;
  wire n_345, n_346, n_348, n_349, n_350, n_351, n_352, n_354;
  wire n_355, n_356, n_357, n_358, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_367, n_368, n_369, n_370, n_371, n_372;
  wire n_374, n_376, n_378, n_379, n_381, n_382, n_384, n_386;
  wire n_388, n_389, n_391, n_392, n_394, n_396, n_398, n_399;
  wire n_401, n_402, n_404, n_406, n_408, n_409, n_411, n_412;
  wire n_414, n_416, n_418, n_419, n_421, n_422, n_424, n_426;
  wire n_428, n_429, n_430, n_432, n_433, n_434, n_436, n_437;
  wire n_438, n_439, n_441, n_443, n_445, n_446, n_447, n_449;
  wire n_450, n_451, n_453, n_454, n_456, n_458, n_460, n_461;
  wire n_462, n_464, n_465, n_466, n_468, n_470, n_471, n_472;
  wire n_474, n_475, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_493, n_496, n_498, n_499, n_500, n_503, n_505;
  wire n_506, n_507, n_509, n_510, n_512, n_513, n_514, n_515;
  wire n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523;
  wire n_525, n_526, n_527, n_529, n_530, n_531, n_533, n_534;
  wire n_535, n_536, n_538, n_539, n_540, n_542, n_543, n_544;
  wire n_545, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_556, n_557, n_559, n_560, n_562, n_563, n_564, n_565;
  wire n_567, n_568, n_569, n_571, n_572, n_573, n_574, n_576;
  wire n_577, n_579, n_580, n_582, n_583, n_584, n_585, n_587;
  wire n_588, n_589, n_590, n_592, n_593, n_594, n_595, n_597;
  wire n_598, n_599;
  xor g31 (n_168, in_0[1], in_2[1]);
  and g2 (n_139, in_0[1], in_2[1]);
  xor g32 (n_177, in_0[2], in_2[2]);
  xor g33 (n_167, n_177, in_1[2]);
  nand g3 (n_178, in_0[2], in_2[2]);
  nand g34 (n_179, in_1[2], in_2[2]);
  nand g35 (n_180, in_0[2], in_1[2]);
  nand g36 (n_138, n_178, n_179, n_180);
  xor g37 (n_181, in_0[3], in_2[3]);
  xor g38 (n_166, n_181, in_1[3]);
  nand g39 (n_182, in_0[3], in_2[3]);
  nand g4 (n_183, in_1[3], in_2[3]);
  nand g40 (n_184, in_0[3], in_1[3]);
  nand g41 (n_137, n_182, n_183, n_184);
  xor g42 (n_185, in_0[4], in_2[4]);
  xor g43 (n_165, n_185, in_1[4]);
  nand g44 (n_186, in_0[4], in_2[4]);
  nand g45 (n_187, in_1[4], in_2[4]);
  nand g5 (n_188, in_0[4], in_1[4]);
  nand g46 (n_136, n_186, n_187, n_188);
  xor g47 (n_189, in_0[5], in_2[5]);
  xor g48 (n_164, n_189, in_1[5]);
  nand g49 (n_190, in_0[5], in_2[5]);
  nand g50 (n_191, in_1[5], in_2[5]);
  nand g51 (n_192, in_0[5], in_1[5]);
  nand g6 (n_135, n_190, n_191, n_192);
  xor g52 (n_193, in_0[6], in_2[6]);
  xor g53 (n_163, n_193, in_1[6]);
  nand g54 (n_194, in_0[6], in_2[6]);
  nand g55 (n_195, in_1[6], in_2[6]);
  nand g56 (n_196, in_0[6], in_1[6]);
  nand g57 (n_134, n_194, n_195, n_196);
  xor g58 (n_197, in_0[7], in_2[7]);
  xor g59 (n_162, n_197, in_1[7]);
  nand g60 (n_198, in_0[7], in_2[7]);
  nand g61 (n_199, in_1[7], in_2[7]);
  nand g62 (n_200, in_0[7], in_1[7]);
  nand g63 (n_133, n_198, n_199, n_200);
  xor g64 (n_201, in_0[8], in_2[8]);
  xor g65 (n_161, n_201, in_1[8]);
  nand g66 (n_202, in_0[8], in_2[8]);
  nand g67 (n_169, in_1[8], in_2[8]);
  nand g68 (n_170, in_0[8], in_1[8]);
  nand g69 (n_132, n_202, n_169, n_170);
  xor g70 (n_203, in_0[9], in_2[9]);
  xor g71 (n_160, n_203, in_1[9]);
  nand g72 (n_204, in_0[9], in_2[9]);
  nand g73 (n_205, in_1[9], in_2[9]);
  nand g74 (n_206, in_0[9], in_1[9]);
  nand g75 (n_131, n_204, n_205, n_206);
  xor g76 (n_207, in_0[10], in_2[10]);
  xor g77 (n_159, n_207, in_1[10]);
  nand g78 (n_208, in_0[10], in_2[10]);
  nand g79 (n_209, in_1[10], in_2[10]);
  nand g80 (n_210, in_0[10], in_1[10]);
  nand g81 (n_130, n_208, n_209, n_210);
  xor g82 (n_211, in_0[11], in_2[11]);
  xor g83 (n_158, n_211, in_1[11]);
  nand g84 (n_212, in_0[11], in_2[11]);
  nand g85 (n_213, in_1[11], in_2[11]);
  nand g86 (n_214, in_0[11], in_1[11]);
  nand g87 (n_129, n_212, n_213, n_214);
  xor g88 (n_215, in_0[12], in_2[12]);
  xor g89 (n_157, n_215, in_1[12]);
  nand g90 (n_216, in_0[12], in_2[12]);
  nand g91 (n_217, in_1[12], in_2[12]);
  nand g92 (n_218, in_0[12], in_1[12]);
  nand g93 (n_128, n_216, n_217, n_218);
  xor g94 (n_219, in_0[13], in_2[13]);
  xor g95 (n_156, n_219, in_1[13]);
  nand g96 (n_220, in_0[13], in_2[13]);
  nand g97 (n_221, in_1[13], in_2[13]);
  nand g98 (n_222, in_0[13], in_1[13]);
  nand g99 (n_127, n_220, n_221, n_222);
  xor g100 (n_223, in_0[14], in_2[14]);
  xor g101 (n_155, n_223, in_1[14]);
  nand g102 (n_224, in_0[14], in_2[14]);
  nand g103 (n_225, in_1[14], in_2[14]);
  nand g104 (n_226, in_0[14], in_1[14]);
  nand g105 (n_126, n_224, n_225, n_226);
  xor g106 (n_227, in_0[15], in_2[15]);
  xor g107 (n_154, n_227, in_1[15]);
  nand g108 (n_228, in_0[15], in_2[15]);
  nand g109 (n_229, in_1[15], in_2[15]);
  nand g110 (n_230, in_0[15], in_1[15]);
  nand g111 (n_125, n_228, n_229, n_230);
  xor g112 (n_231, in_0[16], in_2[16]);
  xor g113 (n_153, n_231, in_1[16]);
  nand g114 (n_232, in_0[16], in_2[16]);
  nand g115 (n_233, in_1[16], in_2[16]);
  nand g116 (n_234, in_0[16], in_1[16]);
  nand g117 (n_124, n_232, n_233, n_234);
  xor g118 (n_235, in_0[17], in_2[17]);
  xor g119 (n_152, n_235, in_1[17]);
  nand g120 (n_236, in_0[17], in_2[17]);
  nand g121 (n_237, in_1[17], in_2[17]);
  nand g122 (n_238, in_0[17], in_1[17]);
  nand g123 (n_123, n_236, n_237, n_238);
  xor g124 (n_239, in_0[18], in_2[18]);
  xor g125 (n_151, n_239, in_1[18]);
  nand g126 (n_240, in_0[18], in_2[18]);
  nand g127 (n_241, in_1[18], in_2[18]);
  nand g128 (n_242, in_0[18], in_1[18]);
  nand g129 (n_122, n_240, n_241, n_242);
  xor g130 (n_243, in_0[19], in_2[19]);
  xor g131 (n_150, n_243, in_1[19]);
  nand g132 (n_244, in_0[19], in_2[19]);
  nand g133 (n_245, in_1[19], in_2[19]);
  nand g134 (n_246, in_0[19], in_1[19]);
  nand g135 (n_121, n_244, n_245, n_246);
  xor g136 (n_247, in_0[20], in_2[20]);
  xor g137 (n_149, n_247, in_1[20]);
  nand g138 (n_248, in_0[20], in_2[20]);
  nand g139 (n_249, in_1[20], in_2[20]);
  nand g140 (n_250, in_0[20], in_1[20]);
  nand g141 (n_120, n_248, n_249, n_250);
  xor g142 (n_251, in_0[21], in_2[21]);
  xor g143 (n_148, n_251, in_1[21]);
  nand g144 (n_252, in_0[21], in_2[21]);
  nand g145 (n_253, in_1[21], in_2[21]);
  nand g146 (n_254, in_0[21], in_1[21]);
  nand g147 (n_119, n_252, n_253, n_254);
  xor g148 (n_255, in_0[22], in_2[22]);
  xor g149 (n_147, n_255, in_1[22]);
  nand g150 (n_256, in_0[22], in_2[22]);
  nand g151 (n_257, in_1[22], in_2[22]);
  nand g152 (n_258, in_0[22], in_1[22]);
  nand g153 (n_118, n_256, n_257, n_258);
  xor g154 (n_259, in_0[23], in_2[23]);
  xor g155 (n_146, n_259, in_1[23]);
  nand g156 (n_260, in_0[23], in_2[23]);
  nand g157 (n_261, in_1[23], in_2[23]);
  nand g158 (n_262, in_0[23], in_1[23]);
  nand g159 (n_117, n_260, n_261, n_262);
  xor g160 (n_263, in_0[24], in_2[24]);
  xor g161 (n_145, n_263, in_1[24]);
  nand g162 (n_264, in_0[24], in_2[24]);
  nand g163 (n_265, in_1[24], in_2[24]);
  nand g164 (n_266, in_0[24], in_1[24]);
  nand g165 (n_116, n_264, n_265, n_266);
  xor g166 (n_267, in_0[25], in_2[25]);
  xor g167 (n_144, n_267, in_1[25]);
  nand g168 (n_268, in_0[25], in_2[25]);
  nand g169 (n_269, in_1[25], in_2[25]);
  nand g170 (n_270, in_0[25], in_1[25]);
  nand g171 (n_115, n_268, n_269, n_270);
  nand g179 (n_114, n_272, n_273, n_274);
  xor g183 (n_142, n_276, in_0[26]);
  xor g190 (n_599, in_2[0], in_1[0]);
  nand g191 (n_283, in_2[0], in_1[0]);
  nand g192 (n_284, in_2[0], in_0[0]);
  nand g7 (n_285, in_1[0], in_0[0]);
  nand g8 (n_287, n_283, n_284, n_285);
  nor g9 (n_286, in_1[1], n_168);
  nand g10 (n_289, in_1[1], n_168);
  nor g11 (n_296, n_139, n_167);
  nand g12 (n_291, n_139, n_167);
  nor g13 (n_292, n_138, n_166);
  nand g14 (n_293, n_138, n_166);
  nor g15 (n_302, n_137, n_165);
  nand g16 (n_297, n_137, n_165);
  nor g17 (n_298, n_136, n_164);
  nand g18 (n_299, n_136, n_164);
  nor g19 (n_308, n_135, n_163);
  nand g20 (n_303, n_135, n_163);
  nor g21 (n_304, n_134, n_162);
  nand g22 (n_305, n_134, n_162);
  nor g23 (n_314, n_133, n_161);
  nand g24 (n_309, n_133, n_161);
  nor g25 (n_310, n_132, n_160);
  nand g26 (n_311, n_132, n_160);
  nor g27 (n_320, n_131, n_159);
  nand g28 (n_315, n_131, n_159);
  nor g29 (n_316, n_130, n_158);
  nand g30 (n_317, n_130, n_158);
  nor g193 (n_326, n_129, n_157);
  nand g194 (n_321, n_129, n_157);
  nor g195 (n_322, n_128, n_156);
  nand g196 (n_323, n_128, n_156);
  nor g197 (n_332, n_127, n_155);
  nand g198 (n_327, n_127, n_155);
  nor g199 (n_328, n_126, n_154);
  nand g200 (n_329, n_126, n_154);
  nor g201 (n_336, n_125, n_153);
  nand g202 (n_140, n_125, n_153);
  nor g203 (n_141, n_124, n_152);
  nand g204 (n_333, n_124, n_152);
  nor g205 (n_342, n_123, n_151);
  nand g206 (n_337, n_123, n_151);
  nor g207 (n_338, n_122, n_150);
  nand g208 (n_339, n_122, n_150);
  nor g209 (n_348, n_121, n_149);
  nand g210 (n_343, n_121, n_149);
  nor g211 (n_344, n_120, n_148);
  nand g212 (n_345, n_120, n_148);
  nor g213 (n_354, n_119, n_147);
  nand g214 (n_349, n_119, n_147);
  nor g215 (n_350, n_118, n_146);
  nand g216 (n_351, n_118, n_146);
  nor g217 (n_360, n_117, n_145);
  nand g218 (n_355, n_117, n_145);
  nor g219 (n_356, n_116, n_144);
  nand g220 (n_357, n_116, n_144);
  nor g221 (n_364, n_115, n_143);
  nand g222 (n_361, n_115, n_143);
  nand g227 (n_365, n_289, n_290);
  nor g228 (n_294, n_291, n_292);
  nor g231 (n_368, n_296, n_292);
  nor g232 (n_300, n_297, n_298);
  nor g235 (n_374, n_302, n_298);
  nor g236 (n_306, n_303, n_304);
  nor g239 (n_376, n_308, n_304);
  nor g240 (n_312, n_309, n_310);
  nor g243 (n_384, n_314, n_310);
  nor g244 (n_318, n_315, n_316);
  nor g247 (n_386, n_320, n_316);
  nor g248 (n_324, n_321, n_322);
  nor g251 (n_394, n_326, n_322);
  nor g252 (n_330, n_327, n_328);
  nor g255 (n_396, n_332, n_328);
  nor g256 (n_334, n_140, n_141);
  nor g259 (n_404, n_336, n_141);
  nor g260 (n_340, n_337, n_338);
  nor g263 (n_406, n_342, n_338);
  nor g264 (n_346, n_343, n_344);
  nor g267 (n_414, n_348, n_344);
  nor g268 (n_352, n_349, n_350);
  nor g271 (n_416, n_354, n_350);
  nor g272 (n_358, n_355, n_356);
  nor g275 (n_424, n_360, n_356);
  nand g278 (n_538, n_291, n_367);
  nand g279 (n_370, n_368, n_365);
  nand g280 (n_426, n_369, n_370);
  nor g281 (n_372, n_308, n_371);
  nand g290 (n_434, n_374, n_376);
  nor g291 (n_382, n_320, n_381);
  nand g300 (n_441, n_384, n_386);
  nor g301 (n_392, n_332, n_391);
  nand g310 (n_449, n_394, n_396);
  nor g311 (n_402, n_342, n_401);
  nand g320 (n_456, n_404, n_406);
  nor g321 (n_412, n_354, n_411);
  nand g330 (n_464, n_414, n_416);
  nor g331 (n_422, n_364, n_421);
  nand g338 (n_542, n_297, n_428);
  nand g339 (n_429, n_374, n_426);
  nand g340 (n_544, n_371, n_429);
  nand g343 (n_547, n_432, n_433);
  nand g346 (n_468, n_436, n_437);
  nor g347 (n_439, n_326, n_438);
  nor g350 (n_478, n_326, n_441);
  nor g356 (n_447, n_445, n_438);
  nor g359 (n_484, n_441, n_445);
  nor g360 (n_451, n_449, n_438);
  nor g363 (n_487, n_441, n_449);
  nor g364 (n_454, n_348, n_453);
  nor g367 (n_513, n_348, n_456);
  nor g373 (n_462, n_460, n_453);
  nor g376 (n_519, n_456, n_460);
  nor g377 (n_466, n_464, n_453);
  nor g380 (n_493, n_456, n_464);
  nand g383 (n_551, n_309, n_470);
  nand g384 (n_471, n_384, n_468);
  nand g385 (n_553, n_381, n_471);
  nand g388 (n_556, n_474, n_475);
  nand g391 (n_559, n_438, n_477);
  nand g392 (n_480, n_478, n_468);
  nand g393 (n_562, n_479, n_480);
  nand g394 (n_483, n_481, n_468);
  nand g395 (n_564, n_482, n_483);
  nand g396 (n_486, n_484, n_468);
  nand g397 (n_567, n_485, n_486);
  nand g398 (n_489, n_487, n_468);
  nand g399 (n_503, n_488, n_489);
  nor g400 (n_491, n_360, n_490);
  nand g409 (n_527, n_424, n_493);
  nor g410 (n_500, n_498, n_490);
  nand g417 (n_571, n_140, n_505);
  nand g418 (n_506, n_404, n_503);
  nand g419 (n_573, n_401, n_506);
  nand g422 (n_576, n_509, n_510);
  nand g425 (n_579, n_453, n_512);
  nand g426 (n_515, n_513, n_503);
  nand g427 (n_582, n_514, n_515);
  nand g428 (n_518, n_516, n_503);
  nand g429 (n_584, n_517, n_518);
  nand g430 (n_521, n_519, n_503);
  nand g431 (n_587, n_520, n_521);
  nand g432 (n_522, n_493, n_503);
  nand g433 (n_589, n_490, n_522);
  nand g436 (n_592, n_525, n_526);
  nand g439 (n_594, n_529, n_530);
  nand g442 (n_597, n_533, n_534);
  xnor g444 (out_0[1], n_287, n_535);
  xnor g446 (out_0[2], n_365, n_536);
  xnor g449 (out_0[3], n_538, n_539);
  xnor g451 (out_0[4], n_426, n_540);
  xnor g454 (out_0[5], n_542, n_543);
  xnor g456 (out_0[6], n_544, n_545);
  xnor g459 (out_0[7], n_547, n_548);
  xnor g461 (out_0[8], n_468, n_549);
  xnor g464 (out_0[9], n_551, n_552);
  xnor g466 (out_0[10], n_553, n_554);
  xnor g469 (out_0[11], n_556, n_557);
  xnor g472 (out_0[12], n_559, n_560);
  xnor g475 (out_0[13], n_562, n_563);
  xnor g477 (out_0[14], n_564, n_565);
  xnor g480 (out_0[15], n_567, n_568);
  xnor g482 (out_0[16], n_503, n_569);
  xnor g485 (out_0[17], n_571, n_572);
  xnor g487 (out_0[18], n_573, n_574);
  xnor g490 (out_0[19], n_576, n_577);
  xnor g493 (out_0[20], n_579, n_580);
  xnor g496 (out_0[21], n_582, n_583);
  xnor g498 (out_0[22], n_584, n_585);
  xnor g501 (out_0[23], n_587, n_588);
  xnor g503 (out_0[24], n_589, n_590);
  xnor g506 (out_0[25], n_592, n_593);
  xnor g508 (out_0[26], n_594, n_595);
  xnor g511 (out_0[27], n_597, n_598);
  xor g512 (out_0[0], in_0[0], n_599);
  xnor g515 (n_271, in_1[26], in_2[26]);
  or g516 (n_272, in_2[26], wc);
  not gc (wc, in_1[26]);
  or g517 (n_273, in_0[26], in_2[26]);
  or g518 (n_274, wc0, in_0[26]);
  not gc0 (wc0, in_1[26]);
  xnor g519 (n_276, in_0[27], in_1[27]);
  xnor g520 (n_143, n_271, in_0[26]);
  or g521 (n_290, n_286, wc1);
  not gc1 (wc1, n_287);
  or g522 (n_535, wc2, n_286);
  not gc2 (wc2, n_289);
  and g523 (n_362, n_114, n_142);
  or g524 (n_363, n_114, n_142);
  and g525 (n_369, wc3, n_293);
  not gc3 (wc3, n_294);
  and g526 (n_371, wc4, n_299);
  not gc4 (wc4, n_300);
  and g527 (n_378, wc5, n_305);
  not gc5 (wc5, n_306);
  and g528 (n_381, wc6, n_311);
  not gc6 (wc6, n_312);
  and g529 (n_388, wc7, n_317);
  not gc7 (wc7, n_318);
  and g530 (n_391, wc8, n_323);
  not gc8 (wc8, n_324);
  and g531 (n_398, wc9, n_329);
  not gc9 (wc9, n_330);
  and g532 (n_401, wc10, n_333);
  not gc10 (wc10, n_334);
  and g533 (n_408, wc11, n_339);
  not gc11 (wc11, n_340);
  and g534 (n_411, wc12, n_345);
  not gc12 (wc12, n_346);
  and g535 (n_418, wc13, n_351);
  not gc13 (wc13, n_352);
  and g536 (n_421, wc14, n_357);
  not gc14 (wc14, n_358);
  or g537 (n_430, wc15, n_308);
  not gc15 (wc15, n_374);
  or g538 (n_472, wc16, n_320);
  not gc16 (wc16, n_384);
  or g539 (n_445, wc17, n_332);
  not gc17 (wc17, n_394);
  or g540 (n_507, wc18, n_342);
  not gc18 (wc18, n_404);
  or g541 (n_460, wc19, n_354);
  not gc19 (wc19, n_414);
  or g542 (n_536, wc20, n_296);
  not gc20 (wc20, n_291);
  or g543 (n_539, wc21, n_292);
  not gc21 (wc21, n_293);
  or g544 (n_540, wc22, n_302);
  not gc22 (wc22, n_297);
  or g545 (n_543, wc23, n_298);
  not gc23 (wc23, n_299);
  or g546 (n_545, wc24, n_308);
  not gc24 (wc24, n_303);
  or g547 (n_548, wc25, n_304);
  not gc25 (wc25, n_305);
  or g548 (n_549, wc26, n_314);
  not gc26 (wc26, n_309);
  or g549 (n_552, wc27, n_310);
  not gc27 (wc27, n_311);
  or g550 (n_554, wc28, n_320);
  not gc28 (wc28, n_315);
  or g551 (n_557, wc29, n_316);
  not gc29 (wc29, n_317);
  or g552 (n_560, wc30, n_326);
  not gc30 (wc30, n_321);
  or g553 (n_563, wc31, n_322);
  not gc31 (wc31, n_323);
  or g554 (n_565, wc32, n_332);
  not gc32 (wc32, n_327);
  or g555 (n_568, wc33, n_328);
  not gc33 (wc33, n_329);
  or g556 (n_569, wc34, n_336);
  not gc34 (wc34, n_140);
  or g557 (n_572, wc35, n_141);
  not gc35 (wc35, n_333);
  or g558 (n_574, wc36, n_342);
  not gc36 (wc36, n_337);
  or g559 (n_577, wc37, n_338);
  not gc37 (wc37, n_339);
  or g560 (n_580, wc38, n_348);
  not gc38 (wc38, n_343);
  or g561 (n_583, wc39, n_344);
  not gc39 (wc39, n_345);
  or g562 (n_585, wc40, n_354);
  not gc40 (wc40, n_349);
  or g563 (n_588, wc41, n_350);
  not gc41 (wc41, n_351);
  or g564 (n_590, wc42, n_360);
  not gc42 (wc42, n_355);
  or g565 (n_593, wc43, n_356);
  not gc43 (wc43, n_357);
  or g566 (n_367, wc44, n_296);
  not gc44 (wc44, n_365);
  and g567 (n_379, wc45, n_376);
  not gc45 (wc45, n_371);
  and g568 (n_389, wc46, n_386);
  not gc46 (wc46, n_381);
  and g569 (n_399, wc47, n_396);
  not gc47 (wc47, n_391);
  and g570 (n_409, wc48, n_406);
  not gc48 (wc48, n_401);
  and g571 (n_419, wc49, n_416);
  not gc49 (wc49, n_411);
  or g572 (n_498, wc50, n_364);
  not gc50 (wc50, n_424);
  and g573 (n_481, wc51, n_394);
  not gc51 (wc51, n_441);
  and g574 (n_516, wc52, n_414);
  not gc52 (wc52, n_456);
  or g575 (n_595, wc53, n_364);
  not gc53 (wc53, n_361);
  and g576 (n_432, wc54, n_303);
  not gc54 (wc54, n_372);
  and g577 (n_436, wc55, n_378);
  not gc55 (wc55, n_379);
  and g578 (n_474, wc56, n_315);
  not gc56 (wc56, n_382);
  and g579 (n_438, wc57, n_388);
  not gc57 (wc57, n_389);
  and g580 (n_446, wc58, n_327);
  not gc58 (wc58, n_392);
  and g581 (n_450, wc59, n_398);
  not gc59 (wc59, n_399);
  and g582 (n_509, wc60, n_337);
  not gc60 (wc60, n_402);
  and g583 (n_453, wc61, n_408);
  not gc61 (wc61, n_409);
  and g584 (n_461, wc62, n_349);
  not gc62 (wc62, n_412);
  and g585 (n_465, wc63, n_418);
  not gc63 (wc63, n_419);
  and g586 (n_499, wc64, n_361);
  not gc64 (wc64, n_422);
  or g587 (n_523, wc65, n_360);
  not gc65 (wc65, n_493);
  or g588 (n_598, wc66, n_362);
  not gc66 (wc66, n_363);
  or g589 (n_428, wc67, n_302);
  not gc67 (wc67, n_426);
  or g590 (n_433, n_430, wc68);
  not gc68 (wc68, n_426);
  or g591 (n_437, n_434, wc69);
  not gc69 (wc69, n_426);
  and g592 (n_443, wc70, n_394);
  not gc70 (wc70, n_438);
  and g593 (n_458, wc71, n_414);
  not gc71 (wc71, n_453);
  or g594 (n_531, n_498, wc72);
  not gc72 (wc72, n_493);
  and g595 (n_479, wc73, n_321);
  not gc73 (wc73, n_439);
  and g596 (n_482, wc74, n_391);
  not gc74 (wc74, n_443);
  and g597 (n_485, n_446, wc75);
  not gc75 (wc75, n_447);
  and g598 (n_488, n_450, wc76);
  not gc76 (wc76, n_451);
  and g599 (n_514, wc77, n_343);
  not gc77 (wc77, n_454);
  and g600 (n_517, wc78, n_411);
  not gc78 (wc78, n_458);
  and g601 (n_520, n_461, wc79);
  not gc79 (wc79, n_462);
  and g602 (n_490, n_465, wc80);
  not gc80 (wc80, n_466);
  or g603 (n_470, wc81, n_314);
  not gc81 (wc81, n_468);
  or g604 (n_475, n_472, wc82);
  not gc82 (wc82, n_468);
  or g605 (n_477, wc83, n_441);
  not gc83 (wc83, n_468);
  and g606 (n_496, wc84, n_424);
  not gc84 (wc84, n_490);
  and g607 (n_525, wc85, n_355);
  not gc85 (wc85, n_491);
  and g608 (n_529, wc86, n_421);
  not gc86 (wc86, n_496);
  and g609 (n_533, n_499, wc87);
  not gc87 (wc87, n_500);
  or g610 (n_505, wc88, n_336);
  not gc88 (wc88, n_503);
  or g611 (n_510, n_507, wc89);
  not gc89 (wc89, n_503);
  or g612 (n_512, wc90, n_456);
  not gc90 (wc90, n_503);
  or g613 (n_526, n_523, wc91);
  not gc91 (wc91, n_503);
  or g614 (n_530, n_527, wc92);
  not gc92 (wc92, n_503);
  or g615 (n_534, n_531, wc93);
  not gc93 (wc93, n_503);
endmodule

module csa_tree_add_449_42_group_16912_GENERIC(in_0, in_1, in_2, out_0);
  input [28:0] in_0, in_1;
  input [26:0] in_2;
  output [27:0] out_0;
  wire [28:0] in_0, in_1;
  wire [26:0] in_2;
  wire [27:0] out_0;
  csa_tree_add_449_42_group_16912_GENERIC_REAL g1(.in_0 ({in_0[28],
       in_0[23], in_0[23], in_0[23], in_0[23], in_0[23:0]}), .in_1
       ({in_1[28], in_1[23], in_1[23], in_1[23], in_1[23],
       in_1[23:0]}), .in_2 ({in_2[25], in_2[25:0]}), .out_0 (out_0));
endmodule

module csa_tree_add_559_42_group_16914_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [32:0] in_0, in_1;
  input [30:0] in_2;
  output [31:0] out_0;
  wire [32:0] in_0, in_1;
  wire [30:0] in_2;
  wire [31:0] out_0;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_235, n_236, n_237, n_238, n_239;
  wire n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_254, n_255;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_316, n_323, n_324, n_325, n_326;
  wire n_327, n_329, n_330, n_331, n_332, n_333, n_334, n_336;
  wire n_337, n_338, n_339, n_340, n_342, n_343, n_344, n_345;
  wire n_346, n_348, n_349, n_350, n_351, n_352, n_354, n_355;
  wire n_356, n_357, n_358, n_360, n_361, n_362, n_363, n_364;
  wire n_366, n_367, n_368, n_369, n_370, n_372, n_373, n_374;
  wire n_375, n_376, n_378, n_379, n_380, n_382, n_383, n_384;
  wire n_385, n_386, n_388, n_389, n_390, n_391, n_392, n_394;
  wire n_395, n_396, n_397, n_398, n_400, n_401, n_402, n_403;
  wire n_404, n_406, n_407, n_408, n_409, n_410, n_412, n_413;
  wire n_414, n_415, n_416, n_417, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_426, n_428, n_430, n_431, n_433, n_434;
  wire n_436, n_438, n_440, n_441, n_443, n_444, n_446, n_448;
  wire n_450, n_451, n_453, n_454, n_456, n_458, n_460, n_461;
  wire n_463, n_464, n_466, n_468, n_470, n_471, n_473, n_474;
  wire n_476, n_478, n_480, n_481, n_483, n_484, n_486, n_488;
  wire n_490, n_491, n_492, n_494, n_495, n_496, n_498, n_499;
  wire n_500, n_501, n_503, n_505, n_507, n_508, n_509, n_511;
  wire n_512, n_513, n_515, n_516, n_518, n_520, n_522, n_523;
  wire n_524, n_526, n_527, n_528, n_530, n_531, n_533, n_535;
  wire n_537, n_538, n_539, n_541, n_543, n_544, n_545, n_547;
  wire n_548, n_550, n_551, n_552, n_553, n_554, n_555, n_556;
  wire n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564;
  wire n_566, n_569, n_571, n_572, n_573, n_576, n_579, n_581;
  wire n_582, n_584, n_586, n_587, n_589, n_591, n_592, n_594;
  wire n_596, n_597, n_598, n_600, n_601, n_603, n_604, n_605;
  wire n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613;
  wire n_614, n_616, n_617, n_618, n_620, n_621, n_622, n_624;
  wire n_625, n_626, n_628, n_629, n_630, n_632, n_633, n_634;
  wire n_636, n_637, n_638, n_640, n_641, n_642, n_643, n_645;
  wire n_646, n_647, n_649, n_650, n_651, n_652, n_654, n_655;
  wire n_656, n_658, n_659, n_660, n_661, n_663, n_664, n_666;
  wire n_667, n_669, n_670, n_671, n_672, n_674, n_675, n_676;
  wire n_678, n_679, n_680, n_681, n_683, n_684, n_686, n_687;
  wire n_689, n_690, n_691, n_692, n_694, n_695, n_696, n_697;
  wire n_699, n_700, n_701, n_702, n_704, n_705, n_707, n_708;
  wire n_710, n_711, n_712, n_713, n_715, n_716, n_717;
  xor g35 (n_192, in_0[1], in_2[1]);
  and g2 (n_159, in_0[1], in_2[1]);
  xor g36 (n_201, in_0[2], in_2[2]);
  xor g37 (n_191, n_201, in_1[2]);
  nand g3 (n_202, in_0[2], in_2[2]);
  nand g38 (n_203, in_1[2], in_2[2]);
  nand g39 (n_204, in_0[2], in_1[2]);
  nand g40 (n_158, n_202, n_203, n_204);
  xor g41 (n_205, in_0[3], in_2[3]);
  xor g42 (n_190, n_205, in_1[3]);
  nand g43 (n_206, in_0[3], in_2[3]);
  nand g4 (n_207, in_1[3], in_2[3]);
  nand g44 (n_208, in_0[3], in_1[3]);
  nand g45 (n_157, n_206, n_207, n_208);
  xor g46 (n_209, in_0[4], in_2[4]);
  xor g47 (n_189, n_209, in_1[4]);
  nand g48 (n_210, in_0[4], in_2[4]);
  nand g49 (n_211, in_1[4], in_2[4]);
  nand g5 (n_212, in_0[4], in_1[4]);
  nand g50 (n_156, n_210, n_211, n_212);
  xor g51 (n_213, in_0[5], in_2[5]);
  xor g52 (n_188, n_213, in_1[5]);
  nand g53 (n_214, in_0[5], in_2[5]);
  nand g54 (n_215, in_1[5], in_2[5]);
  nand g55 (n_216, in_0[5], in_1[5]);
  nand g6 (n_155, n_214, n_215, n_216);
  xor g56 (n_217, in_0[6], in_2[6]);
  xor g57 (n_187, n_217, in_1[6]);
  nand g58 (n_218, in_0[6], in_2[6]);
  nand g59 (n_219, in_1[6], in_2[6]);
  nand g60 (n_220, in_0[6], in_1[6]);
  nand g61 (n_154, n_218, n_219, n_220);
  xor g62 (n_221, in_0[7], in_2[7]);
  xor g63 (n_186, n_221, in_1[7]);
  nand g64 (n_222, in_0[7], in_2[7]);
  nand g65 (n_223, in_1[7], in_2[7]);
  nand g66 (n_224, in_0[7], in_1[7]);
  nand g67 (n_153, n_222, n_223, n_224);
  xor g68 (n_225, in_0[8], in_2[8]);
  xor g69 (n_185, n_225, in_1[8]);
  nand g70 (n_226, in_0[8], in_2[8]);
  nand g71 (n_227, in_1[8], in_2[8]);
  nand g72 (n_228, in_0[8], in_1[8]);
  nand g73 (n_152, n_226, n_227, n_228);
  xor g74 (n_229, in_0[9], in_2[9]);
  xor g75 (n_184, n_229, in_1[9]);
  nand g76 (n_230, in_0[9], in_2[9]);
  nand g77 (n_193, in_1[9], in_2[9]);
  nand g78 (n_194, in_0[9], in_1[9]);
  nand g79 (n_151, n_230, n_193, n_194);
  xor g80 (n_231, in_0[10], in_2[10]);
  xor g81 (n_183, n_231, in_1[10]);
  nand g82 (n_232, in_0[10], in_2[10]);
  nand g83 (n_233, in_1[10], in_2[10]);
  nand g84 (n_234, in_0[10], in_1[10]);
  nand g85 (n_150, n_232, n_233, n_234);
  xor g86 (n_235, in_0[11], in_2[11]);
  xor g87 (n_182, n_235, in_1[11]);
  nand g88 (n_236, in_0[11], in_2[11]);
  nand g89 (n_237, in_1[11], in_2[11]);
  nand g90 (n_238, in_0[11], in_1[11]);
  nand g91 (n_149, n_236, n_237, n_238);
  xor g92 (n_239, in_0[12], in_2[12]);
  xor g93 (n_181, n_239, in_1[12]);
  nand g94 (n_240, in_0[12], in_2[12]);
  nand g95 (n_241, in_1[12], in_2[12]);
  nand g96 (n_242, in_0[12], in_1[12]);
  nand g97 (n_148, n_240, n_241, n_242);
  xor g98 (n_243, in_0[13], in_2[13]);
  xor g99 (n_180, n_243, in_1[13]);
  nand g100 (n_244, in_0[13], in_2[13]);
  nand g101 (n_245, in_1[13], in_2[13]);
  nand g102 (n_246, in_0[13], in_1[13]);
  nand g103 (n_147, n_244, n_245, n_246);
  xor g104 (n_247, in_0[14], in_2[14]);
  xor g105 (n_179, n_247, in_1[14]);
  nand g106 (n_248, in_0[14], in_2[14]);
  nand g107 (n_249, in_1[14], in_2[14]);
  nand g108 (n_250, in_0[14], in_1[14]);
  nand g109 (n_146, n_248, n_249, n_250);
  xor g110 (n_251, in_0[15], in_2[15]);
  xor g111 (n_178, n_251, in_1[15]);
  nand g112 (n_252, in_0[15], in_2[15]);
  nand g113 (n_253, in_1[15], in_2[15]);
  nand g114 (n_254, in_0[15], in_1[15]);
  nand g115 (n_145, n_252, n_253, n_254);
  xor g116 (n_255, in_0[16], in_2[16]);
  xor g117 (n_177, n_255, in_1[16]);
  nand g118 (n_256, in_0[16], in_2[16]);
  nand g119 (n_257, in_1[16], in_2[16]);
  nand g120 (n_258, in_0[16], in_1[16]);
  nand g121 (n_144, n_256, n_257, n_258);
  xor g122 (n_259, in_0[17], in_2[17]);
  xor g123 (n_176, n_259, in_1[17]);
  nand g124 (n_260, in_0[17], in_2[17]);
  nand g125 (n_261, in_1[17], in_2[17]);
  nand g126 (n_262, in_0[17], in_1[17]);
  nand g127 (n_143, n_260, n_261, n_262);
  xor g128 (n_263, in_0[18], in_2[18]);
  xor g129 (n_175, n_263, in_1[18]);
  nand g130 (n_264, in_0[18], in_2[18]);
  nand g131 (n_265, in_1[18], in_2[18]);
  nand g132 (n_266, in_0[18], in_1[18]);
  nand g133 (n_142, n_264, n_265, n_266);
  xor g134 (n_267, in_0[19], in_2[19]);
  xor g135 (n_174, n_267, in_1[19]);
  nand g136 (n_268, in_0[19], in_2[19]);
  nand g137 (n_269, in_1[19], in_2[19]);
  nand g138 (n_270, in_0[19], in_1[19]);
  nand g139 (n_141, n_268, n_269, n_270);
  xor g140 (n_271, in_0[20], in_2[20]);
  xor g141 (n_173, n_271, in_1[20]);
  nand g142 (n_272, in_0[20], in_2[20]);
  nand g143 (n_273, in_1[20], in_2[20]);
  nand g144 (n_274, in_0[20], in_1[20]);
  nand g145 (n_140, n_272, n_273, n_274);
  xor g146 (n_275, in_0[21], in_2[21]);
  xor g147 (n_172, n_275, in_1[21]);
  nand g148 (n_276, in_0[21], in_2[21]);
  nand g149 (n_277, in_1[21], in_2[21]);
  nand g150 (n_278, in_0[21], in_1[21]);
  nand g151 (n_139, n_276, n_277, n_278);
  xor g152 (n_279, in_0[22], in_2[22]);
  xor g153 (n_171, n_279, in_1[22]);
  nand g154 (n_280, in_0[22], in_2[22]);
  nand g155 (n_281, in_1[22], in_2[22]);
  nand g156 (n_282, in_0[22], in_1[22]);
  nand g157 (n_138, n_280, n_281, n_282);
  xor g158 (n_283, in_0[23], in_2[23]);
  xor g159 (n_170, n_283, in_1[23]);
  nand g160 (n_284, in_0[23], in_2[23]);
  nand g161 (n_285, in_1[23], in_2[23]);
  nand g162 (n_286, in_0[23], in_1[23]);
  nand g163 (n_137, n_284, n_285, n_286);
  xor g164 (n_287, in_0[24], in_2[24]);
  xor g165 (n_169, n_287, in_1[24]);
  nand g166 (n_288, in_0[24], in_2[24]);
  nand g167 (n_289, in_1[24], in_2[24]);
  nand g168 (n_290, in_0[24], in_1[24]);
  nand g169 (n_136, n_288, n_289, n_290);
  xor g170 (n_291, in_0[25], in_2[25]);
  xor g171 (n_168, n_291, in_1[25]);
  nand g172 (n_292, in_0[25], in_2[25]);
  nand g173 (n_293, in_1[25], in_2[25]);
  nand g174 (n_294, in_0[25], in_1[25]);
  nand g175 (n_135, n_292, n_293, n_294);
  xor g176 (n_295, in_0[26], in_2[26]);
  xor g177 (n_167, n_295, in_1[26]);
  nand g178 (n_296, in_0[26], in_2[26]);
  nand g179 (n_297, in_1[26], in_2[26]);
  nand g180 (n_298, in_0[26], in_1[26]);
  nand g181 (n_134, n_296, n_297, n_298);
  xor g182 (n_299, in_0[27], in_2[27]);
  xor g183 (n_166, n_299, in_1[27]);
  nand g184 (n_300, in_0[27], in_2[27]);
  nand g185 (n_301, in_1[27], in_2[27]);
  nand g186 (n_302, in_0[27], in_1[27]);
  nand g187 (n_133, n_300, n_301, n_302);
  xor g188 (n_303, in_0[28], in_2[28]);
  xor g189 (n_165, n_303, in_1[28]);
  nand g190 (n_304, in_0[28], in_2[28]);
  nand g191 (n_305, in_1[28], in_2[28]);
  nand g192 (n_306, in_0[28], in_1[28]);
  nand g193 (n_132, n_304, n_305, n_306);
  xor g194 (n_307, in_0[29], in_2[29]);
  xor g195 (n_164, n_307, in_1[29]);
  nand g196 (n_308, in_0[29], in_2[29]);
  nand g197 (n_309, in_1[29], in_2[29]);
  nand g198 (n_310, in_0[29], in_1[29]);
  nand g199 (n_131, n_308, n_309, n_310);
  nand g207 (n_130, n_312, n_313, n_314);
  xor g211 (n_162, n_316, in_0[30]);
  xor g218 (n_717, in_2[0], in_1[0]);
  nand g219 (n_323, in_2[0], in_1[0]);
  nand g220 (n_324, in_2[0], in_0[0]);
  nand g7 (n_325, in_1[0], in_0[0]);
  nand g8 (n_327, n_323, n_324, n_325);
  nor g9 (n_326, in_1[1], n_192);
  nand g10 (n_329, in_1[1], n_192);
  nor g11 (n_336, n_159, n_191);
  nand g12 (n_331, n_159, n_191);
  nor g13 (n_332, n_158, n_190);
  nand g14 (n_333, n_158, n_190);
  nor g15 (n_342, n_157, n_189);
  nand g16 (n_337, n_157, n_189);
  nor g17 (n_338, n_156, n_188);
  nand g18 (n_339, n_156, n_188);
  nor g19 (n_348, n_155, n_187);
  nand g20 (n_343, n_155, n_187);
  nor g21 (n_344, n_154, n_186);
  nand g22 (n_345, n_154, n_186);
  nor g23 (n_354, n_153, n_185);
  nand g24 (n_349, n_153, n_185);
  nor g25 (n_350, n_152, n_184);
  nand g26 (n_351, n_152, n_184);
  nor g27 (n_360, n_151, n_183);
  nand g28 (n_355, n_151, n_183);
  nor g29 (n_356, n_150, n_182);
  nand g30 (n_357, n_150, n_182);
  nor g31 (n_366, n_149, n_181);
  nand g32 (n_361, n_149, n_181);
  nor g33 (n_362, n_148, n_180);
  nand g34 (n_363, n_148, n_180);
  nor g221 (n_372, n_147, n_179);
  nand g222 (n_367, n_147, n_179);
  nor g223 (n_368, n_146, n_178);
  nand g224 (n_369, n_146, n_178);
  nor g225 (n_378, n_145, n_177);
  nand g226 (n_373, n_145, n_177);
  nor g227 (n_374, n_144, n_176);
  nand g228 (n_375, n_144, n_176);
  nor g229 (n_382, n_143, n_175);
  nand g230 (n_379, n_143, n_175);
  nor g231 (n_380, n_142, n_174);
  nand g232 (n_160, n_142, n_174);
  nor g233 (n_388, n_141, n_173);
  nand g234 (n_383, n_141, n_173);
  nor g235 (n_384, n_140, n_172);
  nand g236 (n_385, n_140, n_172);
  nor g237 (n_394, n_139, n_171);
  nand g238 (n_389, n_139, n_171);
  nor g239 (n_390, n_138, n_170);
  nand g240 (n_391, n_138, n_170);
  nor g241 (n_400, n_137, n_169);
  nand g242 (n_395, n_137, n_169);
  nor g243 (n_396, n_136, n_168);
  nand g244 (n_397, n_136, n_168);
  nor g245 (n_406, n_135, n_167);
  nand g246 (n_401, n_135, n_167);
  nor g247 (n_402, n_134, n_166);
  nand g248 (n_403, n_134, n_166);
  nor g249 (n_412, n_133, n_165);
  nand g250 (n_407, n_133, n_165);
  nor g251 (n_408, n_132, n_164);
  nand g252 (n_409, n_132, n_164);
  nor g253 (n_416, n_131, n_163);
  nand g254 (n_413, n_131, n_163);
  nand g259 (n_417, n_329, n_330);
  nor g260 (n_334, n_331, n_332);
  nor g263 (n_420, n_336, n_332);
  nor g264 (n_340, n_337, n_338);
  nor g267 (n_426, n_342, n_338);
  nor g268 (n_346, n_343, n_344);
  nor g271 (n_428, n_348, n_344);
  nor g272 (n_352, n_349, n_350);
  nor g275 (n_436, n_354, n_350);
  nor g276 (n_358, n_355, n_356);
  nor g279 (n_438, n_360, n_356);
  nor g280 (n_364, n_361, n_362);
  nor g283 (n_446, n_366, n_362);
  nor g284 (n_370, n_367, n_368);
  nor g287 (n_448, n_372, n_368);
  nor g288 (n_376, n_373, n_374);
  nor g291 (n_456, n_378, n_374);
  nor g292 (n_161, n_379, n_380);
  nor g295 (n_458, n_382, n_380);
  nor g296 (n_386, n_383, n_384);
  nor g299 (n_466, n_388, n_384);
  nor g300 (n_392, n_389, n_390);
  nor g303 (n_468, n_394, n_390);
  nor g304 (n_398, n_395, n_396);
  nor g307 (n_476, n_400, n_396);
  nor g308 (n_404, n_401, n_402);
  nor g311 (n_478, n_406, n_402);
  nor g312 (n_410, n_407, n_408);
  nor g315 (n_486, n_412, n_408);
  nand g318 (n_645, n_331, n_419);
  nand g319 (n_422, n_420, n_417);
  nand g320 (n_488, n_421, n_422);
  nor g321 (n_424, n_348, n_423);
  nand g330 (n_496, n_426, n_428);
  nor g331 (n_434, n_360, n_433);
  nand g340 (n_503, n_436, n_438);
  nor g341 (n_444, n_372, n_443);
  nand g350 (n_511, n_446, n_448);
  nor g351 (n_454, n_382, n_453);
  nand g360 (n_518, n_456, n_458);
  nor g361 (n_464, n_394, n_463);
  nand g370 (n_526, n_466, n_468);
  nor g371 (n_474, n_406, n_473);
  nand g380 (n_533, n_476, n_478);
  nor g381 (n_484, n_416, n_483);
  nand g388 (n_649, n_337, n_490);
  nand g389 (n_491, n_426, n_488);
  nand g390 (n_651, n_423, n_491);
  nand g393 (n_654, n_494, n_495);
  nand g396 (n_541, n_498, n_499);
  nor g397 (n_501, n_366, n_500);
  nor g400 (n_551, n_366, n_503);
  nor g406 (n_509, n_507, n_500);
  nor g409 (n_557, n_503, n_507);
  nor g410 (n_513, n_511, n_500);
  nor g413 (n_560, n_503, n_511);
  nor g414 (n_516, n_388, n_515);
  nor g417 (n_604, n_388, n_518);
  nor g423 (n_524, n_522, n_515);
  nor g426 (n_610, n_518, n_522);
  nor g427 (n_528, n_526, n_515);
  nor g430 (n_566, n_518, n_526);
  nor g431 (n_531, n_412, n_530);
  nor g434 (n_579, n_412, n_533);
  nor g440 (n_539, n_537, n_530);
  nor g443 (n_589, n_533, n_537);
  nand g446 (n_658, n_349, n_543);
  nand g447 (n_544, n_436, n_541);
  nand g448 (n_660, n_433, n_544);
  nand g451 (n_663, n_547, n_548);
  nand g454 (n_666, n_500, n_550);
  nand g455 (n_553, n_551, n_541);
  nand g456 (n_669, n_552, n_553);
  nand g457 (n_556, n_554, n_541);
  nand g458 (n_671, n_555, n_556);
  nand g459 (n_559, n_557, n_541);
  nand g460 (n_674, n_558, n_559);
  nand g461 (n_562, n_560, n_541);
  nand g462 (n_594, n_561, n_562);
  nor g463 (n_564, n_400, n_563);
  nand g472 (n_618, n_476, n_566);
  nor g473 (n_573, n_571, n_563);
  nor g478 (n_576, n_533, n_563);
  nand g487 (n_630, n_566, n_579);
  nand g492 (n_634, n_566, n_584);
  nand g497 (n_638, n_566, n_589);
  nand g500 (n_678, n_373, n_596);
  nand g501 (n_597, n_456, n_594);
  nand g502 (n_680, n_453, n_597);
  nand g505 (n_683, n_600, n_601);
  nand g508 (n_686, n_515, n_603);
  nand g509 (n_606, n_604, n_594);
  nand g510 (n_689, n_605, n_606);
  nand g511 (n_609, n_607, n_594);
  nand g512 (n_691, n_608, n_609);
  nand g513 (n_612, n_610, n_594);
  nand g514 (n_694, n_611, n_612);
  nand g515 (n_613, n_566, n_594);
  nand g516 (n_696, n_563, n_613);
  nand g519 (n_699, n_616, n_617);
  nand g522 (n_701, n_620, n_621);
  nand g525 (n_704, n_624, n_625);
  nand g528 (n_707, n_628, n_629);
  nand g531 (n_710, n_632, n_633);
  nand g534 (n_712, n_636, n_637);
  nand g537 (n_715, n_640, n_641);
  xnor g539 (out_0[1], n_327, n_642);
  xnor g541 (out_0[2], n_417, n_643);
  xnor g544 (out_0[3], n_645, n_646);
  xnor g546 (out_0[4], n_488, n_647);
  xnor g549 (out_0[5], n_649, n_650);
  xnor g551 (out_0[6], n_651, n_652);
  xnor g554 (out_0[7], n_654, n_655);
  xnor g556 (out_0[8], n_541, n_656);
  xnor g559 (out_0[9], n_658, n_659);
  xnor g561 (out_0[10], n_660, n_661);
  xnor g564 (out_0[11], n_663, n_664);
  xnor g567 (out_0[12], n_666, n_667);
  xnor g570 (out_0[13], n_669, n_670);
  xnor g572 (out_0[14], n_671, n_672);
  xnor g575 (out_0[15], n_674, n_675);
  xnor g577 (out_0[16], n_594, n_676);
  xnor g580 (out_0[17], n_678, n_679);
  xnor g582 (out_0[18], n_680, n_681);
  xnor g585 (out_0[19], n_683, n_684);
  xnor g588 (out_0[20], n_686, n_687);
  xnor g591 (out_0[21], n_689, n_690);
  xnor g593 (out_0[22], n_691, n_692);
  xnor g596 (out_0[23], n_694, n_695);
  xnor g598 (out_0[24], n_696, n_697);
  xnor g601 (out_0[25], n_699, n_700);
  xnor g603 (out_0[26], n_701, n_702);
  xnor g606 (out_0[27], n_704, n_705);
  xnor g609 (out_0[28], n_707, n_708);
  xnor g612 (out_0[29], n_710, n_711);
  xnor g614 (out_0[30], n_712, n_713);
  xnor g617 (out_0[31], n_715, n_716);
  xor g618 (out_0[0], in_0[0], n_717);
  xnor g621 (n_311, in_1[30], in_2[30]);
  or g622 (n_312, in_2[30], wc);
  not gc (wc, in_1[30]);
  or g623 (n_313, in_0[30], in_2[30]);
  or g624 (n_314, wc0, in_0[30]);
  not gc0 (wc0, in_1[30]);
  xnor g625 (n_316, in_0[31], in_1[31]);
  xnor g626 (n_163, n_311, in_0[30]);
  or g627 (n_330, n_326, wc1);
  not gc1 (wc1, n_327);
  or g628 (n_642, wc2, n_326);
  not gc2 (wc2, n_329);
  and g629 (n_414, n_130, n_162);
  or g630 (n_415, n_130, n_162);
  and g631 (n_421, wc3, n_333);
  not gc3 (wc3, n_334);
  and g632 (n_423, wc4, n_339);
  not gc4 (wc4, n_340);
  and g633 (n_430, wc5, n_345);
  not gc5 (wc5, n_346);
  and g634 (n_433, wc6, n_351);
  not gc6 (wc6, n_352);
  and g635 (n_440, wc7, n_357);
  not gc7 (wc7, n_358);
  and g636 (n_443, wc8, n_363);
  not gc8 (wc8, n_364);
  and g637 (n_450, wc9, n_369);
  not gc9 (wc9, n_370);
  and g638 (n_453, wc10, n_375);
  not gc10 (wc10, n_376);
  and g639 (n_460, wc11, n_160);
  not gc11 (wc11, n_161);
  and g640 (n_463, wc12, n_385);
  not gc12 (wc12, n_386);
  and g641 (n_470, wc13, n_391);
  not gc13 (wc13, n_392);
  and g642 (n_473, wc14, n_397);
  not gc14 (wc14, n_398);
  and g643 (n_480, wc15, n_403);
  not gc15 (wc15, n_404);
  and g644 (n_483, wc16, n_409);
  not gc16 (wc16, n_410);
  or g645 (n_492, wc17, n_348);
  not gc17 (wc17, n_426);
  or g646 (n_545, wc18, n_360);
  not gc18 (wc18, n_436);
  or g647 (n_507, wc19, n_372);
  not gc19 (wc19, n_446);
  or g648 (n_598, wc20, n_382);
  not gc20 (wc20, n_456);
  or g649 (n_522, wc21, n_394);
  not gc21 (wc21, n_466);
  or g650 (n_571, wc22, n_406);
  not gc22 (wc22, n_476);
  or g651 (n_643, wc23, n_336);
  not gc23 (wc23, n_331);
  or g652 (n_646, wc24, n_332);
  not gc24 (wc24, n_333);
  or g653 (n_647, wc25, n_342);
  not gc25 (wc25, n_337);
  or g654 (n_650, wc26, n_338);
  not gc26 (wc26, n_339);
  or g655 (n_652, wc27, n_348);
  not gc27 (wc27, n_343);
  or g656 (n_655, wc28, n_344);
  not gc28 (wc28, n_345);
  or g657 (n_656, wc29, n_354);
  not gc29 (wc29, n_349);
  or g658 (n_659, wc30, n_350);
  not gc30 (wc30, n_351);
  or g659 (n_661, wc31, n_360);
  not gc31 (wc31, n_355);
  or g660 (n_664, wc32, n_356);
  not gc32 (wc32, n_357);
  or g661 (n_667, wc33, n_366);
  not gc33 (wc33, n_361);
  or g662 (n_670, wc34, n_362);
  not gc34 (wc34, n_363);
  or g663 (n_672, wc35, n_372);
  not gc35 (wc35, n_367);
  or g664 (n_675, wc36, n_368);
  not gc36 (wc36, n_369);
  or g665 (n_676, wc37, n_378);
  not gc37 (wc37, n_373);
  or g666 (n_679, wc38, n_374);
  not gc38 (wc38, n_375);
  or g667 (n_681, wc39, n_382);
  not gc39 (wc39, n_379);
  or g668 (n_684, wc40, n_380);
  not gc40 (wc40, n_160);
  or g669 (n_687, wc41, n_388);
  not gc41 (wc41, n_383);
  or g670 (n_690, wc42, n_384);
  not gc42 (wc42, n_385);
  or g671 (n_692, wc43, n_394);
  not gc43 (wc43, n_389);
  or g672 (n_695, wc44, n_390);
  not gc44 (wc44, n_391);
  or g673 (n_697, wc45, n_400);
  not gc45 (wc45, n_395);
  or g674 (n_700, wc46, n_396);
  not gc46 (wc46, n_397);
  or g675 (n_702, wc47, n_406);
  not gc47 (wc47, n_401);
  or g676 (n_705, wc48, n_402);
  not gc48 (wc48, n_403);
  or g677 (n_708, wc49, n_412);
  not gc49 (wc49, n_407);
  or g678 (n_711, wc50, n_408);
  not gc50 (wc50, n_409);
  or g679 (n_419, wc51, n_336);
  not gc51 (wc51, n_417);
  and g680 (n_431, wc52, n_428);
  not gc52 (wc52, n_423);
  and g681 (n_441, wc53, n_438);
  not gc53 (wc53, n_433);
  and g682 (n_451, wc54, n_448);
  not gc54 (wc54, n_443);
  and g683 (n_461, wc55, n_458);
  not gc55 (wc55, n_453);
  and g684 (n_471, wc56, n_468);
  not gc56 (wc56, n_463);
  and g685 (n_481, wc57, n_478);
  not gc57 (wc57, n_473);
  or g686 (n_537, wc58, n_416);
  not gc58 (wc58, n_486);
  and g687 (n_554, wc59, n_446);
  not gc59 (wc59, n_503);
  and g688 (n_607, wc60, n_466);
  not gc60 (wc60, n_518);
  and g689 (n_584, wc61, n_486);
  not gc61 (wc61, n_533);
  or g690 (n_713, wc62, n_416);
  not gc62 (wc62, n_413);
  and g691 (n_494, wc63, n_343);
  not gc63 (wc63, n_424);
  and g692 (n_498, wc64, n_430);
  not gc64 (wc64, n_431);
  and g693 (n_547, wc65, n_355);
  not gc65 (wc65, n_434);
  and g694 (n_500, wc66, n_440);
  not gc66 (wc66, n_441);
  and g695 (n_508, wc67, n_367);
  not gc67 (wc67, n_444);
  and g696 (n_512, wc68, n_450);
  not gc68 (wc68, n_451);
  and g697 (n_600, wc69, n_379);
  not gc69 (wc69, n_454);
  and g698 (n_515, wc70, n_460);
  not gc70 (wc70, n_461);
  and g699 (n_523, wc71, n_389);
  not gc71 (wc71, n_464);
  and g700 (n_527, wc72, n_470);
  not gc72 (wc72, n_471);
  and g701 (n_572, wc73, n_401);
  not gc73 (wc73, n_474);
  and g702 (n_530, wc74, n_480);
  not gc74 (wc74, n_481);
  and g703 (n_538, wc75, n_413);
  not gc75 (wc75, n_484);
  or g704 (n_614, wc76, n_400);
  not gc76 (wc76, n_566);
  or g705 (n_622, n_571, wc77);
  not gc77 (wc77, n_566);
  or g706 (n_626, wc78, n_533);
  not gc78 (wc78, n_566);
  or g707 (n_716, wc79, n_414);
  not gc79 (wc79, n_415);
  or g708 (n_490, wc80, n_342);
  not gc80 (wc80, n_488);
  or g709 (n_495, n_492, wc81);
  not gc81 (wc81, n_488);
  or g710 (n_499, n_496, wc82);
  not gc82 (wc82, n_488);
  and g711 (n_505, wc83, n_446);
  not gc83 (wc83, n_500);
  and g712 (n_520, wc84, n_466);
  not gc84 (wc84, n_515);
  and g713 (n_535, wc85, n_486);
  not gc85 (wc85, n_530);
  and g714 (n_552, wc86, n_361);
  not gc86 (wc86, n_501);
  and g715 (n_555, wc87, n_443);
  not gc87 (wc87, n_505);
  and g716 (n_558, n_508, wc88);
  not gc88 (wc88, n_509);
  and g717 (n_561, n_512, wc89);
  not gc89 (wc89, n_513);
  and g718 (n_605, wc90, n_383);
  not gc90 (wc90, n_516);
  and g719 (n_608, wc91, n_463);
  not gc91 (wc91, n_520);
  and g720 (n_611, n_523, wc92);
  not gc92 (wc92, n_524);
  and g721 (n_563, n_527, wc93);
  not gc93 (wc93, n_528);
  and g722 (n_581, wc94, n_407);
  not gc94 (wc94, n_531);
  and g723 (n_586, wc95, n_483);
  not gc95 (wc95, n_535);
  and g724 (n_591, n_538, wc96);
  not gc96 (wc96, n_539);
  or g725 (n_543, wc97, n_354);
  not gc97 (wc97, n_541);
  or g726 (n_548, n_545, wc98);
  not gc98 (wc98, n_541);
  or g727 (n_550, wc99, n_503);
  not gc99 (wc99, n_541);
  and g728 (n_569, wc100, n_476);
  not gc100 (wc100, n_563);
  and g729 (n_582, wc101, n_579);
  not gc101 (wc101, n_563);
  and g730 (n_587, wc102, n_584);
  not gc102 (wc102, n_563);
  and g731 (n_592, wc103, n_589);
  not gc103 (wc103, n_563);
  and g732 (n_616, wc104, n_395);
  not gc104 (wc104, n_564);
  and g733 (n_620, wc105, n_473);
  not gc105 (wc105, n_569);
  and g734 (n_624, n_572, wc106);
  not gc106 (wc106, n_573);
  and g735 (n_628, n_530, wc107);
  not gc107 (wc107, n_576);
  and g736 (n_632, wc108, n_581);
  not gc108 (wc108, n_582);
  and g737 (n_636, wc109, n_586);
  not gc109 (wc109, n_587);
  and g738 (n_640, wc110, n_591);
  not gc110 (wc110, n_592);
  or g739 (n_596, wc111, n_378);
  not gc111 (wc111, n_594);
  or g740 (n_601, n_598, wc112);
  not gc112 (wc112, n_594);
  or g741 (n_603, wc113, n_518);
  not gc113 (wc113, n_594);
  or g742 (n_617, n_614, wc114);
  not gc114 (wc114, n_594);
  or g743 (n_621, n_618, wc115);
  not gc115 (wc115, n_594);
  or g744 (n_625, n_622, wc116);
  not gc116 (wc116, n_594);
  or g745 (n_629, n_626, wc117);
  not gc117 (wc117, n_594);
  or g746 (n_633, n_630, wc118);
  not gc118 (wc118, n_594);
  or g747 (n_637, n_634, wc119);
  not gc119 (wc119, n_594);
  or g748 (n_641, n_638, wc120);
  not gc120 (wc120, n_594);
endmodule

module csa_tree_add_559_42_group_16914_GENERIC(in_0, in_1, in_2, out_0);
  input [32:0] in_0, in_1;
  input [30:0] in_2;
  output [31:0] out_0;
  wire [32:0] in_0, in_1;
  wire [30:0] in_2;
  wire [31:0] out_0;
  csa_tree_add_559_42_group_16914_GENERIC_REAL g1(.in_0 ({in_0[32],
       in_0[28], in_0[28], in_0[28], in_0[28:0]}), .in_1 ({in_1[32],
       in_1[28], in_1[28], in_1[28], in_1[28:0]}), .in_2 ({in_2[29],
       in_2[29:0]}), .out_0 (out_0));
endmodule

module csa_tree_add_607_44_group_16902_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_1) + $signed(in_2) )  + $signed(in_0) )  ;"
  input [55:0] in_0, in_1, in_2;
  output [57:0] out_0;
  wire [55:0] in_0, in_1, in_2;
  wire [57:0] out_0;
  wire n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_241, n_242, n_243, n_244;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268;
  wire n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276;
  wire n_277, n_278, n_279, n_280, n_281, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560;
  wire n_571, n_572, n_573, n_574, n_576, n_577, n_578, n_579;
  wire n_580, n_582, n_583, n_584, n_585, n_586, n_588, n_589;
  wire n_590, n_591, n_592, n_594, n_595, n_596, n_597, n_598;
  wire n_600, n_601, n_602, n_603, n_604, n_606, n_607, n_608;
  wire n_609, n_610, n_612, n_613, n_614, n_615, n_616, n_618;
  wire n_619, n_620, n_621, n_622, n_624, n_625, n_626, n_627;
  wire n_628, n_630, n_631, n_632, n_633, n_634, n_636, n_637;
  wire n_638, n_639, n_640, n_642, n_643, n_644, n_645, n_646;
  wire n_648, n_649, n_650, n_651, n_652, n_654, n_655, n_656;
  wire n_657, n_658, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_666, n_667, n_668, n_669, n_671, n_672, n_673, n_674;
  wire n_675, n_677, n_678, n_679, n_680, n_681, n_683, n_684;
  wire n_685, n_686, n_687, n_689, n_690, n_691, n_692, n_693;
  wire n_695, n_696, n_697, n_698, n_699, n_701, n_702, n_703;
  wire n_704, n_705, n_707, n_708, n_709, n_710, n_711, n_713;
  wire n_714, n_715, n_716, n_717, n_719, n_720, n_721, n_722;
  wire n_723, n_725, n_726, n_727, n_728, n_729, n_731, n_732;
  wire n_735, n_740, n_742, n_743, n_745, n_747, n_749, n_750;
  wire n_752, n_753, n_755, n_757, n_759, n_760, n_762, n_763;
  wire n_765, n_767, n_769, n_770, n_772, n_773, n_775, n_777;
  wire n_779, n_780, n_782, n_783, n_785, n_787, n_789, n_790;
  wire n_792, n_793, n_795, n_797, n_799, n_800, n_802, n_803;
  wire n_805, n_807, n_809, n_810, n_812, n_813, n_815, n_817;
  wire n_819, n_820, n_822, n_823, n_825, n_827, n_829, n_830;
  wire n_832, n_833, n_835, n_837, n_839, n_840, n_842, n_843;
  wire n_845, n_847, n_849, n_850, n_852, n_853, n_855, n_857;
  wire n_859, n_860, n_862, n_863, n_865, n_867, n_869, n_870;
  wire n_874, n_875, n_876, n_878, n_879, n_880, n_882, n_883;
  wire n_884, n_885, n_887, n_889, n_891, n_892, n_893, n_895;
  wire n_896, n_897, n_899, n_900, n_902, n_904, n_906, n_907;
  wire n_908, n_910, n_911, n_912, n_914, n_915, n_917, n_919;
  wire n_921, n_922, n_923, n_925, n_926, n_927, n_929, n_930;
  wire n_932, n_934, n_936, n_937, n_938, n_940, n_941, n_942;
  wire n_944, n_945, n_947, n_949, n_951, n_952, n_953, n_955;
  wire n_956, n_957, n_959, n_960, n_962, n_964, n_966, n_967;
  wire n_968, n_970, n_971, n_972, n_974, n_976, n_977, n_978;
  wire n_980, n_981, n_983, n_984, n_985, n_986, n_987, n_988;
  wire n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996;
  wire n_997, n_999, n_1002, n_1004, n_1005, n_1006, n_1009, n_1012;
  wire n_1014, n_1015, n_1017, n_1019, n_1020, n_1022, n_1024, n_1025;
  wire n_1027, n_1029, n_1030, n_1032, n_1033, n_1035, n_1038, n_1040;
  wire n_1041, n_1042, n_1045, n_1048, n_1050, n_1051, n_1053, n_1055;
  wire n_1056, n_1058, n_1060, n_1061, n_1063, n_1065, n_1066, n_1068;
  wire n_1069, n_1071, n_1073, n_1075, n_1076, n_1077, n_1079, n_1080;
  wire n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089;
  wire n_1090, n_1091, n_1092, n_1093, n_1095, n_1096, n_1097, n_1099;
  wire n_1100, n_1101, n_1103, n_1104, n_1105, n_1107, n_1108, n_1109;
  wire n_1111, n_1112, n_1113, n_1115, n_1116, n_1117, n_1119, n_1120;
  wire n_1121, n_1123, n_1124, n_1125, n_1126, n_1128, n_1130, n_1132;
  wire n_1133, n_1134, n_1136, n_1138, n_1140, n_1141, n_1143, n_1145;
  wire n_1146, n_1148, n_1150, n_1151, n_1154, n_1156, n_1157, n_1158;
  wire n_1160, n_1162, n_1163, n_1164, n_1166, n_1167, n_1169, n_1170;
  wire n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178;
  wire n_1179, n_1180, n_1182, n_1183, n_1184, n_1186, n_1187, n_1188;
  wire n_1190, n_1191, n_1192, n_1194, n_1195, n_1196, n_1198, n_1199;
  wire n_1200, n_1202, n_1203, n_1204, n_1206, n_1207, n_1209, n_1210;
  wire n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218;
  wire n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226;
  wire n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234;
  wire n_1235, n_1236, n_1238, n_1241, n_1242, n_1244, n_1245, n_1246;
  wire n_1247, n_1249, n_1250, n_1251, n_1253, n_1254, n_1255, n_1256;
  wire n_1258, n_1259, n_1261, n_1262, n_1264, n_1265, n_1266, n_1267;
  wire n_1269, n_1270, n_1271, n_1273, n_1274, n_1275, n_1276, n_1278;
  wire n_1279, n_1281, n_1282, n_1284, n_1285, n_1286, n_1287, n_1289;
  wire n_1290, n_1291, n_1292, n_1294, n_1295, n_1296, n_1297, n_1299;
  wire n_1300, n_1302, n_1303, n_1305, n_1306, n_1307, n_1308, n_1310;
  wire n_1311, n_1312, n_1314, n_1315, n_1316, n_1317, n_1319, n_1320;
  wire n_1322, n_1323, n_1325, n_1326, n_1327, n_1328, n_1330, n_1331;
  wire n_1332, n_1333, n_1335, n_1336, n_1337, n_1338, n_1340, n_1341;
  wire n_1343, n_1344, n_1346, n_1347, n_1348, n_1349, n_1351, n_1352;
  wire n_1354, n_1355, n_1357, n_1358, n_1359, n_1360, n_1362, n_1363;
  wire n_1365, n_1366, n_1368, n_1369, n_1370, n_1371, n_1373, n_1374;
  wire n_1375, n_1376, n_1378;
  assign out_0[0] = 1'b0;
  assign out_0[1] = 1'b0;
  xor g59 (n_340, in_0[2], in_2[2]);
  and g60 (n_281, in_0[2], in_2[2]);
  xor g61 (n_349, in_0[3], in_2[3]);
  xor g62 (n_339, n_349, in_1[3]);
  nand g63 (n_350, in_0[3], in_2[3]);
  nand g4 (n_351, in_1[3], in_2[3]);
  nand g5 (n_352, in_0[3], in_1[3]);
  nand g64 (n_280, n_350, n_351, n_352);
  xor g65 (n_353, in_0[4], in_2[4]);
  xor g66 (n_338, n_353, in_1[4]);
  nand g67 (n_354, in_0[4], in_2[4]);
  nand g68 (n_355, in_1[4], in_2[4]);
  nand g69 (n_356, in_0[4], in_1[4]);
  nand g6 (n_279, n_354, n_355, n_356);
  xor g70 (n_357, in_0[5], in_2[5]);
  xor g71 (n_337, n_357, in_1[5]);
  nand g72 (n_358, in_0[5], in_2[5]);
  nand g73 (n_359, in_1[5], in_2[5]);
  nand g74 (n_360, in_0[5], in_1[5]);
  nand g75 (n_278, n_358, n_359, n_360);
  xor g76 (n_361, in_0[6], in_2[6]);
  xor g77 (n_336, n_361, in_1[6]);
  nand g78 (n_362, in_0[6], in_2[6]);
  nand g79 (n_363, in_1[6], in_2[6]);
  nand g80 (n_364, in_0[6], in_1[6]);
  nand g81 (n_277, n_362, n_363, n_364);
  xor g82 (n_365, in_0[7], in_2[7]);
  xor g83 (n_335, n_365, in_1[7]);
  nand g84 (n_366, in_0[7], in_2[7]);
  nand g85 (n_367, in_1[7], in_2[7]);
  nand g86 (n_368, in_0[7], in_1[7]);
  nand g87 (n_276, n_366, n_367, n_368);
  xor g88 (n_369, in_0[8], in_2[8]);
  xor g89 (n_334, n_369, in_1[8]);
  nand g90 (n_370, in_0[8], in_2[8]);
  nand g91 (n_371, in_1[8], in_2[8]);
  nand g92 (n_372, in_0[8], in_1[8]);
  nand g93 (n_275, n_370, n_371, n_372);
  xor g94 (n_373, in_0[9], in_2[9]);
  xor g95 (n_333, n_373, in_1[9]);
  nand g96 (n_374, in_0[9], in_2[9]);
  nand g97 (n_375, in_1[9], in_2[9]);
  nand g98 (n_376, in_0[9], in_1[9]);
  nand g99 (n_274, n_374, n_375, n_376);
  xor g100 (n_377, in_0[10], in_2[10]);
  xor g101 (n_332, n_377, in_1[10]);
  nand g102 (n_378, in_0[10], in_2[10]);
  nand g103 (n_379, in_1[10], in_2[10]);
  nand g104 (n_380, in_0[10], in_1[10]);
  nand g105 (n_273, n_378, n_379, n_380);
  xor g106 (n_381, in_0[11], in_2[11]);
  xor g107 (n_331, n_381, in_1[11]);
  nand g108 (n_382, in_0[11], in_2[11]);
  nand g109 (n_383, in_1[11], in_2[11]);
  nand g110 (n_384, in_0[11], in_1[11]);
  nand g111 (n_272, n_382, n_383, n_384);
  xor g112 (n_385, in_0[12], in_2[12]);
  xor g113 (n_330, n_385, in_1[12]);
  nand g114 (n_386, in_0[12], in_2[12]);
  nand g115 (n_387, in_1[12], in_2[12]);
  nand g116 (n_388, in_0[12], in_1[12]);
  nand g117 (n_271, n_386, n_387, n_388);
  xor g118 (n_389, in_0[13], in_2[13]);
  xor g119 (n_329, n_389, in_1[13]);
  nand g120 (n_390, in_0[13], in_2[13]);
  nand g121 (n_391, in_1[13], in_2[13]);
  nand g122 (n_392, in_0[13], in_1[13]);
  nand g123 (n_270, n_390, n_391, n_392);
  xor g124 (n_393, in_0[14], in_2[14]);
  xor g125 (n_328, n_393, in_1[14]);
  nand g126 (n_394, in_0[14], in_2[14]);
  nand g127 (n_395, in_1[14], in_2[14]);
  nand g128 (n_396, in_0[14], in_1[14]);
  nand g129 (n_269, n_394, n_395, n_396);
  xor g130 (n_397, in_0[15], in_2[15]);
  xor g131 (n_327, n_397, in_1[15]);
  nand g132 (n_398, in_0[15], in_2[15]);
  nand g133 (n_399, in_1[15], in_2[15]);
  nand g134 (n_400, in_0[15], in_1[15]);
  nand g135 (n_268, n_398, n_399, n_400);
  xor g136 (n_401, in_0[16], in_2[16]);
  xor g137 (n_326, n_401, in_1[16]);
  nand g138 (n_402, in_0[16], in_2[16]);
  nand g139 (n_403, in_1[16], in_2[16]);
  nand g140 (n_404, in_0[16], in_1[16]);
  nand g141 (n_267, n_402, n_403, n_404);
  xor g142 (n_405, in_0[17], in_2[17]);
  xor g143 (n_325, n_405, in_1[17]);
  nand g144 (n_406, in_0[17], in_2[17]);
  nand g145 (n_407, in_1[17], in_2[17]);
  nand g146 (n_408, in_0[17], in_1[17]);
  nand g147 (n_266, n_406, n_407, n_408);
  xor g148 (n_409, in_0[18], in_2[18]);
  xor g149 (n_324, n_409, in_1[18]);
  nand g150 (n_410, in_0[18], in_2[18]);
  nand g151 (n_411, in_1[18], in_2[18]);
  nand g152 (n_412, in_0[18], in_1[18]);
  nand g153 (n_265, n_410, n_411, n_412);
  xor g154 (n_413, in_0[19], in_2[19]);
  xor g155 (n_323, n_413, in_1[19]);
  nand g156 (n_414, in_0[19], in_2[19]);
  nand g157 (n_415, in_1[19], in_2[19]);
  nand g158 (n_416, in_0[19], in_1[19]);
  nand g159 (n_264, n_414, n_415, n_416);
  xor g160 (n_417, in_0[20], in_2[20]);
  xor g161 (n_322, n_417, in_1[20]);
  nand g162 (n_418, in_0[20], in_2[20]);
  nand g163 (n_419, in_1[20], in_2[20]);
  nand g164 (n_420, in_0[20], in_1[20]);
  nand g165 (n_263, n_418, n_419, n_420);
  xor g166 (n_421, in_0[21], in_2[21]);
  xor g167 (n_321, n_421, in_1[21]);
  nand g168 (n_422, in_0[21], in_2[21]);
  nand g169 (n_423, in_1[21], in_2[21]);
  nand g170 (n_424, in_0[21], in_1[21]);
  nand g171 (n_262, n_422, n_423, n_424);
  xor g172 (n_425, in_0[22], in_2[22]);
  xor g173 (n_320, n_425, in_1[22]);
  nand g174 (n_426, in_0[22], in_2[22]);
  nand g175 (n_427, in_1[22], in_2[22]);
  nand g176 (n_428, in_0[22], in_1[22]);
  nand g177 (n_261, n_426, n_427, n_428);
  xor g178 (n_429, in_0[23], in_2[23]);
  xor g179 (n_319, n_429, in_1[23]);
  nand g180 (n_430, in_0[23], in_2[23]);
  nand g181 (n_431, in_1[23], in_2[23]);
  nand g182 (n_432, in_0[23], in_1[23]);
  nand g183 (n_260, n_430, n_431, n_432);
  xor g184 (n_433, in_0[24], in_2[24]);
  xor g185 (n_318, n_433, in_1[24]);
  nand g186 (n_434, in_0[24], in_2[24]);
  nand g187 (n_435, in_1[24], in_2[24]);
  nand g188 (n_436, in_0[24], in_1[24]);
  nand g189 (n_259, n_434, n_435, n_436);
  xor g190 (n_437, in_0[25], in_2[25]);
  xor g191 (n_317, n_437, in_1[25]);
  nand g192 (n_438, in_0[25], in_2[25]);
  nand g193 (n_439, in_1[25], in_2[25]);
  nand g194 (n_440, in_0[25], in_1[25]);
  nand g195 (n_258, n_438, n_439, n_440);
  xor g196 (n_441, in_0[26], in_2[26]);
  xor g197 (n_316, n_441, in_1[26]);
  nand g198 (n_442, in_0[26], in_2[26]);
  nand g199 (n_443, in_1[26], in_2[26]);
  nand g200 (n_444, in_0[26], in_1[26]);
  nand g201 (n_257, n_442, n_443, n_444);
  xor g202 (n_445, in_0[27], in_2[27]);
  xor g203 (n_315, n_445, in_1[27]);
  nand g204 (n_446, in_0[27], in_2[27]);
  nand g205 (n_447, in_1[27], in_2[27]);
  nand g206 (n_448, in_0[27], in_1[27]);
  nand g207 (n_256, n_446, n_447, n_448);
  xor g208 (n_449, in_0[28], in_2[28]);
  xor g209 (n_314, n_449, in_1[28]);
  nand g210 (n_450, in_0[28], in_2[28]);
  nand g211 (n_451, in_1[28], in_2[28]);
  nand g212 (n_452, in_0[28], in_1[28]);
  nand g213 (n_255, n_450, n_451, n_452);
  xor g214 (n_453, in_0[29], in_2[29]);
  xor g215 (n_313, n_453, in_1[29]);
  nand g216 (n_454, in_0[29], in_2[29]);
  nand g217 (n_455, in_1[29], in_2[29]);
  nand g218 (n_456, in_0[29], in_1[29]);
  nand g219 (n_254, n_454, n_455, n_456);
  xor g220 (n_457, in_0[30], in_2[30]);
  xor g221 (n_312, n_457, in_1[30]);
  nand g222 (n_458, in_0[30], in_2[30]);
  nand g223 (n_459, in_1[30], in_2[30]);
  nand g224 (n_460, in_0[30], in_1[30]);
  nand g225 (n_253, n_458, n_459, n_460);
  xor g226 (n_461, in_0[31], in_2[31]);
  xor g227 (n_311, n_461, in_1[31]);
  nand g228 (n_462, in_0[31], in_2[31]);
  nand g229 (n_463, in_1[31], in_2[31]);
  nand g230 (n_464, in_0[31], in_1[31]);
  nand g231 (n_252, n_462, n_463, n_464);
  xor g232 (n_465, in_0[32], in_2[32]);
  xor g233 (n_310, n_465, in_1[32]);
  nand g234 (n_466, in_0[32], in_2[32]);
  nand g235 (n_467, in_1[32], in_2[32]);
  nand g236 (n_468, in_0[32], in_1[32]);
  nand g237 (n_251, n_466, n_467, n_468);
  xor g238 (n_469, in_0[33], in_2[33]);
  xor g239 (n_309, n_469, in_1[33]);
  nand g240 (n_470, in_0[33], in_2[33]);
  nand g241 (n_471, in_1[33], in_2[33]);
  nand g242 (n_472, in_0[33], in_1[33]);
  nand g243 (n_250, n_470, n_471, n_472);
  xor g244 (n_473, in_0[34], in_2[34]);
  xor g245 (n_308, n_473, in_1[34]);
  nand g246 (n_474, in_0[34], in_2[34]);
  nand g247 (n_475, in_1[34], in_2[34]);
  nand g248 (n_476, in_0[34], in_1[34]);
  nand g249 (n_249, n_474, n_475, n_476);
  xor g250 (n_477, in_0[35], in_2[35]);
  xor g251 (n_307, n_477, in_1[35]);
  nand g252 (n_478, in_0[35], in_2[35]);
  nand g253 (n_479, in_1[35], in_2[35]);
  nand g254 (n_480, in_0[35], in_1[35]);
  nand g255 (n_248, n_478, n_479, n_480);
  xor g256 (n_481, in_0[36], in_2[36]);
  xor g257 (n_306, n_481, in_1[36]);
  nand g258 (n_482, in_0[36], in_2[36]);
  nand g259 (n_483, in_1[36], in_2[36]);
  nand g260 (n_484, in_0[36], in_1[36]);
  nand g261 (n_247, n_482, n_483, n_484);
  xor g262 (n_485, in_0[37], in_2[37]);
  xor g263 (n_305, n_485, in_1[37]);
  nand g264 (n_486, in_0[37], in_2[37]);
  nand g265 (n_487, in_1[37], in_2[37]);
  nand g266 (n_488, in_0[37], in_1[37]);
  nand g267 (n_246, n_486, n_487, n_488);
  xor g268 (n_489, in_0[38], in_2[38]);
  xor g269 (n_304, n_489, in_1[38]);
  nand g270 (n_490, in_0[38], in_2[38]);
  nand g271 (n_491, in_1[38], in_2[38]);
  nand g272 (n_492, in_0[38], in_1[38]);
  nand g273 (n_245, n_490, n_491, n_492);
  xor g274 (n_493, in_0[39], in_2[39]);
  xor g275 (n_303, n_493, in_1[39]);
  nand g276 (n_494, in_0[39], in_2[39]);
  nand g277 (n_495, in_1[39], in_2[39]);
  nand g278 (n_496, in_0[39], in_1[39]);
  nand g279 (n_244, n_494, n_495, n_496);
  xor g280 (n_497, in_0[40], in_2[40]);
  xor g281 (n_302, n_497, in_1[40]);
  nand g282 (n_498, in_0[40], in_2[40]);
  nand g283 (n_499, in_1[40], in_2[40]);
  nand g284 (n_500, in_0[40], in_1[40]);
  nand g285 (n_243, n_498, n_499, n_500);
  xor g286 (n_501, in_0[41], in_2[41]);
  xor g287 (n_301, n_501, in_1[41]);
  nand g288 (n_502, in_0[41], in_2[41]);
  nand g289 (n_503, in_1[41], in_2[41]);
  nand g290 (n_504, in_0[41], in_1[41]);
  nand g291 (n_242, n_502, n_503, n_504);
  xor g292 (n_505, in_0[42], in_2[42]);
  xor g293 (n_300, n_505, in_1[42]);
  nand g294 (n_506, in_0[42], in_2[42]);
  nand g295 (n_507, in_1[42], in_2[42]);
  nand g296 (n_508, in_0[42], in_1[42]);
  nand g297 (n_241, n_506, n_507, n_508);
  xor g298 (n_509, in_0[43], in_2[43]);
  xor g299 (n_299, n_509, in_1[43]);
  nand g300 (n_510, in_0[43], in_2[43]);
  nand g301 (n_511, in_1[43], in_2[43]);
  nand g302 (n_512, in_0[43], in_1[43]);
  nand g303 (n_240, n_510, n_511, n_512);
  xor g304 (n_513, in_0[44], in_2[44]);
  xor g305 (n_298, n_513, in_1[44]);
  nand g306 (n_514, in_0[44], in_2[44]);
  nand g307 (n_515, in_1[44], in_2[44]);
  nand g308 (n_516, in_0[44], in_1[44]);
  nand g309 (n_239, n_514, n_515, n_516);
  xor g310 (n_517, in_0[45], in_2[45]);
  xor g311 (n_297, n_517, in_1[45]);
  nand g312 (n_518, in_0[45], in_2[45]);
  nand g313 (n_519, in_1[45], in_2[45]);
  nand g314 (n_520, in_0[45], in_1[45]);
  nand g315 (n_238, n_518, n_519, n_520);
  xor g316 (n_521, in_0[46], in_2[46]);
  xor g317 (n_296, n_521, in_1[46]);
  nand g318 (n_522, in_0[46], in_2[46]);
  nand g319 (n_523, in_1[46], in_2[46]);
  nand g320 (n_524, in_0[46], in_1[46]);
  nand g321 (n_237, n_522, n_523, n_524);
  xor g322 (n_525, in_0[47], in_2[47]);
  xor g323 (n_295, n_525, in_1[47]);
  nand g324 (n_526, in_0[47], in_2[47]);
  nand g325 (n_527, in_1[47], in_2[47]);
  nand g326 (n_528, in_0[47], in_1[47]);
  nand g327 (n_236, n_526, n_527, n_528);
  xor g328 (n_529, in_0[48], in_2[48]);
  xor g329 (n_294, n_529, in_1[48]);
  nand g330 (n_530, in_0[48], in_2[48]);
  nand g331 (n_531, in_1[48], in_2[48]);
  nand g332 (n_532, in_0[48], in_1[48]);
  nand g333 (n_235, n_530, n_531, n_532);
  xor g334 (n_533, in_0[49], in_2[49]);
  xor g335 (n_293, n_533, in_1[49]);
  nand g336 (n_534, in_0[49], in_2[49]);
  nand g337 (n_535, in_1[49], in_2[49]);
  nand g338 (n_536, in_0[49], in_1[49]);
  nand g339 (n_234, n_534, n_535, n_536);
  xor g340 (n_537, in_0[50], in_2[50]);
  xor g341 (n_292, n_537, in_1[50]);
  nand g342 (n_538, in_0[50], in_2[50]);
  nand g343 (n_539, in_1[50], in_2[50]);
  nand g344 (n_540, in_0[50], in_1[50]);
  nand g345 (n_233, n_538, n_539, n_540);
  xor g346 (n_541, in_0[51], in_2[51]);
  xor g347 (n_291, n_541, in_1[51]);
  nand g348 (n_542, in_0[51], in_2[51]);
  nand g349 (n_543, in_1[51], in_2[51]);
  nand g350 (n_544, in_0[51], in_1[51]);
  nand g351 (n_232, n_542, n_543, n_544);
  xor g352 (n_545, in_0[52], in_2[52]);
  xor g353 (n_290, n_545, in_1[52]);
  nand g354 (n_546, in_0[52], in_2[52]);
  nand g355 (n_547, in_1[52], in_2[52]);
  nand g356 (n_548, in_0[52], in_1[52]);
  nand g357 (n_231, n_546, n_547, n_548);
  xor g358 (n_549, in_0[53], in_2[53]);
  xor g359 (n_289, n_549, in_1[53]);
  nand g360 (n_550, in_0[53], in_2[53]);
  nand g361 (n_551, in_1[53], in_2[53]);
  nand g362 (n_552, in_0[53], in_1[53]);
  nand g363 (n_230, n_550, n_551, n_552);
  xor g364 (n_553, in_0[54], in_2[54]);
  xor g365 (n_288, n_553, in_1[54]);
  nand g366 (n_554, in_0[54], in_2[54]);
  nand g367 (n_555, in_1[54], in_2[54]);
  nand g368 (n_556, in_0[54], in_1[54]);
  nand g369 (n_229, n_554, n_555, n_556);
  xor g373 (n_287, n_557, in_0[55]);
  nand g377 (n_286, n_558, n_559, n_560);
  nor g11 (n_576, in_1[2], n_340);
  nand g12 (n_571, in_1[2], n_340);
  nor g13 (n_572, n_281, n_339);
  nand g14 (n_573, n_281, n_339);
  nor g15 (n_582, n_280, n_338);
  nand g16 (n_577, n_280, n_338);
  nor g17 (n_578, n_279, n_337);
  nand g18 (n_579, n_279, n_337);
  nor g19 (n_588, n_278, n_336);
  nand g20 (n_583, n_278, n_336);
  nor g21 (n_584, n_277, n_335);
  nand g22 (n_585, n_277, n_335);
  nor g23 (n_594, n_276, n_334);
  nand g24 (n_589, n_276, n_334);
  nor g25 (n_590, n_275, n_333);
  nand g26 (n_591, n_275, n_333);
  nor g27 (n_600, n_274, n_332);
  nand g28 (n_595, n_274, n_332);
  nor g29 (n_596, n_273, n_331);
  nand g30 (n_597, n_273, n_331);
  nor g31 (n_606, n_272, n_330);
  nand g32 (n_601, n_272, n_330);
  nor g33 (n_602, n_271, n_329);
  nand g34 (n_603, n_271, n_329);
  nor g35 (n_612, n_270, n_328);
  nand g36 (n_607, n_270, n_328);
  nor g37 (n_608, n_269, n_327);
  nand g38 (n_609, n_269, n_327);
  nor g39 (n_618, n_268, n_326);
  nand g40 (n_613, n_268, n_326);
  nor g41 (n_614, n_267, n_325);
  nand g42 (n_615, n_267, n_325);
  nor g43 (n_624, n_266, n_324);
  nand g44 (n_619, n_266, n_324);
  nor g45 (n_620, n_265, n_323);
  nand g46 (n_621, n_265, n_323);
  nor g47 (n_630, n_264, n_322);
  nand g48 (n_625, n_264, n_322);
  nor g49 (n_626, n_263, n_321);
  nand g50 (n_627, n_263, n_321);
  nor g51 (n_636, n_262, n_320);
  nand g52 (n_631, n_262, n_320);
  nor g53 (n_632, n_261, n_319);
  nand g54 (n_633, n_261, n_319);
  nor g55 (n_642, n_260, n_318);
  nand g56 (n_637, n_260, n_318);
  nor g57 (n_638, n_259, n_317);
  nand g58 (n_639, n_259, n_317);
  nor g383 (n_648, n_258, n_316);
  nand g384 (n_643, n_258, n_316);
  nor g385 (n_644, n_257, n_315);
  nand g386 (n_645, n_257, n_315);
  nor g387 (n_654, n_256, n_314);
  nand g388 (n_649, n_256, n_314);
  nor g389 (n_650, n_255, n_313);
  nand g390 (n_651, n_255, n_313);
  nor g391 (n_660, n_254, n_312);
  nand g392 (n_655, n_254, n_312);
  nor g393 (n_656, n_253, n_311);
  nand g394 (n_657, n_253, n_311);
  nor g395 (n_665, n_252, n_310);
  nand g396 (n_661, n_252, n_310);
  nor g397 (n_662, n_251, n_309);
  nand g398 (n_663, n_251, n_309);
  nor g399 (n_671, n_250, n_308);
  nand g400 (n_666, n_250, n_308);
  nor g401 (n_667, n_249, n_307);
  nand g402 (n_668, n_249, n_307);
  nor g403 (n_677, n_248, n_306);
  nand g404 (n_672, n_248, n_306);
  nor g405 (n_673, n_247, n_305);
  nand g406 (n_674, n_247, n_305);
  nor g407 (n_683, n_246, n_304);
  nand g408 (n_678, n_246, n_304);
  nor g409 (n_679, n_245, n_303);
  nand g410 (n_680, n_245, n_303);
  nor g411 (n_689, n_244, n_302);
  nand g412 (n_684, n_244, n_302);
  nor g413 (n_685, n_243, n_301);
  nand g414 (n_686, n_243, n_301);
  nor g415 (n_695, n_242, n_300);
  nand g416 (n_690, n_242, n_300);
  nor g417 (n_691, n_241, n_299);
  nand g418 (n_692, n_241, n_299);
  nor g419 (n_701, n_240, n_298);
  nand g420 (n_696, n_240, n_298);
  nor g421 (n_697, n_239, n_297);
  nand g422 (n_698, n_239, n_297);
  nor g423 (n_707, n_238, n_296);
  nand g424 (n_702, n_238, n_296);
  nor g425 (n_703, n_237, n_295);
  nand g426 (n_704, n_237, n_295);
  nor g427 (n_713, n_236, n_294);
  nand g428 (n_708, n_236, n_294);
  nor g429 (n_709, n_235, n_293);
  nand g430 (n_710, n_235, n_293);
  nor g431 (n_719, n_234, n_292);
  nand g432 (n_714, n_234, n_292);
  nor g433 (n_715, n_233, n_291);
  nand g434 (n_716, n_233, n_291);
  nor g435 (n_725, n_232, n_290);
  nand g436 (n_720, n_232, n_290);
  nor g437 (n_721, n_231, n_289);
  nand g438 (n_722, n_231, n_289);
  nor g439 (n_731, n_230, n_288);
  nand g440 (n_726, n_230, n_288);
  nor g441 (n_727, n_229, n_287);
  nand g442 (n_728, n_229, n_287);
  nor g450 (n_574, n_571, n_572);
  nor g454 (n_580, n_577, n_578);
  nor g457 (n_745, n_582, n_578);
  nor g458 (n_586, n_583, n_584);
  nor g461 (n_747, n_588, n_584);
  nor g462 (n_592, n_589, n_590);
  nor g465 (n_755, n_594, n_590);
  nor g466 (n_598, n_595, n_596);
  nor g469 (n_757, n_600, n_596);
  nor g470 (n_604, n_601, n_602);
  nor g473 (n_765, n_606, n_602);
  nor g474 (n_610, n_607, n_608);
  nor g477 (n_767, n_612, n_608);
  nor g478 (n_616, n_613, n_614);
  nor g481 (n_775, n_618, n_614);
  nor g482 (n_622, n_619, n_620);
  nor g485 (n_777, n_624, n_620);
  nor g486 (n_628, n_625, n_626);
  nor g489 (n_785, n_630, n_626);
  nor g490 (n_634, n_631, n_632);
  nor g493 (n_787, n_636, n_632);
  nor g494 (n_640, n_637, n_638);
  nor g497 (n_795, n_642, n_638);
  nor g498 (n_646, n_643, n_644);
  nor g501 (n_797, n_648, n_644);
  nor g502 (n_652, n_649, n_650);
  nor g505 (n_805, n_654, n_650);
  nor g506 (n_658, n_655, n_656);
  nor g509 (n_807, n_660, n_656);
  nor g510 (n_664, n_661, n_662);
  nor g513 (n_815, n_665, n_662);
  nor g514 (n_669, n_666, n_667);
  nor g517 (n_817, n_671, n_667);
  nor g518 (n_675, n_672, n_673);
  nor g521 (n_825, n_677, n_673);
  nor g522 (n_681, n_678, n_679);
  nor g525 (n_827, n_683, n_679);
  nor g526 (n_687, n_684, n_685);
  nor g529 (n_835, n_689, n_685);
  nor g530 (n_693, n_690, n_691);
  nor g533 (n_837, n_695, n_691);
  nor g534 (n_699, n_696, n_697);
  nor g537 (n_845, n_701, n_697);
  nor g538 (n_705, n_702, n_703);
  nor g541 (n_847, n_707, n_703);
  nor g542 (n_711, n_708, n_709);
  nor g545 (n_855, n_713, n_709);
  nor g546 (n_717, n_714, n_715);
  nor g549 (n_857, n_719, n_715);
  nor g550 (n_723, n_720, n_721);
  nor g553 (n_865, n_725, n_721);
  nor g554 (n_729, n_726, n_727);
  nor g557 (n_867, n_731, n_727);
  nor g563 (n_743, n_588, n_742);
  nand g572 (n_880, n_745, n_747);
  nor g573 (n_753, n_600, n_752);
  nand g582 (n_887, n_755, n_757);
  nor g583 (n_763, n_612, n_762);
  nand g592 (n_895, n_765, n_767);
  nor g593 (n_773, n_624, n_772);
  nand g602 (n_902, n_775, n_777);
  nor g603 (n_783, n_636, n_782);
  nand g612 (n_910, n_785, n_787);
  nor g613 (n_793, n_648, n_792);
  nand g622 (n_917, n_795, n_797);
  nor g623 (n_803, n_660, n_802);
  nand g632 (n_925, n_805, n_807);
  nor g633 (n_813, n_671, n_812);
  nand g642 (n_932, n_815, n_817);
  nor g643 (n_823, n_683, n_822);
  nand g652 (n_940, n_825, n_827);
  nor g653 (n_833, n_695, n_832);
  nand g662 (n_947, n_835, n_837);
  nor g663 (n_843, n_707, n_842);
  nand g672 (n_955, n_845, n_847);
  nor g673 (n_853, n_719, n_852);
  nand g682 (n_962, n_855, n_857);
  nor g683 (n_863, n_731, n_862);
  nand g692 (n_970, n_865, n_867);
  nand g695 (n_1244, n_577, n_874);
  nand g697 (n_1246, n_742, n_875);
  nand g700 (n_1249, n_878, n_879);
  nand g703 (n_974, n_882, n_883);
  nor g704 (n_885, n_606, n_884);
  nor g707 (n_984, n_606, n_887);
  nor g713 (n_893, n_891, n_884);
  nor g716 (n_990, n_887, n_891);
  nor g717 (n_897, n_895, n_884);
  nor g720 (n_993, n_887, n_895);
  nor g721 (n_900, n_630, n_899);
  nor g724 (n_1083, n_630, n_902);
  nor g730 (n_908, n_906, n_899);
  nor g733 (n_1089, n_902, n_906);
  nor g734 (n_912, n_910, n_899);
  nor g737 (n_999, n_902, n_910);
  nor g738 (n_915, n_654, n_914);
  nor g741 (n_1012, n_654, n_917);
  nor g747 (n_923, n_921, n_914);
  nor g750 (n_1022, n_917, n_921);
  nor g751 (n_927, n_925, n_914);
  nor g754 (n_1027, n_917, n_925);
  nor g755 (n_930, n_677, n_929);
  nor g758 (n_1170, n_677, n_932);
  nor g764 (n_938, n_936, n_929);
  nor g767 (n_1176, n_932, n_936);
  nor g768 (n_942, n_940, n_929);
  nor g771 (n_1035, n_932, n_940);
  nor g772 (n_945, n_701, n_944);
  nor g775 (n_1048, n_701, n_947);
  nor g781 (n_953, n_951, n_944);
  nor g784 (n_1058, n_947, n_951);
  nor g785 (n_957, n_955, n_944);
  nor g788 (n_1063, n_947, n_955);
  nor g789 (n_960, n_725, n_959);
  nor g792 (n_1138, n_725, n_962);
  nor g798 (n_968, n_966, n_959);
  nor g801 (n_1148, n_962, n_966);
  nor g802 (n_972, n_970, n_959);
  nor g805 (n_1071, n_962, n_970);
  nand g808 (n_1253, n_589, n_976);
  nand g809 (n_977, n_755, n_974);
  nand g810 (n_1255, n_752, n_977);
  nand g813 (n_1258, n_980, n_981);
  nand g816 (n_1261, n_884, n_983);
  nand g817 (n_986, n_984, n_974);
  nand g818 (n_1264, n_985, n_986);
  nand g819 (n_989, n_987, n_974);
  nand g820 (n_1266, n_988, n_989);
  nand g821 (n_992, n_990, n_974);
  nand g822 (n_1269, n_991, n_992);
  nand g823 (n_995, n_993, n_974);
  nand g824 (n_1073, n_994, n_995);
  nor g825 (n_997, n_642, n_996);
  nand g834 (n_1097, n_795, n_999);
  nor g835 (n_1006, n_1004, n_996);
  nor g840 (n_1009, n_917, n_996);
  nand g849 (n_1109, n_999, n_1012);
  nand g854 (n_1113, n_999, n_1017);
  nand g859 (n_1117, n_999, n_1022);
  nand g864 (n_1121, n_999, n_1027);
  nor g865 (n_1033, n_689, n_1032);
  nand g874 (n_1184, n_835, n_1035);
  nor g875 (n_1042, n_1040, n_1032);
  nor g880 (n_1045, n_947, n_1032);
  nand g889 (n_1196, n_1035, n_1048);
  nand g894 (n_1200, n_1035, n_1053);
  nand g899 (n_1204, n_1035, n_1058);
  nand g904 (n_1128, n_1035, n_1063);
  nor g905 (n_1069, n_735, n_1068);
  nand g912 (n_1273, n_613, n_1075);
  nand g913 (n_1076, n_775, n_1073);
  nand g914 (n_1275, n_772, n_1076);
  nand g917 (n_1278, n_1079, n_1080);
  nand g920 (n_1281, n_899, n_1082);
  nand g921 (n_1085, n_1083, n_1073);
  nand g922 (n_1284, n_1084, n_1085);
  nand g923 (n_1088, n_1086, n_1073);
  nand g924 (n_1286, n_1087, n_1088);
  nand g925 (n_1091, n_1089, n_1073);
  nand g926 (n_1289, n_1090, n_1091);
  nand g927 (n_1092, n_999, n_1073);
  nand g928 (n_1291, n_996, n_1092);
  nand g931 (n_1294, n_1095, n_1096);
  nand g934 (n_1296, n_1099, n_1100);
  nand g937 (n_1299, n_1103, n_1104);
  nand g940 (n_1302, n_1107, n_1108);
  nand g943 (n_1305, n_1111, n_1112);
  nand g946 (n_1307, n_1115, n_1116);
  nand g949 (n_1310, n_1119, n_1120);
  nand g952 (n_1160, n_1123, n_1124);
  nor g953 (n_1126, n_713, n_1125);
  nor g956 (n_1210, n_713, n_1128);
  nor g962 (n_1134, n_1132, n_1125);
  nor g965 (n_1216, n_1132, n_1128);
  nor g966 (n_1136, n_962, n_1125);
  nor g969 (n_1219, n_962, n_1128);
  nor g990 (n_1158, n_1156, n_1125);
  nor g993 (n_1234, n_1128, n_1156);
  nand g996 (n_1314, n_661, n_1162);
  nand g997 (n_1163, n_815, n_1160);
  nand g998 (n_1316, n_812, n_1163);
  nand g1001 (n_1319, n_1166, n_1167);
  nand g1004 (n_1322, n_929, n_1169);
  nand g1005 (n_1172, n_1170, n_1160);
  nand g1006 (n_1325, n_1171, n_1172);
  nand g1007 (n_1175, n_1173, n_1160);
  nand g1008 (n_1327, n_1174, n_1175);
  nand g1009 (n_1178, n_1176, n_1160);
  nand g1010 (n_1330, n_1177, n_1178);
  nand g1011 (n_1179, n_1035, n_1160);
  nand g1012 (n_1332, n_1032, n_1179);
  nand g1015 (n_1335, n_1182, n_1183);
  nand g1018 (n_1337, n_1186, n_1187);
  nand g1021 (n_1340, n_1190, n_1191);
  nand g1024 (n_1343, n_1194, n_1195);
  nand g1027 (n_1346, n_1198, n_1199);
  nand g1030 (n_1348, n_1202, n_1203);
  nand g1033 (n_1351, n_1206, n_1207);
  nand g1036 (n_1354, n_1125, n_1209);
  nand g1037 (n_1212, n_1210, n_1160);
  nand g1038 (n_1357, n_1211, n_1212);
  nand g1039 (n_1215, n_1213, n_1160);
  nand g1040 (n_1359, n_1214, n_1215);
  nand g1041 (n_1218, n_1216, n_1160);
  nand g1042 (n_1362, n_1217, n_1218);
  nand g1043 (n_1221, n_1219, n_1160);
  nand g1044 (n_1365, n_1220, n_1221);
  nand g1045 (n_1224, n_1222, n_1160);
  nand g1046 (n_1368, n_1223, n_1224);
  nand g1047 (n_1227, n_1225, n_1160);
  nand g1048 (n_1370, n_1226, n_1227);
  nand g1049 (n_1230, n_1228, n_1160);
  nand g1050 (n_1373, n_1229, n_1230);
  nand g1051 (n_1233, n_1231, n_1160);
  nand g1052 (n_1375, n_1232, n_1233);
  nand g1053 (n_1236, n_1234, n_1160);
  nand g1054 (n_1378, n_1235, n_1236);
  xnor g1066 (out_0[5], n_1244, n_1245);
  xnor g1068 (out_0[6], n_1246, n_1247);
  xnor g1071 (out_0[7], n_1249, n_1250);
  xnor g1073 (out_0[8], n_974, n_1251);
  xnor g1076 (out_0[9], n_1253, n_1254);
  xnor g1078 (out_0[10], n_1255, n_1256);
  xnor g1081 (out_0[11], n_1258, n_1259);
  xnor g1084 (out_0[12], n_1261, n_1262);
  xnor g1087 (out_0[13], n_1264, n_1265);
  xnor g1089 (out_0[14], n_1266, n_1267);
  xnor g1092 (out_0[15], n_1269, n_1270);
  xnor g1094 (out_0[16], n_1073, n_1271);
  xnor g1097 (out_0[17], n_1273, n_1274);
  xnor g1099 (out_0[18], n_1275, n_1276);
  xnor g1102 (out_0[19], n_1278, n_1279);
  xnor g1105 (out_0[20], n_1281, n_1282);
  xnor g1108 (out_0[21], n_1284, n_1285);
  xnor g1110 (out_0[22], n_1286, n_1287);
  xnor g1113 (out_0[23], n_1289, n_1290);
  xnor g1115 (out_0[24], n_1291, n_1292);
  xnor g1118 (out_0[25], n_1294, n_1295);
  xnor g1120 (out_0[26], n_1296, n_1297);
  xnor g1123 (out_0[27], n_1299, n_1300);
  xnor g1126 (out_0[28], n_1302, n_1303);
  xnor g1129 (out_0[29], n_1305, n_1306);
  xnor g1131 (out_0[30], n_1307, n_1308);
  xnor g1134 (out_0[31], n_1310, n_1311);
  xnor g1136 (out_0[32], n_1160, n_1312);
  xnor g1139 (out_0[33], n_1314, n_1315);
  xnor g1141 (out_0[34], n_1316, n_1317);
  xnor g1144 (out_0[35], n_1319, n_1320);
  xnor g1147 (out_0[36], n_1322, n_1323);
  xnor g1150 (out_0[37], n_1325, n_1326);
  xnor g1152 (out_0[38], n_1327, n_1328);
  xnor g1155 (out_0[39], n_1330, n_1331);
  xnor g1157 (out_0[40], n_1332, n_1333);
  xnor g1160 (out_0[41], n_1335, n_1336);
  xnor g1162 (out_0[42], n_1337, n_1338);
  xnor g1165 (out_0[43], n_1340, n_1341);
  xnor g1168 (out_0[44], n_1343, n_1344);
  xnor g1171 (out_0[45], n_1346, n_1347);
  xnor g1173 (out_0[46], n_1348, n_1349);
  xnor g1176 (out_0[47], n_1351, n_1352);
  xnor g1179 (out_0[48], n_1354, n_1355);
  xnor g1182 (out_0[49], n_1357, n_1358);
  xnor g1184 (out_0[50], n_1359, n_1360);
  xnor g1187 (out_0[51], n_1362, n_1363);
  xnor g1190 (out_0[52], n_1365, n_1366);
  xnor g1193 (out_0[53], n_1368, n_1369);
  xnor g1195 (out_0[54], n_1370, n_1371);
  xnor g1198 (out_0[55], n_1373, n_1374);
  xnor g1200 (out_0[56], n_1375, n_1376);
  xor g1205 (n_557, in_1[55], in_2[55]);
  or g1206 (n_558, in_1[55], in_2[55]);
  or g1207 (n_559, in_2[55], wc);
  not gc (wc, in_0[55]);
  or g1208 (n_560, in_1[55], wc0);
  not gc0 (wc0, in_0[55]);
  or g1209 (n_1238, wc1, n_576);
  not gc1 (wc1, n_571);
  and g1210 (n_735, in_0[55], wc2);
  not gc2 (wc2, n_286);
  or g1211 (n_732, in_0[55], wc3);
  not gc3 (wc3, n_286);
  and g1212 (n_740, wc4, n_573);
  not gc4 (wc4, n_574);
  and g1213 (n_742, wc5, n_579);
  not gc5 (wc5, n_580);
  and g1214 (n_749, wc6, n_585);
  not gc6 (wc6, n_586);
  and g1215 (n_752, wc7, n_591);
  not gc7 (wc7, n_592);
  and g1216 (n_759, wc8, n_597);
  not gc8 (wc8, n_598);
  and g1217 (n_762, wc9, n_603);
  not gc9 (wc9, n_604);
  and g1218 (n_769, wc10, n_609);
  not gc10 (wc10, n_610);
  and g1219 (n_772, wc11, n_615);
  not gc11 (wc11, n_616);
  and g1220 (n_779, wc12, n_621);
  not gc12 (wc12, n_622);
  and g1221 (n_782, wc13, n_627);
  not gc13 (wc13, n_628);
  and g1222 (n_789, wc14, n_633);
  not gc14 (wc14, n_634);
  and g1223 (n_792, wc15, n_639);
  not gc15 (wc15, n_640);
  and g1224 (n_799, wc16, n_645);
  not gc16 (wc16, n_646);
  and g1225 (n_802, wc17, n_651);
  not gc17 (wc17, n_652);
  and g1226 (n_809, wc18, n_657);
  not gc18 (wc18, n_658);
  and g1227 (n_812, wc19, n_663);
  not gc19 (wc19, n_664);
  and g1228 (n_819, wc20, n_668);
  not gc20 (wc20, n_669);
  and g1229 (n_822, wc21, n_674);
  not gc21 (wc21, n_675);
  and g1230 (n_829, wc22, n_680);
  not gc22 (wc22, n_681);
  and g1231 (n_832, wc23, n_686);
  not gc23 (wc23, n_687);
  and g1232 (n_839, wc24, n_692);
  not gc24 (wc24, n_693);
  and g1233 (n_842, wc25, n_698);
  not gc25 (wc25, n_699);
  and g1234 (n_849, wc26, n_704);
  not gc26 (wc26, n_705);
  and g1235 (n_852, wc27, n_710);
  not gc27 (wc27, n_711);
  and g1236 (n_859, wc28, n_716);
  not gc28 (wc28, n_717);
  and g1237 (n_862, wc29, n_722);
  not gc29 (wc29, n_723);
  or g1238 (n_876, wc30, n_588);
  not gc30 (wc30, n_745);
  or g1239 (n_978, wc31, n_600);
  not gc31 (wc31, n_755);
  or g1240 (n_891, wc32, n_612);
  not gc32 (wc32, n_765);
  or g1241 (n_1077, wc33, n_624);
  not gc33 (wc33, n_775);
  or g1242 (n_906, wc34, n_636);
  not gc34 (wc34, n_785);
  or g1243 (n_1004, wc35, n_648);
  not gc35 (wc35, n_795);
  or g1244 (n_921, wc36, n_660);
  not gc36 (wc36, n_805);
  or g1245 (n_1164, wc37, n_671);
  not gc37 (wc37, n_815);
  or g1246 (n_936, wc38, n_683);
  not gc38 (wc38, n_825);
  or g1247 (n_1040, wc39, n_695);
  not gc39 (wc39, n_835);
  or g1248 (n_951, wc40, n_707);
  not gc40 (wc40, n_845);
  or g1249 (n_1132, wc41, n_719);
  not gc41 (wc41, n_855);
  or g1250 (n_966, wc42, n_731);
  not gc42 (wc42, n_865);
  not g1251 (out_0[2], n_1238);
  or g1252 (n_1241, wc43, n_572);
  not gc43 (wc43, n_573);
  or g1253 (n_1242, wc44, n_582);
  not gc44 (wc44, n_577);
  or g1254 (n_1245, wc45, n_578);
  not gc45 (wc45, n_579);
  or g1255 (n_1247, wc46, n_588);
  not gc46 (wc46, n_583);
  or g1256 (n_1250, wc47, n_584);
  not gc47 (wc47, n_585);
  or g1257 (n_1251, wc48, n_594);
  not gc48 (wc48, n_589);
  or g1258 (n_1254, wc49, n_590);
  not gc49 (wc49, n_591);
  or g1259 (n_1256, wc50, n_600);
  not gc50 (wc50, n_595);
  or g1260 (n_1259, wc51, n_596);
  not gc51 (wc51, n_597);
  or g1261 (n_1262, wc52, n_606);
  not gc52 (wc52, n_601);
  or g1262 (n_1265, wc53, n_602);
  not gc53 (wc53, n_603);
  or g1263 (n_1267, wc54, n_612);
  not gc54 (wc54, n_607);
  or g1264 (n_1270, wc55, n_608);
  not gc55 (wc55, n_609);
  or g1265 (n_1271, wc56, n_618);
  not gc56 (wc56, n_613);
  or g1266 (n_1274, wc57, n_614);
  not gc57 (wc57, n_615);
  or g1267 (n_1276, wc58, n_624);
  not gc58 (wc58, n_619);
  or g1268 (n_1279, wc59, n_620);
  not gc59 (wc59, n_621);
  or g1269 (n_1282, wc60, n_630);
  not gc60 (wc60, n_625);
  or g1270 (n_1285, wc61, n_626);
  not gc61 (wc61, n_627);
  or g1271 (n_1287, wc62, n_636);
  not gc62 (wc62, n_631);
  or g1272 (n_1290, wc63, n_632);
  not gc63 (wc63, n_633);
  or g1273 (n_1292, wc64, n_642);
  not gc64 (wc64, n_637);
  or g1274 (n_1295, wc65, n_638);
  not gc65 (wc65, n_639);
  or g1275 (n_1297, wc66, n_648);
  not gc66 (wc66, n_643);
  or g1276 (n_1300, wc67, n_644);
  not gc67 (wc67, n_645);
  or g1277 (n_1303, wc68, n_654);
  not gc68 (wc68, n_649);
  or g1278 (n_1306, wc69, n_650);
  not gc69 (wc69, n_651);
  or g1279 (n_1308, wc70, n_660);
  not gc70 (wc70, n_655);
  or g1280 (n_1311, wc71, n_656);
  not gc71 (wc71, n_657);
  or g1281 (n_1312, wc72, n_665);
  not gc72 (wc72, n_661);
  or g1282 (n_1315, wc73, n_662);
  not gc73 (wc73, n_663);
  or g1283 (n_1317, wc74, n_671);
  not gc74 (wc74, n_666);
  or g1284 (n_1320, wc75, n_667);
  not gc75 (wc75, n_668);
  or g1285 (n_1323, wc76, n_677);
  not gc76 (wc76, n_672);
  or g1286 (n_1326, wc77, n_673);
  not gc77 (wc77, n_674);
  or g1287 (n_1328, wc78, n_683);
  not gc78 (wc78, n_678);
  or g1288 (n_1331, wc79, n_679);
  not gc79 (wc79, n_680);
  or g1289 (n_1333, wc80, n_689);
  not gc80 (wc80, n_684);
  or g1290 (n_1336, wc81, n_685);
  not gc81 (wc81, n_686);
  or g1291 (n_1338, wc82, n_695);
  not gc82 (wc82, n_690);
  or g1292 (n_1341, wc83, n_691);
  not gc83 (wc83, n_692);
  or g1293 (n_1344, wc84, n_701);
  not gc84 (wc84, n_696);
  or g1294 (n_1347, wc85, n_697);
  not gc85 (wc85, n_698);
  or g1295 (n_1349, wc86, n_707);
  not gc86 (wc86, n_702);
  or g1296 (n_1352, wc87, n_703);
  not gc87 (wc87, n_704);
  or g1297 (n_1355, wc88, n_713);
  not gc88 (wc88, n_708);
  or g1298 (n_1358, wc89, n_709);
  not gc89 (wc89, n_710);
  or g1299 (n_1360, wc90, n_719);
  not gc90 (wc90, n_714);
  or g1300 (n_1363, wc91, n_715);
  not gc91 (wc91, n_716);
  or g1301 (n_1366, wc92, n_725);
  not gc92 (wc92, n_720);
  or g1302 (n_1369, wc93, n_721);
  not gc93 (wc93, n_722);
  or g1303 (n_1371, wc94, n_731);
  not gc94 (wc94, n_726);
  and g1304 (n_869, wc95, n_728);
  not gc95 (wc95, n_729);
  and g1307 (n_750, wc96, n_747);
  not gc96 (wc96, n_742);
  and g1308 (n_760, wc97, n_757);
  not gc97 (wc97, n_752);
  and g1309 (n_770, wc98, n_767);
  not gc98 (wc98, n_762);
  and g1310 (n_780, wc99, n_777);
  not gc99 (wc99, n_772);
  and g1311 (n_790, wc100, n_787);
  not gc100 (wc100, n_782);
  and g1312 (n_800, wc101, n_797);
  not gc101 (wc101, n_792);
  and g1313 (n_810, wc102, n_807);
  not gc102 (wc102, n_802);
  and g1314 (n_820, wc103, n_817);
  not gc103 (wc103, n_812);
  and g1315 (n_830, wc104, n_827);
  not gc104 (wc104, n_822);
  and g1316 (n_840, wc105, n_837);
  not gc105 (wc105, n_832);
  and g1317 (n_850, wc106, n_847);
  not gc106 (wc106, n_842);
  and g1318 (n_860, wc107, n_857);
  not gc107 (wc107, n_852);
  and g1319 (n_987, wc108, n_765);
  not gc108 (wc108, n_887);
  and g1320 (n_1086, wc109, n_785);
  not gc109 (wc109, n_902);
  and g1321 (n_1017, wc110, n_805);
  not gc110 (wc110, n_917);
  and g1322 (n_1173, wc111, n_825);
  not gc111 (wc111, n_932);
  and g1323 (n_1053, wc112, n_845);
  not gc112 (wc112, n_947);
  and g1324 (n_1143, wc113, n_865);
  not gc113 (wc113, n_962);
  or g1325 (n_1374, wc114, n_727);
  not gc114 (wc114, n_728);
  and g1326 (n_878, wc115, n_583);
  not gc115 (wc115, n_743);
  and g1327 (n_882, wc116, n_749);
  not gc116 (wc116, n_750);
  and g1328 (n_980, wc117, n_595);
  not gc117 (wc117, n_753);
  and g1329 (n_884, wc118, n_759);
  not gc118 (wc118, n_760);
  and g1330 (n_892, wc119, n_607);
  not gc119 (wc119, n_763);
  and g1331 (n_896, wc120, n_769);
  not gc120 (wc120, n_770);
  and g1332 (n_1079, wc121, n_619);
  not gc121 (wc121, n_773);
  and g1333 (n_899, wc122, n_779);
  not gc122 (wc122, n_780);
  and g1334 (n_907, wc123, n_631);
  not gc123 (wc123, n_783);
  and g1335 (n_911, wc124, n_789);
  not gc124 (wc124, n_790);
  and g1336 (n_1005, wc125, n_643);
  not gc125 (wc125, n_793);
  and g1337 (n_914, wc126, n_799);
  not gc126 (wc126, n_800);
  and g1338 (n_922, wc127, n_655);
  not gc127 (wc127, n_803);
  and g1339 (n_926, wc128, n_809);
  not gc128 (wc128, n_810);
  and g1340 (n_1166, wc129, n_666);
  not gc129 (wc129, n_813);
  and g1341 (n_929, wc130, n_819);
  not gc130 (wc130, n_820);
  and g1342 (n_937, wc131, n_678);
  not gc131 (wc131, n_823);
  and g1343 (n_941, wc132, n_829);
  not gc132 (wc132, n_830);
  and g1344 (n_1041, wc133, n_690);
  not gc133 (wc133, n_833);
  and g1345 (n_944, wc134, n_839);
  not gc134 (wc134, n_840);
  and g1346 (n_952, wc135, n_702);
  not gc135 (wc135, n_843);
  and g1347 (n_956, wc136, n_849);
  not gc136 (wc136, n_850);
  and g1348 (n_1133, wc137, n_714);
  not gc137 (wc137, n_853);
  and g1349 (n_959, wc138, n_859);
  not gc138 (wc138, n_860);
  and g1350 (n_967, wc139, n_726);
  not gc139 (wc139, n_863);
  and g1351 (n_870, wc140, n_867);
  not gc140 (wc140, n_862);
  or g1352 (n_874, n_582, n_740);
  or g1353 (n_875, n_740, wc141);
  not gc141 (wc141, n_745);
  or g1354 (n_879, n_740, n_876);
  or g1355 (n_883, n_880, n_740);
  or g1356 (n_1093, wc142, n_642);
  not gc142 (wc142, n_999);
  or g1357 (n_1101, n_1004, wc143);
  not gc143 (wc143, n_999);
  or g1358 (n_1105, wc144, n_917);
  not gc144 (wc144, n_999);
  or g1359 (n_1180, wc145, n_689);
  not gc145 (wc145, n_1035);
  or g1360 (n_1188, n_1040, wc146);
  not gc146 (wc146, n_1035);
  or g1361 (n_1192, wc147, n_947);
  not gc147 (wc147, n_1035);
  xor g1362 (out_0[3], n_571, n_1241);
  xor g1363 (out_0[4], n_740, n_1242);
  or g1364 (n_1376, wc148, n_735);
  not gc148 (wc148, n_732);
  and g1365 (n_971, wc149, n_869);
  not gc149 (wc149, n_870);
  and g1366 (n_889, wc150, n_765);
  not gc150 (wc150, n_884);
  and g1367 (n_904, wc151, n_785);
  not gc151 (wc151, n_899);
  and g1368 (n_919, wc152, n_805);
  not gc152 (wc152, n_914);
  and g1369 (n_934, wc153, n_825);
  not gc153 (wc153, n_929);
  and g1370 (n_949, wc154, n_845);
  not gc154 (wc154, n_944);
  and g1371 (n_964, wc155, n_865);
  not gc155 (wc155, n_959);
  or g1372 (n_1156, n_735, wc156);
  not gc156 (wc156, n_1071);
  and g1373 (n_1213, wc157, n_855);
  not gc157 (wc157, n_1128);
  and g1374 (n_1222, wc158, n_1138);
  not gc158 (wc158, n_1128);
  and g1375 (n_1225, n_1143, wc159);
  not gc159 (wc159, n_1128);
  and g1376 (n_1228, wc160, n_1148);
  not gc160 (wc160, n_1128);
  and g1377 (n_985, wc161, n_601);
  not gc161 (wc161, n_885);
  and g1378 (n_988, wc162, n_762);
  not gc162 (wc162, n_889);
  and g1379 (n_991, n_892, wc163);
  not gc163 (wc163, n_893);
  and g1380 (n_994, n_896, wc164);
  not gc164 (wc164, n_897);
  and g1381 (n_1084, wc165, n_625);
  not gc165 (wc165, n_900);
  and g1382 (n_1087, wc166, n_782);
  not gc166 (wc166, n_904);
  and g1383 (n_1090, n_907, wc167);
  not gc167 (wc167, n_908);
  and g1384 (n_996, n_911, wc168);
  not gc168 (wc168, n_912);
  and g1385 (n_1014, wc169, n_649);
  not gc169 (wc169, n_915);
  and g1386 (n_1019, wc170, n_802);
  not gc170 (wc170, n_919);
  and g1387 (n_1024, n_922, wc171);
  not gc171 (wc171, n_923);
  and g1388 (n_1029, n_926, wc172);
  not gc172 (wc172, n_927);
  and g1389 (n_1171, wc173, n_672);
  not gc173 (wc173, n_930);
  and g1390 (n_1174, wc174, n_822);
  not gc174 (wc174, n_934);
  and g1391 (n_1177, n_937, wc175);
  not gc175 (wc175, n_938);
  and g1392 (n_1032, n_941, wc176);
  not gc176 (wc176, n_942);
  and g1393 (n_1050, wc177, n_696);
  not gc177 (wc177, n_945);
  and g1394 (n_1055, wc178, n_842);
  not gc178 (wc178, n_949);
  and g1395 (n_1060, n_952, wc179);
  not gc179 (wc179, n_953);
  and g1396 (n_1065, n_956, wc180);
  not gc180 (wc180, n_957);
  and g1397 (n_1140, wc181, n_720);
  not gc181 (wc181, n_960);
  and g1398 (n_1145, wc182, n_862);
  not gc182 (wc182, n_964);
  and g1399 (n_1150, n_967, wc183);
  not gc183 (wc183, n_968);
  or g1400 (n_976, wc184, n_594);
  not gc184 (wc184, n_974);
  or g1401 (n_981, n_978, wc185);
  not gc185 (wc185, n_974);
  or g1402 (n_983, wc186, n_887);
  not gc186 (wc186, n_974);
  and g1403 (n_1231, wc187, n_1071);
  not gc187 (wc187, n_1128);
  and g1404 (n_1068, n_971, wc188);
  not gc188 (wc188, n_972);
  and g1405 (n_1002, wc189, n_795);
  not gc189 (wc189, n_996);
  and g1406 (n_1015, wc190, n_1012);
  not gc190 (wc190, n_996);
  and g1407 (n_1020, wc191, n_1017);
  not gc191 (wc191, n_996);
  and g1408 (n_1025, wc192, n_1022);
  not gc192 (wc192, n_996);
  and g1409 (n_1030, wc193, n_1027);
  not gc193 (wc193, n_996);
  and g1410 (n_1038, wc194, n_835);
  not gc194 (wc194, n_1032);
  and g1411 (n_1051, wc195, n_1048);
  not gc195 (wc195, n_1032);
  and g1412 (n_1056, wc196, n_1053);
  not gc196 (wc196, n_1032);
  and g1413 (n_1061, wc197, n_1058);
  not gc197 (wc197, n_1032);
  and g1414 (n_1066, wc198, n_1063);
  not gc198 (wc198, n_1032);
  and g1415 (n_1095, wc199, n_637);
  not gc199 (wc199, n_997);
  and g1416 (n_1099, wc200, n_792);
  not gc200 (wc200, n_1002);
  and g1417 (n_1103, n_1005, wc201);
  not gc201 (wc201, n_1006);
  and g1418 (n_1107, n_914, wc202);
  not gc202 (wc202, n_1009);
  and g1419 (n_1111, wc203, n_1014);
  not gc203 (wc203, n_1015);
  and g1420 (n_1115, wc204, n_1019);
  not gc204 (wc204, n_1020);
  and g1421 (n_1119, wc205, n_1024);
  not gc205 (wc205, n_1025);
  and g1422 (n_1123, wc206, n_1029);
  not gc206 (wc206, n_1030);
  and g1423 (n_1182, wc207, n_684);
  not gc207 (wc207, n_1033);
  and g1424 (n_1186, wc208, n_832);
  not gc208 (wc208, n_1038);
  and g1425 (n_1190, n_1041, wc209);
  not gc209 (wc209, n_1042);
  and g1426 (n_1194, n_944, wc210);
  not gc210 (wc210, n_1045);
  and g1427 (n_1198, wc211, n_1050);
  not gc211 (wc211, n_1051);
  and g1428 (n_1202, wc212, n_1055);
  not gc212 (wc212, n_1056);
  and g1429 (n_1206, wc213, n_1060);
  not gc213 (wc213, n_1061);
  and g1430 (n_1125, wc214, n_1065);
  not gc214 (wc214, n_1066);
  or g1431 (n_1075, wc215, n_618);
  not gc215 (wc215, n_1073);
  or g1432 (n_1080, n_1077, wc216);
  not gc216 (wc216, n_1073);
  or g1433 (n_1082, wc217, n_902);
  not gc217 (wc217, n_1073);
  or g1434 (n_1096, n_1093, wc218);
  not gc218 (wc218, n_1073);
  or g1435 (n_1100, n_1097, wc219);
  not gc219 (wc219, n_1073);
  or g1436 (n_1104, n_1101, wc220);
  not gc220 (wc220, n_1073);
  or g1437 (n_1108, n_1105, wc221);
  not gc221 (wc221, n_1073);
  or g1438 (n_1112, n_1109, wc222);
  not gc222 (wc222, n_1073);
  or g1439 (n_1116, n_1113, wc223);
  not gc223 (wc223, n_1073);
  or g1440 (n_1120, n_1117, wc224);
  not gc224 (wc224, n_1073);
  or g1441 (n_1124, n_1121, wc225);
  not gc225 (wc225, n_1073);
  and g1442 (n_1157, n_732, wc226);
  not gc226 (wc226, n_1069);
  and g1443 (n_1130, wc227, n_855);
  not gc227 (wc227, n_1125);
  and g1444 (n_1141, wc228, n_1138);
  not gc228 (wc228, n_1125);
  and g1445 (n_1146, wc229, n_1143);
  not gc229 (wc229, n_1125);
  and g1446 (n_1151, wc230, n_1148);
  not gc230 (wc230, n_1125);
  and g1447 (n_1154, wc231, n_1071);
  not gc231 (wc231, n_1125);
  and g1448 (n_1211, wc232, n_708);
  not gc232 (wc232, n_1126);
  and g1449 (n_1214, wc233, n_852);
  not gc233 (wc233, n_1130);
  and g1450 (n_1217, n_1133, wc234);
  not gc234 (wc234, n_1134);
  and g1451 (n_1220, n_959, wc235);
  not gc235 (wc235, n_1136);
  and g1452 (n_1223, wc236, n_1140);
  not gc236 (wc236, n_1141);
  and g1453 (n_1226, wc237, n_1145);
  not gc237 (wc237, n_1146);
  and g1454 (n_1229, wc238, n_1150);
  not gc238 (wc238, n_1151);
  and g1455 (n_1232, wc239, n_1068);
  not gc239 (wc239, n_1154);
  or g1456 (n_1162, wc240, n_665);
  not gc240 (wc240, n_1160);
  or g1457 (n_1167, n_1164, wc241);
  not gc241 (wc241, n_1160);
  or g1458 (n_1169, wc242, n_932);
  not gc242 (wc242, n_1160);
  or g1459 (n_1183, n_1180, wc243);
  not gc243 (wc243, n_1160);
  or g1460 (n_1187, wc244, n_1184);
  not gc244 (wc244, n_1160);
  or g1461 (n_1191, n_1188, wc245);
  not gc245 (wc245, n_1160);
  or g1462 (n_1195, n_1192, wc246);
  not gc246 (wc246, n_1160);
  or g1463 (n_1199, wc247, n_1196);
  not gc247 (wc247, n_1160);
  or g1464 (n_1203, wc248, n_1200);
  not gc248 (wc248, n_1160);
  or g1465 (n_1207, wc249, n_1204);
  not gc249 (wc249, n_1160);
  or g1466 (n_1209, wc250, n_1128);
  not gc250 (wc250, n_1160);
  and g1467 (n_1235, n_1157, wc251);
  not gc251 (wc251, n_1158);
  not g1468 (out_0[57], n_1378);
endmodule

module csa_tree_add_607_44_group_16902_GENERIC(in_0, in_1, in_2, out_0);
  input [55:0] in_0, in_1, in_2;
  output [57:0] out_0;
  wire [55:0] in_0, in_1, in_2;
  wire [57:0] out_0;
  csa_tree_add_607_44_group_16902_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module increment_unsigned_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [18:0] A;
  input CI;
  output [18:0] Z;
  wire [18:0] A;
  wire CI;
  wire [18:0] Z;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_40, A[0], CI);
  xor g19 (Z[1], A[1], n_40);
  and g20 (n_41, A[1], n_40);
  xor g21 (Z[2], A[2], n_41);
  and g22 (n_42, A[2], n_41);
  xor g23 (Z[3], A[3], n_42);
  and g24 (n_43, A[3], n_42);
  xor g25 (Z[4], A[4], n_43);
  and g26 (n_44, A[4], n_43);
  xor g27 (Z[5], A[5], n_44);
  and g28 (n_45, A[5], n_44);
  xor g29 (Z[6], A[6], n_45);
  and g30 (n_46, A[6], n_45);
  xor g31 (Z[7], A[7], n_46);
  and g32 (n_47, A[7], n_46);
  xor g33 (Z[8], A[8], n_47);
  and g34 (n_48, A[8], n_47);
  xor g35 (Z[9], A[9], n_48);
  and g36 (n_49, A[9], n_48);
  xor g37 (Z[10], A[10], n_49);
  and g38 (n_50, A[10], n_49);
  xor g39 (Z[11], A[11], n_50);
  and g40 (n_51, A[11], n_50);
  xor g41 (Z[12], A[12], n_51);
  and g42 (n_52, A[12], n_51);
  xor g43 (Z[13], A[13], n_52);
  and g44 (n_53, A[13], n_52);
  xor g45 (Z[14], A[14], n_53);
  and g46 (n_54, A[14], n_53);
  xor g47 (Z[15], A[15], n_54);
  and g48 (n_55, A[15], n_54);
  xor g49 (Z[16], A[16], n_55);
  and g50 (n_56, A[16], n_55);
  xor g51 (Z[17], A[17], n_56);
  and g52 (n_57, A[17], n_56);
  xor g53 (Z[18], A[18], n_57);
endmodule

module increment_unsigned_GENERIC(A, CI, Z);
  input [18:0] A;
  input CI;
  output [18:0] Z;
  wire [18:0] A;
  wire CI;
  wire [18:0] Z;
  increment_unsigned_GENERIC_REAL g1(.A (A), .CI (CI), .Z (Z));
endmodule

module increment_unsigned_1_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [18:0] A;
  input CI;
  output [18:0] Z;
  wire [18:0] A;
  wire CI;
  wire [18:0] Z;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_40, A[0], CI);
  xor g19 (Z[1], A[1], n_40);
  and g20 (n_41, A[1], n_40);
  xor g21 (Z[2], A[2], n_41);
  and g22 (n_42, A[2], n_41);
  xor g23 (Z[3], A[3], n_42);
  and g24 (n_43, A[3], n_42);
  xor g25 (Z[4], A[4], n_43);
  and g26 (n_44, A[4], n_43);
  xor g27 (Z[5], A[5], n_44);
  and g28 (n_45, A[5], n_44);
  xor g29 (Z[6], A[6], n_45);
  and g30 (n_46, A[6], n_45);
  xor g31 (Z[7], A[7], n_46);
  and g32 (n_47, A[7], n_46);
  xor g33 (Z[8], A[8], n_47);
  and g34 (n_48, A[8], n_47);
  xor g35 (Z[9], A[9], n_48);
  and g36 (n_49, A[9], n_48);
  xor g37 (Z[10], A[10], n_49);
  and g38 (n_50, A[10], n_49);
  xor g39 (Z[11], A[11], n_50);
  and g40 (n_51, A[11], n_50);
  xor g41 (Z[12], A[12], n_51);
  and g42 (n_52, A[12], n_51);
  xor g43 (Z[13], A[13], n_52);
  and g44 (n_53, A[13], n_52);
  xor g45 (Z[14], A[14], n_53);
  and g46 (n_54, A[14], n_53);
  xor g47 (Z[15], A[15], n_54);
  and g48 (n_55, A[15], n_54);
  xor g49 (Z[16], A[16], n_55);
  and g50 (n_56, A[16], n_55);
  xor g51 (Z[17], A[17], n_56);
  and g52 (n_57, A[17], n_56);
  xor g53 (Z[18], A[18], n_57);
endmodule

module increment_unsigned_1_GENERIC(A, CI, Z);
  input [18:0] A;
  input CI;
  output [18:0] Z;
  wire [18:0] A;
  wire CI;
  wire [18:0] Z;
  increment_unsigned_1_GENERIC_REAL g1(.A ({A[16], A[16], A[16:0]}),
       .CI (CI), .Z (Z));
endmodule

module increment_unsigned_16827_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [60:0] A;
  input CI;
  output [60:0] Z;
  wire [60:0] A;
  wire CI;
  wire [60:0] Z;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163;
  wire n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171;
  wire n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179;
  wire n_180, n_181, n_182, n_183;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_124, A[0], CI);
  xor g61 (Z[1], A[1], n_124);
  and g62 (n_125, A[1], n_124);
  xor g63 (Z[2], A[2], n_125);
  and g64 (n_126, A[2], n_125);
  xor g65 (Z[3], A[3], n_126);
  and g66 (n_127, A[3], n_126);
  xor g67 (Z[4], A[4], n_127);
  and g68 (n_128, A[4], n_127);
  xor g69 (Z[5], A[5], n_128);
  and g70 (n_129, A[5], n_128);
  xor g71 (Z[6], A[6], n_129);
  and g72 (n_130, A[6], n_129);
  xor g73 (Z[7], A[7], n_130);
  and g74 (n_131, A[7], n_130);
  xor g75 (Z[8], A[8], n_131);
  and g76 (n_132, A[8], n_131);
  xor g77 (Z[9], A[9], n_132);
  and g78 (n_133, A[9], n_132);
  xor g79 (Z[10], A[10], n_133);
  and g80 (n_134, A[10], n_133);
  xor g81 (Z[11], A[11], n_134);
  and g82 (n_135, A[11], n_134);
  xor g83 (Z[12], A[12], n_135);
  and g84 (n_136, A[12], n_135);
  xor g85 (Z[13], A[13], n_136);
  and g86 (n_137, A[13], n_136);
  xor g87 (Z[14], A[14], n_137);
  and g88 (n_138, A[14], n_137);
  xor g89 (Z[15], A[15], n_138);
  and g90 (n_139, A[15], n_138);
  xor g91 (Z[16], A[16], n_139);
  and g92 (n_140, A[16], n_139);
  xor g93 (Z[17], A[17], n_140);
  and g94 (n_141, A[17], n_140);
  xor g95 (Z[18], A[18], n_141);
  and g96 (n_142, A[18], n_141);
  xor g97 (Z[19], A[19], n_142);
  and g98 (n_143, A[19], n_142);
  xor g99 (Z[20], A[20], n_143);
  and g100 (n_144, A[20], n_143);
  xor g101 (Z[21], A[21], n_144);
  and g102 (n_145, A[21], n_144);
  xor g103 (Z[22], A[22], n_145);
  and g104 (n_146, A[22], n_145);
  xor g105 (Z[23], A[23], n_146);
  and g106 (n_147, A[23], n_146);
  xor g107 (Z[24], A[24], n_147);
  and g108 (n_148, A[24], n_147);
  xor g109 (Z[25], A[25], n_148);
  and g110 (n_149, A[25], n_148);
  xor g111 (Z[26], A[26], n_149);
  and g112 (n_150, A[26], n_149);
  xor g113 (Z[27], A[27], n_150);
  and g114 (n_151, A[27], n_150);
  xor g115 (Z[28], A[28], n_151);
  and g116 (n_152, A[28], n_151);
  xor g117 (Z[29], A[29], n_152);
  and g118 (n_153, A[29], n_152);
  xor g119 (Z[30], A[30], n_153);
  and g120 (n_154, A[30], n_153);
  xor g121 (Z[31], A[31], n_154);
  and g122 (n_155, A[31], n_154);
  xor g123 (Z[32], A[32], n_155);
  and g124 (n_156, A[32], n_155);
  xor g125 (Z[33], A[33], n_156);
  and g126 (n_157, A[33], n_156);
  xor g127 (Z[34], A[34], n_157);
  and g128 (n_158, A[34], n_157);
  xor g129 (Z[35], A[35], n_158);
  and g130 (n_159, A[35], n_158);
  xor g131 (Z[36], A[36], n_159);
  and g132 (n_160, A[36], n_159);
  xor g133 (Z[37], A[37], n_160);
  and g134 (n_161, A[37], n_160);
  xor g135 (Z[38], A[38], n_161);
  and g136 (n_162, A[38], n_161);
  xor g137 (Z[39], A[39], n_162);
  and g138 (n_163, A[39], n_162);
  xor g139 (Z[40], A[40], n_163);
  and g140 (n_164, A[40], n_163);
  xor g141 (Z[41], A[41], n_164);
  and g142 (n_165, A[41], n_164);
  xor g143 (Z[42], A[42], n_165);
  and g144 (n_166, A[42], n_165);
  xor g145 (Z[43], A[43], n_166);
  and g146 (n_167, A[43], n_166);
  xor g147 (Z[44], A[44], n_167);
  and g148 (n_168, A[44], n_167);
  xor g149 (Z[45], A[45], n_168);
  and g150 (n_169, A[45], n_168);
  xor g151 (Z[46], A[46], n_169);
  and g152 (n_170, A[46], n_169);
  xor g153 (Z[47], A[47], n_170);
  and g154 (n_171, A[47], n_170);
  xor g155 (Z[48], A[48], n_171);
  and g156 (n_172, A[48], n_171);
  xor g157 (Z[49], A[49], n_172);
  and g158 (n_173, A[49], n_172);
  xor g159 (Z[50], A[50], n_173);
  and g160 (n_174, A[50], n_173);
  xor g161 (Z[51], A[51], n_174);
  and g162 (n_175, A[51], n_174);
  xor g163 (Z[52], A[52], n_175);
  and g164 (n_176, A[52], n_175);
  xor g165 (Z[53], A[53], n_176);
  and g166 (n_177, A[53], n_176);
  xor g167 (Z[54], A[54], n_177);
  and g168 (n_178, A[54], n_177);
  xor g169 (Z[55], A[55], n_178);
  and g170 (n_179, A[55], n_178);
  xor g171 (Z[56], A[56], n_179);
  and g172 (n_180, A[56], n_179);
  xor g173 (Z[57], A[57], n_180);
  and g174 (n_181, A[57], n_180);
  xor g175 (Z[58], A[58], n_181);
  and g176 (n_182, A[58], n_181);
  xor g177 (Z[59], A[59], n_182);
  and g178 (n_183, A[59], n_182);
  xor g179 (Z[60], A[60], n_183);
endmodule

module increment_unsigned_16827_GENERIC(A, CI, Z);
  input [60:0] A;
  input CI;
  output [60:0] Z;
  wire [60:0] A;
  wire CI;
  wire [60:0] Z;
  increment_unsigned_16827_GENERIC_REAL g1(.A ({A[59], A[59:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16828_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [66:0] A;
  input CI;
  output [66:0] Z;
  wire [66:0] A;
  wire CI;
  wire [66:0] Z;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_136, A[0], CI);
  xor g67 (Z[1], A[1], n_136);
  and g68 (n_137, A[1], n_136);
  xor g69 (Z[2], A[2], n_137);
  and g70 (n_138, A[2], n_137);
  xor g71 (Z[3], A[3], n_138);
  and g72 (n_139, A[3], n_138);
  xor g73 (Z[4], A[4], n_139);
  and g74 (n_140, A[4], n_139);
  xor g75 (Z[5], A[5], n_140);
  and g76 (n_141, A[5], n_140);
  xor g77 (Z[6], A[6], n_141);
  and g78 (n_142, A[6], n_141);
  xor g79 (Z[7], A[7], n_142);
  and g80 (n_143, A[7], n_142);
  xor g81 (Z[8], A[8], n_143);
  and g82 (n_144, A[8], n_143);
  xor g83 (Z[9], A[9], n_144);
  and g84 (n_145, A[9], n_144);
  xor g85 (Z[10], A[10], n_145);
  and g86 (n_146, A[10], n_145);
  xor g87 (Z[11], A[11], n_146);
  and g88 (n_147, A[11], n_146);
  xor g89 (Z[12], A[12], n_147);
  and g90 (n_148, A[12], n_147);
  xor g91 (Z[13], A[13], n_148);
  and g92 (n_149, A[13], n_148);
  xor g93 (Z[14], A[14], n_149);
  and g94 (n_150, A[14], n_149);
  xor g95 (Z[15], A[15], n_150);
  and g96 (n_151, A[15], n_150);
  xor g97 (Z[16], A[16], n_151);
  and g98 (n_152, A[16], n_151);
  xor g99 (Z[17], A[17], n_152);
  and g100 (n_153, A[17], n_152);
  xor g101 (Z[18], A[18], n_153);
  and g102 (n_154, A[18], n_153);
  xor g103 (Z[19], A[19], n_154);
  and g104 (n_155, A[19], n_154);
  xor g105 (Z[20], A[20], n_155);
  and g106 (n_156, A[20], n_155);
  xor g107 (Z[21], A[21], n_156);
  and g108 (n_157, A[21], n_156);
  xor g109 (Z[22], A[22], n_157);
  and g110 (n_158, A[22], n_157);
  xor g111 (Z[23], A[23], n_158);
  and g112 (n_159, A[23], n_158);
  xor g113 (Z[24], A[24], n_159);
  and g114 (n_160, A[24], n_159);
  xor g115 (Z[25], A[25], n_160);
  and g116 (n_161, A[25], n_160);
  xor g117 (Z[26], A[26], n_161);
  and g118 (n_162, A[26], n_161);
  xor g119 (Z[27], A[27], n_162);
  and g120 (n_163, A[27], n_162);
  xor g121 (Z[28], A[28], n_163);
  and g122 (n_164, A[28], n_163);
  xor g123 (Z[29], A[29], n_164);
  and g124 (n_165, A[29], n_164);
  xor g125 (Z[30], A[30], n_165);
  and g126 (n_166, A[30], n_165);
  xor g127 (Z[31], A[31], n_166);
  and g128 (n_167, A[31], n_166);
  xor g129 (Z[32], A[32], n_167);
  and g130 (n_168, A[32], n_167);
  xor g131 (Z[33], A[33], n_168);
  and g132 (n_169, A[33], n_168);
  xor g133 (Z[34], A[34], n_169);
  and g134 (n_170, A[34], n_169);
  xor g135 (Z[35], A[35], n_170);
  and g136 (n_171, A[35], n_170);
  xor g137 (Z[36], A[36], n_171);
  and g138 (n_172, A[36], n_171);
  xor g139 (Z[37], A[37], n_172);
  and g140 (n_173, A[37], n_172);
  xor g141 (Z[38], A[38], n_173);
  and g142 (n_174, A[38], n_173);
  xor g143 (Z[39], A[39], n_174);
  and g144 (n_175, A[39], n_174);
  xor g145 (Z[40], A[40], n_175);
  and g146 (n_176, A[40], n_175);
  xor g147 (Z[41], A[41], n_176);
  and g148 (n_177, A[41], n_176);
  xor g149 (Z[42], A[42], n_177);
  and g150 (n_178, A[42], n_177);
  xor g151 (Z[43], A[43], n_178);
  and g152 (n_179, A[43], n_178);
  xor g153 (Z[44], A[44], n_179);
  and g154 (n_180, A[44], n_179);
  xor g155 (Z[45], A[45], n_180);
  and g156 (n_181, A[45], n_180);
  xor g157 (Z[46], A[46], n_181);
  and g158 (n_182, A[46], n_181);
  xor g159 (Z[47], A[47], n_182);
  and g160 (n_183, A[47], n_182);
  xor g161 (Z[48], A[48], n_183);
  and g162 (n_184, A[48], n_183);
  xor g163 (Z[49], A[49], n_184);
  and g164 (n_185, A[49], n_184);
  xor g165 (Z[50], A[50], n_185);
  and g166 (n_186, A[50], n_185);
  xor g167 (Z[51], A[51], n_186);
  and g168 (n_187, A[51], n_186);
  xor g169 (Z[52], A[52], n_187);
  and g170 (n_188, A[52], n_187);
  xor g171 (Z[53], A[53], n_188);
  and g172 (n_189, A[53], n_188);
  xor g173 (Z[54], A[54], n_189);
  and g174 (n_190, A[54], n_189);
  xor g175 (Z[55], A[55], n_190);
  and g176 (n_191, A[55], n_190);
  xor g177 (Z[56], A[56], n_191);
  and g178 (n_192, A[56], n_191);
  xor g179 (Z[57], A[57], n_192);
  and g180 (n_193, A[57], n_192);
  xor g181 (Z[58], A[58], n_193);
  and g182 (n_194, A[58], n_193);
  xor g183 (Z[59], A[59], n_194);
  and g184 (n_195, A[59], n_194);
  xor g185 (Z[60], A[60], n_195);
  and g186 (n_196, A[60], n_195);
  xor g187 (Z[61], A[61], n_196);
  and g188 (n_197, A[61], n_196);
  xor g189 (Z[62], A[62], n_197);
  and g190 (n_198, A[62], n_197);
  xor g191 (Z[63], A[63], n_198);
  and g192 (n_199, A[63], n_198);
  xor g193 (Z[64], A[64], n_199);
  and g194 (n_200, A[64], n_199);
  xor g195 (Z[65], A[65], n_200);
  and g196 (n_201, A[65], n_200);
  xor g197 (Z[66], A[66], n_201);
endmodule

module increment_unsigned_16828_GENERIC(A, CI, Z);
  input [66:0] A;
  input CI;
  output [66:0] Z;
  wire [66:0] A;
  wire CI;
  wire [66:0] Z;
  increment_unsigned_16828_GENERIC_REAL g1(.A ({A[65], A[65:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16830_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [58:0] A;
  input CI;
  output [58:0] Z;
  wire [58:0] A;
  wire CI;
  wire [58:0] Z;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_120, A[0], CI);
  xor g59 (Z[1], A[1], n_120);
  and g60 (n_121, A[1], n_120);
  xor g61 (Z[2], A[2], n_121);
  and g62 (n_122, A[2], n_121);
  xor g63 (Z[3], A[3], n_122);
  and g64 (n_123, A[3], n_122);
  xor g65 (Z[4], A[4], n_123);
  and g66 (n_124, A[4], n_123);
  xor g67 (Z[5], A[5], n_124);
  and g68 (n_125, A[5], n_124);
  xor g69 (Z[6], A[6], n_125);
  and g70 (n_126, A[6], n_125);
  xor g71 (Z[7], A[7], n_126);
  and g72 (n_127, A[7], n_126);
  xor g73 (Z[8], A[8], n_127);
  and g74 (n_128, A[8], n_127);
  xor g75 (Z[9], A[9], n_128);
  and g76 (n_129, A[9], n_128);
  xor g77 (Z[10], A[10], n_129);
  and g78 (n_130, A[10], n_129);
  xor g79 (Z[11], A[11], n_130);
  and g80 (n_131, A[11], n_130);
  xor g81 (Z[12], A[12], n_131);
  and g82 (n_132, A[12], n_131);
  xor g83 (Z[13], A[13], n_132);
  and g84 (n_133, A[13], n_132);
  xor g85 (Z[14], A[14], n_133);
  and g86 (n_134, A[14], n_133);
  xor g87 (Z[15], A[15], n_134);
  and g88 (n_135, A[15], n_134);
  xor g89 (Z[16], A[16], n_135);
  and g90 (n_136, A[16], n_135);
  xor g91 (Z[17], A[17], n_136);
  and g92 (n_137, A[17], n_136);
  xor g93 (Z[18], A[18], n_137);
  and g94 (n_138, A[18], n_137);
  xor g95 (Z[19], A[19], n_138);
  and g96 (n_139, A[19], n_138);
  xor g97 (Z[20], A[20], n_139);
  and g98 (n_140, A[20], n_139);
  xor g99 (Z[21], A[21], n_140);
  and g100 (n_141, A[21], n_140);
  xor g101 (Z[22], A[22], n_141);
  and g102 (n_142, A[22], n_141);
  xor g103 (Z[23], A[23], n_142);
  and g104 (n_143, A[23], n_142);
  xor g105 (Z[24], A[24], n_143);
  and g106 (n_144, A[24], n_143);
  xor g107 (Z[25], A[25], n_144);
  and g108 (n_145, A[25], n_144);
  xor g109 (Z[26], A[26], n_145);
  and g110 (n_146, A[26], n_145);
  xor g111 (Z[27], A[27], n_146);
  and g112 (n_147, A[27], n_146);
  xor g113 (Z[28], A[28], n_147);
  and g114 (n_148, A[28], n_147);
  xor g115 (Z[29], A[29], n_148);
  and g116 (n_149, A[29], n_148);
  xor g117 (Z[30], A[30], n_149);
  and g118 (n_150, A[30], n_149);
  xor g119 (Z[31], A[31], n_150);
  and g120 (n_151, A[31], n_150);
  xor g121 (Z[32], A[32], n_151);
  and g122 (n_152, A[32], n_151);
  xor g123 (Z[33], A[33], n_152);
  and g124 (n_153, A[33], n_152);
  xor g125 (Z[34], A[34], n_153);
  and g126 (n_154, A[34], n_153);
  xor g127 (Z[35], A[35], n_154);
  and g128 (n_155, A[35], n_154);
  xor g129 (Z[36], A[36], n_155);
  and g130 (n_156, A[36], n_155);
  xor g131 (Z[37], A[37], n_156);
  and g132 (n_157, A[37], n_156);
  xor g133 (Z[38], A[38], n_157);
  and g134 (n_158, A[38], n_157);
  xor g135 (Z[39], A[39], n_158);
  and g136 (n_159, A[39], n_158);
  xor g137 (Z[40], A[40], n_159);
  and g138 (n_160, A[40], n_159);
  xor g139 (Z[41], A[41], n_160);
  and g140 (n_161, A[41], n_160);
  xor g141 (Z[42], A[42], n_161);
  and g142 (n_162, A[42], n_161);
  xor g143 (Z[43], A[43], n_162);
  and g144 (n_163, A[43], n_162);
  xor g145 (Z[44], A[44], n_163);
  and g146 (n_164, A[44], n_163);
  xor g147 (Z[45], A[45], n_164);
  and g148 (n_165, A[45], n_164);
  xor g149 (Z[46], A[46], n_165);
  and g150 (n_166, A[46], n_165);
  xor g151 (Z[47], A[47], n_166);
  and g152 (n_167, A[47], n_166);
  xor g153 (Z[48], A[48], n_167);
  and g154 (n_168, A[48], n_167);
  xor g155 (Z[49], A[49], n_168);
  and g156 (n_169, A[49], n_168);
  xor g157 (Z[50], A[50], n_169);
  and g158 (n_170, A[50], n_169);
  xor g159 (Z[51], A[51], n_170);
  and g160 (n_171, A[51], n_170);
  xor g161 (Z[52], A[52], n_171);
  and g162 (n_172, A[52], n_171);
  xor g163 (Z[53], A[53], n_172);
  and g164 (n_173, A[53], n_172);
  xor g165 (Z[54], A[54], n_173);
  and g166 (n_174, A[54], n_173);
  xor g167 (Z[55], A[55], n_174);
  and g168 (n_175, A[55], n_174);
  xor g169 (Z[56], A[56], n_175);
  and g170 (n_176, A[56], n_175);
  xor g171 (Z[57], A[57], n_176);
  and g172 (n_177, A[57], n_176);
  xor g173 (Z[58], A[58], n_177);
endmodule

module increment_unsigned_16830_GENERIC(A, CI, Z);
  input [58:0] A;
  input CI;
  output [58:0] Z;
  wire [58:0] A;
  wire CI;
  wire [58:0] Z;
  increment_unsigned_16830_GENERIC_REAL g1(.A ({A[57], A[57:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16830_1_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [58:0] A;
  input CI;
  output [58:0] Z;
  wire [58:0] A;
  wire CI;
  wire [58:0] Z;
  wire n_120, n_122, n_123, n_125, n_127, n_128, n_130, n_131;
  wire n_133, n_134, n_136, n_137, n_139, n_140, n_142, n_143;
  wire n_145, n_146, n_148, n_149, n_151, n_152, n_154, n_155;
  wire n_157, n_158, n_160, n_161, n_163, n_164, n_166, n_168;
  wire n_170, n_172, n_174, n_175, n_176, n_178, n_179, n_180;
  wire n_182, n_183, n_184, n_186, n_187, n_188, n_190, n_191;
  wire n_192, n_194, n_195, n_196, n_198, n_199, n_201, n_203;
  wire n_205, n_207, n_209, n_212, n_213, n_214, n_215, n_216;
  wire n_218, n_221, n_222, n_223, n_224, n_225, n_229, n_231;
  wire n_234, n_235, n_236, n_237, n_239, n_241, n_243, n_245;
  wire n_247, n_249, n_251, n_253, n_255, n_256, n_258, n_260;
  wire n_263, n_264, n_266, n_268, n_269, n_271, n_273, n_276;
  wire n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_285;
  wire n_287, n_289, n_291, n_293, n_295, n_297, n_299, n_301;
  wire n_306, n_309, n_310, n_311, n_312, n_314, n_316, n_318;
  wire n_320, n_322, n_324, n_327, n_328, n_329, n_330, n_331;
  wire n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339;
  wire n_340, n_341, n_342, n_344, n_346, n_348, n_350, n_352;
  wire n_354, n_356, n_358, n_360, n_362, n_364, n_366, n_368;
  wire n_370, n_372, n_374, n_376, n_378, n_380, n_382, n_384;
  wire n_386, n_388, n_390, n_392;
  nand g1 (n_120, A[0], CI);
  nand g4 (n_123, A[2], A[3]);
  nand g5 (n_125, A[4], A[5]);
  nand g6 (n_127, A[6], A[7]);
  nand g7 (n_128, A[8], A[9]);
  nand g8 (n_130, A[10], A[11]);
  nand g9 (n_131, A[12], A[13]);
  nand g10 (n_133, A[14], A[15]);
  nand g11 (n_134, A[16], A[17]);
  nand g12 (n_136, A[18], A[19]);
  nand g13 (n_137, A[20], A[21]);
  nand g14 (n_139, A[22], A[23]);
  nand g15 (n_140, A[24], A[25]);
  nand g16 (n_142, A[26], A[27]);
  nand g17 (n_143, A[28], A[29]);
  nand g18 (n_145, A[30], A[31]);
  nand g19 (n_146, A[32], A[33]);
  nand g20 (n_148, A[34], A[35]);
  nand g21 (n_149, A[36], A[37]);
  nand g22 (n_151, A[38], A[39]);
  nand g23 (n_152, A[40], A[41]);
  nand g24 (n_154, A[42], A[43]);
  nand g25 (n_155, A[44], A[45]);
  nand g26 (n_157, A[46], A[47]);
  nand g27 (n_158, A[48], A[49]);
  nand g28 (n_160, A[50], A[51]);
  nand g29 (n_161, A[52], A[53]);
  nand g30 (n_163, A[54], A[55]);
  nand g31 (n_164, A[56], A[57]);
  nand g32 (n_306, A[2], n_122);
  nor g37 (n_170, n_125, n_127);
  nor g40 (n_172, n_128, n_130);
  nor g43 (n_175, n_131, n_133);
  nor g46 (n_176, n_134, n_136);
  nor g49 (n_179, n_137, n_139);
  nor g52 (n_180, n_140, n_142);
  nor g55 (n_183, n_143, n_145);
  nor g58 (n_184, n_146, n_148);
  nor g61 (n_187, n_149, n_151);
  nor g64 (n_188, n_152, n_154);
  nor g67 (n_191, n_155, n_157);
  nor g70 (n_192, n_158, n_160);
  nor g73 (n_195, n_161, n_163);
  nor g78 (n_310, n_125, n_166);
  nand g83 (n_199, A[12], n_172);
  nand g86 (n_203, n_172, n_174);
  nand g87 (n_205, n_172, n_175);
  nand g88 (n_234, A[20], n_176);
  nand g91 (n_236, n_176, n_178);
  nand g92 (n_207, n_176, n_179);
  nand g93 (n_212, A[28], n_180);
  nand g96 (n_214, n_180, n_182);
  nand g97 (n_215, n_180, n_183);
  nand g98 (n_269, A[36], n_184);
  nand g101 (n_273, n_184, n_186);
  nand g102 (n_216, n_184, n_187);
  nand g103 (n_221, A[44], n_188);
  nand g106 (n_223, n_188, n_190);
  nand g107 (n_224, n_188, n_191);
  nand g108 (n_256, A[52], n_192);
  nand g111 (n_260, n_192, n_194);
  nand g112 (n_225, n_192, n_195);
  nand g113 (n_312, A[8], n_196);
  nand g116 (n_316, n_198, n_196);
  nand g117 (n_318, n_172, n_196);
  nor g128 (n_239, n_140, n_207);
  nor g133 (n_245, n_207, n_212);
  nor g134 (n_247, n_207, n_213);
  nor g135 (n_249, n_207, n_214);
  nor g136 (n_251, n_207, n_215);
  nor g139 (n_277, n_152, n_216);
  nor g144 (n_280, n_216, n_221);
  nor g145 (n_281, n_216, n_222);
  nor g146 (n_282, n_216, n_223);
  nor g147 (n_253, n_216, n_224);
  nor g150 (n_264, n_164, n_225);
  nor g155 (n_328, n_134, n_229);
  nor g160 (n_331, n_234, n_229);
  nor g161 (n_332, n_235, n_229);
  nor g162 (n_333, n_236, n_229);
  nor g163 (n_334, n_207, n_229);
  nand g180 (n_283, A[48], n_253);
  nand g183 (n_287, n_255, n_253);
  nand g184 (n_289, n_192, n_253);
  nand g193 (n_299, n_253, n_263);
  nand g194 (n_301, n_253, n_264);
  nand g196 (n_342, A[32], n_266);
  nand g199 (n_346, n_268, n_266);
  nand g200 (n_348, n_184, n_266);
  nand g209 (n_358, n_276, n_266);
  nand g210 (n_360, n_277, n_266);
  nand g211 (n_362, n_278, n_266);
  nand g212 (n_364, n_279, n_266);
  nand g213 (n_366, n_280, n_266);
  nand g214 (n_368, n_281, n_266);
  nand g215 (n_370, n_282, n_266);
  nand g216 (n_372, n_253, n_266);
  xor g239 (Z[0], A[0], CI);
  xor g242 (Z[2], A[2], n_122);
  xor g247 (Z[5], A[5], n_309);
  xor g248 (Z[6], A[6], n_310);
  xor g249 (Z[7], A[7], n_311);
  xor g250 (Z[8], A[8], n_196);
  xor g267 (Z[17], A[17], n_327);
  xor g268 (Z[18], A[18], n_328);
  xor g269 (Z[19], A[19], n_329);
  xor g270 (Z[20], A[20], n_330);
  xor g271 (Z[21], A[21], n_331);
  xor g272 (Z[22], A[22], n_332);
  xor g273 (Z[23], A[23], n_333);
  xor g274 (Z[24], A[24], n_334);
  xor g275 (Z[25], A[25], n_335);
  xor g276 (Z[26], A[26], n_336);
  xor g277 (Z[27], A[27], n_337);
  xor g278 (Z[28], A[28], n_338);
  xor g279 (Z[29], A[29], n_339);
  xor g280 (Z[30], A[30], n_340);
  xor g281 (Z[31], A[31], n_341);
  xor g282 (Z[32], A[32], n_266);
  and g336 (n_122, A[1], wc);
  not gc (wc, n_120);
  and g337 (n_168, A[6], wc0);
  not gc0 (wc0, n_125);
  and g338 (n_198, A[10], wc1);
  not gc1 (wc1, n_128);
  and g339 (n_174, A[14], wc2);
  not gc2 (wc2, n_131);
  and g340 (n_231, A[18], wc3);
  not gc3 (wc3, n_134);
  and g341 (n_178, A[22], wc4);
  not gc4 (wc4, n_137);
  and g342 (n_209, A[26], wc5);
  not gc5 (wc5, n_140);
  and g343 (n_182, A[30], wc6);
  not gc6 (wc6, n_143);
  and g344 (n_268, A[34], wc7);
  not gc7 (wc7, n_146);
  and g345 (n_186, A[38], wc8);
  not gc8 (wc8, n_149);
  and g346 (n_218, A[42], wc9);
  not gc9 (wc9, n_152);
  and g347 (n_190, A[46], wc10);
  not gc10 (wc10, n_155);
  and g348 (n_255, A[50], wc11);
  not gc11 (wc11, n_158);
  and g349 (n_194, A[54], wc12);
  not gc12 (wc12, n_161);
  or g350 (n_166, wc13, n_123);
  not gc13 (wc13, n_122);
  or g351 (n_201, wc14, n_131);
  not gc14 (wc14, n_172);
  or g352 (n_235, wc15, n_137);
  not gc15 (wc15, n_176);
  or g353 (n_213, wc16, n_143);
  not gc16 (wc16, n_180);
  or g354 (n_271, wc17, n_149);
  not gc17 (wc17, n_184);
  or g355 (n_222, wc18, n_155);
  not gc18 (wc18, n_188);
  or g356 (n_258, wc19, n_161);
  not gc19 (wc19, n_192);
  xnor g357 (Z[1], n_120, A[1]);
  and g358 (n_309, A[4], wc20);
  not gc20 (wc20, n_166);
  and g359 (n_311, wc21, n_168);
  not gc21 (wc21, n_166);
  and g360 (n_196, wc22, n_170);
  not gc22 (wc22, n_166);
  and g361 (n_237, A[24], wc23);
  not gc23 (wc23, n_207);
  and g362 (n_241, n_209, wc24);
  not gc24 (wc24, n_207);
  and g363 (n_243, wc25, n_180);
  not gc25 (wc25, n_207);
  and g364 (n_276, A[40], wc26);
  not gc26 (wc26, n_216);
  and g365 (n_278, n_218, wc27);
  not gc27 (wc27, n_216);
  and g366 (n_279, wc28, n_188);
  not gc28 (wc28, n_216);
  and g367 (n_263, A[56], wc29);
  not gc29 (wc29, n_225);
  or g368 (n_314, wc30, n_128);
  not gc30 (wc30, n_196);
  or g369 (n_320, wc31, n_199);
  not gc31 (wc31, n_196);
  or g370 (n_322, wc32, n_201);
  not gc32 (wc32, n_196);
  or g371 (n_324, wc33, n_203);
  not gc33 (wc33, n_196);
  or g372 (n_229, wc34, n_205);
  not gc34 (wc34, n_196);
  or g373 (n_285, wc35, n_158);
  not gc35 (wc35, n_253);
  or g374 (n_291, wc36, n_256);
  not gc36 (wc36, n_253);
  or g375 (n_293, n_258, wc37);
  not gc37 (wc37, n_253);
  or g376 (n_295, wc38, n_260);
  not gc38 (wc38, n_253);
  or g377 (n_297, wc39, n_225);
  not gc39 (wc39, n_253);
  xnor g378 (Z[3], n_306, A[3]);
  xnor g379 (Z[4], n_166, A[4]);
  and g380 (n_327, A[16], wc40);
  not gc40 (wc40, n_229);
  and g381 (n_329, wc41, n_231);
  not gc41 (wc41, n_229);
  and g382 (n_330, wc42, n_176);
  not gc42 (wc42, n_229);
  and g383 (n_335, wc43, n_237);
  not gc43 (wc43, n_229);
  and g384 (n_336, wc44, n_239);
  not gc44 (wc44, n_229);
  and g385 (n_337, wc45, n_241);
  not gc45 (wc45, n_229);
  and g386 (n_338, wc46, n_243);
  not gc46 (wc46, n_229);
  and g387 (n_339, wc47, n_245);
  not gc47 (wc47, n_229);
  and g388 (n_340, wc48, n_247);
  not gc48 (wc48, n_229);
  and g389 (n_341, wc49, n_249);
  not gc49 (wc49, n_229);
  and g390 (n_266, wc50, n_251);
  not gc50 (wc50, n_229);
  or g391 (n_344, wc51, n_146);
  not gc51 (wc51, n_266);
  or g392 (n_350, wc52, n_269);
  not gc52 (wc52, n_266);
  or g393 (n_352, wc53, n_271);
  not gc53 (wc53, n_266);
  or g394 (n_354, wc54, n_273);
  not gc54 (wc54, n_266);
  or g395 (n_356, wc55, n_216);
  not gc55 (wc55, n_266);
  or g396 (n_374, wc56, n_283);
  not gc56 (wc56, n_266);
  or g397 (n_376, wc57, n_285);
  not gc57 (wc57, n_266);
  or g398 (n_378, wc58, n_287);
  not gc58 (wc58, n_266);
  or g399 (n_380, wc59, n_289);
  not gc59 (wc59, n_266);
  or g400 (n_382, wc60, n_291);
  not gc60 (wc60, n_266);
  or g401 (n_384, wc61, n_293);
  not gc61 (wc61, n_266);
  or g402 (n_386, wc62, n_295);
  not gc62 (wc62, n_266);
  or g403 (n_388, wc63, n_297);
  not gc63 (wc63, n_266);
  or g404 (n_390, wc64, n_299);
  not gc64 (wc64, n_266);
  or g405 (n_392, wc65, n_301);
  not gc65 (wc65, n_266);
  xnor g406 (Z[9], n_312, A[9]);
  xnor g407 (Z[10], n_314, A[10]);
  xnor g408 (Z[11], n_316, A[11]);
  xnor g409 (Z[12], n_318, A[12]);
  xnor g410 (Z[13], n_320, A[13]);
  xnor g411 (Z[14], n_322, A[14]);
  xnor g412 (Z[15], n_324, A[15]);
  xnor g413 (Z[16], n_229, A[16]);
  xnor g414 (Z[33], n_342, A[33]);
  xnor g415 (Z[34], n_344, A[34]);
  xnor g416 (Z[35], n_346, A[35]);
  xnor g417 (Z[36], n_348, A[36]);
  xnor g418 (Z[37], n_350, A[37]);
  xnor g419 (Z[38], n_352, A[38]);
  xnor g420 (Z[39], n_354, A[39]);
  xnor g421 (Z[40], n_356, A[40]);
  xnor g422 (Z[41], n_358, A[41]);
  xnor g423 (Z[42], n_360, A[42]);
  xnor g424 (Z[43], n_362, A[43]);
  xnor g425 (Z[44], n_364, A[44]);
  xnor g426 (Z[45], n_366, A[45]);
  xnor g427 (Z[46], n_368, A[46]);
  xnor g428 (Z[47], n_370, A[47]);
  xnor g429 (Z[48], n_372, A[48]);
  xnor g430 (Z[49], n_374, A[49]);
  xnor g431 (Z[50], n_376, A[50]);
  xnor g432 (Z[51], n_378, A[51]);
  xnor g433 (Z[52], n_380, A[52]);
  xnor g434 (Z[53], n_382, A[53]);
  xnor g435 (Z[54], n_384, A[54]);
  xnor g436 (Z[55], n_386, A[55]);
  xnor g437 (Z[56], n_388, A[56]);
  xnor g438 (Z[57], n_390, A[57]);
  xnor g439 (Z[58], n_392, A[58]);
endmodule

module increment_unsigned_16830_1_GENERIC(A, CI, Z);
  input [58:0] A;
  input CI;
  output [58:0] Z;
  wire [58:0] A;
  wire CI;
  wire [58:0] Z;
  increment_unsigned_16830_1_GENERIC_REAL g1(.A ({A[57], A[57:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16832_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [56:0] A;
  input CI;
  output [56:0] Z;
  wire [56:0] A;
  wire CI;
  wire [56:0] Z;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163;
  wire n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_116, A[0], CI);
  xor g57 (Z[1], A[1], n_116);
  and g58 (n_117, A[1], n_116);
  xor g59 (Z[2], A[2], n_117);
  and g60 (n_118, A[2], n_117);
  xor g61 (Z[3], A[3], n_118);
  and g62 (n_119, A[3], n_118);
  xor g63 (Z[4], A[4], n_119);
  and g64 (n_120, A[4], n_119);
  xor g65 (Z[5], A[5], n_120);
  and g66 (n_121, A[5], n_120);
  xor g67 (Z[6], A[6], n_121);
  and g68 (n_122, A[6], n_121);
  xor g69 (Z[7], A[7], n_122);
  and g70 (n_123, A[7], n_122);
  xor g71 (Z[8], A[8], n_123);
  and g72 (n_124, A[8], n_123);
  xor g73 (Z[9], A[9], n_124);
  and g74 (n_125, A[9], n_124);
  xor g75 (Z[10], A[10], n_125);
  and g76 (n_126, A[10], n_125);
  xor g77 (Z[11], A[11], n_126);
  and g78 (n_127, A[11], n_126);
  xor g79 (Z[12], A[12], n_127);
  and g80 (n_128, A[12], n_127);
  xor g81 (Z[13], A[13], n_128);
  and g82 (n_129, A[13], n_128);
  xor g83 (Z[14], A[14], n_129);
  and g84 (n_130, A[14], n_129);
  xor g85 (Z[15], A[15], n_130);
  and g86 (n_131, A[15], n_130);
  xor g87 (Z[16], A[16], n_131);
  and g88 (n_132, A[16], n_131);
  xor g89 (Z[17], A[17], n_132);
  and g90 (n_133, A[17], n_132);
  xor g91 (Z[18], A[18], n_133);
  and g92 (n_134, A[18], n_133);
  xor g93 (Z[19], A[19], n_134);
  and g94 (n_135, A[19], n_134);
  xor g95 (Z[20], A[20], n_135);
  and g96 (n_136, A[20], n_135);
  xor g97 (Z[21], A[21], n_136);
  and g98 (n_137, A[21], n_136);
  xor g99 (Z[22], A[22], n_137);
  and g100 (n_138, A[22], n_137);
  xor g101 (Z[23], A[23], n_138);
  and g102 (n_139, A[23], n_138);
  xor g103 (Z[24], A[24], n_139);
  and g104 (n_140, A[24], n_139);
  xor g105 (Z[25], A[25], n_140);
  and g106 (n_141, A[25], n_140);
  xor g107 (Z[26], A[26], n_141);
  and g108 (n_142, A[26], n_141);
  xor g109 (Z[27], A[27], n_142);
  and g110 (n_143, A[27], n_142);
  xor g111 (Z[28], A[28], n_143);
  and g112 (n_144, A[28], n_143);
  xor g113 (Z[29], A[29], n_144);
  and g114 (n_145, A[29], n_144);
  xor g115 (Z[30], A[30], n_145);
  and g116 (n_146, A[30], n_145);
  xor g117 (Z[31], A[31], n_146);
  and g118 (n_147, A[31], n_146);
  xor g119 (Z[32], A[32], n_147);
  and g120 (n_148, A[32], n_147);
  xor g121 (Z[33], A[33], n_148);
  and g122 (n_149, A[33], n_148);
  xor g123 (Z[34], A[34], n_149);
  and g124 (n_150, A[34], n_149);
  xor g125 (Z[35], A[35], n_150);
  and g126 (n_151, A[35], n_150);
  xor g127 (Z[36], A[36], n_151);
  and g128 (n_152, A[36], n_151);
  xor g129 (Z[37], A[37], n_152);
  and g130 (n_153, A[37], n_152);
  xor g131 (Z[38], A[38], n_153);
  and g132 (n_154, A[38], n_153);
  xor g133 (Z[39], A[39], n_154);
  and g134 (n_155, A[39], n_154);
  xor g135 (Z[40], A[40], n_155);
  and g136 (n_156, A[40], n_155);
  xor g137 (Z[41], A[41], n_156);
  and g138 (n_157, A[41], n_156);
  xor g139 (Z[42], A[42], n_157);
  and g140 (n_158, A[42], n_157);
  xor g141 (Z[43], A[43], n_158);
  and g142 (n_159, A[43], n_158);
  xor g143 (Z[44], A[44], n_159);
  and g144 (n_160, A[44], n_159);
  xor g145 (Z[45], A[45], n_160);
  and g146 (n_161, A[45], n_160);
  xor g147 (Z[46], A[46], n_161);
  and g148 (n_162, A[46], n_161);
  xor g149 (Z[47], A[47], n_162);
  and g150 (n_163, A[47], n_162);
  xor g151 (Z[48], A[48], n_163);
  and g152 (n_164, A[48], n_163);
  xor g153 (Z[49], A[49], n_164);
  and g154 (n_165, A[49], n_164);
  xor g155 (Z[50], A[50], n_165);
  and g156 (n_166, A[50], n_165);
  xor g157 (Z[51], A[51], n_166);
  and g158 (n_167, A[51], n_166);
  xor g159 (Z[52], A[52], n_167);
  and g160 (n_168, A[52], n_167);
  xor g161 (Z[53], A[53], n_168);
  and g162 (n_169, A[53], n_168);
  xor g163 (Z[54], A[54], n_169);
  and g164 (n_170, A[54], n_169);
  xor g165 (Z[55], A[55], n_170);
  and g166 (n_171, A[55], n_170);
  xor g167 (Z[56], A[56], n_171);
endmodule

module increment_unsigned_16832_GENERIC(A, CI, Z);
  input [56:0] A;
  input CI;
  output [56:0] Z;
  wire [56:0] A;
  wire CI;
  wire [56:0] Z;
  increment_unsigned_16832_GENERIC_REAL g1(.A ({A[55], A[55:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16833_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [61:0] A;
  input CI;
  output [61:0] Z;
  wire [61:0] A;
  wire CI;
  wire [61:0] Z;
  wire n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133;
  wire n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_126, A[0], CI);
  xor g62 (Z[1], A[1], n_126);
  and g63 (n_127, A[1], n_126);
  xor g64 (Z[2], A[2], n_127);
  and g65 (n_128, A[2], n_127);
  xor g66 (Z[3], A[3], n_128);
  and g67 (n_129, A[3], n_128);
  xor g68 (Z[4], A[4], n_129);
  and g69 (n_130, A[4], n_129);
  xor g70 (Z[5], A[5], n_130);
  and g71 (n_131, A[5], n_130);
  xor g72 (Z[6], A[6], n_131);
  and g73 (n_132, A[6], n_131);
  xor g74 (Z[7], A[7], n_132);
  and g75 (n_133, A[7], n_132);
  xor g76 (Z[8], A[8], n_133);
  and g77 (n_134, A[8], n_133);
  xor g78 (Z[9], A[9], n_134);
  and g79 (n_135, A[9], n_134);
  xor g80 (Z[10], A[10], n_135);
  and g81 (n_136, A[10], n_135);
  xor g82 (Z[11], A[11], n_136);
  and g83 (n_137, A[11], n_136);
  xor g84 (Z[12], A[12], n_137);
  and g85 (n_138, A[12], n_137);
  xor g86 (Z[13], A[13], n_138);
  and g87 (n_139, A[13], n_138);
  xor g88 (Z[14], A[14], n_139);
  and g89 (n_140, A[14], n_139);
  xor g90 (Z[15], A[15], n_140);
  and g91 (n_141, A[15], n_140);
  xor g92 (Z[16], A[16], n_141);
  and g93 (n_142, A[16], n_141);
  xor g94 (Z[17], A[17], n_142);
  and g95 (n_143, A[17], n_142);
  xor g96 (Z[18], A[18], n_143);
  and g97 (n_144, A[18], n_143);
  xor g98 (Z[19], A[19], n_144);
  and g99 (n_145, A[19], n_144);
  xor g100 (Z[20], A[20], n_145);
  and g101 (n_146, A[20], n_145);
  xor g102 (Z[21], A[21], n_146);
  and g103 (n_147, A[21], n_146);
  xor g104 (Z[22], A[22], n_147);
  and g105 (n_148, A[22], n_147);
  xor g106 (Z[23], A[23], n_148);
  and g107 (n_149, A[23], n_148);
  xor g108 (Z[24], A[24], n_149);
  and g109 (n_150, A[24], n_149);
  xor g110 (Z[25], A[25], n_150);
  and g111 (n_151, A[25], n_150);
  xor g112 (Z[26], A[26], n_151);
  and g113 (n_152, A[26], n_151);
  xor g114 (Z[27], A[27], n_152);
  and g115 (n_153, A[27], n_152);
  xor g116 (Z[28], A[28], n_153);
  and g117 (n_154, A[28], n_153);
  xor g118 (Z[29], A[29], n_154);
  and g119 (n_155, A[29], n_154);
  xor g120 (Z[30], A[30], n_155);
  and g121 (n_156, A[30], n_155);
  xor g122 (Z[31], A[31], n_156);
  and g123 (n_157, A[31], n_156);
  xor g124 (Z[32], A[32], n_157);
  and g125 (n_158, A[32], n_157);
  xor g126 (Z[33], A[33], n_158);
  and g127 (n_159, A[33], n_158);
  xor g128 (Z[34], A[34], n_159);
  and g129 (n_160, A[34], n_159);
  xor g130 (Z[35], A[35], n_160);
  and g131 (n_161, A[35], n_160);
  xor g132 (Z[36], A[36], n_161);
  and g133 (n_162, A[36], n_161);
  xor g134 (Z[37], A[37], n_162);
  and g135 (n_163, A[37], n_162);
  xor g136 (Z[38], A[38], n_163);
  and g137 (n_164, A[38], n_163);
  xor g138 (Z[39], A[39], n_164);
  and g139 (n_165, A[39], n_164);
  xor g140 (Z[40], A[40], n_165);
  and g141 (n_166, A[40], n_165);
  xor g142 (Z[41], A[41], n_166);
  and g143 (n_167, A[41], n_166);
  xor g144 (Z[42], A[42], n_167);
  and g145 (n_168, A[42], n_167);
  xor g146 (Z[43], A[43], n_168);
  and g147 (n_169, A[43], n_168);
  xor g148 (Z[44], A[44], n_169);
  and g149 (n_170, A[44], n_169);
  xor g150 (Z[45], A[45], n_170);
  and g151 (n_171, A[45], n_170);
  xor g152 (Z[46], A[46], n_171);
  and g153 (n_172, A[46], n_171);
  xor g154 (Z[47], A[47], n_172);
  and g155 (n_173, A[47], n_172);
  xor g156 (Z[48], A[48], n_173);
  and g157 (n_174, A[48], n_173);
  xor g158 (Z[49], A[49], n_174);
  and g159 (n_175, A[49], n_174);
  xor g160 (Z[50], A[50], n_175);
  and g161 (n_176, A[50], n_175);
  xor g162 (Z[51], A[51], n_176);
  and g163 (n_177, A[51], n_176);
  xor g164 (Z[52], A[52], n_177);
  and g165 (n_178, A[52], n_177);
  xor g166 (Z[53], A[53], n_178);
  and g167 (n_179, A[53], n_178);
  xor g168 (Z[54], A[54], n_179);
  and g169 (n_180, A[54], n_179);
  xor g170 (Z[55], A[55], n_180);
  and g171 (n_181, A[55], n_180);
  xor g172 (Z[56], A[56], n_181);
  and g173 (n_182, A[56], n_181);
  xor g174 (Z[57], A[57], n_182);
  and g175 (n_183, A[57], n_182);
  xor g176 (Z[58], A[58], n_183);
  and g177 (n_184, A[58], n_183);
  xor g178 (Z[59], A[59], n_184);
  and g179 (n_185, A[59], n_184);
  xor g180 (Z[60], A[60], n_185);
  and g181 (n_186, A[60], n_185);
  xor g182 (Z[61], A[61], n_186);
endmodule

module increment_unsigned_16833_GENERIC(A, CI, Z);
  input [61:0] A;
  input CI;
  output [61:0] Z;
  wire [61:0] A;
  wire CI;
  wire [61:0] Z;
  increment_unsigned_16833_GENERIC_REAL g1(.A ({A[60], A[60:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16834_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [53:0] A;
  input CI;
  output [53:0] Z;
  wire [53:0] A;
  wire CI;
  wire [53:0] Z;
  wire n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117;
  wire n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125;
  wire n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133;
  wire n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_159, n_160, n_161, n_162;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_110, A[0], CI);
  xor g54 (Z[1], A[1], n_110);
  and g55 (n_111, A[1], n_110);
  xor g56 (Z[2], A[2], n_111);
  and g57 (n_112, A[2], n_111);
  xor g58 (Z[3], A[3], n_112);
  and g59 (n_113, A[3], n_112);
  xor g60 (Z[4], A[4], n_113);
  and g61 (n_114, A[4], n_113);
  xor g62 (Z[5], A[5], n_114);
  and g63 (n_115, A[5], n_114);
  xor g64 (Z[6], A[6], n_115);
  and g65 (n_116, A[6], n_115);
  xor g66 (Z[7], A[7], n_116);
  and g67 (n_117, A[7], n_116);
  xor g68 (Z[8], A[8], n_117);
  and g69 (n_118, A[8], n_117);
  xor g70 (Z[9], A[9], n_118);
  and g71 (n_119, A[9], n_118);
  xor g72 (Z[10], A[10], n_119);
  and g73 (n_120, A[10], n_119);
  xor g74 (Z[11], A[11], n_120);
  and g75 (n_121, A[11], n_120);
  xor g76 (Z[12], A[12], n_121);
  and g77 (n_122, A[12], n_121);
  xor g78 (Z[13], A[13], n_122);
  and g79 (n_123, A[13], n_122);
  xor g80 (Z[14], A[14], n_123);
  and g81 (n_124, A[14], n_123);
  xor g82 (Z[15], A[15], n_124);
  and g83 (n_125, A[15], n_124);
  xor g84 (Z[16], A[16], n_125);
  and g85 (n_126, A[16], n_125);
  xor g86 (Z[17], A[17], n_126);
  and g87 (n_127, A[17], n_126);
  xor g88 (Z[18], A[18], n_127);
  and g89 (n_128, A[18], n_127);
  xor g90 (Z[19], A[19], n_128);
  and g91 (n_129, A[19], n_128);
  xor g92 (Z[20], A[20], n_129);
  and g93 (n_130, A[20], n_129);
  xor g94 (Z[21], A[21], n_130);
  and g95 (n_131, A[21], n_130);
  xor g96 (Z[22], A[22], n_131);
  and g97 (n_132, A[22], n_131);
  xor g98 (Z[23], A[23], n_132);
  and g99 (n_133, A[23], n_132);
  xor g100 (Z[24], A[24], n_133);
  and g101 (n_134, A[24], n_133);
  xor g102 (Z[25], A[25], n_134);
  and g103 (n_135, A[25], n_134);
  xor g104 (Z[26], A[26], n_135);
  and g105 (n_136, A[26], n_135);
  xor g106 (Z[27], A[27], n_136);
  and g107 (n_137, A[27], n_136);
  xor g108 (Z[28], A[28], n_137);
  and g109 (n_138, A[28], n_137);
  xor g110 (Z[29], A[29], n_138);
  and g111 (n_139, A[29], n_138);
  xor g112 (Z[30], A[30], n_139);
  and g113 (n_140, A[30], n_139);
  xor g114 (Z[31], A[31], n_140);
  and g115 (n_141, A[31], n_140);
  xor g116 (Z[32], A[32], n_141);
  and g117 (n_142, A[32], n_141);
  xor g118 (Z[33], A[33], n_142);
  and g119 (n_143, A[33], n_142);
  xor g120 (Z[34], A[34], n_143);
  and g121 (n_144, A[34], n_143);
  xor g122 (Z[35], A[35], n_144);
  and g123 (n_145, A[35], n_144);
  xor g124 (Z[36], A[36], n_145);
  and g125 (n_146, A[36], n_145);
  xor g126 (Z[37], A[37], n_146);
  and g127 (n_147, A[37], n_146);
  xor g128 (Z[38], A[38], n_147);
  and g129 (n_148, A[38], n_147);
  xor g130 (Z[39], A[39], n_148);
  and g131 (n_149, A[39], n_148);
  xor g132 (Z[40], A[40], n_149);
  and g133 (n_150, A[40], n_149);
  xor g134 (Z[41], A[41], n_150);
  and g135 (n_151, A[41], n_150);
  xor g136 (Z[42], A[42], n_151);
  and g137 (n_152, A[42], n_151);
  xor g138 (Z[43], A[43], n_152);
  and g139 (n_153, A[43], n_152);
  xor g140 (Z[44], A[44], n_153);
  and g141 (n_154, A[44], n_153);
  xor g142 (Z[45], A[45], n_154);
  and g143 (n_155, A[45], n_154);
  xor g144 (Z[46], A[46], n_155);
  and g145 (n_156, A[46], n_155);
  xor g146 (Z[47], A[47], n_156);
  and g147 (n_157, A[47], n_156);
  xor g148 (Z[48], A[48], n_157);
  and g149 (n_158, A[48], n_157);
  xor g150 (Z[49], A[49], n_158);
  and g151 (n_159, A[49], n_158);
  xor g152 (Z[50], A[50], n_159);
  and g153 (n_160, A[50], n_159);
  xor g154 (Z[51], A[51], n_160);
  and g155 (n_161, A[51], n_160);
  xor g156 (Z[52], A[52], n_161);
  and g157 (n_162, A[52], n_161);
  xor g158 (Z[53], A[53], n_162);
endmodule

module increment_unsigned_16834_GENERIC(A, CI, Z);
  input [53:0] A;
  input CI;
  output [53:0] Z;
  wire [53:0] A;
  wire CI;
  wire [53:0] Z;
  increment_unsigned_16834_GENERIC_REAL g1(.A ({A[52], A[52:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16835_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [52:0] A;
  input CI;
  output [52:0] Z;
  wire [52:0] A;
  wire CI;
  wire [52:0] Z;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_157, n_158, n_159;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_108, A[0], CI);
  xor g53 (Z[1], A[1], n_108);
  and g54 (n_109, A[1], n_108);
  xor g55 (Z[2], A[2], n_109);
  and g56 (n_110, A[2], n_109);
  xor g57 (Z[3], A[3], n_110);
  and g58 (n_111, A[3], n_110);
  xor g59 (Z[4], A[4], n_111);
  and g60 (n_112, A[4], n_111);
  xor g61 (Z[5], A[5], n_112);
  and g62 (n_113, A[5], n_112);
  xor g63 (Z[6], A[6], n_113);
  and g64 (n_114, A[6], n_113);
  xor g65 (Z[7], A[7], n_114);
  and g66 (n_115, A[7], n_114);
  xor g67 (Z[8], A[8], n_115);
  and g68 (n_116, A[8], n_115);
  xor g69 (Z[9], A[9], n_116);
  and g70 (n_117, A[9], n_116);
  xor g71 (Z[10], A[10], n_117);
  and g72 (n_118, A[10], n_117);
  xor g73 (Z[11], A[11], n_118);
  and g74 (n_119, A[11], n_118);
  xor g75 (Z[12], A[12], n_119);
  and g76 (n_120, A[12], n_119);
  xor g77 (Z[13], A[13], n_120);
  and g78 (n_121, A[13], n_120);
  xor g79 (Z[14], A[14], n_121);
  and g80 (n_122, A[14], n_121);
  xor g81 (Z[15], A[15], n_122);
  and g82 (n_123, A[15], n_122);
  xor g83 (Z[16], A[16], n_123);
  and g84 (n_124, A[16], n_123);
  xor g85 (Z[17], A[17], n_124);
  and g86 (n_125, A[17], n_124);
  xor g87 (Z[18], A[18], n_125);
  and g88 (n_126, A[18], n_125);
  xor g89 (Z[19], A[19], n_126);
  and g90 (n_127, A[19], n_126);
  xor g91 (Z[20], A[20], n_127);
  and g92 (n_128, A[20], n_127);
  xor g93 (Z[21], A[21], n_128);
  and g94 (n_129, A[21], n_128);
  xor g95 (Z[22], A[22], n_129);
  and g96 (n_130, A[22], n_129);
  xor g97 (Z[23], A[23], n_130);
  and g98 (n_131, A[23], n_130);
  xor g99 (Z[24], A[24], n_131);
  and g100 (n_132, A[24], n_131);
  xor g101 (Z[25], A[25], n_132);
  and g102 (n_133, A[25], n_132);
  xor g103 (Z[26], A[26], n_133);
  and g104 (n_134, A[26], n_133);
  xor g105 (Z[27], A[27], n_134);
  and g106 (n_135, A[27], n_134);
  xor g107 (Z[28], A[28], n_135);
  and g108 (n_136, A[28], n_135);
  xor g109 (Z[29], A[29], n_136);
  and g110 (n_137, A[29], n_136);
  xor g111 (Z[30], A[30], n_137);
  and g112 (n_138, A[30], n_137);
  xor g113 (Z[31], A[31], n_138);
  and g114 (n_139, A[31], n_138);
  xor g115 (Z[32], A[32], n_139);
  and g116 (n_140, A[32], n_139);
  xor g117 (Z[33], A[33], n_140);
  and g118 (n_141, A[33], n_140);
  xor g119 (Z[34], A[34], n_141);
  and g120 (n_142, A[34], n_141);
  xor g121 (Z[35], A[35], n_142);
  and g122 (n_143, A[35], n_142);
  xor g123 (Z[36], A[36], n_143);
  and g124 (n_144, A[36], n_143);
  xor g125 (Z[37], A[37], n_144);
  and g126 (n_145, A[37], n_144);
  xor g127 (Z[38], A[38], n_145);
  and g128 (n_146, A[38], n_145);
  xor g129 (Z[39], A[39], n_146);
  and g130 (n_147, A[39], n_146);
  xor g131 (Z[40], A[40], n_147);
  and g132 (n_148, A[40], n_147);
  xor g133 (Z[41], A[41], n_148);
  and g134 (n_149, A[41], n_148);
  xor g135 (Z[42], A[42], n_149);
  and g136 (n_150, A[42], n_149);
  xor g137 (Z[43], A[43], n_150);
  and g138 (n_151, A[43], n_150);
  xor g139 (Z[44], A[44], n_151);
  and g140 (n_152, A[44], n_151);
  xor g141 (Z[45], A[45], n_152);
  and g142 (n_153, A[45], n_152);
  xor g143 (Z[46], A[46], n_153);
  and g144 (n_154, A[46], n_153);
  xor g145 (Z[47], A[47], n_154);
  and g146 (n_155, A[47], n_154);
  xor g147 (Z[48], A[48], n_155);
  and g148 (n_156, A[48], n_155);
  xor g149 (Z[49], A[49], n_156);
  and g150 (n_157, A[49], n_156);
  xor g151 (Z[50], A[50], n_157);
  and g152 (n_158, A[50], n_157);
  xor g153 (Z[51], A[51], n_158);
  and g154 (n_159, A[51], n_158);
  xor g155 (Z[52], A[52], n_159);
endmodule

module increment_unsigned_16835_GENERIC(A, CI, Z);
  input [52:0] A;
  input CI;
  output [52:0] Z;
  wire [52:0] A;
  wire CI;
  wire [52:0] Z;
  increment_unsigned_16835_GENERIC_REAL g1(.A ({A[51], A[51:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16836_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [50:0] A;
  input CI;
  output [50:0] Z;
  wire [50:0] A;
  wire CI;
  wire [50:0] Z;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_104, A[0], CI);
  xor g51 (Z[1], A[1], n_104);
  and g52 (n_105, A[1], n_104);
  xor g53 (Z[2], A[2], n_105);
  and g54 (n_106, A[2], n_105);
  xor g55 (Z[3], A[3], n_106);
  and g56 (n_107, A[3], n_106);
  xor g57 (Z[4], A[4], n_107);
  and g58 (n_108, A[4], n_107);
  xor g59 (Z[5], A[5], n_108);
  and g60 (n_109, A[5], n_108);
  xor g61 (Z[6], A[6], n_109);
  and g62 (n_110, A[6], n_109);
  xor g63 (Z[7], A[7], n_110);
  and g64 (n_111, A[7], n_110);
  xor g65 (Z[8], A[8], n_111);
  and g66 (n_112, A[8], n_111);
  xor g67 (Z[9], A[9], n_112);
  and g68 (n_113, A[9], n_112);
  xor g69 (Z[10], A[10], n_113);
  and g70 (n_114, A[10], n_113);
  xor g71 (Z[11], A[11], n_114);
  and g72 (n_115, A[11], n_114);
  xor g73 (Z[12], A[12], n_115);
  and g74 (n_116, A[12], n_115);
  xor g75 (Z[13], A[13], n_116);
  and g76 (n_117, A[13], n_116);
  xor g77 (Z[14], A[14], n_117);
  and g78 (n_118, A[14], n_117);
  xor g79 (Z[15], A[15], n_118);
  and g80 (n_119, A[15], n_118);
  xor g81 (Z[16], A[16], n_119);
  and g82 (n_120, A[16], n_119);
  xor g83 (Z[17], A[17], n_120);
  and g84 (n_121, A[17], n_120);
  xor g85 (Z[18], A[18], n_121);
  and g86 (n_122, A[18], n_121);
  xor g87 (Z[19], A[19], n_122);
  and g88 (n_123, A[19], n_122);
  xor g89 (Z[20], A[20], n_123);
  and g90 (n_124, A[20], n_123);
  xor g91 (Z[21], A[21], n_124);
  and g92 (n_125, A[21], n_124);
  xor g93 (Z[22], A[22], n_125);
  and g94 (n_126, A[22], n_125);
  xor g95 (Z[23], A[23], n_126);
  and g96 (n_127, A[23], n_126);
  xor g97 (Z[24], A[24], n_127);
  and g98 (n_128, A[24], n_127);
  xor g99 (Z[25], A[25], n_128);
  and g100 (n_129, A[25], n_128);
  xor g101 (Z[26], A[26], n_129);
  and g102 (n_130, A[26], n_129);
  xor g103 (Z[27], A[27], n_130);
  and g104 (n_131, A[27], n_130);
  xor g105 (Z[28], A[28], n_131);
  and g106 (n_132, A[28], n_131);
  xor g107 (Z[29], A[29], n_132);
  and g108 (n_133, A[29], n_132);
  xor g109 (Z[30], A[30], n_133);
  and g110 (n_134, A[30], n_133);
  xor g111 (Z[31], A[31], n_134);
  and g112 (n_135, A[31], n_134);
  xor g113 (Z[32], A[32], n_135);
  and g114 (n_136, A[32], n_135);
  xor g115 (Z[33], A[33], n_136);
  and g116 (n_137, A[33], n_136);
  xor g117 (Z[34], A[34], n_137);
  and g118 (n_138, A[34], n_137);
  xor g119 (Z[35], A[35], n_138);
  and g120 (n_139, A[35], n_138);
  xor g121 (Z[36], A[36], n_139);
  and g122 (n_140, A[36], n_139);
  xor g123 (Z[37], A[37], n_140);
  and g124 (n_141, A[37], n_140);
  xor g125 (Z[38], A[38], n_141);
  and g126 (n_142, A[38], n_141);
  xor g127 (Z[39], A[39], n_142);
  and g128 (n_143, A[39], n_142);
  xor g129 (Z[40], A[40], n_143);
  and g130 (n_144, A[40], n_143);
  xor g131 (Z[41], A[41], n_144);
  and g132 (n_145, A[41], n_144);
  xor g133 (Z[42], A[42], n_145);
  and g134 (n_146, A[42], n_145);
  xor g135 (Z[43], A[43], n_146);
  and g136 (n_147, A[43], n_146);
  xor g137 (Z[44], A[44], n_147);
  and g138 (n_148, A[44], n_147);
  xor g139 (Z[45], A[45], n_148);
  and g140 (n_149, A[45], n_148);
  xor g141 (Z[46], A[46], n_149);
  and g142 (n_150, A[46], n_149);
  xor g143 (Z[47], A[47], n_150);
  and g144 (n_151, A[47], n_150);
  xor g145 (Z[48], A[48], n_151);
  and g146 (n_152, A[48], n_151);
  xor g147 (Z[49], A[49], n_152);
  and g148 (n_153, A[49], n_152);
  xor g149 (Z[50], A[50], n_153);
endmodule

module increment_unsigned_16836_GENERIC(A, CI, Z);
  input [50:0] A;
  input CI;
  output [50:0] Z;
  wire [50:0] A;
  wire CI;
  wire [50:0] Z;
  increment_unsigned_16836_GENERIC_REAL g1(.A ({A[49], A[49:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16837_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [49:0] A;
  input CI;
  output [49:0] Z;
  wire [49:0] A;
  wire CI;
  wire [49:0] Z;
  wire n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109;
  wire n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117;
  wire n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125;
  wire n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133;
  wire n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_102, A[0], CI);
  xor g50 (Z[1], A[1], n_102);
  and g51 (n_103, A[1], n_102);
  xor g52 (Z[2], A[2], n_103);
  and g53 (n_104, A[2], n_103);
  xor g54 (Z[3], A[3], n_104);
  and g55 (n_105, A[3], n_104);
  xor g56 (Z[4], A[4], n_105);
  and g57 (n_106, A[4], n_105);
  xor g58 (Z[5], A[5], n_106);
  and g59 (n_107, A[5], n_106);
  xor g60 (Z[6], A[6], n_107);
  and g61 (n_108, A[6], n_107);
  xor g62 (Z[7], A[7], n_108);
  and g63 (n_109, A[7], n_108);
  xor g64 (Z[8], A[8], n_109);
  and g65 (n_110, A[8], n_109);
  xor g66 (Z[9], A[9], n_110);
  and g67 (n_111, A[9], n_110);
  xor g68 (Z[10], A[10], n_111);
  and g69 (n_112, A[10], n_111);
  xor g70 (Z[11], A[11], n_112);
  and g71 (n_113, A[11], n_112);
  xor g72 (Z[12], A[12], n_113);
  and g73 (n_114, A[12], n_113);
  xor g74 (Z[13], A[13], n_114);
  and g75 (n_115, A[13], n_114);
  xor g76 (Z[14], A[14], n_115);
  and g77 (n_116, A[14], n_115);
  xor g78 (Z[15], A[15], n_116);
  and g79 (n_117, A[15], n_116);
  xor g80 (Z[16], A[16], n_117);
  and g81 (n_118, A[16], n_117);
  xor g82 (Z[17], A[17], n_118);
  and g83 (n_119, A[17], n_118);
  xor g84 (Z[18], A[18], n_119);
  and g85 (n_120, A[18], n_119);
  xor g86 (Z[19], A[19], n_120);
  and g87 (n_121, A[19], n_120);
  xor g88 (Z[20], A[20], n_121);
  and g89 (n_122, A[20], n_121);
  xor g90 (Z[21], A[21], n_122);
  and g91 (n_123, A[21], n_122);
  xor g92 (Z[22], A[22], n_123);
  and g93 (n_124, A[22], n_123);
  xor g94 (Z[23], A[23], n_124);
  and g95 (n_125, A[23], n_124);
  xor g96 (Z[24], A[24], n_125);
  and g97 (n_126, A[24], n_125);
  xor g98 (Z[25], A[25], n_126);
  and g99 (n_127, A[25], n_126);
  xor g100 (Z[26], A[26], n_127);
  and g101 (n_128, A[26], n_127);
  xor g102 (Z[27], A[27], n_128);
  and g103 (n_129, A[27], n_128);
  xor g104 (Z[28], A[28], n_129);
  and g105 (n_130, A[28], n_129);
  xor g106 (Z[29], A[29], n_130);
  and g107 (n_131, A[29], n_130);
  xor g108 (Z[30], A[30], n_131);
  and g109 (n_132, A[30], n_131);
  xor g110 (Z[31], A[31], n_132);
  and g111 (n_133, A[31], n_132);
  xor g112 (Z[32], A[32], n_133);
  and g113 (n_134, A[32], n_133);
  xor g114 (Z[33], A[33], n_134);
  and g115 (n_135, A[33], n_134);
  xor g116 (Z[34], A[34], n_135);
  and g117 (n_136, A[34], n_135);
  xor g118 (Z[35], A[35], n_136);
  and g119 (n_137, A[35], n_136);
  xor g120 (Z[36], A[36], n_137);
  and g121 (n_138, A[36], n_137);
  xor g122 (Z[37], A[37], n_138);
  and g123 (n_139, A[37], n_138);
  xor g124 (Z[38], A[38], n_139);
  and g125 (n_140, A[38], n_139);
  xor g126 (Z[39], A[39], n_140);
  and g127 (n_141, A[39], n_140);
  xor g128 (Z[40], A[40], n_141);
  and g129 (n_142, A[40], n_141);
  xor g130 (Z[41], A[41], n_142);
  and g131 (n_143, A[41], n_142);
  xor g132 (Z[42], A[42], n_143);
  and g133 (n_144, A[42], n_143);
  xor g134 (Z[43], A[43], n_144);
  and g135 (n_145, A[43], n_144);
  xor g136 (Z[44], A[44], n_145);
  and g137 (n_146, A[44], n_145);
  xor g138 (Z[45], A[45], n_146);
  and g139 (n_147, A[45], n_146);
  xor g140 (Z[46], A[46], n_147);
  and g141 (n_148, A[46], n_147);
  xor g142 (Z[47], A[47], n_148);
  and g143 (n_149, A[47], n_148);
  xor g144 (Z[48], A[48], n_149);
  and g145 (n_150, A[48], n_149);
  xor g146 (Z[49], A[49], n_150);
endmodule

module increment_unsigned_16837_GENERIC(A, CI, Z);
  input [49:0] A;
  input CI;
  output [49:0] Z;
  wire [49:0] A;
  wire CI;
  wire [49:0] Z;
  increment_unsigned_16837_GENERIC_REAL g1(.A ({A[48], A[48:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16838_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [47:0] A;
  input CI;
  output [47:0] Z;
  wire [47:0] A;
  wire CI;
  wire [47:0] Z;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_98, A[0], CI);
  xor g48 (Z[1], A[1], n_98);
  and g49 (n_99, A[1], n_98);
  xor g50 (Z[2], A[2], n_99);
  and g51 (n_100, A[2], n_99);
  xor g52 (Z[3], A[3], n_100);
  and g53 (n_101, A[3], n_100);
  xor g54 (Z[4], A[4], n_101);
  and g55 (n_102, A[4], n_101);
  xor g56 (Z[5], A[5], n_102);
  and g57 (n_103, A[5], n_102);
  xor g58 (Z[6], A[6], n_103);
  and g59 (n_104, A[6], n_103);
  xor g60 (Z[7], A[7], n_104);
  and g61 (n_105, A[7], n_104);
  xor g62 (Z[8], A[8], n_105);
  and g63 (n_106, A[8], n_105);
  xor g64 (Z[9], A[9], n_106);
  and g65 (n_107, A[9], n_106);
  xor g66 (Z[10], A[10], n_107);
  and g67 (n_108, A[10], n_107);
  xor g68 (Z[11], A[11], n_108);
  and g69 (n_109, A[11], n_108);
  xor g70 (Z[12], A[12], n_109);
  and g71 (n_110, A[12], n_109);
  xor g72 (Z[13], A[13], n_110);
  and g73 (n_111, A[13], n_110);
  xor g74 (Z[14], A[14], n_111);
  and g75 (n_112, A[14], n_111);
  xor g76 (Z[15], A[15], n_112);
  and g77 (n_113, A[15], n_112);
  xor g78 (Z[16], A[16], n_113);
  and g79 (n_114, A[16], n_113);
  xor g80 (Z[17], A[17], n_114);
  and g81 (n_115, A[17], n_114);
  xor g82 (Z[18], A[18], n_115);
  and g83 (n_116, A[18], n_115);
  xor g84 (Z[19], A[19], n_116);
  and g85 (n_117, A[19], n_116);
  xor g86 (Z[20], A[20], n_117);
  and g87 (n_118, A[20], n_117);
  xor g88 (Z[21], A[21], n_118);
  and g89 (n_119, A[21], n_118);
  xor g90 (Z[22], A[22], n_119);
  and g91 (n_120, A[22], n_119);
  xor g92 (Z[23], A[23], n_120);
  and g93 (n_121, A[23], n_120);
  xor g94 (Z[24], A[24], n_121);
  and g95 (n_122, A[24], n_121);
  xor g96 (Z[25], A[25], n_122);
  and g97 (n_123, A[25], n_122);
  xor g98 (Z[26], A[26], n_123);
  and g99 (n_124, A[26], n_123);
  xor g100 (Z[27], A[27], n_124);
  and g101 (n_125, A[27], n_124);
  xor g102 (Z[28], A[28], n_125);
  and g103 (n_126, A[28], n_125);
  xor g104 (Z[29], A[29], n_126);
  and g105 (n_127, A[29], n_126);
  xor g106 (Z[30], A[30], n_127);
  and g107 (n_128, A[30], n_127);
  xor g108 (Z[31], A[31], n_128);
  and g109 (n_129, A[31], n_128);
  xor g110 (Z[32], A[32], n_129);
  and g111 (n_130, A[32], n_129);
  xor g112 (Z[33], A[33], n_130);
  and g113 (n_131, A[33], n_130);
  xor g114 (Z[34], A[34], n_131);
  and g115 (n_132, A[34], n_131);
  xor g116 (Z[35], A[35], n_132);
  and g117 (n_133, A[35], n_132);
  xor g118 (Z[36], A[36], n_133);
  and g119 (n_134, A[36], n_133);
  xor g120 (Z[37], A[37], n_134);
  and g121 (n_135, A[37], n_134);
  xor g122 (Z[38], A[38], n_135);
  and g123 (n_136, A[38], n_135);
  xor g124 (Z[39], A[39], n_136);
  and g125 (n_137, A[39], n_136);
  xor g126 (Z[40], A[40], n_137);
  and g127 (n_138, A[40], n_137);
  xor g128 (Z[41], A[41], n_138);
  and g129 (n_139, A[41], n_138);
  xor g130 (Z[42], A[42], n_139);
  and g131 (n_140, A[42], n_139);
  xor g132 (Z[43], A[43], n_140);
  and g133 (n_141, A[43], n_140);
  xor g134 (Z[44], A[44], n_141);
  and g135 (n_142, A[44], n_141);
  xor g136 (Z[45], A[45], n_142);
  and g137 (n_143, A[45], n_142);
  xor g138 (Z[46], A[46], n_143);
  and g139 (n_144, A[46], n_143);
  xor g140 (Z[47], A[47], n_144);
endmodule

module increment_unsigned_16838_GENERIC(A, CI, Z);
  input [47:0] A;
  input CI;
  output [47:0] Z;
  wire [47:0] A;
  wire CI;
  wire [47:0] Z;
  increment_unsigned_16838_GENERIC_REAL g1(.A ({A[46], A[46:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16839_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [46:0] A;
  input CI;
  output [46:0] Z;
  wire [46:0] A;
  wire CI;
  wire [46:0] Z;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_96, A[0], CI);
  xor g47 (Z[1], A[1], n_96);
  and g48 (n_97, A[1], n_96);
  xor g49 (Z[2], A[2], n_97);
  and g50 (n_98, A[2], n_97);
  xor g51 (Z[3], A[3], n_98);
  and g52 (n_99, A[3], n_98);
  xor g53 (Z[4], A[4], n_99);
  and g54 (n_100, A[4], n_99);
  xor g55 (Z[5], A[5], n_100);
  and g56 (n_101, A[5], n_100);
  xor g57 (Z[6], A[6], n_101);
  and g58 (n_102, A[6], n_101);
  xor g59 (Z[7], A[7], n_102);
  and g60 (n_103, A[7], n_102);
  xor g61 (Z[8], A[8], n_103);
  and g62 (n_104, A[8], n_103);
  xor g63 (Z[9], A[9], n_104);
  and g64 (n_105, A[9], n_104);
  xor g65 (Z[10], A[10], n_105);
  and g66 (n_106, A[10], n_105);
  xor g67 (Z[11], A[11], n_106);
  and g68 (n_107, A[11], n_106);
  xor g69 (Z[12], A[12], n_107);
  and g70 (n_108, A[12], n_107);
  xor g71 (Z[13], A[13], n_108);
  and g72 (n_109, A[13], n_108);
  xor g73 (Z[14], A[14], n_109);
  and g74 (n_110, A[14], n_109);
  xor g75 (Z[15], A[15], n_110);
  and g76 (n_111, A[15], n_110);
  xor g77 (Z[16], A[16], n_111);
  and g78 (n_112, A[16], n_111);
  xor g79 (Z[17], A[17], n_112);
  and g80 (n_113, A[17], n_112);
  xor g81 (Z[18], A[18], n_113);
  and g82 (n_114, A[18], n_113);
  xor g83 (Z[19], A[19], n_114);
  and g84 (n_115, A[19], n_114);
  xor g85 (Z[20], A[20], n_115);
  and g86 (n_116, A[20], n_115);
  xor g87 (Z[21], A[21], n_116);
  and g88 (n_117, A[21], n_116);
  xor g89 (Z[22], A[22], n_117);
  and g90 (n_118, A[22], n_117);
  xor g91 (Z[23], A[23], n_118);
  and g92 (n_119, A[23], n_118);
  xor g93 (Z[24], A[24], n_119);
  and g94 (n_120, A[24], n_119);
  xor g95 (Z[25], A[25], n_120);
  and g96 (n_121, A[25], n_120);
  xor g97 (Z[26], A[26], n_121);
  and g98 (n_122, A[26], n_121);
  xor g99 (Z[27], A[27], n_122);
  and g100 (n_123, A[27], n_122);
  xor g101 (Z[28], A[28], n_123);
  and g102 (n_124, A[28], n_123);
  xor g103 (Z[29], A[29], n_124);
  and g104 (n_125, A[29], n_124);
  xor g105 (Z[30], A[30], n_125);
  and g106 (n_126, A[30], n_125);
  xor g107 (Z[31], A[31], n_126);
  and g108 (n_127, A[31], n_126);
  xor g109 (Z[32], A[32], n_127);
  and g110 (n_128, A[32], n_127);
  xor g111 (Z[33], A[33], n_128);
  and g112 (n_129, A[33], n_128);
  xor g113 (Z[34], A[34], n_129);
  and g114 (n_130, A[34], n_129);
  xor g115 (Z[35], A[35], n_130);
  and g116 (n_131, A[35], n_130);
  xor g117 (Z[36], A[36], n_131);
  and g118 (n_132, A[36], n_131);
  xor g119 (Z[37], A[37], n_132);
  and g120 (n_133, A[37], n_132);
  xor g121 (Z[38], A[38], n_133);
  and g122 (n_134, A[38], n_133);
  xor g123 (Z[39], A[39], n_134);
  and g124 (n_135, A[39], n_134);
  xor g125 (Z[40], A[40], n_135);
  and g126 (n_136, A[40], n_135);
  xor g127 (Z[41], A[41], n_136);
  and g128 (n_137, A[41], n_136);
  xor g129 (Z[42], A[42], n_137);
  and g130 (n_138, A[42], n_137);
  xor g131 (Z[43], A[43], n_138);
  and g132 (n_139, A[43], n_138);
  xor g133 (Z[44], A[44], n_139);
  and g134 (n_140, A[44], n_139);
  xor g135 (Z[45], A[45], n_140);
  and g136 (n_141, A[45], n_140);
  xor g137 (Z[46], A[46], n_141);
endmodule

module increment_unsigned_16839_GENERIC(A, CI, Z);
  input [46:0] A;
  input CI;
  output [46:0] Z;
  wire [46:0] A;
  wire CI;
  wire [46:0] Z;
  increment_unsigned_16839_GENERIC_REAL g1(.A ({A[45], A[45:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16840_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [44:0] A;
  input CI;
  output [44:0] Z;
  wire [44:0] A;
  wire CI;
  wire [44:0] Z;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_92, A[0], CI);
  xor g45 (Z[1], A[1], n_92);
  and g46 (n_93, A[1], n_92);
  xor g47 (Z[2], A[2], n_93);
  and g48 (n_94, A[2], n_93);
  xor g49 (Z[3], A[3], n_94);
  and g50 (n_95, A[3], n_94);
  xor g51 (Z[4], A[4], n_95);
  and g52 (n_96, A[4], n_95);
  xor g53 (Z[5], A[5], n_96);
  and g54 (n_97, A[5], n_96);
  xor g55 (Z[6], A[6], n_97);
  and g56 (n_98, A[6], n_97);
  xor g57 (Z[7], A[7], n_98);
  and g58 (n_99, A[7], n_98);
  xor g59 (Z[8], A[8], n_99);
  and g60 (n_100, A[8], n_99);
  xor g61 (Z[9], A[9], n_100);
  and g62 (n_101, A[9], n_100);
  xor g63 (Z[10], A[10], n_101);
  and g64 (n_102, A[10], n_101);
  xor g65 (Z[11], A[11], n_102);
  and g66 (n_103, A[11], n_102);
  xor g67 (Z[12], A[12], n_103);
  and g68 (n_104, A[12], n_103);
  xor g69 (Z[13], A[13], n_104);
  and g70 (n_105, A[13], n_104);
  xor g71 (Z[14], A[14], n_105);
  and g72 (n_106, A[14], n_105);
  xor g73 (Z[15], A[15], n_106);
  and g74 (n_107, A[15], n_106);
  xor g75 (Z[16], A[16], n_107);
  and g76 (n_108, A[16], n_107);
  xor g77 (Z[17], A[17], n_108);
  and g78 (n_109, A[17], n_108);
  xor g79 (Z[18], A[18], n_109);
  and g80 (n_110, A[18], n_109);
  xor g81 (Z[19], A[19], n_110);
  and g82 (n_111, A[19], n_110);
  xor g83 (Z[20], A[20], n_111);
  and g84 (n_112, A[20], n_111);
  xor g85 (Z[21], A[21], n_112);
  and g86 (n_113, A[21], n_112);
  xor g87 (Z[22], A[22], n_113);
  and g88 (n_114, A[22], n_113);
  xor g89 (Z[23], A[23], n_114);
  and g90 (n_115, A[23], n_114);
  xor g91 (Z[24], A[24], n_115);
  and g92 (n_116, A[24], n_115);
  xor g93 (Z[25], A[25], n_116);
  and g94 (n_117, A[25], n_116);
  xor g95 (Z[26], A[26], n_117);
  and g96 (n_118, A[26], n_117);
  xor g97 (Z[27], A[27], n_118);
  and g98 (n_119, A[27], n_118);
  xor g99 (Z[28], A[28], n_119);
  and g100 (n_120, A[28], n_119);
  xor g101 (Z[29], A[29], n_120);
  and g102 (n_121, A[29], n_120);
  xor g103 (Z[30], A[30], n_121);
  and g104 (n_122, A[30], n_121);
  xor g105 (Z[31], A[31], n_122);
  and g106 (n_123, A[31], n_122);
  xor g107 (Z[32], A[32], n_123);
  and g108 (n_124, A[32], n_123);
  xor g109 (Z[33], A[33], n_124);
  and g110 (n_125, A[33], n_124);
  xor g111 (Z[34], A[34], n_125);
  and g112 (n_126, A[34], n_125);
  xor g113 (Z[35], A[35], n_126);
  and g114 (n_127, A[35], n_126);
  xor g115 (Z[36], A[36], n_127);
  and g116 (n_128, A[36], n_127);
  xor g117 (Z[37], A[37], n_128);
  and g118 (n_129, A[37], n_128);
  xor g119 (Z[38], A[38], n_129);
  and g120 (n_130, A[38], n_129);
  xor g121 (Z[39], A[39], n_130);
  and g122 (n_131, A[39], n_130);
  xor g123 (Z[40], A[40], n_131);
  and g124 (n_132, A[40], n_131);
  xor g125 (Z[41], A[41], n_132);
  and g126 (n_133, A[41], n_132);
  xor g127 (Z[42], A[42], n_133);
  and g128 (n_134, A[42], n_133);
  xor g129 (Z[43], A[43], n_134);
  and g130 (n_135, A[43], n_134);
  xor g131 (Z[44], A[44], n_135);
endmodule

module increment_unsigned_16840_GENERIC(A, CI, Z);
  input [44:0] A;
  input CI;
  output [44:0] Z;
  wire [44:0] A;
  wire CI;
  wire [44:0] Z;
  increment_unsigned_16840_GENERIC_REAL g1(.A ({A[43], A[43:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16842_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [65:0] A;
  input CI;
  output [65:0] Z;
  wire [65:0] A;
  wire CI;
  wire [65:0] Z;
  wire n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_134, A[0], CI);
  xor g66 (Z[1], A[1], n_134);
  and g67 (n_135, A[1], n_134);
  xor g68 (Z[2], A[2], n_135);
  and g69 (n_136, A[2], n_135);
  xor g70 (Z[3], A[3], n_136);
  and g71 (n_137, A[3], n_136);
  xor g72 (Z[4], A[4], n_137);
  and g73 (n_138, A[4], n_137);
  xor g74 (Z[5], A[5], n_138);
  and g75 (n_139, A[5], n_138);
  xor g76 (Z[6], A[6], n_139);
  and g77 (n_140, A[6], n_139);
  xor g78 (Z[7], A[7], n_140);
  and g79 (n_141, A[7], n_140);
  xor g80 (Z[8], A[8], n_141);
  and g81 (n_142, A[8], n_141);
  xor g82 (Z[9], A[9], n_142);
  and g83 (n_143, A[9], n_142);
  xor g84 (Z[10], A[10], n_143);
  and g85 (n_144, A[10], n_143);
  xor g86 (Z[11], A[11], n_144);
  and g87 (n_145, A[11], n_144);
  xor g88 (Z[12], A[12], n_145);
  and g89 (n_146, A[12], n_145);
  xor g90 (Z[13], A[13], n_146);
  and g91 (n_147, A[13], n_146);
  xor g92 (Z[14], A[14], n_147);
  and g93 (n_148, A[14], n_147);
  xor g94 (Z[15], A[15], n_148);
  and g95 (n_149, A[15], n_148);
  xor g96 (Z[16], A[16], n_149);
  and g97 (n_150, A[16], n_149);
  xor g98 (Z[17], A[17], n_150);
  and g99 (n_151, A[17], n_150);
  xor g100 (Z[18], A[18], n_151);
  and g101 (n_152, A[18], n_151);
  xor g102 (Z[19], A[19], n_152);
  and g103 (n_153, A[19], n_152);
  xor g104 (Z[20], A[20], n_153);
  and g105 (n_154, A[20], n_153);
  xor g106 (Z[21], A[21], n_154);
  and g107 (n_155, A[21], n_154);
  xor g108 (Z[22], A[22], n_155);
  and g109 (n_156, A[22], n_155);
  xor g110 (Z[23], A[23], n_156);
  and g111 (n_157, A[23], n_156);
  xor g112 (Z[24], A[24], n_157);
  and g113 (n_158, A[24], n_157);
  xor g114 (Z[25], A[25], n_158);
  and g115 (n_159, A[25], n_158);
  xor g116 (Z[26], A[26], n_159);
  and g117 (n_160, A[26], n_159);
  xor g118 (Z[27], A[27], n_160);
  and g119 (n_161, A[27], n_160);
  xor g120 (Z[28], A[28], n_161);
  and g121 (n_162, A[28], n_161);
  xor g122 (Z[29], A[29], n_162);
  and g123 (n_163, A[29], n_162);
  xor g124 (Z[30], A[30], n_163);
  and g125 (n_164, A[30], n_163);
  xor g126 (Z[31], A[31], n_164);
  and g127 (n_165, A[31], n_164);
  xor g128 (Z[32], A[32], n_165);
  and g129 (n_166, A[32], n_165);
  xor g130 (Z[33], A[33], n_166);
  and g131 (n_167, A[33], n_166);
  xor g132 (Z[34], A[34], n_167);
  and g133 (n_168, A[34], n_167);
  xor g134 (Z[35], A[35], n_168);
  and g135 (n_169, A[35], n_168);
  xor g136 (Z[36], A[36], n_169);
  and g137 (n_170, A[36], n_169);
  xor g138 (Z[37], A[37], n_170);
  and g139 (n_171, A[37], n_170);
  xor g140 (Z[38], A[38], n_171);
  and g141 (n_172, A[38], n_171);
  xor g142 (Z[39], A[39], n_172);
  and g143 (n_173, A[39], n_172);
  xor g144 (Z[40], A[40], n_173);
  and g145 (n_174, A[40], n_173);
  xor g146 (Z[41], A[41], n_174);
  and g147 (n_175, A[41], n_174);
  xor g148 (Z[42], A[42], n_175);
  and g149 (n_176, A[42], n_175);
  xor g150 (Z[43], A[43], n_176);
  and g151 (n_177, A[43], n_176);
  xor g152 (Z[44], A[44], n_177);
  and g153 (n_178, A[44], n_177);
  xor g154 (Z[45], A[45], n_178);
  and g155 (n_179, A[45], n_178);
  xor g156 (Z[46], A[46], n_179);
  and g157 (n_180, A[46], n_179);
  xor g158 (Z[47], A[47], n_180);
  and g159 (n_181, A[47], n_180);
  xor g160 (Z[48], A[48], n_181);
  and g161 (n_182, A[48], n_181);
  xor g162 (Z[49], A[49], n_182);
  and g163 (n_183, A[49], n_182);
  xor g164 (Z[50], A[50], n_183);
  and g165 (n_184, A[50], n_183);
  xor g166 (Z[51], A[51], n_184);
  and g167 (n_185, A[51], n_184);
  xor g168 (Z[52], A[52], n_185);
  and g169 (n_186, A[52], n_185);
  xor g170 (Z[53], A[53], n_186);
  and g171 (n_187, A[53], n_186);
  xor g172 (Z[54], A[54], n_187);
  and g173 (n_188, A[54], n_187);
  xor g174 (Z[55], A[55], n_188);
  and g175 (n_189, A[55], n_188);
  xor g176 (Z[56], A[56], n_189);
  and g177 (n_190, A[56], n_189);
  xor g178 (Z[57], A[57], n_190);
  and g179 (n_191, A[57], n_190);
  xor g180 (Z[58], A[58], n_191);
  and g181 (n_192, A[58], n_191);
  xor g182 (Z[59], A[59], n_192);
  and g183 (n_193, A[59], n_192);
  xor g184 (Z[60], A[60], n_193);
  and g185 (n_194, A[60], n_193);
  xor g186 (Z[61], A[61], n_194);
  and g187 (n_195, A[61], n_194);
  xor g188 (Z[62], A[62], n_195);
  and g189 (n_196, A[62], n_195);
  xor g190 (Z[63], A[63], n_196);
  and g191 (n_197, A[63], n_196);
  xor g192 (Z[64], A[64], n_197);
  and g193 (n_198, A[64], n_197);
  xor g194 (Z[65], A[65], n_198);
endmodule

module increment_unsigned_16842_GENERIC(A, CI, Z);
  input [65:0] A;
  input CI;
  output [65:0] Z;
  wire [65:0] A;
  wire CI;
  wire [65:0] Z;
  increment_unsigned_16842_GENERIC_REAL g1(.A ({A[64], A[64:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_16843_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [63:0] A;
  input CI;
  output [63:0] Z;
  wire [63:0] A;
  wire CI;
  wire [63:0] Z;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_130, A[0], CI);
  xor g64 (Z[1], A[1], n_130);
  and g65 (n_131, A[1], n_130);
  xor g66 (Z[2], A[2], n_131);
  and g67 (n_132, A[2], n_131);
  xor g68 (Z[3], A[3], n_132);
  and g69 (n_133, A[3], n_132);
  xor g70 (Z[4], A[4], n_133);
  and g71 (n_134, A[4], n_133);
  xor g72 (Z[5], A[5], n_134);
  and g73 (n_135, A[5], n_134);
  xor g74 (Z[6], A[6], n_135);
  and g75 (n_136, A[6], n_135);
  xor g76 (Z[7], A[7], n_136);
  and g77 (n_137, A[7], n_136);
  xor g78 (Z[8], A[8], n_137);
  and g79 (n_138, A[8], n_137);
  xor g80 (Z[9], A[9], n_138);
  and g81 (n_139, A[9], n_138);
  xor g82 (Z[10], A[10], n_139);
  and g83 (n_140, A[10], n_139);
  xor g84 (Z[11], A[11], n_140);
  and g85 (n_141, A[11], n_140);
  xor g86 (Z[12], A[12], n_141);
  and g87 (n_142, A[12], n_141);
  xor g88 (Z[13], A[13], n_142);
  and g89 (n_143, A[13], n_142);
  xor g90 (Z[14], A[14], n_143);
  and g91 (n_144, A[14], n_143);
  xor g92 (Z[15], A[15], n_144);
  and g93 (n_145, A[15], n_144);
  xor g94 (Z[16], A[16], n_145);
  and g95 (n_146, A[16], n_145);
  xor g96 (Z[17], A[17], n_146);
  and g97 (n_147, A[17], n_146);
  xor g98 (Z[18], A[18], n_147);
  and g99 (n_148, A[18], n_147);
  xor g100 (Z[19], A[19], n_148);
  and g101 (n_149, A[19], n_148);
  xor g102 (Z[20], A[20], n_149);
  and g103 (n_150, A[20], n_149);
  xor g104 (Z[21], A[21], n_150);
  and g105 (n_151, A[21], n_150);
  xor g106 (Z[22], A[22], n_151);
  and g107 (n_152, A[22], n_151);
  xor g108 (Z[23], A[23], n_152);
  and g109 (n_153, A[23], n_152);
  xor g110 (Z[24], A[24], n_153);
  and g111 (n_154, A[24], n_153);
  xor g112 (Z[25], A[25], n_154);
  and g113 (n_155, A[25], n_154);
  xor g114 (Z[26], A[26], n_155);
  and g115 (n_156, A[26], n_155);
  xor g116 (Z[27], A[27], n_156);
  and g117 (n_157, A[27], n_156);
  xor g118 (Z[28], A[28], n_157);
  and g119 (n_158, A[28], n_157);
  xor g120 (Z[29], A[29], n_158);
  and g121 (n_159, A[29], n_158);
  xor g122 (Z[30], A[30], n_159);
  and g123 (n_160, A[30], n_159);
  xor g124 (Z[31], A[31], n_160);
  and g125 (n_161, A[31], n_160);
  xor g126 (Z[32], A[32], n_161);
  and g127 (n_162, A[32], n_161);
  xor g128 (Z[33], A[33], n_162);
  and g129 (n_163, A[33], n_162);
  xor g130 (Z[34], A[34], n_163);
  and g131 (n_164, A[34], n_163);
  xor g132 (Z[35], A[35], n_164);
  and g133 (n_165, A[35], n_164);
  xor g134 (Z[36], A[36], n_165);
  and g135 (n_166, A[36], n_165);
  xor g136 (Z[37], A[37], n_166);
  and g137 (n_167, A[37], n_166);
  xor g138 (Z[38], A[38], n_167);
  and g139 (n_168, A[38], n_167);
  xor g140 (Z[39], A[39], n_168);
  and g141 (n_169, A[39], n_168);
  xor g142 (Z[40], A[40], n_169);
  and g143 (n_170, A[40], n_169);
  xor g144 (Z[41], A[41], n_170);
  and g145 (n_171, A[41], n_170);
  xor g146 (Z[42], A[42], n_171);
  and g147 (n_172, A[42], n_171);
  xor g148 (Z[43], A[43], n_172);
  and g149 (n_173, A[43], n_172);
  xor g150 (Z[44], A[44], n_173);
  and g151 (n_174, A[44], n_173);
  xor g152 (Z[45], A[45], n_174);
  and g153 (n_175, A[45], n_174);
  xor g154 (Z[46], A[46], n_175);
  and g155 (n_176, A[46], n_175);
  xor g156 (Z[47], A[47], n_176);
  and g157 (n_177, A[47], n_176);
  xor g158 (Z[48], A[48], n_177);
  and g159 (n_178, A[48], n_177);
  xor g160 (Z[49], A[49], n_178);
  and g161 (n_179, A[49], n_178);
  xor g162 (Z[50], A[50], n_179);
  and g163 (n_180, A[50], n_179);
  xor g164 (Z[51], A[51], n_180);
  and g165 (n_181, A[51], n_180);
  xor g166 (Z[52], A[52], n_181);
  and g167 (n_182, A[52], n_181);
  xor g168 (Z[53], A[53], n_182);
  and g169 (n_183, A[53], n_182);
  xor g170 (Z[54], A[54], n_183);
  and g171 (n_184, A[54], n_183);
  xor g172 (Z[55], A[55], n_184);
  and g173 (n_185, A[55], n_184);
  xor g174 (Z[56], A[56], n_185);
  and g175 (n_186, A[56], n_185);
  xor g176 (Z[57], A[57], n_186);
  and g177 (n_187, A[57], n_186);
  xor g178 (Z[58], A[58], n_187);
  and g179 (n_188, A[58], n_187);
  xor g180 (Z[59], A[59], n_188);
  and g181 (n_189, A[59], n_188);
  xor g182 (Z[60], A[60], n_189);
  and g183 (n_190, A[60], n_189);
  xor g184 (Z[61], A[61], n_190);
  and g185 (n_191, A[61], n_190);
  xor g186 (Z[62], A[62], n_191);
  and g187 (n_192, A[62], n_191);
  xor g188 (Z[63], A[63], n_192);
endmodule

module increment_unsigned_16843_GENERIC(A, CI, Z);
  input [63:0] A;
  input CI;
  output [63:0] Z;
  wire [63:0] A;
  wire CI;
  wire [63:0] Z;
  increment_unsigned_16843_GENERIC_REAL g1(.A ({A[62], A[62:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_9286_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [42:0] A;
  input CI;
  output [42:0] Z;
  wire [42:0] A;
  wire CI;
  wire [42:0] Z;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_88, A[0], CI);
  xor g43 (Z[1], A[1], n_88);
  and g44 (n_89, A[1], n_88);
  xor g45 (Z[2], A[2], n_89);
  and g46 (n_90, A[2], n_89);
  xor g47 (Z[3], A[3], n_90);
  and g48 (n_91, A[3], n_90);
  xor g49 (Z[4], A[4], n_91);
  and g50 (n_92, A[4], n_91);
  xor g51 (Z[5], A[5], n_92);
  and g52 (n_93, A[5], n_92);
  xor g53 (Z[6], A[6], n_93);
  and g54 (n_94, A[6], n_93);
  xor g55 (Z[7], A[7], n_94);
  and g56 (n_95, A[7], n_94);
  xor g57 (Z[8], A[8], n_95);
  and g58 (n_96, A[8], n_95);
  xor g59 (Z[9], A[9], n_96);
  and g60 (n_97, A[9], n_96);
  xor g61 (Z[10], A[10], n_97);
  and g62 (n_98, A[10], n_97);
  xor g63 (Z[11], A[11], n_98);
  and g64 (n_99, A[11], n_98);
  xor g65 (Z[12], A[12], n_99);
  and g66 (n_100, A[12], n_99);
  xor g67 (Z[13], A[13], n_100);
  and g68 (n_101, A[13], n_100);
  xor g69 (Z[14], A[14], n_101);
  and g70 (n_102, A[14], n_101);
  xor g71 (Z[15], A[15], n_102);
  and g72 (n_103, A[15], n_102);
  xor g73 (Z[16], A[16], n_103);
  and g74 (n_104, A[16], n_103);
  xor g75 (Z[17], A[17], n_104);
  and g76 (n_105, A[17], n_104);
  xor g77 (Z[18], A[18], n_105);
  and g78 (n_106, A[18], n_105);
  xor g79 (Z[19], A[19], n_106);
  and g80 (n_107, A[19], n_106);
  xor g81 (Z[20], A[20], n_107);
  and g82 (n_108, A[20], n_107);
  xor g83 (Z[21], A[21], n_108);
  and g84 (n_109, A[21], n_108);
  xor g85 (Z[22], A[22], n_109);
  and g86 (n_110, A[22], n_109);
  xor g87 (Z[23], A[23], n_110);
  and g88 (n_111, A[23], n_110);
  xor g89 (Z[24], A[24], n_111);
  and g90 (n_112, A[24], n_111);
  xor g91 (Z[25], A[25], n_112);
  and g92 (n_113, A[25], n_112);
  xor g93 (Z[26], A[26], n_113);
  and g94 (n_114, A[26], n_113);
  xor g95 (Z[27], A[27], n_114);
  and g96 (n_115, A[27], n_114);
  xor g97 (Z[28], A[28], n_115);
  and g98 (n_116, A[28], n_115);
  xor g99 (Z[29], A[29], n_116);
  and g100 (n_117, A[29], n_116);
  xor g101 (Z[30], A[30], n_117);
  and g102 (n_118, A[30], n_117);
  xor g103 (Z[31], A[31], n_118);
  and g104 (n_119, A[31], n_118);
  xor g105 (Z[32], A[32], n_119);
  and g106 (n_120, A[32], n_119);
  xor g107 (Z[33], A[33], n_120);
  and g108 (n_121, A[33], n_120);
  xor g109 (Z[34], A[34], n_121);
  and g110 (n_122, A[34], n_121);
  xor g111 (Z[35], A[35], n_122);
  and g112 (n_123, A[35], n_122);
  xor g113 (Z[36], A[36], n_123);
  and g114 (n_124, A[36], n_123);
  xor g115 (Z[37], A[37], n_124);
  and g116 (n_125, A[37], n_124);
  xor g117 (Z[38], A[38], n_125);
  and g118 (n_126, A[38], n_125);
  xor g119 (Z[39], A[39], n_126);
  and g120 (n_127, A[39], n_126);
  xor g121 (Z[40], A[40], n_127);
  and g122 (n_128, A[40], n_127);
  xor g123 (Z[41], A[41], n_128);
  and g124 (n_129, A[41], n_128);
  xor g125 (Z[42], A[42], n_129);
endmodule

module increment_unsigned_9286_GENERIC(A, CI, Z);
  input [42:0] A;
  input CI;
  output [42:0] Z;
  wire [42:0] A;
  wire CI;
  wire [42:0] Z;
  increment_unsigned_9286_GENERIC_REAL g1(.A ({A[41], A[41:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_9286_1_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [42:0] A;
  input CI;
  output [42:0] Z;
  wire [42:0] A;
  wire CI;
  wire [42:0] Z;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129;
  xor g1 (Z[0], A[0], CI);
  and g2 (n_88, A[0], CI);
  xor g43 (Z[1], A[1], n_88);
  and g44 (n_89, A[1], n_88);
  xor g45 (Z[2], A[2], n_89);
  and g46 (n_90, A[2], n_89);
  xor g47 (Z[3], A[3], n_90);
  and g48 (n_91, A[3], n_90);
  xor g49 (Z[4], A[4], n_91);
  and g50 (n_92, A[4], n_91);
  xor g51 (Z[5], A[5], n_92);
  and g52 (n_93, A[5], n_92);
  xor g53 (Z[6], A[6], n_93);
  and g54 (n_94, A[6], n_93);
  xor g55 (Z[7], A[7], n_94);
  and g56 (n_95, A[7], n_94);
  xor g57 (Z[8], A[8], n_95);
  and g58 (n_96, A[8], n_95);
  xor g59 (Z[9], A[9], n_96);
  and g60 (n_97, A[9], n_96);
  xor g61 (Z[10], A[10], n_97);
  and g62 (n_98, A[10], n_97);
  xor g63 (Z[11], A[11], n_98);
  and g64 (n_99, A[11], n_98);
  xor g65 (Z[12], A[12], n_99);
  and g66 (n_100, A[12], n_99);
  xor g67 (Z[13], A[13], n_100);
  and g68 (n_101, A[13], n_100);
  xor g69 (Z[14], A[14], n_101);
  and g70 (n_102, A[14], n_101);
  xor g71 (Z[15], A[15], n_102);
  and g72 (n_103, A[15], n_102);
  xor g73 (Z[16], A[16], n_103);
  and g74 (n_104, A[16], n_103);
  xor g75 (Z[17], A[17], n_104);
  and g76 (n_105, A[17], n_104);
  xor g77 (Z[18], A[18], n_105);
  and g78 (n_106, A[18], n_105);
  xor g79 (Z[19], A[19], n_106);
  and g80 (n_107, A[19], n_106);
  xor g81 (Z[20], A[20], n_107);
  and g82 (n_108, A[20], n_107);
  xor g83 (Z[21], A[21], n_108);
  and g84 (n_109, A[21], n_108);
  xor g85 (Z[22], A[22], n_109);
  and g86 (n_110, A[22], n_109);
  xor g87 (Z[23], A[23], n_110);
  and g88 (n_111, A[23], n_110);
  xor g89 (Z[24], A[24], n_111);
  and g90 (n_112, A[24], n_111);
  xor g91 (Z[25], A[25], n_112);
  and g92 (n_113, A[25], n_112);
  xor g93 (Z[26], A[26], n_113);
  and g94 (n_114, A[26], n_113);
  xor g95 (Z[27], A[27], n_114);
  and g96 (n_115, A[27], n_114);
  xor g97 (Z[28], A[28], n_115);
  and g98 (n_116, A[28], n_115);
  xor g99 (Z[29], A[29], n_116);
  and g100 (n_117, A[29], n_116);
  xor g101 (Z[30], A[30], n_117);
  and g102 (n_118, A[30], n_117);
  xor g103 (Z[31], A[31], n_118);
  and g104 (n_119, A[31], n_118);
  xor g105 (Z[32], A[32], n_119);
  and g106 (n_120, A[32], n_119);
  xor g107 (Z[33], A[33], n_120);
  and g108 (n_121, A[33], n_120);
  xor g109 (Z[34], A[34], n_121);
  and g110 (n_122, A[34], n_121);
  xor g111 (Z[35], A[35], n_122);
  and g112 (n_123, A[35], n_122);
  xor g113 (Z[36], A[36], n_123);
  and g114 (n_124, A[36], n_123);
  xor g115 (Z[37], A[37], n_124);
  and g116 (n_125, A[37], n_124);
  xor g117 (Z[38], A[38], n_125);
  and g118 (n_126, A[38], n_125);
  xor g119 (Z[39], A[39], n_126);
  and g120 (n_127, A[39], n_126);
  xor g121 (Z[40], A[40], n_127);
  and g122 (n_128, A[40], n_127);
  xor g123 (Z[41], A[41], n_128);
  and g124 (n_129, A[41], n_128);
  xor g125 (Z[42], A[42], n_129);
endmodule

module increment_unsigned_9286_1_GENERIC(A, CI, Z);
  input [42:0] A;
  input CI;
  output [42:0] Z;
  wire [42:0] A;
  wire CI;
  wire [42:0] Z;
  increment_unsigned_9286_1_GENERIC_REAL g1(.A ({A[41], A[41:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_9286_2_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [42:0] A;
  input CI;
  output [42:0] Z;
  wire [42:0] A;
  wire CI;
  wire [42:0] Z;
  wire n_88, n_90, n_91, n_93, n_95, n_96, n_98, n_99;
  wire n_101, n_102, n_104, n_105, n_107, n_108, n_110, n_111;
  wire n_113, n_114, n_116, n_117, n_119, n_120, n_122, n_124;
  wire n_126, n_128, n_130, n_131, n_132, n_134, n_135, n_136;
  wire n_138, n_139, n_140, n_142, n_143, n_144, n_146, n_147;
  wire n_149, n_151, n_153, n_155, n_157, n_160, n_161, n_162;
  wire n_163, n_164, n_168, n_170, n_173, n_174, n_175, n_176;
  wire n_178, n_180, n_182, n_184, n_186, n_188, n_190, n_192;
  wire n_194, n_195, n_197, n_199, n_202, n_203, n_206, n_209;
  wire n_210, n_211, n_212, n_214, n_216, n_218, n_220, n_222;
  wire n_224, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_244, n_246, n_248, n_250, n_252, n_254, n_256;
  wire n_258, n_260;
  nand g1 (n_88, A[0], CI);
  nand g4 (n_91, A[2], A[3]);
  nand g5 (n_93, A[4], A[5]);
  nand g6 (n_95, A[6], A[7]);
  nand g7 (n_96, A[8], A[9]);
  nand g8 (n_98, A[10], A[11]);
  nand g9 (n_99, A[12], A[13]);
  nand g10 (n_101, A[14], A[15]);
  nand g11 (n_102, A[16], A[17]);
  nand g12 (n_104, A[18], A[19]);
  nand g13 (n_105, A[20], A[21]);
  nand g14 (n_107, A[22], A[23]);
  nand g15 (n_108, A[24], A[25]);
  nand g16 (n_110, A[26], A[27]);
  nand g17 (n_111, A[28], A[29]);
  nand g18 (n_113, A[30], A[31]);
  nand g19 (n_114, A[32], A[33]);
  nand g20 (n_116, A[34], A[35]);
  nand g21 (n_117, A[36], A[37]);
  nand g22 (n_119, A[38], A[39]);
  nand g23 (n_120, A[40], A[41]);
  nand g24 (n_206, A[2], n_90);
  nor g29 (n_126, n_93, n_95);
  nor g32 (n_128, n_96, n_98);
  nor g35 (n_131, n_99, n_101);
  nor g38 (n_132, n_102, n_104);
  nor g41 (n_135, n_105, n_107);
  nor g44 (n_136, n_108, n_110);
  nor g47 (n_139, n_111, n_113);
  nor g50 (n_140, n_114, n_116);
  nor g53 (n_143, n_117, n_119);
  nor g58 (n_210, n_93, n_122);
  nand g63 (n_147, A[12], n_128);
  nand g66 (n_151, n_128, n_130);
  nand g67 (n_153, n_128, n_131);
  nand g68 (n_173, A[20], n_132);
  nand g71 (n_175, n_132, n_134);
  nand g72 (n_155, n_132, n_135);
  nand g73 (n_160, A[28], n_136);
  nand g76 (n_162, n_136, n_138);
  nand g77 (n_163, n_136, n_139);
  nand g78 (n_195, A[36], n_140);
  nand g81 (n_199, n_140, n_142);
  nand g82 (n_164, n_140, n_143);
  nand g83 (n_212, A[8], n_144);
  nand g86 (n_216, n_146, n_144);
  nand g87 (n_218, n_128, n_144);
  nor g98 (n_178, n_108, n_155);
  nor g103 (n_184, n_155, n_160);
  nor g104 (n_186, n_155, n_161);
  nor g105 (n_188, n_155, n_162);
  nor g106 (n_190, n_155, n_163);
  nor g109 (n_203, n_120, n_164);
  nor g114 (n_228, n_102, n_168);
  nor g119 (n_231, n_173, n_168);
  nor g120 (n_232, n_174, n_168);
  nor g121 (n_233, n_175, n_168);
  nor g122 (n_234, n_155, n_168);
  nand g139 (n_242, A[32], n_192);
  nand g142 (n_246, n_194, n_192);
  nand g143 (n_248, n_140, n_192);
  nand g152 (n_258, n_202, n_192);
  nand g153 (n_260, n_203, n_192);
  xor g155 (Z[0], A[0], CI);
  xor g158 (Z[2], A[2], n_90);
  xor g163 (Z[5], A[5], n_209);
  xor g164 (Z[6], A[6], n_210);
  xor g165 (Z[7], A[7], n_211);
  xor g166 (Z[8], A[8], n_144);
  xor g183 (Z[17], A[17], n_227);
  xor g184 (Z[18], A[18], n_228);
  xor g185 (Z[19], A[19], n_229);
  xor g186 (Z[20], A[20], n_230);
  xor g187 (Z[21], A[21], n_231);
  xor g188 (Z[22], A[22], n_232);
  xor g189 (Z[23], A[23], n_233);
  xor g190 (Z[24], A[24], n_234);
  xor g191 (Z[25], A[25], n_235);
  xor g192 (Z[26], A[26], n_236);
  xor g193 (Z[27], A[27], n_237);
  xor g194 (Z[28], A[28], n_238);
  xor g195 (Z[29], A[29], n_239);
  xor g196 (Z[30], A[30], n_240);
  xor g197 (Z[31], A[31], n_241);
  xor g198 (Z[32], A[32], n_192);
  and g220 (n_90, A[1], wc);
  not gc (wc, n_88);
  and g221 (n_124, A[6], wc0);
  not gc0 (wc0, n_93);
  and g222 (n_146, A[10], wc1);
  not gc1 (wc1, n_96);
  and g223 (n_130, A[14], wc2);
  not gc2 (wc2, n_99);
  and g224 (n_170, A[18], wc3);
  not gc3 (wc3, n_102);
  and g225 (n_134, A[22], wc4);
  not gc4 (wc4, n_105);
  and g226 (n_157, A[26], wc5);
  not gc5 (wc5, n_108);
  and g227 (n_138, A[30], wc6);
  not gc6 (wc6, n_111);
  and g228 (n_194, A[34], wc7);
  not gc7 (wc7, n_114);
  and g229 (n_142, A[38], wc8);
  not gc8 (wc8, n_117);
  or g230 (n_122, wc9, n_91);
  not gc9 (wc9, n_90);
  or g231 (n_149, wc10, n_99);
  not gc10 (wc10, n_128);
  or g232 (n_174, wc11, n_105);
  not gc11 (wc11, n_132);
  or g233 (n_161, wc12, n_111);
  not gc12 (wc12, n_136);
  or g234 (n_197, wc13, n_117);
  not gc13 (wc13, n_140);
  xnor g235 (Z[1], n_88, A[1]);
  and g236 (n_209, A[4], wc14);
  not gc14 (wc14, n_122);
  and g237 (n_211, wc15, n_124);
  not gc15 (wc15, n_122);
  and g238 (n_144, wc16, n_126);
  not gc16 (wc16, n_122);
  and g239 (n_176, A[24], wc17);
  not gc17 (wc17, n_155);
  and g240 (n_180, n_157, wc18);
  not gc18 (wc18, n_155);
  and g241 (n_182, wc19, n_136);
  not gc19 (wc19, n_155);
  and g242 (n_202, A[40], wc20);
  not gc20 (wc20, n_164);
  or g243 (n_214, wc21, n_96);
  not gc21 (wc21, n_144);
  or g244 (n_220, wc22, n_147);
  not gc22 (wc22, n_144);
  or g245 (n_222, wc23, n_149);
  not gc23 (wc23, n_144);
  or g246 (n_224, wc24, n_151);
  not gc24 (wc24, n_144);
  or g247 (n_168, wc25, n_153);
  not gc25 (wc25, n_144);
  xnor g248 (Z[3], n_206, A[3]);
  xnor g249 (Z[4], n_122, A[4]);
  and g250 (n_227, A[16], wc26);
  not gc26 (wc26, n_168);
  and g251 (n_229, wc27, n_170);
  not gc27 (wc27, n_168);
  and g252 (n_230, wc28, n_132);
  not gc28 (wc28, n_168);
  and g253 (n_235, wc29, n_176);
  not gc29 (wc29, n_168);
  and g254 (n_236, wc30, n_178);
  not gc30 (wc30, n_168);
  and g255 (n_237, wc31, n_180);
  not gc31 (wc31, n_168);
  and g256 (n_238, wc32, n_182);
  not gc32 (wc32, n_168);
  and g257 (n_239, wc33, n_184);
  not gc33 (wc33, n_168);
  and g258 (n_240, wc34, n_186);
  not gc34 (wc34, n_168);
  and g259 (n_241, wc35, n_188);
  not gc35 (wc35, n_168);
  and g260 (n_192, wc36, n_190);
  not gc36 (wc36, n_168);
  or g261 (n_244, wc37, n_114);
  not gc37 (wc37, n_192);
  or g262 (n_250, wc38, n_195);
  not gc38 (wc38, n_192);
  or g263 (n_252, wc39, n_197);
  not gc39 (wc39, n_192);
  or g264 (n_254, wc40, n_199);
  not gc40 (wc40, n_192);
  or g265 (n_256, wc41, n_164);
  not gc41 (wc41, n_192);
  xnor g266 (Z[9], n_212, A[9]);
  xnor g267 (Z[10], n_214, A[10]);
  xnor g268 (Z[11], n_216, A[11]);
  xnor g269 (Z[12], n_218, A[12]);
  xnor g270 (Z[13], n_220, A[13]);
  xnor g271 (Z[14], n_222, A[14]);
  xnor g272 (Z[15], n_224, A[15]);
  xnor g273 (Z[16], n_168, A[16]);
  xnor g274 (Z[33], n_242, A[33]);
  xnor g275 (Z[34], n_244, A[34]);
  xnor g276 (Z[35], n_246, A[35]);
  xnor g277 (Z[36], n_248, A[36]);
  xnor g278 (Z[37], n_250, A[37]);
  xnor g279 (Z[38], n_252, A[38]);
  xnor g280 (Z[39], n_254, A[39]);
  xnor g281 (Z[40], n_256, A[40]);
  xnor g282 (Z[41], n_258, A[41]);
  xnor g283 (Z[42], n_260, A[42]);
endmodule

module increment_unsigned_9286_2_GENERIC(A, CI, Z);
  input [42:0] A;
  input CI;
  output [42:0] Z;
  wire [42:0] A;
  wire CI;
  wire [42:0] Z;
  increment_unsigned_9286_2_GENERIC_REAL g1(.A ({A[41], A[41:0]}), .CI
       (CI), .Z (Z));
endmodule

module increment_unsigned_9286_3_GENERIC_REAL(A, CI, Z);
// synthesis_equation increment_unsigned
  input [42:0] A;
  input CI;
  output [42:0] Z;
  wire [42:0] A;
  wire CI;
  wire [42:0] Z;
  wire n_88, n_90, n_91, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_125, n_126, n_127, n_128, n_130, n_131, n_134;
  wire n_136, n_137, n_140, n_142, n_143, n_144, n_146, n_147;
  wire n_150, n_152, n_153, n_155, n_158, n_159, n_162, n_164;
  wire n_166, n_169, n_170, n_172, n_175, n_177, n_178, n_181;
  wire n_182, n_184, n_187, n_188, n_191, n_193, n_194, n_196;
  wire n_199, n_201, n_202, n_205;
  nand g1 (n_88, A[0], CI);
  nand g4 (n_90, A[2], A[3]);
  nand g5 (n_93, A[4], A[5]);
  nand g6 (n_94, A[6], A[7]);
  nand g7 (n_95, A[8], A[9]);
  nand g8 (n_96, A[10], A[11]);
  nand g9 (n_97, A[12], A[13]);
  nand g10 (n_98, A[14], A[15]);
  nand g11 (n_99, A[16], A[17]);
  nand g12 (n_100, A[18], A[19]);
  nand g13 (n_101, A[20], A[21]);
  nand g14 (n_102, A[22], A[23]);
  nand g15 (n_103, A[24], A[25]);
  nand g16 (n_104, A[26], A[27]);
  nand g17 (n_105, A[28], A[29]);
  nand g18 (n_106, A[30], A[31]);
  nand g19 (n_107, A[32], A[33]);
  nand g20 (n_108, A[34], A[35]);
  nand g21 (n_109, A[36], A[37]);
  nand g22 (n_110, A[38], A[39]);
  nand g23 (n_143, A[40], A[41]);
  nor g26 (n_111, n_93, n_94);
  nor g27 (n_114, n_95, n_96);
  nor g28 (n_115, n_97, n_98);
  nor g29 (n_116, n_99, n_100);
  nor g30 (n_117, n_101, n_102);
  nor g31 (n_118, n_103, n_104);
  nor g32 (n_119, n_105, n_106);
  nor g33 (n_120, n_107, n_108);
  nor g34 (n_121, n_109, n_110);
  nand g37 (n_122, n_114, n_115);
  nand g38 (n_125, n_116, n_117);
  nand g39 (n_126, n_118, n_119);
  nand g40 (n_130, n_120, n_121);
  nor g43 (n_127, n_125, n_126);
  nor g46 (n_134, n_125, n_128);
  nand g49 (n_136, n_114, n_123);
  nand g52 (n_140, n_118, n_134);
  nand g53 (n_142, n_120, n_131);
  nor g54 (n_146, n_93, n_112);
  nor g57 (n_150, n_97, n_136);
  nor g58 (n_152, n_99, n_128);
  nor g63 (n_158, n_105, n_140);
  nor g66 (n_162, n_109, n_142);
  nor g67 (n_164, n_143, n_144);
  nand g68 (n_166, A[2], n_91);
  nand g71 (n_170, A[6], n_146);
  nand g72 (n_172, A[8], n_123);
  nand g77 (n_178, A[14], n_150);
  nand g80 (n_182, A[18], n_152);
  nand g81 (n_184, A[20], n_137);
  nand g84 (n_188, A[24], n_134);
  nand g89 (n_194, A[30], n_158);
  nand g90 (n_196, A[32], n_131);
  nand g95 (n_202, A[38], n_162);
  xor g99 (Z[0], A[0], CI);
  xor g102 (Z[2], A[2], n_91);
  xor g107 (Z[5], A[5], n_169);
  xor g108 (Z[6], A[6], n_146);
  xor g111 (Z[8], A[8], n_123);
  xor g116 (Z[11], A[11], n_175);
  xor g119 (Z[13], A[13], n_177);
  xor g120 (Z[14], A[14], n_150);
  xor g125 (Z[17], A[17], n_181);
  xor g126 (Z[18], A[18], n_152);
  xor g129 (Z[20], A[20], n_137);
  xor g134 (Z[23], A[23], n_187);
  xor g135 (Z[24], A[24], n_134);
  xor g140 (Z[27], A[27], n_191);
  xor g143 (Z[29], A[29], n_193);
  xor g144 (Z[30], A[30], n_158);
  xor g147 (Z[32], A[32], n_131);
  xor g152 (Z[35], A[35], n_199);
  xor g155 (Z[37], A[37], n_201);
  xor g156 (Z[38], A[38], n_162);
  xor g161 (Z[41], A[41], n_205);
  xor g162 (Z[42], A[42], n_164);
  and g164 (n_91, A[1], wc);
  not gc (wc, n_88);
  or g165 (n_112, wc0, n_90);
  not gc0 (wc0, n_91);
  xnor g166 (Z[1], n_88, A[1]);
  and g167 (n_123, wc1, n_111);
  not gc1 (wc1, n_112);
  and g168 (n_169, A[4], wc2);
  not gc2 (wc2, n_112);
  or g169 (n_128, wc3, n_122);
  not gc3 (wc3, n_123);
  or g170 (n_147, wc4, n_95);
  not gc4 (wc4, n_123);
  xnor g171 (Z[3], n_166, A[3]);
  xnor g172 (Z[4], n_112, A[4]);
  and g173 (n_131, wc5, n_127);
  not gc5 (wc5, n_128);
  and g174 (n_137, wc6, n_116);
  not gc6 (wc6, n_128);
  and g175 (n_175, A[10], wc7);
  not gc7 (wc7, n_147);
  and g176 (n_177, A[12], wc8);
  not gc8 (wc8, n_136);
  and g177 (n_181, A[16], wc9);
  not gc9 (wc9, n_128);
  or g178 (n_144, wc10, n_130);
  not gc10 (wc10, n_131);
  or g179 (n_153, wc11, n_101);
  not gc11 (wc11, n_137);
  or g180 (n_155, wc12, n_103);
  not gc12 (wc12, n_134);
  or g181 (n_159, wc13, n_107);
  not gc13 (wc13, n_131);
  xnor g182 (Z[7], n_170, A[7]);
  xnor g183 (Z[9], n_172, A[9]);
  xnor g184 (Z[10], n_147, A[10]);
  xnor g185 (Z[12], n_136, A[12]);
  xnor g186 (Z[16], n_128, A[16]);
  and g187 (n_187, A[22], wc14);
  not gc14 (wc14, n_153);
  and g188 (n_191, A[26], wc15);
  not gc15 (wc15, n_155);
  and g189 (n_193, A[28], wc16);
  not gc16 (wc16, n_140);
  and g190 (n_199, A[34], wc17);
  not gc17 (wc17, n_159);
  and g191 (n_201, A[36], wc18);
  not gc18 (wc18, n_142);
  and g192 (n_205, A[40], wc19);
  not gc19 (wc19, n_144);
  xnor g193 (Z[15], n_178, A[15]);
  xnor g194 (Z[19], n_182, A[19]);
  xnor g195 (Z[21], n_184, A[21]);
  xnor g196 (Z[22], n_153, A[22]);
  xnor g197 (Z[25], n_188, A[25]);
  xnor g198 (Z[26], n_155, A[26]);
  xnor g199 (Z[28], n_140, A[28]);
  xnor g200 (Z[33], n_196, A[33]);
  xnor g201 (Z[34], n_159, A[34]);
  xnor g202 (Z[36], n_142, A[36]);
  xnor g203 (Z[40], n_144, A[40]);
  xnor g204 (Z[31], n_194, A[31]);
  xnor g205 (Z[39], n_202, A[39]);
endmodule

module increment_unsigned_9286_3_GENERIC(A, CI, Z);
  input [42:0] A;
  input CI;
  output [42:0] Z;
  wire [42:0] A;
  wire CI;
  wire [42:0] Z;
  increment_unsigned_9286_3_GENERIC_REAL g1(.A ({A[41], A[41:0]}), .CI
       (CI), .Z (Z));
endmodule

module mult_signed_const_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [42:0] A;
  output [61:0] Z;
  wire [42:0] A;
  wire [61:0] Z;
  wire n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54;
  wire n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62;
  wire n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78;
  wire n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241;
  wire n_242, n_243, n_244, n_245, n_246, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257;
  wire n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538;
  wire n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562;
  wire n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578;
  wire n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586;
  wire n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594;
  wire n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602;
  wire n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_611;
  wire n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619;
  wire n_620, n_621, n_622, n_623, n_625, n_626, n_627, n_628;
  wire n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636;
  wire n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646;
  wire n_647, n_648, n_649, n_650, n_651, n_652, n_656, n_657;
  wire n_658, n_659, n_660, n_662, n_663, n_664, n_665, n_666;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_677;
  wire n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_687;
  wire n_688, n_692, n_693, n_694, n_695, n_696, n_697, n_698;
  wire n_699, n_704, n_705, n_706, n_707, n_708, n_709, n_710;
  wire n_711, n_712, n_716, n_717, n_718, n_719, n_720, n_721;
  wire n_722, n_723, n_724, n_725, n_727, n_728, n_729, n_731;
  wire n_732, n_733, n_734, n_735, n_736, n_739, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_749, n_750, n_751;
  wire n_753, n_754, n_755, n_756, n_760, n_762, n_763, n_764;
  wire n_765, n_769, n_770, n_771, n_772, n_776, n_777, n_778;
  wire n_779, n_782, n_783, n_784, n_788, n_789, n_791, n_792;
  wire n_795, n_798, n_799, n_800, n_801, n_802, n_803, n_804;
  wire n_805, n_806, n_807, n_809, n_810, n_811, n_812, n_813;
  wire n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824;
  wire n_825, n_826, n_828, n_829, n_830, n_831, n_832, n_833;
  wire n_834, n_836, n_838, n_839, n_840, n_841, n_842, n_843;
  wire n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_854;
  wire n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_864;
  wire n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875;
  wire n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_886;
  wire n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894;
  wire n_895, n_896, n_897, n_898, n_899, n_900, n_902, n_903;
  wire n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_912;
  wire n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920;
  wire n_921, n_922, n_925, n_928, n_929, n_930, n_931, n_932;
  wire n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940;
  wire n_941, n_942, n_945, n_946, n_947, n_948, n_950, n_951;
  wire n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959;
  wire n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967;
  wire n_968, n_969, n_970, n_972, n_974, n_977, n_978, n_979;
  wire n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_997, n_998, n_1000, n_1001, n_1004, n_1005, n_1006, n_1007;
  wire n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015;
  wire n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023;
  wire n_1024, n_1025, n_1028, n_1030, n_1031, n_1034, n_1035, n_1036;
  wire n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044;
  wire n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052;
  wire n_1053, n_1054, n_1055, n_1056, n_1057, n_1062, n_1063, n_1064;
  wire n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073;
  wire n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081;
  wire n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089;
  wire n_1094, n_1095, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103;
  wire n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111;
  wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119;
  wire n_1120, n_1121, n_1124, n_1125, n_1126, n_1127, n_1128, n_1130;
  wire n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138;
  wire n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146;
  wire n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1156;
  wire n_1158, n_1159, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167;
  wire n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175;
  wire n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183;
  wire n_1184, n_1185, n_1188, n_1190, n_1191, n_1194, n_1195, n_1196;
  wire n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204;
  wire n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212;
  wire n_1213, n_1214, n_1215, n_1216, n_1217, n_1220, n_1222, n_1223;
  wire n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233;
  wire n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241;
  wire n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249;
  wire n_1252, n_1254, n_1255, n_1258, n_1259, n_1260, n_1261, n_1262;
  wire n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270;
  wire n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278;
  wire n_1279, n_1280, n_1281, n_1284, n_1286, n_1287, n_1290, n_1291;
  wire n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299;
  wire n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307;
  wire n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1316, n_1318;
  wire n_1319, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328;
  wire n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336;
  wire n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344;
  wire n_1345, n_1348, n_1350, n_1351, n_1354, n_1355, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1380, n_1382, n_1383, n_1386;
  wire n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394;
  wire n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402;
  wire n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1412;
  wire n_1414, n_1415, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423;
  wire n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431;
  wire n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439;
  wire n_1440, n_1441, n_1442, n_1443, n_1444, n_1446, n_1449, n_1450;
  wire n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458;
  wire n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466;
  wire n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474;
  wire n_1475, n_1476, n_1478, n_1481, n_1482, n_1483, n_1484, n_1485;
  wire n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493;
  wire n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501;
  wire n_1505, n_1506, n_1508, n_1512, n_1513, n_1514, n_1515, n_1516;
  wire n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524;
  wire n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532;
  wire n_1533, n_1534, n_1535, n_1537, n_1538, n_1540, n_1542, n_1545;
  wire n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553;
  wire n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561;
  wire n_1562, n_1563, n_1564, n_1565, n_1569, n_1574, n_1575, n_1576;
  wire n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584;
  wire n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592;
  wire n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1601;
  wire n_1602, n_1604, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613;
  wire n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621;
  wire n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629;
  wire n_1630, n_1634, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643;
  wire n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651;
  wire n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659;
  wire n_1660, n_1661, n_1665, n_1670, n_1671, n_1672, n_1674, n_1675;
  wire n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683;
  wire n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691;
  wire n_1692, n_1693, n_1694, n_1695, n_1697, n_1698, n_1702, n_1703;
  wire n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712;
  wire n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720;
  wire n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1730;
  wire n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741;
  wire n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749;
  wire n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757;
  wire n_1758, n_1759, n_1761, n_1762, n_1765, n_1766, n_1770, n_1771;
  wire n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779;
  wire n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787;
  wire n_1788, n_1789, n_1790, n_1792, n_1793, n_1802, n_1803, n_1804;
  wire n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812;
  wire n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820;
  wire n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
  wire n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841;
  wire n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849;
  wire n_1850, n_1851, n_1852, n_1853, n_1862, n_1863, n_1864, n_1865;
  wire n_1866, n_1867, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874;
  wire n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1886;
  wire n_1887, n_1889, n_1892, n_1893, n_1894, n_1895, n_1897, n_1898;
  wire n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906;
  wire n_1907, n_1908, n_1909, n_1912, n_1913, n_1914, n_1917, n_1918;
  wire n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927;
  wire n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1942, n_1944;
  wire n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952;
  wire n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1961, n_1962;
  wire n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972;
  wire n_1973, n_1974, n_1975, n_1976, n_1977, n_1980, n_1981, n_1986;
  wire n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994;
  wire n_1995, n_1996, n_1997, n_2004, n_2005, n_2006, n_2007, n_2008;
  wire n_2009, n_2010, n_2011, n_2012, n_2013, n_2021, n_2022, n_2023;
  wire n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2032, n_2034;
  wire n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2049;
  wire n_2050, n_2051, n_2052, n_2053, n_2054, n_2056, n_2057, n_2058;
  wire n_2059, n_2060, n_2061, n_2064, n_2065, n_2066, n_2067, n_2068;
  wire n_2069, n_2071, n_2072, n_2073, n_2076, n_2077, n_2089, n_2091;
  wire n_2093, n_2094, n_2095, n_2096, n_2097, n_2099, n_2100, n_2101;
  wire n_2102, n_2103, n_2105, n_2106, n_2107, n_2108, n_2109, n_2111;
  wire n_2112, n_2113, n_2114, n_2115, n_2117, n_2118, n_2119, n_2120;
  wire n_2121, n_2123, n_2124, n_2125, n_2126, n_2127, n_2129, n_2130;
  wire n_2131, n_2132, n_2133, n_2135, n_2136, n_2137, n_2138, n_2139;
  wire n_2141, n_2142, n_2143, n_2144, n_2145, n_2147, n_2148, n_2149;
  wire n_2150, n_2151, n_2153, n_2154, n_2155, n_2156, n_2157, n_2159;
  wire n_2160, n_2161, n_2162, n_2163, n_2165, n_2166, n_2167, n_2168;
  wire n_2169, n_2171, n_2172, n_2173, n_2174, n_2175, n_2177, n_2178;
  wire n_2179, n_2180, n_2181, n_2183, n_2184, n_2185, n_2186, n_2187;
  wire n_2189, n_2190, n_2191, n_2192, n_2193, n_2195, n_2196, n_2197;
  wire n_2198, n_2199, n_2201, n_2202, n_2203, n_2204, n_2205, n_2207;
  wire n_2208, n_2209, n_2210, n_2211, n_2213, n_2214, n_2215, n_2216;
  wire n_2217, n_2219, n_2220, n_2221, n_2222, n_2223, n_2225, n_2226;
  wire n_2227, n_2228, n_2229, n_2231, n_2232, n_2233, n_2234, n_2235;
  wire n_2237, n_2238, n_2239, n_2240, n_2241, n_2243, n_2244, n_2245;
  wire n_2246, n_2247, n_2249, n_2250, n_2251, n_2252, n_2253, n_2255;
  wire n_2256, n_2257, n_2258, n_2259, n_2261, n_2262, n_2265, n_2270;
  wire n_2272, n_2273, n_2275, n_2277, n_2279, n_2280, n_2282, n_2283;
  wire n_2285, n_2287, n_2289, n_2290, n_2292, n_2293, n_2295, n_2297;
  wire n_2299, n_2300, n_2302, n_2303, n_2305, n_2307, n_2309, n_2310;
  wire n_2312, n_2313, n_2315, n_2317, n_2319, n_2320, n_2322, n_2323;
  wire n_2325, n_2327, n_2329, n_2330, n_2332, n_2333, n_2335, n_2337;
  wire n_2339, n_2340, n_2342, n_2343, n_2345, n_2347, n_2349, n_2350;
  wire n_2352, n_2353, n_2355, n_2357, n_2359, n_2360, n_2362, n_2363;
  wire n_2365, n_2367, n_2369, n_2370, n_2372, n_2373, n_2375, n_2377;
  wire n_2379, n_2380, n_2382, n_2383, n_2385, n_2387, n_2389, n_2390;
  wire n_2392, n_2393, n_2395, n_2397, n_2399, n_2400, n_2402, n_2403;
  wire n_2405, n_2407, n_2409, n_2410, n_2414, n_2415, n_2416, n_2418;
  wire n_2419, n_2420, n_2422, n_2423, n_2424, n_2425, n_2427, n_2429;
  wire n_2431, n_2432, n_2433, n_2435, n_2436, n_2437, n_2439, n_2440;
  wire n_2442, n_2444, n_2446, n_2447, n_2448, n_2450, n_2451, n_2452;
  wire n_2454, n_2455, n_2457, n_2459, n_2461, n_2462, n_2463, n_2465;
  wire n_2466, n_2467, n_2469, n_2470, n_2472, n_2474, n_2476, n_2477;
  wire n_2478, n_2480, n_2481, n_2482, n_2484, n_2485, n_2487, n_2489;
  wire n_2491, n_2492, n_2493, n_2495, n_2496, n_2497, n_2499, n_2500;
  wire n_2502, n_2504, n_2506, n_2507, n_2508, n_2510, n_2511, n_2512;
  wire n_2514, n_2515, n_2517, n_2518, n_2520, n_2521, n_2522, n_2524;
  wire n_2525, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533;
  wire n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541;
  wire n_2543, n_2546, n_2548, n_2549, n_2550, n_2553, n_2556, n_2558;
  wire n_2559, n_2561, n_2563, n_2564, n_2566, n_2568, n_2569, n_2571;
  wire n_2573, n_2574, n_2576, n_2577, n_2579, n_2582, n_2584, n_2585;
  wire n_2586, n_2589, n_2592, n_2594, n_2595, n_2597, n_2599, n_2600;
  wire n_2602, n_2604, n_2605, n_2607, n_2609, n_2610, n_2612, n_2613;
  wire n_2615, n_2618, n_2620, n_2621, n_2622, n_2625, n_2628, n_2630;
  wire n_2631, n_2633, n_2635, n_2636, n_2637, n_2639, n_2640, n_2642;
  wire n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650;
  wire n_2651, n_2652, n_2653, n_2655, n_2656, n_2657, n_2659, n_2660;
  wire n_2661, n_2663, n_2664, n_2665, n_2667, n_2668, n_2669, n_2671;
  wire n_2672, n_2673, n_2675, n_2676, n_2677, n_2679, n_2680, n_2681;
  wire n_2683, n_2684, n_2685, n_2686, n_2688, n_2690, n_2692, n_2693;
  wire n_2694, n_2696, n_2698, n_2700, n_2701, n_2703, n_2705, n_2706;
  wire n_2708, n_2710, n_2711, n_2714, n_2716, n_2717, n_2718, n_2720;
  wire n_2721, n_2722, n_2724, n_2725, n_2726, n_2728, n_2729, n_2730;
  wire n_2732, n_2733, n_2734, n_2736, n_2738, n_2739, n_2740, n_2742;
  wire n_2743, n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751;
  wire n_2752, n_2753, n_2754, n_2755, n_2756, n_2758, n_2759, n_2760;
  wire n_2762, n_2763, n_2764, n_2766, n_2767, n_2768, n_2770, n_2771;
  wire n_2772, n_2774, n_2775, n_2776, n_2778, n_2779, n_2780, n_2782;
  wire n_2783, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791;
  wire n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799;
  wire n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807;
  wire n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815;
  wire n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823;
  wire n_2824, n_2826, n_2829, n_2830, n_2832, n_2833, n_2834, n_2835;
  wire n_2837, n_2838, n_2839, n_2841, n_2842, n_2843, n_2844, n_2846;
  wire n_2847, n_2849, n_2850, n_2852, n_2853, n_2854, n_2855, n_2857;
  wire n_2858, n_2859, n_2861, n_2862, n_2863, n_2864, n_2866, n_2867;
  wire n_2869, n_2870, n_2872, n_2873, n_2874, n_2875, n_2877, n_2878;
  wire n_2879, n_2880, n_2882, n_2883, n_2884, n_2885, n_2887, n_2888;
  wire n_2890, n_2891, n_2893, n_2894, n_2895, n_2896, n_2898, n_2899;
  wire n_2900, n_2902, n_2903, n_2904, n_2905, n_2907, n_2908, n_2910;
  wire n_2911, n_2913, n_2914, n_2915, n_2916, n_2918, n_2919, n_2920;
  wire n_2921, n_2923, n_2924, n_2925, n_2926, n_2928, n_2929, n_2931;
  wire n_2932, n_2934, n_2935, n_2936, n_2937, n_2939, n_2940, n_2942;
  wire n_2943, n_2945, n_2946, n_2947, n_2948, n_2950, n_2951, n_2953;
  wire n_2954, n_2956, n_2957, n_2958, n_2959, n_2961, n_2962, n_2963;
  wire n_2964, n_2966, n_2967, n_2968, n_2969, n_2971, n_2972, n_2974;
  wire n_2975, n_2977;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g340 (n_163, A[4], A[0]);
  and g2 (n_100, A[4], A[0]);
  xor g341 (n_798, A[5], A[3]);
  xor g342 (n_162, n_798, A[1]);
  nand g3 (n_799, A[5], A[3]);
  nand g343 (n_800, A[1], A[3]);
  nand g344 (n_801, A[5], A[1]);
  nand g345 (n_99, n_799, n_800, n_801);
  xor g346 (n_231, A[6], A[4]);
  and g347 (n_232, A[6], A[4]);
  xor g348 (n_802, A[0], A[2]);
  xor g349 (n_161, n_802, n_231);
  nand g350 (n_803, A[0], A[2]);
  nand g4 (n_804, n_231, A[2]);
  nand g5 (n_805, A[0], n_231);
  nand g351 (n_98, n_803, n_804, n_805);
  xor g352 (n_806, A[7], A[5]);
  xor g353 (n_233, n_806, A[1]);
  nand g354 (n_807, A[7], A[5]);
  nand g356 (n_809, A[7], A[1]);
  nand g6 (n_235, n_807, n_801, n_809);
  xor g357 (n_810, A[3], n_232);
  xor g358 (n_160, n_810, n_233);
  nand g359 (n_811, A[3], n_232);
  nand g360 (n_812, n_233, n_232);
  nand g361 (n_813, A[3], n_233);
  nand g362 (n_97, n_811, n_812, n_813);
  xor g363 (n_234, A[8], A[6]);
  and g364 (n_237, A[8], A[6]);
  xor g366 (n_236, n_802, A[4]);
  nand g369 (n_817, A[2], A[4]);
  xor g371 (n_818, n_234, n_235);
  xor g372 (n_159, n_818, n_236);
  nand g373 (n_819, n_234, n_235);
  nand g374 (n_820, n_236, n_235);
  nand g375 (n_821, n_234, n_236);
  nand g376 (n_96, n_819, n_820, n_821);
  xor g377 (n_822, A[9], A[7]);
  xor g378 (n_239, n_822, A[3]);
  nand g379 (n_823, A[9], A[7]);
  nand g380 (n_824, A[3], A[7]);
  nand g381 (n_825, A[9], A[3]);
  nand g382 (n_242, n_823, n_824, n_825);
  xor g383 (n_826, A[1], A[5]);
  xor g384 (n_240, n_826, n_237);
  nand g386 (n_828, n_237, A[5]);
  nand g387 (n_829, A[1], n_237);
  nand g388 (n_244, n_801, n_828, n_829);
  xor g389 (n_830, n_238, n_239);
  xor g390 (n_158, n_830, n_240);
  nand g391 (n_831, n_238, n_239);
  nand g392 (n_832, n_240, n_239);
  nand g393 (n_833, n_238, n_240);
  nand g394 (n_95, n_831, n_832, n_833);
  xor g395 (n_241, A[10], A[8]);
  and g396 (n_246, A[10], A[8]);
  xor g397 (n_834, A[4], A[2]);
  xor g398 (n_243, n_834, A[6]);
  nand g400 (n_836, A[6], A[2]);
  xor g403 (n_838, A[0], n_241);
  xor g404 (n_245, n_838, n_242);
  nand g405 (n_839, A[0], n_241);
  nand g406 (n_840, n_242, n_241);
  nand g407 (n_841, A[0], n_242);
  nand g408 (n_250, n_839, n_840, n_841);
  xor g409 (n_842, n_243, n_244);
  xor g410 (n_157, n_842, n_245);
  nand g411 (n_843, n_243, n_244);
  nand g412 (n_844, n_245, n_244);
  nand g413 (n_845, n_243, n_245);
  nand g414 (n_94, n_843, n_844, n_845);
  xor g415 (n_846, A[11], A[9]);
  xor g416 (n_248, n_846, A[5]);
  nand g417 (n_847, A[11], A[9]);
  nand g418 (n_848, A[5], A[9]);
  nand g419 (n_849, A[11], A[5]);
  nand g420 (n_253, n_847, n_848, n_849);
  xor g421 (n_850, A[3], A[7]);
  xor g422 (n_249, n_850, A[1]);
  nand g426 (n_254, n_824, n_809, n_800);
  xor g427 (n_854, n_246, n_247);
  xor g428 (n_251, n_854, n_248);
  nand g429 (n_855, n_246, n_247);
  nand g430 (n_856, n_248, n_247);
  nand g431 (n_857, n_246, n_248);
  nand g432 (n_258, n_855, n_856, n_857);
  xor g433 (n_858, n_249, n_250);
  xor g434 (n_156, n_858, n_251);
  nand g435 (n_859, n_249, n_250);
  nand g436 (n_860, n_251, n_250);
  nand g437 (n_861, n_249, n_251);
  nand g438 (n_93, n_859, n_860, n_861);
  xor g439 (n_252, A[12], A[10]);
  and g440 (n_259, A[12], A[10]);
  xor g442 (n_255, n_231, A[8]);
  nand g444 (n_864, A[8], A[4]);
  xor g448 (n_256, n_802, n_252);
  nand g450 (n_868, n_252, A[0]);
  nand g451 (n_869, A[2], n_252);
  nand g452 (n_263, n_803, n_868, n_869);
  xor g453 (n_870, n_253, n_254);
  xor g454 (n_257, n_870, n_255);
  nand g455 (n_871, n_253, n_254);
  nand g456 (n_872, n_255, n_254);
  nand g457 (n_873, n_253, n_255);
  nand g458 (n_265, n_871, n_872, n_873);
  xor g459 (n_874, n_256, n_257);
  xor g460 (n_155, n_874, n_258);
  nand g461 (n_875, n_256, n_257);
  nand g462 (n_876, n_258, n_257);
  nand g463 (n_877, n_256, n_258);
  nand g464 (n_92, n_875, n_876, n_877);
  xor g465 (n_878, A[13], A[11]);
  xor g466 (n_262, n_878, A[7]);
  nand g467 (n_879, A[13], A[11]);
  nand g468 (n_880, A[7], A[11]);
  nand g469 (n_881, A[13], A[7]);
  nand g470 (n_268, n_879, n_880, n_881);
  xor g471 (n_882, A[5], A[9]);
  xor g472 (n_261, n_882, A[3]);
  nand g476 (n_269, n_848, n_825, n_799);
  xor g477 (n_886, A[1], n_259);
  xor g478 (n_264, n_886, n_260);
  nand g479 (n_887, A[1], n_259);
  nand g480 (n_888, n_260, n_259);
  nand g481 (n_889, A[1], n_260);
  nand g482 (n_272, n_887, n_888, n_889);
  xor g483 (n_890, n_261, n_262);
  xor g484 (n_266, n_890, n_263);
  nand g485 (n_891, n_261, n_262);
  nand g486 (n_892, n_263, n_262);
  nand g487 (n_893, n_261, n_263);
  nand g488 (n_274, n_891, n_892, n_893);
  xor g489 (n_894, n_264, n_265);
  xor g490 (n_154, n_894, n_266);
  nand g491 (n_895, n_264, n_265);
  nand g492 (n_896, n_266, n_265);
  nand g493 (n_897, n_264, n_266);
  nand g494 (n_91, n_895, n_896, n_897);
  xor g495 (n_267, A[14], A[12]);
  and g496 (n_276, A[14], A[12]);
  xor g497 (n_898, A[8], A[0]);
  xor g498 (n_271, n_898, A[6]);
  nand g499 (n_899, A[8], A[0]);
  nand g500 (n_900, A[6], A[0]);
  xor g503 (n_902, A[10], A[4]);
  xor g504 (n_270, n_902, A[2]);
  nand g505 (n_903, A[10], A[4]);
  nand g507 (n_905, A[10], A[2]);
  nand g508 (n_278, n_903, n_817, n_905);
  xor g509 (n_906, n_267, n_268);
  xor g510 (n_273, n_906, n_269);
  nand g511 (n_907, n_267, n_268);
  nand g512 (n_908, n_269, n_268);
  nand g513 (n_909, n_267, n_269);
  nand g514 (n_282, n_907, n_908, n_909);
  xor g515 (n_910, n_270, n_271);
  xor g516 (n_275, n_910, n_272);
  nand g517 (n_911, n_270, n_271);
  nand g518 (n_912, n_272, n_271);
  nand g519 (n_913, n_270, n_272);
  nand g520 (n_285, n_911, n_912, n_913);
  xor g521 (n_914, n_273, n_274);
  xor g522 (n_153, n_914, n_275);
  nand g523 (n_915, n_273, n_274);
  nand g524 (n_916, n_275, n_274);
  nand g525 (n_917, n_273, n_275);
  nand g526 (n_90, n_915, n_916, n_917);
  xor g527 (n_918, A[15], A[13]);
  xor g528 (n_279, n_918, A[9]);
  nand g529 (n_919, A[15], A[13]);
  nand g530 (n_920, A[9], A[13]);
  nand g531 (n_921, A[15], A[9]);
  nand g532 (n_287, n_919, n_920, n_921);
  xor g533 (n_922, A[1], A[7]);
  xor g534 (n_280, n_922, A[11]);
  nand g537 (n_925, A[1], A[11]);
  nand g538 (n_288, n_809, n_880, n_925);
  xor g540 (n_281, n_798, n_276);
  nand g542 (n_928, n_276, A[3]);
  nand g543 (n_929, A[5], n_276);
  nand g544 (n_291, n_799, n_928, n_929);
  xor g545 (n_930, n_277, n_278);
  xor g546 (n_283, n_930, n_279);
  nand g547 (n_931, n_277, n_278);
  nand g548 (n_932, n_279, n_278);
  nand g549 (n_933, n_277, n_279);
  nand g550 (n_293, n_931, n_932, n_933);
  xor g551 (n_934, n_280, n_281);
  xor g552 (n_284, n_934, n_282);
  nand g553 (n_935, n_280, n_281);
  nand g554 (n_936, n_282, n_281);
  nand g555 (n_937, n_280, n_282);
  nand g556 (n_295, n_935, n_936, n_937);
  xor g557 (n_938, n_283, n_284);
  xor g558 (n_152, n_938, n_285);
  nand g559 (n_939, n_283, n_284);
  nand g560 (n_940, n_285, n_284);
  nand g561 (n_941, n_283, n_285);
  nand g562 (n_89, n_939, n_940, n_941);
  xor g563 (n_286, A[16], A[14]);
  and g564 (n_297, A[16], A[14]);
  xor g565 (n_942, A[10], A[2]);
  xor g566 (n_290, n_942, A[0]);
  nand g569 (n_945, A[10], A[0]);
  nand g570 (n_298, n_905, n_803, n_945);
  xor g571 (n_946, A[8], A[12]);
  xor g572 (n_289, n_946, A[6]);
  nand g573 (n_947, A[8], A[12]);
  nand g574 (n_948, A[6], A[12]);
  xor g577 (n_950, A[4], n_286);
  xor g578 (n_292, n_950, n_287);
  nand g579 (n_951, A[4], n_286);
  nand g580 (n_952, n_287, n_286);
  nand g581 (n_953, A[4], n_287);
  nand g582 (n_303, n_951, n_952, n_953);
  xor g583 (n_954, n_288, n_289);
  xor g584 (n_294, n_954, n_290);
  nand g585 (n_955, n_288, n_289);
  nand g586 (n_956, n_290, n_289);
  nand g587 (n_957, n_288, n_290);
  nand g588 (n_305, n_955, n_956, n_957);
  xor g589 (n_958, n_291, n_292);
  xor g590 (n_296, n_958, n_293);
  nand g591 (n_959, n_291, n_292);
  nand g592 (n_960, n_293, n_292);
  nand g593 (n_961, n_291, n_293);
  nand g594 (n_307, n_959, n_960, n_961);
  xor g595 (n_962, n_294, n_295);
  xor g596 (n_151, n_962, n_296);
  nand g597 (n_963, n_294, n_295);
  nand g598 (n_964, n_296, n_295);
  nand g599 (n_965, n_294, n_296);
  nand g600 (n_88, n_963, n_964, n_965);
  xor g601 (n_966, A[17], A[15]);
  xor g602 (n_301, n_966, A[11]);
  nand g603 (n_967, A[17], A[15]);
  nand g604 (n_968, A[11], A[15]);
  nand g605 (n_969, A[17], A[11]);
  nand g606 (n_310, n_967, n_968, n_969);
  xor g607 (n_970, A[3], A[1]);
  xor g608 (n_302, n_970, A[9]);
  nand g610 (n_972, A[9], A[1]);
  nand g612 (n_102, n_800, n_972, n_825);
  xor g613 (n_974, A[13], A[7]);
  xor g614 (n_300, n_974, A[5]);
  nand g617 (n_977, A[13], A[5]);
  nand g618 (n_101, n_881, n_807, n_977);
  xor g619 (n_978, n_297, n_298);
  xor g620 (n_304, n_978, n_299);
  nand g621 (n_979, n_297, n_298);
  nand g622 (n_980, n_299, n_298);
  nand g623 (n_981, n_297, n_299);
  nand g624 (n_311, n_979, n_980, n_981);
  xor g625 (n_982, n_300, n_301);
  xor g626 (n_306, n_982, n_302);
  nand g627 (n_983, n_300, n_301);
  nand g628 (n_984, n_302, n_301);
  nand g629 (n_985, n_300, n_302);
  nand g630 (n_313, n_983, n_984, n_985);
  xor g631 (n_986, n_303, n_304);
  xor g632 (n_308, n_986, n_305);
  nand g633 (n_987, n_303, n_304);
  nand g634 (n_988, n_305, n_304);
  nand g635 (n_989, n_303, n_305);
  nand g636 (n_315, n_987, n_988, n_989);
  xor g637 (n_990, n_306, n_307);
  xor g638 (n_150, n_990, n_308);
  nand g639 (n_991, n_306, n_307);
  nand g640 (n_992, n_308, n_307);
  nand g641 (n_993, n_306, n_308);
  nand g642 (n_87, n_991, n_992, n_993);
  xor g643 (n_309, A[18], A[16]);
  and g644 (n_317, A[18], A[16]);
  xor g645 (n_994, A[12], A[4]);
  xor g646 (n_103, n_994, A[2]);
  nand g647 (n_995, A[12], A[4]);
  nand g649 (n_997, A[12], A[2]);
  nand g650 (n_318, n_995, n_817, n_997);
  xor g651 (n_998, A[10], A[0]);
  xor g652 (n_104, n_998, A[14]);
  nand g654 (n_1000, A[14], A[0]);
  nand g655 (n_1001, A[10], A[14]);
  nand g656 (n_319, n_945, n_1000, n_1001);
  xor g658 (n_105, n_234, n_309);
  nand g660 (n_1004, n_309, A[6]);
  nand g661 (n_1005, A[8], n_309);
  xor g663 (n_1006, n_310, n_101);
  xor g664 (n_312, n_1006, n_102);
  nand g665 (n_1007, n_310, n_101);
  nand g666 (n_1008, n_102, n_101);
  nand g667 (n_1009, n_310, n_102);
  nand g668 (n_325, n_1007, n_1008, n_1009);
  xor g669 (n_1010, n_103, n_104);
  xor g670 (n_314, n_1010, n_105);
  nand g671 (n_1011, n_103, n_104);
  nand g672 (n_1012, n_105, n_104);
  nand g673 (n_1013, n_103, n_105);
  nand g674 (n_326, n_1011, n_1012, n_1013);
  xor g675 (n_1014, n_311, n_312);
  xor g676 (n_316, n_1014, n_313);
  nand g677 (n_1015, n_311, n_312);
  nand g678 (n_1016, n_313, n_312);
  nand g679 (n_1017, n_311, n_313);
  nand g680 (n_329, n_1015, n_1016, n_1017);
  xor g681 (n_1018, n_314, n_315);
  xor g682 (n_149, n_1018, n_316);
  nand g683 (n_1019, n_314, n_315);
  nand g684 (n_1020, n_316, n_315);
  nand g685 (n_1021, n_314, n_316);
  nand g686 (n_86, n_1019, n_1020, n_1021);
  xor g687 (n_1022, A[19], A[17]);
  xor g688 (n_321, n_1022, A[13]);
  nand g689 (n_1023, A[19], A[17]);
  nand g690 (n_1024, A[13], A[17]);
  nand g691 (n_1025, A[19], A[13]);
  nand g692 (n_331, n_1023, n_1024, n_1025);
  xor g694 (n_322, n_798, A[11]);
  nand g696 (n_1028, A[11], A[3]);
  nand g698 (n_332, n_799, n_1028, n_849);
  xor g699 (n_1030, A[1], A[15]);
  xor g700 (n_320, n_1030, A[9]);
  nand g701 (n_1031, A[1], A[15]);
  nand g704 (n_333, n_1031, n_921, n_972);
  xor g705 (n_1034, A[7], n_317);
  xor g706 (n_324, n_1034, n_318);
  nand g707 (n_1035, A[7], n_317);
  nand g708 (n_1036, n_318, n_317);
  nand g709 (n_1037, A[7], n_318);
  nand g710 (n_337, n_1035, n_1036, n_1037);
  xor g711 (n_1038, n_319, n_320);
  xor g712 (n_327, n_1038, n_321);
  nand g713 (n_1039, n_319, n_320);
  nand g714 (n_1040, n_321, n_320);
  nand g715 (n_1041, n_319, n_321);
  nand g716 (n_339, n_1039, n_1040, n_1041);
  xor g717 (n_1042, n_322, n_323);
  xor g718 (n_328, n_1042, n_324);
  nand g719 (n_1043, n_322, n_323);
  nand g720 (n_1044, n_324, n_323);
  nand g721 (n_1045, n_322, n_324);
  nand g722 (n_341, n_1043, n_1044, n_1045);
  xor g723 (n_1046, n_325, n_326);
  xor g724 (n_330, n_1046, n_327);
  nand g725 (n_1047, n_325, n_326);
  nand g726 (n_1048, n_327, n_326);
  nand g727 (n_1049, n_325, n_327);
  nand g728 (n_343, n_1047, n_1048, n_1049);
  xor g729 (n_1050, n_328, n_329);
  xor g730 (n_148, n_1050, n_330);
  nand g731 (n_1051, n_328, n_329);
  nand g732 (n_1052, n_330, n_329);
  nand g733 (n_1053, n_328, n_330);
  nand g734 (n_85, n_1051, n_1052, n_1053);
  xor g735 (n_1054, A[20], A[18]);
  xor g736 (n_335, n_1054, A[14]);
  nand g737 (n_1055, A[20], A[18]);
  nand g738 (n_1056, A[14], A[18]);
  nand g739 (n_1057, A[20], A[14]);
  nand g740 (n_345, n_1055, n_1056, n_1057);
  xor g742 (n_336, n_231, A[12]);
  xor g747 (n_1062, A[2], A[16]);
  xor g748 (n_334, n_1062, A[10]);
  nand g749 (n_1063, A[2], A[16]);
  nand g750 (n_1064, A[10], A[16]);
  nand g752 (n_347, n_1063, n_1064, n_905);
  xor g753 (n_1066, A[8], n_331);
  xor g754 (n_338, n_1066, n_332);
  nand g755 (n_1067, A[8], n_331);
  nand g756 (n_1068, n_332, n_331);
  nand g757 (n_1069, A[8], n_332);
  nand g758 (n_351, n_1067, n_1068, n_1069);
  xor g759 (n_1070, n_333, n_334);
  xor g760 (n_340, n_1070, n_335);
  nand g761 (n_1071, n_333, n_334);
  nand g762 (n_1072, n_335, n_334);
  nand g763 (n_1073, n_333, n_335);
  nand g764 (n_353, n_1071, n_1072, n_1073);
  xor g765 (n_1074, n_336, n_337);
  xor g766 (n_342, n_1074, n_338);
  nand g767 (n_1075, n_336, n_337);
  nand g768 (n_1076, n_338, n_337);
  nand g769 (n_1077, n_336, n_338);
  nand g770 (n_355, n_1075, n_1076, n_1077);
  xor g771 (n_1078, n_339, n_340);
  xor g772 (n_344, n_1078, n_341);
  nand g773 (n_1079, n_339, n_340);
  nand g774 (n_1080, n_341, n_340);
  nand g775 (n_1081, n_339, n_341);
  nand g776 (n_357, n_1079, n_1080, n_1081);
  xor g777 (n_1082, n_342, n_343);
  xor g778 (n_147, n_1082, n_344);
  nand g779 (n_1083, n_342, n_343);
  nand g780 (n_1084, n_344, n_343);
  nand g781 (n_1085, n_342, n_344);
  nand g782 (n_84, n_1083, n_1084, n_1085);
  xor g783 (n_1086, A[21], A[19]);
  xor g784 (n_349, n_1086, A[15]);
  nand g785 (n_1087, A[21], A[19]);
  nand g786 (n_1088, A[15], A[19]);
  nand g787 (n_1089, A[21], A[15]);
  nand g788 (n_359, n_1087, n_1088, n_1089);
  xor g790 (n_350, n_806, A[13]);
  xor g795 (n_1094, A[3], A[17]);
  xor g796 (n_348, n_1094, A[11]);
  nand g797 (n_1095, A[3], A[17]);
  nand g800 (n_361, n_1095, n_969, n_1028);
  xor g801 (n_1098, A[9], n_345);
  xor g802 (n_352, n_1098, n_346);
  nand g803 (n_1099, A[9], n_345);
  nand g804 (n_1100, n_346, n_345);
  nand g805 (n_1101, A[9], n_346);
  nand g806 (n_164, n_1099, n_1100, n_1101);
  xor g807 (n_1102, n_347, n_348);
  xor g808 (n_354, n_1102, n_349);
  nand g809 (n_1103, n_347, n_348);
  nand g810 (n_1104, n_349, n_348);
  nand g811 (n_1105, n_347, n_349);
  nand g812 (n_365, n_1103, n_1104, n_1105);
  xor g813 (n_1106, n_350, n_351);
  xor g814 (n_356, n_1106, n_352);
  nand g815 (n_1107, n_350, n_351);
  nand g816 (n_1108, n_352, n_351);
  nand g817 (n_1109, n_350, n_352);
  nand g818 (n_367, n_1107, n_1108, n_1109);
  xor g819 (n_1110, n_353, n_354);
  xor g820 (n_358, n_1110, n_355);
  nand g821 (n_1111, n_353, n_354);
  nand g822 (n_1112, n_355, n_354);
  nand g823 (n_1113, n_353, n_355);
  nand g824 (n_370, n_1111, n_1112, n_1113);
  xor g825 (n_1114, n_356, n_357);
  xor g826 (n_146, n_1114, n_358);
  nand g827 (n_1115, n_356, n_357);
  nand g828 (n_1116, n_358, n_357);
  nand g829 (n_1117, n_356, n_358);
  nand g830 (n_83, n_1115, n_1116, n_1117);
  xor g831 (n_1118, A[22], A[20]);
  xor g832 (n_363, n_1118, A[16]);
  nand g833 (n_1119, A[22], A[20]);
  nand g834 (n_1120, A[16], A[20]);
  nand g835 (n_1121, A[22], A[16]);
  nand g836 (n_371, n_1119, n_1120, n_1121);
  xor g838 (n_364, n_234, A[14]);
  nand g840 (n_1124, A[14], A[6]);
  nand g841 (n_1125, A[8], A[14]);
  xor g843 (n_1126, A[4], A[18]);
  xor g844 (n_362, n_1126, A[12]);
  nand g845 (n_1127, A[4], A[18]);
  nand g846 (n_1128, A[12], A[18]);
  nand g848 (n_373, n_1127, n_1128, n_995);
  xor g849 (n_1130, A[10], n_359);
  xor g850 (n_165, n_1130, n_101);
  nand g851 (n_1131, A[10], n_359);
  nand g852 (n_1132, n_101, n_359);
  nand g853 (n_1133, A[10], n_101);
  nand g854 (n_377, n_1131, n_1132, n_1133);
  xor g855 (n_1134, n_361, n_362);
  xor g856 (n_366, n_1134, n_363);
  nand g857 (n_1135, n_361, n_362);
  nand g858 (n_1136, n_363, n_362);
  nand g859 (n_1137, n_361, n_363);
  nand g860 (n_379, n_1135, n_1136, n_1137);
  xor g861 (n_1138, n_364, n_164);
  xor g862 (n_368, n_1138, n_165);
  nand g863 (n_1139, n_364, n_164);
  nand g864 (n_1140, n_165, n_164);
  nand g865 (n_1141, n_364, n_165);
  nand g866 (n_381, n_1139, n_1140, n_1141);
  xor g867 (n_1142, n_365, n_366);
  xor g868 (n_369, n_1142, n_367);
  nand g869 (n_1143, n_365, n_366);
  nand g870 (n_1144, n_367, n_366);
  nand g871 (n_1145, n_365, n_367);
  nand g872 (n_384, n_1143, n_1144, n_1145);
  xor g873 (n_1146, n_368, n_369);
  xor g874 (n_145, n_1146, n_370);
  nand g875 (n_1147, n_368, n_369);
  nand g876 (n_1148, n_370, n_369);
  nand g877 (n_1149, n_368, n_370);
  nand g878 (n_82, n_1147, n_1148, n_1149);
  xor g879 (n_1150, A[23], A[21]);
  xor g880 (n_375, n_1150, A[17]);
  nand g881 (n_1151, A[23], A[21]);
  nand g882 (n_1152, A[17], A[21]);
  nand g883 (n_1153, A[23], A[17]);
  nand g884 (n_385, n_1151, n_1152, n_1153);
  xor g886 (n_376, n_822, A[15]);
  nand g888 (n_1156, A[15], A[7]);
  nand g890 (n_386, n_823, n_1156, n_921);
  xor g891 (n_1158, A[5], A[19]);
  xor g892 (n_374, n_1158, A[13]);
  nand g893 (n_1159, A[5], A[19]);
  nand g896 (n_387, n_1159, n_1025, n_977);
  xor g897 (n_1162, A[11], n_371);
  xor g898 (n_378, n_1162, n_372);
  nand g899 (n_1163, A[11], n_371);
  nand g900 (n_1164, n_372, n_371);
  nand g901 (n_1165, A[11], n_372);
  nand g902 (n_391, n_1163, n_1164, n_1165);
  xor g903 (n_1166, n_373, n_374);
  xor g904 (n_380, n_1166, n_375);
  nand g905 (n_1167, n_373, n_374);
  nand g906 (n_1168, n_375, n_374);
  nand g907 (n_1169, n_373, n_375);
  nand g908 (n_393, n_1167, n_1168, n_1169);
  xor g909 (n_1170, n_376, n_377);
  xor g910 (n_382, n_1170, n_378);
  nand g911 (n_1171, n_376, n_377);
  nand g912 (n_1172, n_378, n_377);
  nand g913 (n_1173, n_376, n_378);
  nand g914 (n_395, n_1171, n_1172, n_1173);
  xor g915 (n_1174, n_379, n_380);
  xor g916 (n_383, n_1174, n_381);
  nand g917 (n_1175, n_379, n_380);
  nand g918 (n_1176, n_381, n_380);
  nand g919 (n_1177, n_379, n_381);
  nand g920 (n_398, n_1175, n_1176, n_1177);
  xor g921 (n_1178, n_382, n_383);
  xor g922 (n_144, n_1178, n_384);
  nand g923 (n_1179, n_382, n_383);
  nand g924 (n_1180, n_384, n_383);
  nand g925 (n_1181, n_382, n_384);
  nand g926 (n_81, n_1179, n_1180, n_1181);
  xor g927 (n_1182, A[24], A[22]);
  xor g928 (n_389, n_1182, A[18]);
  nand g929 (n_1183, A[24], A[22]);
  nand g930 (n_1184, A[18], A[22]);
  nand g931 (n_1185, A[24], A[18]);
  nand g932 (n_399, n_1183, n_1184, n_1185);
  xor g934 (n_390, n_241, A[16]);
  nand g936 (n_1188, A[16], A[8]);
  xor g939 (n_1190, A[6], A[20]);
  xor g940 (n_388, n_1190, A[14]);
  nand g941 (n_1191, A[6], A[20]);
  nand g944 (n_401, n_1191, n_1057, n_1124);
  xor g945 (n_1194, A[12], n_385);
  xor g946 (n_392, n_1194, n_386);
  nand g947 (n_1195, A[12], n_385);
  nand g948 (n_1196, n_386, n_385);
  nand g949 (n_1197, A[12], n_386);
  nand g950 (n_405, n_1195, n_1196, n_1197);
  xor g951 (n_1198, n_387, n_388);
  xor g952 (n_394, n_1198, n_389);
  nand g953 (n_1199, n_387, n_388);
  nand g954 (n_1200, n_389, n_388);
  nand g955 (n_1201, n_387, n_389);
  nand g956 (n_407, n_1199, n_1200, n_1201);
  xor g957 (n_1202, n_390, n_391);
  xor g958 (n_396, n_1202, n_392);
  nand g959 (n_1203, n_390, n_391);
  nand g960 (n_1204, n_392, n_391);
  nand g961 (n_1205, n_390, n_392);
  nand g962 (n_409, n_1203, n_1204, n_1205);
  xor g963 (n_1206, n_393, n_394);
  xor g964 (n_397, n_1206, n_395);
  nand g965 (n_1207, n_393, n_394);
  nand g966 (n_1208, n_395, n_394);
  nand g967 (n_1209, n_393, n_395);
  nand g968 (n_412, n_1207, n_1208, n_1209);
  xor g969 (n_1210, n_396, n_397);
  xor g970 (n_143, n_1210, n_398);
  nand g971 (n_1211, n_396, n_397);
  nand g972 (n_1212, n_398, n_397);
  nand g973 (n_1213, n_396, n_398);
  nand g974 (n_80, n_1211, n_1212, n_1213);
  xor g975 (n_1214, A[25], A[23]);
  xor g976 (n_403, n_1214, A[19]);
  nand g977 (n_1215, A[25], A[23]);
  nand g978 (n_1216, A[19], A[23]);
  nand g979 (n_1217, A[25], A[19]);
  nand g980 (n_413, n_1215, n_1216, n_1217);
  xor g982 (n_404, n_846, A[17]);
  nand g984 (n_1220, A[17], A[9]);
  nand g986 (n_414, n_847, n_1220, n_969);
  xor g987 (n_1222, A[7], A[21]);
  xor g988 (n_402, n_1222, A[15]);
  nand g989 (n_1223, A[7], A[21]);
  nand g992 (n_415, n_1223, n_1089, n_1156);
  xor g993 (n_1226, A[13], n_399);
  xor g994 (n_406, n_1226, n_400);
  nand g995 (n_1227, A[13], n_399);
  nand g996 (n_1228, n_400, n_399);
  nand g997 (n_1229, A[13], n_400);
  nand g998 (n_419, n_1227, n_1228, n_1229);
  xor g999 (n_1230, n_401, n_402);
  xor g1000 (n_408, n_1230, n_403);
  nand g1001 (n_1231, n_401, n_402);
  nand g1002 (n_1232, n_403, n_402);
  nand g1003 (n_1233, n_401, n_403);
  nand g1004 (n_421, n_1231, n_1232, n_1233);
  xor g1005 (n_1234, n_404, n_405);
  xor g1006 (n_410, n_1234, n_406);
  nand g1007 (n_1235, n_404, n_405);
  nand g1008 (n_1236, n_406, n_405);
  nand g1009 (n_1237, n_404, n_406);
  nand g1010 (n_423, n_1235, n_1236, n_1237);
  xor g1011 (n_1238, n_407, n_408);
  xor g1012 (n_411, n_1238, n_409);
  nand g1013 (n_1239, n_407, n_408);
  nand g1014 (n_1240, n_409, n_408);
  nand g1015 (n_1241, n_407, n_409);
  nand g1016 (n_426, n_1239, n_1240, n_1241);
  xor g1017 (n_1242, n_410, n_411);
  xor g1018 (n_142, n_1242, n_412);
  nand g1019 (n_1243, n_410, n_411);
  nand g1020 (n_1244, n_412, n_411);
  nand g1021 (n_1245, n_410, n_412);
  nand g1022 (n_79, n_1243, n_1244, n_1245);
  xor g1023 (n_1246, A[26], A[24]);
  xor g1024 (n_417, n_1246, A[20]);
  nand g1025 (n_1247, A[26], A[24]);
  nand g1026 (n_1248, A[20], A[24]);
  nand g1027 (n_1249, A[26], A[20]);
  nand g1028 (n_427, n_1247, n_1248, n_1249);
  xor g1030 (n_418, n_252, A[18]);
  nand g1032 (n_1252, A[18], A[10]);
  xor g1035 (n_1254, A[8], A[22]);
  xor g1036 (n_416, n_1254, A[16]);
  nand g1037 (n_1255, A[8], A[22]);
  nand g1040 (n_429, n_1255, n_1121, n_1188);
  xor g1041 (n_1258, A[14], n_413);
  xor g1042 (n_420, n_1258, n_414);
  nand g1043 (n_1259, A[14], n_413);
  nand g1044 (n_1260, n_414, n_413);
  nand g1045 (n_1261, A[14], n_414);
  nand g1046 (n_433, n_1259, n_1260, n_1261);
  xor g1047 (n_1262, n_415, n_416);
  xor g1048 (n_422, n_1262, n_417);
  nand g1049 (n_1263, n_415, n_416);
  nand g1050 (n_1264, n_417, n_416);
  nand g1051 (n_1265, n_415, n_417);
  nand g1052 (n_435, n_1263, n_1264, n_1265);
  xor g1053 (n_1266, n_418, n_419);
  xor g1054 (n_424, n_1266, n_420);
  nand g1055 (n_1267, n_418, n_419);
  nand g1056 (n_1268, n_420, n_419);
  nand g1057 (n_1269, n_418, n_420);
  nand g1058 (n_437, n_1267, n_1268, n_1269);
  xor g1059 (n_1270, n_421, n_422);
  xor g1060 (n_425, n_1270, n_423);
  nand g1061 (n_1271, n_421, n_422);
  nand g1062 (n_1272, n_423, n_422);
  nand g1063 (n_1273, n_421, n_423);
  nand g1064 (n_440, n_1271, n_1272, n_1273);
  xor g1065 (n_1274, n_424, n_425);
  xor g1066 (n_141, n_1274, n_426);
  nand g1067 (n_1275, n_424, n_425);
  nand g1068 (n_1276, n_426, n_425);
  nand g1069 (n_1277, n_424, n_426);
  nand g1070 (n_78, n_1275, n_1276, n_1277);
  xor g1071 (n_1278, A[27], A[25]);
  xor g1072 (n_431, n_1278, A[21]);
  nand g1073 (n_1279, A[27], A[25]);
  nand g1074 (n_1280, A[21], A[25]);
  nand g1075 (n_1281, A[27], A[21]);
  nand g1076 (n_441, n_1279, n_1280, n_1281);
  xor g1078 (n_432, n_878, A[19]);
  nand g1080 (n_1284, A[19], A[11]);
  nand g1082 (n_442, n_879, n_1284, n_1025);
  xor g1083 (n_1286, A[9], A[23]);
  xor g1084 (n_430, n_1286, A[17]);
  nand g1085 (n_1287, A[9], A[23]);
  nand g1088 (n_443, n_1287, n_1153, n_1220);
  xor g1089 (n_1290, A[15], n_427);
  xor g1090 (n_434, n_1290, n_428);
  nand g1091 (n_1291, A[15], n_427);
  nand g1092 (n_1292, n_428, n_427);
  nand g1093 (n_1293, A[15], n_428);
  nand g1094 (n_447, n_1291, n_1292, n_1293);
  xor g1095 (n_1294, n_429, n_430);
  xor g1096 (n_436, n_1294, n_431);
  nand g1097 (n_1295, n_429, n_430);
  nand g1098 (n_1296, n_431, n_430);
  nand g1099 (n_1297, n_429, n_431);
  nand g1100 (n_449, n_1295, n_1296, n_1297);
  xor g1101 (n_1298, n_432, n_433);
  xor g1102 (n_438, n_1298, n_434);
  nand g1103 (n_1299, n_432, n_433);
  nand g1104 (n_1300, n_434, n_433);
  nand g1105 (n_1301, n_432, n_434);
  nand g1106 (n_451, n_1299, n_1300, n_1301);
  xor g1107 (n_1302, n_435, n_436);
  xor g1108 (n_439, n_1302, n_437);
  nand g1109 (n_1303, n_435, n_436);
  nand g1110 (n_1304, n_437, n_436);
  nand g1111 (n_1305, n_435, n_437);
  nand g1112 (n_454, n_1303, n_1304, n_1305);
  xor g1113 (n_1306, n_438, n_439);
  xor g1114 (n_140, n_1306, n_440);
  nand g1115 (n_1307, n_438, n_439);
  nand g1116 (n_1308, n_440, n_439);
  nand g1117 (n_1309, n_438, n_440);
  nand g1118 (n_77, n_1307, n_1308, n_1309);
  xor g1119 (n_1310, A[28], A[26]);
  xor g1120 (n_445, n_1310, A[22]);
  nand g1121 (n_1311, A[28], A[26]);
  nand g1122 (n_1312, A[22], A[26]);
  nand g1123 (n_1313, A[28], A[22]);
  nand g1124 (n_455, n_1311, n_1312, n_1313);
  xor g1126 (n_446, n_267, A[20]);
  nand g1128 (n_1316, A[20], A[12]);
  xor g1131 (n_1318, A[10], A[24]);
  xor g1132 (n_444, n_1318, A[18]);
  nand g1133 (n_1319, A[10], A[24]);
  nand g1136 (n_457, n_1319, n_1185, n_1252);
  xor g1137 (n_1322, A[16], n_441);
  xor g1138 (n_448, n_1322, n_442);
  nand g1139 (n_1323, A[16], n_441);
  nand g1140 (n_1324, n_442, n_441);
  nand g1141 (n_1325, A[16], n_442);
  nand g1142 (n_461, n_1323, n_1324, n_1325);
  xor g1143 (n_1326, n_443, n_444);
  xor g1144 (n_450, n_1326, n_445);
  nand g1145 (n_1327, n_443, n_444);
  nand g1146 (n_1328, n_445, n_444);
  nand g1147 (n_1329, n_443, n_445);
  nand g1148 (n_463, n_1327, n_1328, n_1329);
  xor g1149 (n_1330, n_446, n_447);
  xor g1150 (n_452, n_1330, n_448);
  nand g1151 (n_1331, n_446, n_447);
  nand g1152 (n_1332, n_448, n_447);
  nand g1153 (n_1333, n_446, n_448);
  nand g1154 (n_465, n_1331, n_1332, n_1333);
  xor g1155 (n_1334, n_449, n_450);
  xor g1156 (n_453, n_1334, n_451);
  nand g1157 (n_1335, n_449, n_450);
  nand g1158 (n_1336, n_451, n_450);
  nand g1159 (n_1337, n_449, n_451);
  nand g1160 (n_468, n_1335, n_1336, n_1337);
  xor g1161 (n_1338, n_452, n_453);
  xor g1162 (n_139, n_1338, n_454);
  nand g1163 (n_1339, n_452, n_453);
  nand g1164 (n_1340, n_454, n_453);
  nand g1165 (n_1341, n_452, n_454);
  nand g1166 (n_76, n_1339, n_1340, n_1341);
  xor g1167 (n_1342, A[29], A[27]);
  xor g1168 (n_459, n_1342, A[23]);
  nand g1169 (n_1343, A[29], A[27]);
  nand g1170 (n_1344, A[23], A[27]);
  nand g1171 (n_1345, A[29], A[23]);
  nand g1172 (n_469, n_1343, n_1344, n_1345);
  xor g1174 (n_460, n_918, A[21]);
  nand g1176 (n_1348, A[21], A[13]);
  nand g1178 (n_470, n_919, n_1348, n_1089);
  xor g1179 (n_1350, A[11], A[25]);
  xor g1180 (n_458, n_1350, A[19]);
  nand g1181 (n_1351, A[11], A[25]);
  nand g1184 (n_471, n_1351, n_1217, n_1284);
  xor g1185 (n_1354, A[17], n_455);
  xor g1186 (n_462, n_1354, n_456);
  nand g1187 (n_1355, A[17], n_455);
  nand g1188 (n_1356, n_456, n_455);
  nand g1189 (n_1357, A[17], n_456);
  nand g1190 (n_475, n_1355, n_1356, n_1357);
  xor g1191 (n_1358, n_457, n_458);
  xor g1192 (n_464, n_1358, n_459);
  nand g1193 (n_1359, n_457, n_458);
  nand g1194 (n_1360, n_459, n_458);
  nand g1195 (n_1361, n_457, n_459);
  nand g1196 (n_477, n_1359, n_1360, n_1361);
  xor g1197 (n_1362, n_460, n_461);
  xor g1198 (n_466, n_1362, n_462);
  nand g1199 (n_1363, n_460, n_461);
  nand g1200 (n_1364, n_462, n_461);
  nand g1201 (n_1365, n_460, n_462);
  nand g1202 (n_479, n_1363, n_1364, n_1365);
  xor g1203 (n_1366, n_463, n_464);
  xor g1204 (n_467, n_1366, n_465);
  nand g1205 (n_1367, n_463, n_464);
  nand g1206 (n_1368, n_465, n_464);
  nand g1207 (n_1369, n_463, n_465);
  nand g1208 (n_482, n_1367, n_1368, n_1369);
  xor g1209 (n_1370, n_466, n_467);
  xor g1210 (n_138, n_1370, n_468);
  nand g1211 (n_1371, n_466, n_467);
  nand g1212 (n_1372, n_468, n_467);
  nand g1213 (n_1373, n_466, n_468);
  nand g1214 (n_75, n_1371, n_1372, n_1373);
  xor g1215 (n_1374, A[30], A[28]);
  xor g1216 (n_473, n_1374, A[24]);
  nand g1217 (n_1375, A[30], A[28]);
  nand g1218 (n_1376, A[24], A[28]);
  nand g1219 (n_1377, A[30], A[24]);
  nand g1220 (n_483, n_1375, n_1376, n_1377);
  xor g1222 (n_474, n_286, A[22]);
  nand g1224 (n_1380, A[22], A[14]);
  xor g1227 (n_1382, A[12], A[26]);
  xor g1228 (n_472, n_1382, A[20]);
  nand g1229 (n_1383, A[12], A[26]);
  nand g1232 (n_485, n_1383, n_1249, n_1316);
  xor g1233 (n_1386, A[18], n_469);
  xor g1234 (n_476, n_1386, n_470);
  nand g1235 (n_1387, A[18], n_469);
  nand g1236 (n_1388, n_470, n_469);
  nand g1237 (n_1389, A[18], n_470);
  nand g1238 (n_489, n_1387, n_1388, n_1389);
  xor g1239 (n_1390, n_471, n_472);
  xor g1240 (n_478, n_1390, n_473);
  nand g1241 (n_1391, n_471, n_472);
  nand g1242 (n_1392, n_473, n_472);
  nand g1243 (n_1393, n_471, n_473);
  nand g1244 (n_491, n_1391, n_1392, n_1393);
  xor g1245 (n_1394, n_474, n_475);
  xor g1246 (n_480, n_1394, n_476);
  nand g1247 (n_1395, n_474, n_475);
  nand g1248 (n_1396, n_476, n_475);
  nand g1249 (n_1397, n_474, n_476);
  nand g1250 (n_493, n_1395, n_1396, n_1397);
  xor g1251 (n_1398, n_477, n_478);
  xor g1252 (n_481, n_1398, n_479);
  nand g1253 (n_1399, n_477, n_478);
  nand g1254 (n_1400, n_479, n_478);
  nand g1255 (n_1401, n_477, n_479);
  nand g1256 (n_496, n_1399, n_1400, n_1401);
  xor g1257 (n_1402, n_480, n_481);
  xor g1258 (n_137, n_1402, n_482);
  nand g1259 (n_1403, n_480, n_481);
  nand g1260 (n_1404, n_482, n_481);
  nand g1261 (n_1405, n_480, n_482);
  nand g1262 (n_74, n_1403, n_1404, n_1405);
  xor g1263 (n_1406, A[31], A[29]);
  xor g1264 (n_487, n_1406, A[25]);
  nand g1265 (n_1407, A[31], A[29]);
  nand g1266 (n_1408, A[25], A[29]);
  nand g1267 (n_1409, A[31], A[25]);
  nand g1268 (n_497, n_1407, n_1408, n_1409);
  xor g1270 (n_488, n_966, A[23]);
  nand g1272 (n_1412, A[23], A[15]);
  nand g1274 (n_499, n_967, n_1412, n_1153);
  xor g1275 (n_1414, A[13], A[27]);
  xor g1276 (n_486, n_1414, A[21]);
  nand g1277 (n_1415, A[13], A[27]);
  nand g1280 (n_498, n_1415, n_1281, n_1348);
  xor g1281 (n_1418, A[19], n_483);
  xor g1282 (n_490, n_1418, n_484);
  nand g1283 (n_1419, A[19], n_483);
  nand g1284 (n_1420, n_484, n_483);
  nand g1285 (n_1421, A[19], n_484);
  nand g1286 (n_503, n_1419, n_1420, n_1421);
  xor g1287 (n_1422, n_485, n_486);
  xor g1288 (n_492, n_1422, n_487);
  nand g1289 (n_1423, n_485, n_486);
  nand g1290 (n_1424, n_487, n_486);
  nand g1291 (n_1425, n_485, n_487);
  nand g1292 (n_505, n_1423, n_1424, n_1425);
  xor g1293 (n_1426, n_488, n_489);
  xor g1294 (n_494, n_1426, n_490);
  nand g1295 (n_1427, n_488, n_489);
  nand g1296 (n_1428, n_490, n_489);
  nand g1297 (n_1429, n_488, n_490);
  nand g1298 (n_508, n_1427, n_1428, n_1429);
  xor g1299 (n_1430, n_491, n_492);
  xor g1300 (n_495, n_1430, n_493);
  nand g1301 (n_1431, n_491, n_492);
  nand g1302 (n_1432, n_493, n_492);
  nand g1303 (n_1433, n_491, n_493);
  nand g1304 (n_510, n_1431, n_1432, n_1433);
  xor g1305 (n_1434, n_494, n_495);
  xor g1306 (n_136, n_1434, n_496);
  nand g1307 (n_1435, n_494, n_495);
  nand g1308 (n_1436, n_496, n_495);
  nand g1309 (n_1437, n_494, n_496);
  nand g1310 (n_73, n_1435, n_1436, n_1437);
  xor g1311 (n_1438, A[30], A[26]);
  xor g1312 (n_501, n_1438, A[18]);
  nand g1313 (n_1439, A[30], A[26]);
  nand g1314 (n_1440, A[18], A[26]);
  nand g1315 (n_1441, A[30], A[18]);
  nand g1316 (n_511, n_1439, n_1440, n_1441);
  xor g1317 (n_1442, A[16], A[24]);
  xor g1318 (n_502, n_1442, A[14]);
  nand g1319 (n_1443, A[16], A[24]);
  nand g1320 (n_1444, A[14], A[24]);
  xor g1323 (n_1446, A[28], A[22]);
  xor g1324 (n_500, n_1446, A[20]);
  nand g1327 (n_1449, A[28], A[20]);
  nand g1328 (n_512, n_1313, n_1119, n_1449);
  xor g1329 (n_1450, A[32], n_497);
  xor g1330 (n_504, n_1450, n_498);
  nand g1331 (n_1451, A[32], n_497);
  nand g1332 (n_1452, n_498, n_497);
  nand g1333 (n_1453, A[32], n_498);
  nand g1334 (n_517, n_1451, n_1452, n_1453);
  xor g1335 (n_1454, n_499, n_500);
  xor g1336 (n_506, n_1454, n_501);
  nand g1337 (n_1455, n_499, n_500);
  nand g1338 (n_1456, n_501, n_500);
  nand g1339 (n_1457, n_499, n_501);
  nand g1340 (n_519, n_1455, n_1456, n_1457);
  xor g1341 (n_1458, n_502, n_503);
  xor g1342 (n_507, n_1458, n_504);
  nand g1343 (n_1459, n_502, n_503);
  nand g1344 (n_1460, n_504, n_503);
  nand g1345 (n_1461, n_502, n_504);
  nand g1346 (n_522, n_1459, n_1460, n_1461);
  xor g1347 (n_1462, n_505, n_506);
  xor g1348 (n_509, n_1462, n_507);
  nand g1349 (n_1463, n_505, n_506);
  nand g1350 (n_1464, n_507, n_506);
  nand g1351 (n_1465, n_505, n_507);
  nand g1352 (n_524, n_1463, n_1464, n_1465);
  xor g1353 (n_1466, n_508, n_509);
  xor g1354 (n_135, n_1466, n_510);
  nand g1355 (n_1467, n_508, n_509);
  nand g1356 (n_1468, n_510, n_509);
  nand g1357 (n_1469, n_508, n_510);
  nand g1358 (n_72, n_1467, n_1468, n_1469);
  xor g1359 (n_1470, A[31], A[27]);
  xor g1360 (n_515, n_1470, A[19]);
  nand g1361 (n_1471, A[31], A[27]);
  nand g1362 (n_1472, A[19], A[27]);
  nand g1363 (n_1473, A[31], A[19]);
  nand g1364 (n_526, n_1471, n_1472, n_1473);
  xor g1365 (n_1474, A[17], A[25]);
  xor g1366 (n_516, n_1474, A[15]);
  nand g1367 (n_1475, A[17], A[25]);
  nand g1368 (n_1476, A[15], A[25]);
  nand g1370 (n_527, n_1475, n_1476, n_967);
  xor g1371 (n_1478, A[29], A[23]);
  xor g1372 (n_514, n_1478, A[21]);
  nand g1375 (n_1481, A[29], A[21]);
  nand g1376 (n_525, n_1345, n_1151, n_1481);
  xor g1377 (n_1482, A[33], n_511);
  xor g1378 (n_518, n_1482, n_512);
  nand g1379 (n_1483, A[33], n_511);
  nand g1380 (n_1484, n_512, n_511);
  nand g1381 (n_1485, A[33], n_512);
  nand g1382 (n_531, n_1483, n_1484, n_1485);
  xor g1383 (n_1486, n_513, n_514);
  xor g1384 (n_520, n_1486, n_515);
  nand g1385 (n_1487, n_513, n_514);
  nand g1386 (n_1488, n_515, n_514);
  nand g1387 (n_1489, n_513, n_515);
  nand g1388 (n_532, n_1487, n_1488, n_1489);
  xor g1389 (n_1490, n_516, n_517);
  xor g1390 (n_521, n_1490, n_518);
  nand g1391 (n_1491, n_516, n_517);
  nand g1392 (n_1492, n_518, n_517);
  nand g1393 (n_1493, n_516, n_518);
  nand g1394 (n_536, n_1491, n_1492, n_1493);
  xor g1395 (n_1494, n_519, n_520);
  xor g1396 (n_523, n_1494, n_521);
  nand g1397 (n_1495, n_519, n_520);
  nand g1398 (n_1496, n_521, n_520);
  nand g1399 (n_1497, n_519, n_521);
  nand g1400 (n_538, n_1495, n_1496, n_1497);
  xor g1401 (n_1498, n_522, n_523);
  xor g1402 (n_134, n_1498, n_524);
  nand g1403 (n_1499, n_522, n_523);
  nand g1404 (n_1500, n_524, n_523);
  nand g1405 (n_1501, n_522, n_524);
  nand g1406 (n_71, n_1499, n_1500, n_1501);
  xor g1408 (n_528, n_1374, A[20]);
  nand g1411 (n_1505, A[30], A[20]);
  nand g1412 (n_539, n_1375, n_1449, n_1505);
  xor g1413 (n_1506, A[18], A[26]);
  xor g1414 (n_530, n_1506, A[16]);
  nand g1416 (n_1508, A[16], A[26]);
  xor g1420 (n_529, n_1182, A[32]);
  nand g1422 (n_1512, A[32], A[22]);
  nand g1423 (n_1513, A[24], A[32]);
  nand g1424 (n_543, n_1183, n_1512, n_1513);
  xor g1425 (n_1514, A[34], n_525);
  xor g1426 (n_533, n_1514, n_526);
  nand g1427 (n_1515, A[34], n_525);
  nand g1428 (n_1516, n_526, n_525);
  nand g1429 (n_1517, A[34], n_526);
  nand g1430 (n_545, n_1515, n_1516, n_1517);
  xor g1431 (n_1518, n_527, n_528);
  xor g1432 (n_534, n_1518, n_529);
  nand g1433 (n_1519, n_527, n_528);
  nand g1434 (n_1520, n_529, n_528);
  nand g1435 (n_1521, n_527, n_529);
  nand g1436 (n_546, n_1519, n_1520, n_1521);
  xor g1437 (n_1522, n_530, n_531);
  xor g1438 (n_535, n_1522, n_532);
  nand g1439 (n_1523, n_530, n_531);
  nand g1440 (n_1524, n_532, n_531);
  nand g1441 (n_1525, n_530, n_532);
  nand g1442 (n_550, n_1523, n_1524, n_1525);
  xor g1443 (n_1526, n_533, n_534);
  xor g1444 (n_537, n_1526, n_535);
  nand g1445 (n_1527, n_533, n_534);
  nand g1446 (n_1528, n_535, n_534);
  nand g1447 (n_1529, n_533, n_535);
  nand g1448 (n_552, n_1527, n_1528, n_1529);
  xor g1449 (n_1530, n_536, n_537);
  xor g1450 (n_133, n_1530, n_538);
  nand g1451 (n_1531, n_536, n_537);
  nand g1452 (n_1532, n_538, n_537);
  nand g1453 (n_1533, n_536, n_538);
  nand g1454 (n_70, n_1531, n_1532, n_1533);
  xor g1455 (n_1534, A[35], A[29]);
  xor g1456 (n_542, n_1534, A[21]);
  nand g1457 (n_1535, A[35], A[29]);
  nand g1459 (n_1537, A[35], A[21]);
  nand g1460 (n_554, n_1535, n_1481, n_1537);
  xor g1461 (n_1538, A[19], A[27]);
  xor g1462 (n_544, n_1538, A[17]);
  nand g1464 (n_1540, A[17], A[27]);
  nand g1466 (n_555, n_1472, n_1540, n_1023);
  xor g1467 (n_1542, A[31], A[25]);
  xor g1468 (n_541, n_1542, A[23]);
  nand g1471 (n_1545, A[31], A[23]);
  nand g1472 (n_553, n_1409, n_1215, n_1545);
  xor g1473 (n_1546, A[33], n_539);
  xor g1474 (n_547, n_1546, n_540);
  nand g1475 (n_1547, A[33], n_539);
  nand g1476 (n_1548, n_540, n_539);
  nand g1477 (n_1549, A[33], n_540);
  nand g1478 (n_559, n_1547, n_1548, n_1549);
  xor g1479 (n_1550, n_541, n_542);
  xor g1480 (n_548, n_1550, n_543);
  nand g1481 (n_1551, n_541, n_542);
  nand g1482 (n_1552, n_543, n_542);
  nand g1483 (n_1553, n_541, n_543);
  nand g1484 (n_560, n_1551, n_1552, n_1553);
  xor g1485 (n_1554, n_544, n_545);
  xor g1486 (n_549, n_1554, n_546);
  nand g1487 (n_1555, n_544, n_545);
  nand g1488 (n_1556, n_546, n_545);
  nand g1489 (n_1557, n_544, n_546);
  nand g1490 (n_564, n_1555, n_1556, n_1557);
  xor g1491 (n_1558, n_547, n_548);
  xor g1492 (n_551, n_1558, n_549);
  nand g1493 (n_1559, n_547, n_548);
  nand g1494 (n_1560, n_549, n_548);
  nand g1495 (n_1561, n_547, n_549);
  nand g1496 (n_566, n_1559, n_1560, n_1561);
  xor g1497 (n_1562, n_550, n_551);
  xor g1498 (n_132, n_1562, n_552);
  nand g1499 (n_1563, n_550, n_551);
  nand g1500 (n_1564, n_552, n_551);
  nand g1501 (n_1565, n_550, n_552);
  nand g1502 (n_69, n_1563, n_1564, n_1565);
  xor g1504 (n_556, n_1374, A[22]);
  nand g1507 (n_1569, A[30], A[22]);
  nand g1508 (n_567, n_1375, n_1313, n_1569);
  xor g1510 (n_557, n_1054, A[26]);
  nand g1514 (n_568, n_1055, n_1440, n_1249);
  xor g1515 (n_1574, A[24], A[34]);
  xor g1516 (n_558, n_1574, A[36]);
  nand g1517 (n_1575, A[24], A[34]);
  nand g1518 (n_1576, A[36], A[34]);
  nand g1519 (n_1577, A[24], A[36]);
  nand g1520 (n_570, n_1575, n_1576, n_1577);
  xor g1521 (n_1578, A[32], n_553);
  xor g1522 (n_561, n_1578, n_554);
  nand g1523 (n_1579, A[32], n_553);
  nand g1524 (n_1580, n_554, n_553);
  nand g1525 (n_1581, A[32], n_554);
  nand g1526 (n_573, n_1579, n_1580, n_1581);
  xor g1527 (n_1582, n_555, n_556);
  xor g1528 (n_562, n_1582, n_557);
  nand g1529 (n_1583, n_555, n_556);
  nand g1530 (n_1584, n_557, n_556);
  nand g1531 (n_1585, n_555, n_557);
  nand g1532 (n_574, n_1583, n_1584, n_1585);
  xor g1533 (n_1586, n_558, n_559);
  xor g1534 (n_563, n_1586, n_560);
  nand g1535 (n_1587, n_558, n_559);
  nand g1536 (n_1588, n_560, n_559);
  nand g1537 (n_1589, n_558, n_560);
  nand g1538 (n_578, n_1587, n_1588, n_1589);
  xor g1539 (n_1590, n_561, n_562);
  xor g1540 (n_565, n_1590, n_563);
  nand g1541 (n_1591, n_561, n_562);
  nand g1542 (n_1592, n_563, n_562);
  nand g1543 (n_1593, n_561, n_563);
  nand g1544 (n_580, n_1591, n_1592, n_1593);
  xor g1545 (n_1594, n_564, n_565);
  xor g1546 (n_131, n_1594, n_566);
  nand g1547 (n_1595, n_564, n_565);
  nand g1548 (n_1596, n_566, n_565);
  nand g1549 (n_1597, n_564, n_566);
  nand g1550 (n_68, n_1595, n_1596, n_1597);
  xor g1551 (n_1598, A[35], A[31]);
  xor g1552 (n_569, n_1598, A[23]);
  nand g1553 (n_1599, A[35], A[31]);
  nand g1555 (n_1601, A[35], A[23]);
  nand g1556 (n_581, n_1599, n_1545, n_1601);
  xor g1557 (n_1602, A[21], A[29]);
  xor g1558 (n_572, n_1602, A[19]);
  nand g1560 (n_1604, A[19], A[29]);
  nand g1562 (n_582, n_1481, n_1604, n_1087);
  xor g1564 (n_571, n_1278, A[37]);
  nand g1566 (n_1608, A[37], A[25]);
  nand g1567 (n_1609, A[27], A[37]);
  nand g1568 (n_584, n_1279, n_1608, n_1609);
  xor g1569 (n_1610, A[33], n_567);
  xor g1570 (n_575, n_1610, n_568);
  nand g1571 (n_1611, A[33], n_567);
  nand g1572 (n_1612, n_568, n_567);
  nand g1573 (n_1613, A[33], n_568);
  nand g1574 (n_587, n_1611, n_1612, n_1613);
  xor g1575 (n_1614, n_569, n_570);
  xor g1576 (n_576, n_1614, n_571);
  nand g1577 (n_1615, n_569, n_570);
  nand g1578 (n_1616, n_571, n_570);
  nand g1579 (n_1617, n_569, n_571);
  nand g1580 (n_588, n_1615, n_1616, n_1617);
  xor g1581 (n_1618, n_572, n_573);
  xor g1582 (n_577, n_1618, n_574);
  nand g1583 (n_1619, n_572, n_573);
  nand g1584 (n_1620, n_574, n_573);
  nand g1585 (n_1621, n_572, n_574);
  nand g1586 (n_592, n_1619, n_1620, n_1621);
  xor g1587 (n_1622, n_575, n_576);
  xor g1588 (n_579, n_1622, n_577);
  nand g1589 (n_1623, n_575, n_576);
  nand g1590 (n_1624, n_577, n_576);
  nand g1591 (n_1625, n_575, n_577);
  nand g1592 (n_594, n_1623, n_1624, n_1625);
  xor g1593 (n_1626, n_578, n_579);
  xor g1594 (n_130, n_1626, n_580);
  nand g1595 (n_1627, n_578, n_579);
  nand g1596 (n_1628, n_580, n_579);
  nand g1597 (n_1629, n_578, n_580);
  nand g1598 (n_67, n_1627, n_1628, n_1629);
  xor g1599 (n_1630, A[30], A[24]);
  xor g1600 (n_583, n_1630, A[22]);
  nand g1604 (n_595, n_1377, n_1183, n_1569);
  xor g1605 (n_1634, A[20], A[28]);
  xor g1606 (n_585, n_1634, A[26]);
  nand g1610 (n_596, n_1449, n_1311, n_1249);
  xor g1611 (n_1638, A[32], A[38]);
  xor g1612 (n_586, n_1638, A[36]);
  nand g1613 (n_1639, A[32], A[38]);
  nand g1614 (n_1640, A[36], A[38]);
  nand g1615 (n_1641, A[32], A[36]);
  nand g1616 (n_598, n_1639, n_1640, n_1641);
  xor g1617 (n_1642, A[34], n_581);
  xor g1618 (n_589, n_1642, n_582);
  nand g1619 (n_1643, A[34], n_581);
  nand g1620 (n_1644, n_582, n_581);
  nand g1621 (n_1645, A[34], n_582);
  nand g1622 (n_601, n_1643, n_1644, n_1645);
  xor g1623 (n_1646, n_583, n_584);
  xor g1624 (n_590, n_1646, n_585);
  nand g1625 (n_1647, n_583, n_584);
  nand g1626 (n_1648, n_585, n_584);
  nand g1627 (n_1649, n_583, n_585);
  nand g1628 (n_602, n_1647, n_1648, n_1649);
  xor g1629 (n_1650, n_586, n_587);
  xor g1630 (n_591, n_1650, n_588);
  nand g1631 (n_1651, n_586, n_587);
  nand g1632 (n_1652, n_588, n_587);
  nand g1633 (n_1653, n_586, n_588);
  nand g1634 (n_606, n_1651, n_1652, n_1653);
  xor g1635 (n_1654, n_589, n_590);
  xor g1636 (n_593, n_1654, n_591);
  nand g1637 (n_1655, n_589, n_590);
  nand g1638 (n_1656, n_591, n_590);
  nand g1639 (n_1657, n_589, n_591);
  nand g1640 (n_608, n_1655, n_1656, n_1657);
  xor g1641 (n_1658, n_592, n_593);
  xor g1642 (n_129, n_1658, n_594);
  nand g1643 (n_1659, n_592, n_593);
  nand g1644 (n_1660, n_594, n_593);
  nand g1645 (n_1661, n_592, n_594);
  nand g1646 (n_66, n_1659, n_1660, n_1661);
  xor g1648 (n_597, n_1598, A[25]);
  nand g1651 (n_1665, A[35], A[25]);
  nand g1652 (n_609, n_1599, n_1409, n_1665);
  xor g1654 (n_599, n_1150, A[29]);
  xor g1659 (n_1670, A[27], A[33]);
  xor g1660 (n_600, n_1670, A[37]);
  nand g1661 (n_1671, A[27], A[33]);
  nand g1662 (n_1672, A[37], A[33]);
  nand g1664 (n_612, n_1671, n_1672, n_1609);
  xor g1665 (n_1674, A[39], n_595);
  xor g1666 (n_603, n_1674, n_596);
  nand g1667 (n_1675, A[39], n_595);
  nand g1668 (n_1676, n_596, n_595);
  nand g1669 (n_1677, A[39], n_596);
  nand g1670 (n_615, n_1675, n_1676, n_1677);
  xor g1671 (n_1678, n_597, n_598);
  xor g1672 (n_604, n_1678, n_599);
  nand g1673 (n_1679, n_597, n_598);
  nand g1674 (n_1680, n_599, n_598);
  nand g1675 (n_1681, n_597, n_599);
  nand g1676 (n_616, n_1679, n_1680, n_1681);
  xor g1677 (n_1682, n_600, n_601);
  xor g1678 (n_605, n_1682, n_602);
  nand g1679 (n_1683, n_600, n_601);
  nand g1680 (n_1684, n_602, n_601);
  nand g1681 (n_1685, n_600, n_602);
  nand g1682 (n_620, n_1683, n_1684, n_1685);
  xor g1683 (n_1686, n_603, n_604);
  xor g1684 (n_607, n_1686, n_605);
  nand g1685 (n_1687, n_603, n_604);
  nand g1686 (n_1688, n_605, n_604);
  nand g1687 (n_1689, n_603, n_605);
  nand g1688 (n_622, n_1687, n_1688, n_1689);
  xor g1689 (n_1690, n_606, n_607);
  xor g1690 (n_128, n_1690, n_608);
  nand g1691 (n_1691, n_606, n_607);
  nand g1692 (n_1692, n_608, n_607);
  nand g1693 (n_1693, n_606, n_608);
  nand g1694 (n_65, n_1691, n_1692, n_1693);
  xor g1695 (n_1694, A[40], A[26]);
  xor g1696 (n_611, n_1694, A[24]);
  nand g1697 (n_1695, A[40], A[26]);
  nand g1699 (n_1697, A[40], A[24]);
  nand g1700 (n_623, n_1695, n_1247, n_1697);
  xor g1701 (n_1698, A[22], A[30]);
  xor g1702 (n_613, n_1698, A[28]);
  xor g1707 (n_1702, A[34], A[38]);
  xor g1708 (n_614, n_1702, A[32]);
  nand g1709 (n_1703, A[34], A[38]);
  nand g1711 (n_1705, A[34], A[32]);
  nand g1712 (n_626, n_1703, n_1639, n_1705);
  xor g1713 (n_1706, A[36], n_609);
  xor g1714 (n_617, n_1706, n_525);
  nand g1715 (n_1707, A[36], n_609);
  nand g1716 (n_1708, n_525, n_609);
  nand g1717 (n_1709, A[36], n_525);
  nand g1718 (n_629, n_1707, n_1708, n_1709);
  xor g1719 (n_1710, n_611, n_612);
  xor g1720 (n_618, n_1710, n_613);
  nand g1721 (n_1711, n_611, n_612);
  nand g1722 (n_1712, n_613, n_612);
  nand g1723 (n_1713, n_611, n_613);
  nand g1724 (n_630, n_1711, n_1712, n_1713);
  xor g1725 (n_1714, n_614, n_615);
  xor g1726 (n_619, n_1714, n_616);
  nand g1727 (n_1715, n_614, n_615);
  nand g1728 (n_1716, n_616, n_615);
  nand g1729 (n_1717, n_614, n_616);
  nand g1730 (n_634, n_1715, n_1716, n_1717);
  xor g1731 (n_1718, n_617, n_618);
  xor g1732 (n_621, n_1718, n_619);
  nand g1733 (n_1719, n_617, n_618);
  nand g1734 (n_1720, n_619, n_618);
  nand g1735 (n_1721, n_617, n_619);
  nand g1736 (n_636, n_1719, n_1720, n_1721);
  xor g1737 (n_1722, n_620, n_621);
  xor g1738 (n_127, n_1722, n_622);
  nand g1739 (n_1723, n_620, n_621);
  nand g1740 (n_1724, n_622, n_621);
  nand g1741 (n_1725, n_620, n_622);
  nand g1742 (n_64, n_1723, n_1724, n_1725);
  xor g1743 (n_1726, A[35], A[27]);
  xor g1744 (n_625, n_1726, A[25]);
  nand g1745 (n_1727, A[35], A[27]);
  nand g1748 (n_639, n_1727, n_1279, n_1665);
  xor g1749 (n_1730, A[23], A[31]);
  xor g1750 (n_627, n_1730, A[29]);
  nand g1754 (n_640, n_1545, n_1407, n_1345);
  xor g1755 (n_1734, A[39], A[41]);
  xor g1756 (n_628, n_1734, A[33]);
  nand g1757 (n_1735, A[39], A[41]);
  nand g1758 (n_1736, A[33], A[41]);
  nand g1759 (n_1737, A[39], A[33]);
  nand g1760 (n_643, n_1735, n_1736, n_1737);
  xor g1761 (n_1738, A[37], n_623);
  xor g1762 (n_631, n_1738, n_567);
  nand g1763 (n_1739, A[37], n_623);
  nand g1764 (n_1740, n_567, n_623);
  nand g1765 (n_1741, A[37], n_567);
  nand g1766 (n_645, n_1739, n_1740, n_1741);
  xor g1767 (n_1742, n_625, n_626);
  xor g1768 (n_632, n_1742, n_627);
  nand g1769 (n_1743, n_625, n_626);
  nand g1770 (n_1744, n_627, n_626);
  nand g1771 (n_1745, n_625, n_627);
  nand g1772 (n_646, n_1743, n_1744, n_1745);
  xor g1773 (n_1746, n_628, n_629);
  xor g1774 (n_633, n_1746, n_630);
  nand g1775 (n_1747, n_628, n_629);
  nand g1776 (n_1748, n_630, n_629);
  nand g1777 (n_1749, n_628, n_630);
  nand g1778 (n_650, n_1747, n_1748, n_1749);
  xor g1779 (n_1750, n_631, n_632);
  xor g1780 (n_635, n_1750, n_633);
  nand g1781 (n_1751, n_631, n_632);
  nand g1782 (n_1752, n_633, n_632);
  nand g1783 (n_1753, n_631, n_633);
  nand g1784 (n_652, n_1751, n_1752, n_1753);
  xor g1785 (n_1754, n_634, n_635);
  xor g1786 (n_126, n_1754, n_636);
  nand g1787 (n_1755, n_634, n_635);
  nand g1788 (n_1756, n_636, n_635);
  nand g1789 (n_1757, n_634, n_636);
  nand g1790 (n_63, n_1755, n_1756, n_1757);
  xor g1793 (n_1758, A[42], A[28]);
  xor g1794 (n_642, n_1758, A[26]);
  nand g1795 (n_1759, A[42], A[28]);
  nand g1797 (n_1761, A[42], A[26]);
  nand g1798 (n_657, n_1759, n_1311, n_1761);
  xor g1799 (n_1762, A[40], A[24]);
  xor g1800 (n_641, n_1762, A[30]);
  nand g1803 (n_1765, A[40], A[30]);
  nand g1804 (n_656, n_1697, n_1377, n_1765);
  xor g1805 (n_1766, A[36], A[34]);
  xor g1806 (n_644, n_1766, A[32]);
  nand g1810 (n_660, n_1576, n_1705, n_1641);
  xor g1811 (n_1770, A[38], n_639);
  xor g1812 (n_647, n_1770, n_640);
  nand g1813 (n_1771, A[38], n_639);
  nand g1814 (n_1772, n_640, n_639);
  nand g1815 (n_1773, A[38], n_640);
  nand g1816 (n_662, n_1771, n_1772, n_1773);
  xor g1817 (n_1774, n_641, n_642);
  xor g1818 (n_648, n_1774, n_643);
  nand g1819 (n_1775, n_641, n_642);
  nand g1820 (n_1776, n_643, n_642);
  nand g1821 (n_1777, n_641, n_643);
  nand g1822 (n_663, n_1775, n_1776, n_1777);
  xor g1823 (n_1778, n_644, n_645);
  xor g1824 (n_649, n_1778, n_646);
  nand g1825 (n_1779, n_644, n_645);
  nand g1826 (n_1780, n_646, n_645);
  nand g1827 (n_1781, n_644, n_646);
  nand g1828 (n_667, n_1779, n_1780, n_1781);
  xor g1829 (n_1782, n_647, n_648);
  xor g1830 (n_651, n_1782, n_649);
  nand g1831 (n_1783, n_647, n_648);
  nand g1832 (n_1784, n_649, n_648);
  nand g1833 (n_1785, n_647, n_649);
  nand g1834 (n_669, n_1783, n_1784, n_1785);
  xor g1835 (n_1786, n_650, n_651);
  xor g1836 (n_125, n_1786, n_652);
  nand g1837 (n_1787, n_650, n_651);
  nand g1838 (n_1788, n_652, n_651);
  nand g1839 (n_1789, n_650, n_652);
  nand g1840 (n_62, n_1787, n_1788, n_1789);
  xor g1843 (n_1790, A[25], A[35]);
  xor g1844 (n_658, n_1790, A[42]);
  nand g1846 (n_1792, A[42], A[35]);
  nand g1847 (n_1793, A[25], A[42]);
  nand g1848 (n_671, n_1665, n_1792, n_1793);
  xor g1850 (n_659, n_1470, A[29]);
  nand g1854 (n_672, n_1471, n_1407, n_1343);
  xor g1861 (n_1802, A[37], n_656);
  xor g1862 (n_664, n_1802, n_657);
  nand g1863 (n_1803, A[37], n_656);
  nand g1864 (n_1804, n_657, n_656);
  nand g1865 (n_1805, A[37], n_657);
  nand g1866 (n_677, n_1803, n_1804, n_1805);
  xor g1867 (n_1806, n_658, n_659);
  xor g1868 (n_665, n_1806, n_660);
  nand g1869 (n_1807, n_658, n_659);
  nand g1870 (n_1808, n_660, n_659);
  nand g1871 (n_1809, n_658, n_660);
  nand g1872 (n_678, n_1807, n_1808, n_1809);
  xor g1873 (n_1810, n_628, n_662);
  xor g1874 (n_666, n_1810, n_663);
  nand g1875 (n_1811, n_628, n_662);
  nand g1876 (n_1812, n_663, n_662);
  nand g1877 (n_1813, n_628, n_663);
  nand g1878 (n_682, n_1811, n_1812, n_1813);
  xor g1879 (n_1814, n_664, n_665);
  xor g1880 (n_668, n_1814, n_666);
  nand g1881 (n_1815, n_664, n_665);
  nand g1882 (n_1816, n_666, n_665);
  nand g1883 (n_1817, n_664, n_666);
  nand g1884 (n_684, n_1815, n_1816, n_1817);
  xor g1885 (n_1818, n_667, n_668);
  xor g1886 (n_124, n_1818, n_669);
  nand g1887 (n_1819, n_667, n_668);
  nand g1888 (n_1820, n_669, n_668);
  nand g1889 (n_1821, n_667, n_669);
  nand g1890 (n_61, n_1819, n_1820, n_1821);
  xor g1892 (n_673, n_1822, A[28]);
  nand g1894 (n_1824, A[28], A[40]);
  nand g1896 (n_687, n_1823, n_1824, n_1825);
  xor g1898 (n_674, n_1826, A[30]);
  nand g1902 (n_688, n_1827, n_1828, n_1439);
  xor g1909 (n_1834, A[38], n_671);
  xor g1910 (n_679, n_1834, n_672);
  nand g1911 (n_1835, A[38], n_671);
  nand g1912 (n_1836, n_672, n_671);
  nand g1913 (n_1837, A[38], n_672);
  nand g1914 (n_692, n_1835, n_1836, n_1837);
  xor g1915 (n_1838, n_673, n_674);
  xor g1916 (n_680, n_1838, n_643);
  nand g1917 (n_1839, n_673, n_674);
  nand g1918 (n_1840, n_643, n_674);
  nand g1919 (n_1841, n_673, n_643);
  nand g1920 (n_694, n_1839, n_1840, n_1841);
  xor g1921 (n_1842, n_644, n_677);
  xor g1922 (n_681, n_1842, n_678);
  nand g1923 (n_1843, n_644, n_677);
  nand g1924 (n_1844, n_678, n_677);
  nand g1925 (n_1845, n_644, n_678);
  nand g1926 (n_696, n_1843, n_1844, n_1845);
  xor g1927 (n_1846, n_679, n_680);
  xor g1928 (n_683, n_1846, n_681);
  nand g1929 (n_1847, n_679, n_680);
  nand g1930 (n_1848, n_681, n_680);
  nand g1931 (n_1849, n_679, n_681);
  nand g1932 (n_699, n_1847, n_1848, n_1849);
  xor g1933 (n_1850, n_682, n_683);
  xor g1934 (n_123, n_1850, n_684);
  nand g1935 (n_1851, n_682, n_683);
  nand g1936 (n_1852, n_684, n_683);
  nand g1937 (n_1853, n_682, n_684);
  nand g1938 (n_60, n_1851, n_1852, n_1853);
  xor g1954 (n_693, n_1862, n_687);
  nand g1957 (n_1865, A[37], n_687);
  nand g1958 (n_706, n_1863, n_1864, n_1865);
  xor g1959 (n_1866, n_688, n_660);
  xor g1960 (n_695, n_1866, n_659);
  nand g1961 (n_1867, n_688, n_660);
  nand g1963 (n_1869, n_688, n_659);
  nand g1964 (n_707, n_1867, n_1808, n_1869);
  xor g1965 (n_1870, n_628, n_692);
  xor g1966 (n_697, n_1870, n_693);
  nand g1967 (n_1871, n_628, n_692);
  nand g1968 (n_1872, n_693, n_692);
  nand g1969 (n_1873, n_628, n_693);
  nand g1970 (n_710, n_1871, n_1872, n_1873);
  xor g1971 (n_1874, n_694, n_695);
  xor g1972 (n_698, n_1874, n_696);
  nand g1973 (n_1875, n_694, n_695);
  nand g1974 (n_1876, n_696, n_695);
  nand g1975 (n_1877, n_694, n_696);
  nand g1976 (n_712, n_1875, n_1876, n_1877);
  xor g1977 (n_1878, n_697, n_698);
  xor g1978 (n_122, n_1878, n_699);
  nand g1979 (n_1879, n_697, n_698);
  nand g1980 (n_1880, n_699, n_698);
  nand g1981 (n_1881, n_697, n_699);
  nand g1982 (n_59, n_1879, n_1880, n_1881);
  xor g1989 (n_1886, A[30], A[36]);
  xor g1990 (n_705, n_1886, A[34]);
  nand g1991 (n_1887, A[30], A[36]);
  nand g1993 (n_1889, A[30], A[34]);
  nand g1994 (n_716, n_1887, n_1576, n_1889);
  xor g1996 (n_704, n_1638, A[35]);
  nand g1998 (n_1892, A[35], A[38]);
  nand g1999 (n_1893, A[32], A[35]);
  nand g2000 (n_719, n_1639, n_1892, n_1893);
  xor g2001 (n_1894, n_672, n_673);
  xor g2002 (n_708, n_1894, n_643);
  nand g2003 (n_1895, n_672, n_673);
  nand g2005 (n_1897, n_672, n_643);
  nand g2006 (n_721, n_1895, n_1841, n_1897);
  xor g2007 (n_1898, n_704, n_705);
  xor g2008 (n_709, n_1898, n_706);
  nand g2009 (n_1899, n_704, n_705);
  nand g2010 (n_1900, n_706, n_705);
  nand g2011 (n_1901, n_704, n_706);
  nand g2012 (n_722, n_1899, n_1900, n_1901);
  xor g2013 (n_1902, n_707, n_708);
  xor g2014 (n_711, n_1902, n_709);
  nand g2015 (n_1903, n_707, n_708);
  nand g2016 (n_1904, n_709, n_708);
  nand g2017 (n_1905, n_707, n_709);
  nand g2018 (n_725, n_1903, n_1904, n_1905);
  xor g2019 (n_1906, n_710, n_711);
  xor g2020 (n_121, n_1906, n_712);
  nand g2021 (n_1907, n_710, n_711);
  nand g2022 (n_1908, n_712, n_711);
  nand g2023 (n_1909, n_710, n_712);
  nand g2024 (n_58, n_1907, n_1908, n_1909);
  xor g2028 (n_717, n_1406, A[41]);
  nand g2030 (n_1912, A[41], A[29]);
  nand g2031 (n_1913, A[31], A[41]);
  nand g2032 (n_727, n_1407, n_1912, n_1913);
  xor g2033 (n_1914, A[39], A[33]);
  xor g2034 (n_718, n_1914, A[37]);
  nand g2037 (n_1917, A[39], A[37]);
  nand g2038 (n_728, n_1737, n_1672, n_1917);
  xor g2040 (n_720, n_1918, n_716);
  nand g2042 (n_1920, n_716, n_687);
  nand g2044 (n_732, n_1864, n_1920, n_1921);
  xor g2045 (n_1922, n_717, n_718);
  xor g2046 (n_723, n_1922, n_719);
  nand g2047 (n_1923, n_717, n_718);
  nand g2048 (n_1924, n_719, n_718);
  nand g2049 (n_1925, n_717, n_719);
  nand g2050 (n_733, n_1923, n_1924, n_1925);
  xor g2051 (n_1926, n_720, n_721);
  xor g2052 (n_724, n_1926, n_722);
  nand g2053 (n_1927, n_720, n_721);
  nand g2054 (n_1928, n_722, n_721);
  nand g2055 (n_1929, n_720, n_722);
  nand g2056 (n_736, n_1927, n_1928, n_1929);
  xor g2057 (n_1930, n_723, n_724);
  xor g2058 (n_120, n_1930, n_725);
  nand g2059 (n_1931, n_723, n_724);
  nand g2060 (n_1932, n_725, n_724);
  nand g2061 (n_1933, n_723, n_725);
  nand g2062 (n_57, n_1931, n_1932, n_1933);
  xor g2064 (n_729, n_1822, A[30]);
  nand g2068 (n_739, n_1823, n_1765, n_1828);
  xor g2075 (n_1942, A[38], A[35]);
  xor g2076 (n_731, n_1942, n_727);
  nand g2078 (n_1944, n_727, A[35]);
  nand g2079 (n_1945, A[38], n_727);
  nand g2080 (n_743, n_1892, n_1944, n_1945);
  xor g2081 (n_1946, n_728, n_729);
  xor g2082 (n_734, n_1946, n_644);
  nand g2083 (n_1947, n_728, n_729);
  nand g2084 (n_1948, n_644, n_729);
  nand g2085 (n_1949, n_728, n_644);
  nand g2086 (n_744, n_1947, n_1948, n_1949);
  xor g2087 (n_1950, n_731, n_732);
  xor g2088 (n_735, n_1950, n_733);
  nand g2089 (n_1951, n_731, n_732);
  nand g2090 (n_1952, n_733, n_732);
  nand g2091 (n_1953, n_731, n_733);
  nand g2092 (n_747, n_1951, n_1952, n_1953);
  xor g2093 (n_1954, n_734, n_735);
  xor g2094 (n_119, n_1954, n_736);
  nand g2095 (n_1955, n_734, n_735);
  nand g2096 (n_1956, n_736, n_735);
  nand g2097 (n_1957, n_734, n_736);
  nand g2098 (n_56, n_1955, n_1956, n_1957);
  xor g2101 (n_1958, A[31], A[41]);
  xor g2102 (n_742, n_1958, A[39]);
  nand g2105 (n_1961, A[31], A[39]);
  nand g2106 (n_749, n_1913, n_1735, n_1961);
  xor g2107 (n_1962, A[33], A[37]);
  nand g2112 (n_751, n_1672, n_1863, n_1965);
  xor g2113 (n_1966, n_739, n_660);
  xor g2114 (n_745, n_1966, n_741);
  nand g2115 (n_1967, n_739, n_660);
  nand g2116 (n_1968, n_741, n_660);
  nand g2117 (n_1969, n_739, n_741);
  nand g2118 (n_754, n_1967, n_1968, n_1969);
  xor g2119 (n_1970, n_742, n_743);
  xor g2120 (n_746, n_1970, n_744);
  nand g2121 (n_1971, n_742, n_743);
  nand g2122 (n_1972, n_744, n_743);
  nand g2123 (n_1973, n_742, n_744);
  nand g2124 (n_756, n_1971, n_1972, n_1973);
  xor g2125 (n_1974, n_745, n_746);
  xor g2126 (n_118, n_1974, n_747);
  nand g2127 (n_1975, n_745, n_746);
  nand g2128 (n_1976, n_747, n_746);
  nand g2129 (n_1977, n_745, n_747);
  nand g2130 (n_55, n_1975, n_1976, n_1977);
  xor g2132 (n_750, n_1822, A[36]);
  nand g2134 (n_1980, A[36], A[40]);
  nand g2136 (n_760, n_1823, n_1980, n_1981);
  xor g2143 (n_1986, A[35], n_749);
  xor g2144 (n_753, n_1986, n_750);
  nand g2145 (n_1987, A[35], n_749);
  nand g2146 (n_1988, n_750, n_749);
  nand g2147 (n_1989, A[35], n_750);
  nand g2148 (n_762, n_1987, n_1988, n_1989);
  xor g2149 (n_1990, n_751, n_614);
  xor g2150 (n_755, n_1990, n_753);
  nand g2151 (n_1991, n_751, n_614);
  nand g2152 (n_1992, n_753, n_614);
  nand g2153 (n_1993, n_751, n_753);
  nand g2154 (n_765, n_1991, n_1992, n_1993);
  xor g2155 (n_1994, n_754, n_755);
  xor g2156 (n_117, n_1994, n_756);
  nand g2157 (n_1995, n_754, n_755);
  nand g2158 (n_1996, n_756, n_755);
  nand g2159 (n_1997, n_754, n_756);
  nand g2160 (n_54, n_1995, n_1996, n_1997);
  xor g2170 (n_763, n_1862, n_626);
  nand g2173 (n_2005, A[37], n_626);
  nand g2174 (n_770, n_1863, n_2004, n_2005);
  xor g2175 (n_2006, n_760, n_628);
  xor g2176 (n_764, n_2006, n_762);
  nand g2177 (n_2007, n_760, n_628);
  nand g2178 (n_2008, n_762, n_628);
  nand g2179 (n_2009, n_760, n_762);
  nand g2180 (n_772, n_2007, n_2008, n_2009);
  xor g2181 (n_2010, n_763, n_764);
  xor g2182 (n_116, n_2010, n_765);
  nand g2183 (n_2011, n_763, n_764);
  nand g2184 (n_2012, n_765, n_764);
  nand g2185 (n_2013, n_763, n_765);
  nand g2186 (n_115, n_2011, n_2012, n_2013);
  xor g2194 (n_769, n_1702, A[35]);
  nand g2197 (n_2021, A[34], A[35]);
  nand g2198 (n_776, n_1703, n_1892, n_2021);
  xor g2199 (n_2022, n_750, n_643);
  xor g2200 (n_771, n_2022, n_769);
  nand g2201 (n_2023, n_750, n_643);
  nand g2202 (n_2024, n_769, n_643);
  nand g2203 (n_2025, n_750, n_769);
  nand g2204 (n_779, n_2023, n_2024, n_2025);
  xor g2205 (n_2026, n_770, n_771);
  xor g2206 (n_53, n_2026, n_772);
  nand g2207 (n_2027, n_770, n_771);
  nand g2208 (n_2028, n_772, n_771);
  nand g2209 (n_2029, n_770, n_772);
  nand g2210 (n_114, n_2027, n_2028, n_2029);
  xor g2214 (n_777, n_1734, A[37]);
  nand g2216 (n_2032, A[37], A[41]);
  nand g2218 (n_782, n_1735, n_2032, n_1917);
  xor g2220 (n_778, n_2034, n_776);
  nand g2222 (n_2036, n_776, n_760);
  nand g2224 (n_784, n_2035, n_2036, n_2037);
  xor g2225 (n_2038, n_777, n_778);
  xor g2226 (n_52, n_2038, n_779);
  nand g2227 (n_2039, n_777, n_778);
  nand g2228 (n_2040, n_779, n_778);
  nand g2229 (n_2041, n_777, n_779);
  nand g2230 (n_51, n_2039, n_2040, n_2041);
  xor g2238 (n_783, n_1942, n_750);
  nand g2241 (n_2049, A[38], n_750);
  nand g2242 (n_789, n_1892, n_1989, n_2049);
  xor g2243 (n_2050, n_782, n_783);
  xor g2244 (n_113, n_2050, n_784);
  nand g2245 (n_2051, n_782, n_783);
  nand g2246 (n_2052, n_784, n_783);
  nand g2247 (n_2053, n_782, n_784);
  nand g2248 (n_112, n_2051, n_2052, n_2053);
  xor g2251 (n_2054, A[39], A[37]);
  nand g2256 (n_792, n_1917, n_2056, n_2057);
  xor g2257 (n_2058, n_760, n_788);
  xor g2258 (n_50, n_2058, n_789);
  nand g2259 (n_2059, n_760, n_788);
  nand g2260 (n_2060, n_789, n_788);
  nand g2261 (n_2061, n_760, n_789);
  nand g2262 (n_111, n_2059, n_2060, n_2061);
  xor g2264 (n_791, n_1822, A[38]);
  nand g2266 (n_2064, A[38], A[40]);
  nand g2268 (n_795, n_1823, n_2064, n_2065);
  xor g2269 (n_2066, A[41], n_791);
  xor g2270 (n_49, n_2066, n_792);
  nand g2271 (n_2067, A[41], n_791);
  nand g2272 (n_2068, n_792, n_791);
  nand g2273 (n_2069, A[41], n_792);
  nand g2274 (n_110, n_2067, n_2068, n_2069);
  nand g2281 (n_2073, A[41], n_795);
  nand g2282 (n_109, n_2071, n_2072, n_2073);
  xor g2284 (n_47, n_1822, A[39]);
  nand g2286 (n_2076, A[39], A[40]);
  nand g2288 (n_108, n_1823, n_2076, n_2077);
  nor g11 (n_2093, A[2], A[0]);
  nor g13 (n_2089, A[3], A[1]);
  nor g15 (n_2099, A[2], n_163);
  nand g16 (n_2094, A[2], n_163);
  nor g17 (n_2095, n_100, n_162);
  nand g18 (n_2096, n_100, n_162);
  nor g19 (n_2105, n_99, n_161);
  nand g20 (n_2100, n_99, n_161);
  nor g21 (n_2101, n_98, n_160);
  nand g22 (n_2102, n_98, n_160);
  nor g23 (n_2111, n_97, n_159);
  nand g24 (n_2106, n_97, n_159);
  nor g25 (n_2107, n_96, n_158);
  nand g26 (n_2108, n_96, n_158);
  nor g27 (n_2117, n_95, n_157);
  nand g28 (n_2112, n_95, n_157);
  nor g29 (n_2113, n_94, n_156);
  nand g30 (n_2114, n_94, n_156);
  nor g31 (n_2123, n_93, n_155);
  nand g32 (n_2118, n_93, n_155);
  nor g33 (n_2119, n_92, n_154);
  nand g34 (n_2120, n_92, n_154);
  nor g35 (n_2129, n_91, n_153);
  nand g36 (n_2124, n_91, n_153);
  nor g37 (n_2125, n_90, n_152);
  nand g38 (n_2126, n_90, n_152);
  nor g39 (n_2135, n_89, n_151);
  nand g40 (n_2130, n_89, n_151);
  nor g41 (n_2131, n_88, n_150);
  nand g42 (n_2132, n_88, n_150);
  nor g43 (n_2141, n_87, n_149);
  nand g44 (n_2136, n_87, n_149);
  nor g45 (n_2137, n_86, n_148);
  nand g46 (n_2138, n_86, n_148);
  nor g47 (n_2147, n_85, n_147);
  nand g48 (n_2142, n_85, n_147);
  nor g49 (n_2143, n_84, n_146);
  nand g50 (n_2144, n_84, n_146);
  nor g51 (n_2153, n_83, n_145);
  nand g52 (n_2148, n_83, n_145);
  nor g53 (n_2149, n_82, n_144);
  nand g54 (n_2150, n_82, n_144);
  nor g55 (n_2159, n_81, n_143);
  nand g56 (n_2154, n_81, n_143);
  nor g57 (n_2155, n_80, n_142);
  nand g58 (n_2156, n_80, n_142);
  nor g59 (n_2165, n_79, n_141);
  nand g60 (n_2160, n_79, n_141);
  nor g61 (n_2161, n_78, n_140);
  nand g62 (n_2162, n_78, n_140);
  nor g63 (n_2171, n_77, n_139);
  nand g64 (n_2166, n_77, n_139);
  nor g65 (n_2167, n_76, n_138);
  nand g66 (n_2168, n_76, n_138);
  nor g67 (n_2177, n_75, n_137);
  nand g68 (n_2172, n_75, n_137);
  nor g69 (n_2173, n_74, n_136);
  nand g70 (n_2174, n_74, n_136);
  nor g71 (n_2183, n_73, n_135);
  nand g72 (n_2178, n_73, n_135);
  nor g73 (n_2179, n_72, n_134);
  nand g74 (n_2180, n_72, n_134);
  nor g75 (n_2189, n_71, n_133);
  nand g76 (n_2184, n_71, n_133);
  nor g77 (n_2185, n_70, n_132);
  nand g78 (n_2186, n_70, n_132);
  nor g79 (n_2195, n_69, n_131);
  nand g80 (n_2190, n_69, n_131);
  nor g81 (n_2191, n_68, n_130);
  nand g82 (n_2192, n_68, n_130);
  nor g83 (n_2201, n_67, n_129);
  nand g84 (n_2196, n_67, n_129);
  nor g85 (n_2197, n_66, n_128);
  nand g86 (n_2198, n_66, n_128);
  nor g87 (n_2207, n_65, n_127);
  nand g88 (n_2202, n_65, n_127);
  nor g89 (n_2203, n_64, n_126);
  nand g90 (n_2204, n_64, n_126);
  nor g91 (n_2213, n_63, n_125);
  nand g92 (n_2208, n_63, n_125);
  nor g93 (n_2209, n_62, n_124);
  nand g94 (n_2210, n_62, n_124);
  nor g95 (n_2219, n_61, n_123);
  nand g96 (n_2214, n_61, n_123);
  nor g97 (n_2215, n_60, n_122);
  nand g98 (n_2216, n_60, n_122);
  nor g99 (n_2225, n_59, n_121);
  nand g100 (n_2220, n_59, n_121);
  nor g101 (n_2221, n_58, n_120);
  nand g102 (n_2222, n_58, n_120);
  nor g103 (n_2231, n_57, n_119);
  nand g104 (n_2226, n_57, n_119);
  nor g105 (n_2227, n_56, n_118);
  nand g106 (n_2228, n_56, n_118);
  nor g107 (n_2237, n_55, n_117);
  nand g108 (n_2232, n_55, n_117);
  nor g109 (n_2233, n_54, n_116);
  nand g110 (n_2234, n_54, n_116);
  nor g111 (n_2243, n_53, n_115);
  nand g112 (n_2238, n_53, n_115);
  nor g113 (n_2239, n_52, n_114);
  nand g114 (n_2240, n_52, n_114);
  nor g115 (n_2249, n_51, n_113);
  nand g116 (n_2244, n_51, n_113);
  nor g117 (n_2245, n_50, n_112);
  nand g118 (n_2246, n_50, n_112);
  nor g119 (n_2255, n_49, n_111);
  nand g120 (n_2250, n_49, n_111);
  nor g121 (n_2251, n_48, n_110);
  nand g122 (n_2252, n_48, n_110);
  nor g123 (n_2261, n_47, n_109);
  nand g124 (n_2256, n_47, n_109);
  nor g134 (n_2091, n_803, n_2089);
  nor g138 (n_2097, n_2094, n_2095);
  nor g141 (n_2275, n_2099, n_2095);
  nor g142 (n_2103, n_2100, n_2101);
  nor g145 (n_2277, n_2105, n_2101);
  nor g146 (n_2109, n_2106, n_2107);
  nor g149 (n_2285, n_2111, n_2107);
  nor g150 (n_2115, n_2112, n_2113);
  nor g153 (n_2287, n_2117, n_2113);
  nor g154 (n_2121, n_2118, n_2119);
  nor g157 (n_2295, n_2123, n_2119);
  nor g158 (n_2127, n_2124, n_2125);
  nor g161 (n_2297, n_2129, n_2125);
  nor g162 (n_2133, n_2130, n_2131);
  nor g165 (n_2305, n_2135, n_2131);
  nor g166 (n_2139, n_2136, n_2137);
  nor g169 (n_2307, n_2141, n_2137);
  nor g170 (n_2145, n_2142, n_2143);
  nor g173 (n_2315, n_2147, n_2143);
  nor g174 (n_2151, n_2148, n_2149);
  nor g177 (n_2317, n_2153, n_2149);
  nor g178 (n_2157, n_2154, n_2155);
  nor g181 (n_2325, n_2159, n_2155);
  nor g182 (n_2163, n_2160, n_2161);
  nor g185 (n_2327, n_2165, n_2161);
  nor g186 (n_2169, n_2166, n_2167);
  nor g189 (n_2335, n_2171, n_2167);
  nor g190 (n_2175, n_2172, n_2173);
  nor g193 (n_2337, n_2177, n_2173);
  nor g194 (n_2181, n_2178, n_2179);
  nor g197 (n_2345, n_2183, n_2179);
  nor g198 (n_2187, n_2184, n_2185);
  nor g201 (n_2347, n_2189, n_2185);
  nor g202 (n_2193, n_2190, n_2191);
  nor g205 (n_2355, n_2195, n_2191);
  nor g206 (n_2199, n_2196, n_2197);
  nor g209 (n_2357, n_2201, n_2197);
  nor g210 (n_2205, n_2202, n_2203);
  nor g213 (n_2365, n_2207, n_2203);
  nor g214 (n_2211, n_2208, n_2209);
  nor g217 (n_2367, n_2213, n_2209);
  nor g218 (n_2217, n_2214, n_2215);
  nor g221 (n_2375, n_2219, n_2215);
  nor g222 (n_2223, n_2220, n_2221);
  nor g225 (n_2377, n_2225, n_2221);
  nor g226 (n_2229, n_2226, n_2227);
  nor g229 (n_2385, n_2231, n_2227);
  nor g230 (n_2235, n_2232, n_2233);
  nor g233 (n_2387, n_2237, n_2233);
  nor g234 (n_2241, n_2238, n_2239);
  nor g237 (n_2395, n_2243, n_2239);
  nor g238 (n_2247, n_2244, n_2245);
  nor g241 (n_2397, n_2249, n_2245);
  nor g242 (n_2253, n_2250, n_2251);
  nor g245 (n_2405, n_2255, n_2251);
  nor g246 (n_2259, n_2256, n_2257);
  nor g249 (n_2407, n_2261, n_2257);
  nor g259 (n_2273, n_2105, n_2272);
  nand g268 (n_2420, n_2275, n_2277);
  nor g269 (n_2283, n_2117, n_2282);
  nand g278 (n_2427, n_2285, n_2287);
  nor g279 (n_2293, n_2129, n_2292);
  nand g288 (n_2435, n_2295, n_2297);
  nor g289 (n_2303, n_2141, n_2302);
  nand g298 (n_2442, n_2305, n_2307);
  nor g299 (n_2313, n_2153, n_2312);
  nand g308 (n_2450, n_2315, n_2317);
  nor g309 (n_2323, n_2165, n_2322);
  nand g318 (n_2457, n_2325, n_2327);
  nor g319 (n_2333, n_2177, n_2332);
  nand g328 (n_2465, n_2335, n_2337);
  nor g329 (n_2343, n_2189, n_2342);
  nand g338 (n_2472, n_2345, n_2347);
  nor g339 (n_2353, n_2201, n_2352);
  nand g2304 (n_2480, n_2355, n_2357);
  nor g2305 (n_2363, n_2213, n_2362);
  nand g2314 (n_2487, n_2365, n_2367);
  nor g2315 (n_2373, n_2225, n_2372);
  nand g2324 (n_2495, n_2375, n_2377);
  nor g2325 (n_2383, n_2237, n_2382);
  nand g2334 (n_2502, n_2385, n_2387);
  nor g2335 (n_2393, n_2249, n_2392);
  nand g2344 (n_2510, n_2395, n_2397);
  nor g2345 (n_2403, n_2261, n_2402);
  nand g2354 (n_2517, n_2405, n_2407);
  nand g2357 (n_2832, n_2094, n_2414);
  nand g2359 (n_2834, n_2272, n_2415);
  nand g2362 (n_2837, n_2418, n_2419);
  nand g2365 (n_2518, n_2422, n_2423);
  nor g2366 (n_2425, n_2123, n_2424);
  nor g2369 (n_2528, n_2123, n_2427);
  nor g2375 (n_2433, n_2431, n_2424);
  nor g2378 (n_2534, n_2427, n_2431);
  nor g2379 (n_2437, n_2435, n_2424);
  nor g2382 (n_2537, n_2427, n_2435);
  nor g2383 (n_2440, n_2147, n_2439);
  nor g2386 (n_2643, n_2147, n_2442);
  nor g2392 (n_2448, n_2446, n_2439);
  nor g2395 (n_2649, n_2442, n_2446);
  nor g2396 (n_2452, n_2450, n_2439);
  nor g2399 (n_2543, n_2442, n_2450);
  nor g2400 (n_2455, n_2171, n_2454);
  nor g2403 (n_2556, n_2171, n_2457);
  nor g2409 (n_2463, n_2461, n_2454);
  nor g2412 (n_2566, n_2457, n_2461);
  nor g2413 (n_2467, n_2465, n_2454);
  nor g2416 (n_2571, n_2457, n_2465);
  nor g2417 (n_2470, n_2195, n_2469);
  nor g2420 (n_2746, n_2195, n_2472);
  nor g2426 (n_2478, n_2476, n_2469);
  nor g2429 (n_2752, n_2472, n_2476);
  nor g2430 (n_2482, n_2480, n_2469);
  nor g2433 (n_2579, n_2472, n_2480);
  nor g2434 (n_2485, n_2219, n_2484);
  nor g2437 (n_2592, n_2219, n_2487);
  nor g2443 (n_2493, n_2491, n_2484);
  nor g2446 (n_2602, n_2487, n_2491);
  nor g2447 (n_2497, n_2495, n_2484);
  nor g2450 (n_2607, n_2487, n_2495);
  nor g2451 (n_2500, n_2243, n_2499);
  nor g2454 (n_2698, n_2243, n_2502);
  nor g2460 (n_2508, n_2506, n_2499);
  nor g2463 (n_2708, n_2502, n_2506);
  nor g2464 (n_2512, n_2510, n_2499);
  nor g2467 (n_2615, n_2502, n_2510);
  nor g2468 (n_2515, n_2265, n_2514);
  nor g2471 (n_2628, n_2265, n_2517);
  nand g2474 (n_2841, n_2106, n_2520);
  nand g2475 (n_2521, n_2285, n_2518);
  nand g2476 (n_2843, n_2282, n_2521);
  nand g2479 (n_2846, n_2524, n_2525);
  nand g2482 (n_2849, n_2424, n_2527);
  nand g2483 (n_2530, n_2528, n_2518);
  nand g2484 (n_2852, n_2529, n_2530);
  nand g2485 (n_2533, n_2531, n_2518);
  nand g2486 (n_2854, n_2532, n_2533);
  nand g2487 (n_2536, n_2534, n_2518);
  nand g2488 (n_2857, n_2535, n_2536);
  nand g2489 (n_2539, n_2537, n_2518);
  nand g2490 (n_2633, n_2538, n_2539);
  nor g2491 (n_2541, n_2159, n_2540);
  nand g2500 (n_2657, n_2325, n_2543);
  nor g2501 (n_2550, n_2548, n_2540);
  nor g2506 (n_2553, n_2457, n_2540);
  nand g2515 (n_2669, n_2543, n_2556);
  nand g2520 (n_2673, n_2543, n_2561);
  nand g2525 (n_2677, n_2543, n_2566);
  nand g2530 (n_2681, n_2543, n_2571);
  nor g2531 (n_2577, n_2207, n_2576);
  nand g2540 (n_2760, n_2365, n_2579);
  nor g2541 (n_2586, n_2584, n_2576);
  nor g2546 (n_2589, n_2487, n_2576);
  nand g2555 (n_2772, n_2579, n_2592);
  nand g2560 (n_2776, n_2579, n_2597);
  nand g2565 (n_2780, n_2579, n_2602);
  nand g2570 (n_2688, n_2579, n_2607);
  nor g2571 (n_2613, n_2255, n_2612);
  nand g2580 (n_2720, n_2405, n_2615);
  nor g2581 (n_2622, n_2620, n_2612);
  nor g2586 (n_2625, n_2517, n_2612);
  nand g2595 (n_2732, n_2615, n_2628);
  nand g2598 (n_2861, n_2130, n_2635);
  nand g2599 (n_2636, n_2305, n_2633);
  nand g2600 (n_2863, n_2302, n_2636);
  nand g2603 (n_2866, n_2639, n_2640);
  nand g2606 (n_2869, n_2439, n_2642);
  nand g2607 (n_2645, n_2643, n_2633);
  nand g2608 (n_2872, n_2644, n_2645);
  nand g2609 (n_2648, n_2646, n_2633);
  nand g2610 (n_2874, n_2647, n_2648);
  nand g2611 (n_2651, n_2649, n_2633);
  nand g2612 (n_2877, n_2650, n_2651);
  nand g2613 (n_2652, n_2543, n_2633);
  nand g2614 (n_2879, n_2540, n_2652);
  nand g2617 (n_2882, n_2655, n_2656);
  nand g2620 (n_2884, n_2659, n_2660);
  nand g2623 (n_2887, n_2663, n_2664);
  nand g2626 (n_2890, n_2667, n_2668);
  nand g2629 (n_2893, n_2671, n_2672);
  nand g2632 (n_2895, n_2675, n_2676);
  nand g2635 (n_2898, n_2679, n_2680);
  nand g2638 (n_2736, n_2683, n_2684);
  nor g2639 (n_2686, n_2231, n_2685);
  nor g2642 (n_2786, n_2231, n_2688);
  nor g2648 (n_2694, n_2692, n_2685);
  nor g2651 (n_2792, n_2692, n_2688);
  nor g2652 (n_2696, n_2502, n_2685);
  nor g2655 (n_2795, n_2502, n_2688);
  nor g2676 (n_2718, n_2716, n_2685);
  nor g2679 (n_2810, n_2688, n_2716);
  nor g2680 (n_2722, n_2720, n_2685);
  nor g2683 (n_2813, n_2688, n_2720);
  nor g2684 (n_2726, n_2724, n_2685);
  nor g2687 (n_2816, n_2688, n_2724);
  nor g2688 (n_2730, n_2728, n_2685);
  nor g2691 (n_2819, n_2688, n_2728);
  nor g2692 (n_2734, n_2732, n_2685);
  nor g2695 (n_2822, n_2688, n_2732);
  nand g2698 (n_2902, n_2178, n_2738);
  nand g2699 (n_2739, n_2345, n_2736);
  nand g2700 (n_2904, n_2342, n_2739);
  nand g2703 (n_2907, n_2742, n_2743);
  nand g2706 (n_2910, n_2469, n_2745);
  nand g2707 (n_2748, n_2746, n_2736);
  nand g2708 (n_2913, n_2747, n_2748);
  nand g2709 (n_2751, n_2749, n_2736);
  nand g2710 (n_2915, n_2750, n_2751);
  nand g2711 (n_2754, n_2752, n_2736);
  nand g2712 (n_2918, n_2753, n_2754);
  nand g2713 (n_2755, n_2579, n_2736);
  nand g2714 (n_2920, n_2576, n_2755);
  nand g2717 (n_2923, n_2758, n_2759);
  nand g2720 (n_2925, n_2762, n_2763);
  nand g2723 (n_2928, n_2766, n_2767);
  nand g2726 (n_2931, n_2770, n_2771);
  nand g2729 (n_2934, n_2774, n_2775);
  nand g2732 (n_2936, n_2778, n_2779);
  nand g2735 (n_2939, n_2782, n_2783);
  nand g2738 (n_2942, n_2685, n_2785);
  nand g2739 (n_2788, n_2786, n_2736);
  nand g2740 (n_2945, n_2787, n_2788);
  nand g2741 (n_2791, n_2789, n_2736);
  nand g2742 (n_2947, n_2790, n_2791);
  nand g2743 (n_2794, n_2792, n_2736);
  nand g2744 (n_2950, n_2793, n_2794);
  nand g2745 (n_2797, n_2795, n_2736);
  nand g2746 (n_2953, n_2796, n_2797);
  nand g2747 (n_2800, n_2798, n_2736);
  nand g2748 (n_2956, n_2799, n_2800);
  nand g2749 (n_2803, n_2801, n_2736);
  nand g2750 (n_2958, n_2802, n_2803);
  nand g2751 (n_2806, n_2804, n_2736);
  nand g2752 (n_2961, n_2805, n_2806);
  nand g2753 (n_2809, n_2807, n_2736);
  nand g2754 (n_2963, n_2808, n_2809);
  nand g2755 (n_2812, n_2810, n_2736);
  nand g2756 (n_2966, n_2811, n_2812);
  nand g2757 (n_2815, n_2813, n_2736);
  nand g2758 (n_2968, n_2814, n_2815);
  nand g2759 (n_2818, n_2816, n_2736);
  nand g2760 (n_2971, n_2817, n_2818);
  nand g2761 (n_2821, n_2819, n_2736);
  nand g2762 (n_2974, n_2820, n_2821);
  nand g2763 (n_2824, n_2822, n_2736);
  nand g2764 (n_2977, n_2823, n_2824);
  xnor g2776 (Z[5], n_2832, n_2833);
  xnor g2778 (Z[6], n_2834, n_2835);
  xnor g2781 (Z[7], n_2837, n_2838);
  xnor g2783 (Z[8], n_2518, n_2839);
  xnor g2786 (Z[9], n_2841, n_2842);
  xnor g2788 (Z[10], n_2843, n_2844);
  xnor g2791 (Z[11], n_2846, n_2847);
  xnor g2794 (Z[12], n_2849, n_2850);
  xnor g2797 (Z[13], n_2852, n_2853);
  xnor g2799 (Z[14], n_2854, n_2855);
  xnor g2802 (Z[15], n_2857, n_2858);
  xnor g2804 (Z[16], n_2633, n_2859);
  xnor g2807 (Z[17], n_2861, n_2862);
  xnor g2809 (Z[18], n_2863, n_2864);
  xnor g2812 (Z[19], n_2866, n_2867);
  xnor g2815 (Z[20], n_2869, n_2870);
  xnor g2818 (Z[21], n_2872, n_2873);
  xnor g2820 (Z[22], n_2874, n_2875);
  xnor g2823 (Z[23], n_2877, n_2878);
  xnor g2825 (Z[24], n_2879, n_2880);
  xnor g2828 (Z[25], n_2882, n_2883);
  xnor g2830 (Z[26], n_2884, n_2885);
  xnor g2833 (Z[27], n_2887, n_2888);
  xnor g2836 (Z[28], n_2890, n_2891);
  xnor g2839 (Z[29], n_2893, n_2894);
  xnor g2841 (Z[30], n_2895, n_2896);
  xnor g2844 (Z[31], n_2898, n_2899);
  xnor g2846 (Z[32], n_2736, n_2900);
  xnor g2849 (Z[33], n_2902, n_2903);
  xnor g2851 (Z[34], n_2904, n_2905);
  xnor g2854 (Z[35], n_2907, n_2908);
  xnor g2857 (Z[36], n_2910, n_2911);
  xnor g2860 (Z[37], n_2913, n_2914);
  xnor g2862 (Z[38], n_2915, n_2916);
  xnor g2865 (Z[39], n_2918, n_2919);
  xnor g2867 (Z[40], n_2920, n_2921);
  xnor g2870 (Z[41], n_2923, n_2924);
  xnor g2872 (Z[42], n_2925, n_2926);
  xnor g2875 (Z[43], n_2928, n_2929);
  xnor g2878 (Z[44], n_2931, n_2932);
  xnor g2881 (Z[45], n_2934, n_2935);
  xnor g2883 (Z[46], n_2936, n_2937);
  xnor g2886 (Z[47], n_2939, n_2940);
  xnor g2889 (Z[48], n_2942, n_2943);
  xnor g2892 (Z[49], n_2945, n_2946);
  xnor g2894 (Z[50], n_2947, n_2948);
  xnor g2897 (Z[51], n_2950, n_2951);
  xnor g2900 (Z[52], n_2953, n_2954);
  xnor g2903 (Z[53], n_2956, n_2957);
  xnor g2905 (Z[54], n_2958, n_2959);
  xnor g2908 (Z[55], n_2961, n_2962);
  xnor g2910 (Z[56], n_2963, n_2964);
  xnor g2913 (Z[57], n_2966, n_2967);
  xnor g2915 (Z[58], n_2968, n_2969);
  xnor g2918 (Z[59], n_2971, n_2972);
  xnor g2921 (Z[60], n_2974, n_2975);
  or g2938 (n_238, wc, wc0, n_100);
  not gc0 (wc0, n_803);
  not gc (wc, n_817);
  or g2939 (n_247, wc1, wc2, n_232);
  not gc2 (wc2, n_817);
  not gc1 (wc1, n_836);
  or g2940 (n_260, wc3, n_237, n_232);
  not gc3 (wc3, n_864);
  or g2941 (n_277, wc4, wc5, n_237);
  not gc5 (wc5, n_899);
  not gc4 (wc4, n_900);
  or g2942 (n_299, wc6, wc7, n_237);
  not gc7 (wc7, n_947);
  not gc6 (wc6, n_948);
  or g2943 (n_346, wc8, wc9, n_232);
  not gc9 (wc9, n_948);
  not gc8 (wc8, n_995);
  or g2944 (n_372, wc10, wc11, n_237);
  not gc11 (wc11, n_1124);
  not gc10 (wc10, n_1125);
  or g2945 (n_400, wc12, wc13, n_246);
  not gc13 (wc13, n_1064);
  not gc12 (wc12, n_1188);
  or g2946 (n_428, wc14, wc15, n_259);
  not gc15 (wc15, n_1128);
  not gc14 (wc14, n_1252);
  or g2947 (n_456, wc16, wc17, n_276);
  not gc17 (wc17, n_1057);
  not gc16 (wc16, n_1316);
  or g2948 (n_484, wc18, wc19, n_297);
  not gc19 (wc19, n_1121);
  not gc18 (wc18, n_1380);
  or g2949 (n_513, wc20, wc21, n_297);
  not gc21 (wc21, n_1443);
  not gc20 (wc20, n_1444);
  or g2950 (n_540, wc22, wc23, n_317);
  not gc23 (wc23, n_1440);
  not gc22 (wc22, n_1508);
  xnor g2951 (n_1822, A[42], A[40]);
  or g2952 (n_1823, wc24, A[42]);
  not gc24 (wc24, A[40]);
  or g2953 (n_1825, wc25, A[42]);
  not gc25 (wc25, A[28]);
  xnor g2954 (n_1862, A[37], A[35]);
  or g2955 (n_1863, A[35], wc26);
  not gc26 (wc26, A[37]);
  or g2956 (n_1828, wc27, A[42]);
  not gc27 (wc27, A[30]);
  xnor g2957 (n_741, n_1962, A[35]);
  or g2958 (n_1965, wc28, A[35]);
  not gc28 (wc28, A[33]);
  or g2959 (n_1981, wc29, A[42]);
  not gc29 (wc29, A[36]);
  xnor g2960 (n_788, n_2054, A[41]);
  or g2961 (n_2056, wc30, A[41]);
  not gc30 (wc30, A[37]);
  or g2962 (n_2057, wc31, A[41]);
  not gc31 (wc31, A[39]);
  or g2963 (n_2065, wc32, A[42]);
  not gc32 (wc32, A[38]);
  or g2965 (n_2071, A[39], wc33);
  not gc33 (wc33, A[41]);
  or g2966 (n_2077, wc34, A[42]);
  not gc34 (wc34, A[39]);
  and g2967 (n_2265, wc35, A[42]);
  not gc35 (wc35, A[41]);
  or g2968 (n_2262, wc36, A[42]);
  not gc36 (wc36, A[41]);
  or g2969 (n_323, wc37, wc38, n_237);
  not gc38 (wc38, n_1004);
  not gc37 (wc37, n_1005);
  or g2970 (n_1921, A[35], wc39);
  not gc39 (wc39, n_716);
  or g2971 (n_2004, A[35], wc40);
  not gc40 (wc40, n_626);
  and g2972 (n_2270, wc41, n_800);
  not gc41 (wc41, n_2091);
  or g2974 (n_2826, n_2093, wc42);
  not gc42 (wc42, n_803);
  or g2975 (n_2829, n_2089, wc43);
  not gc43 (wc43, n_800);
  xnor g2976 (n_1826, A[42], A[26]);
  or g2977 (n_1827, wc44, A[42]);
  not gc44 (wc44, A[26]);
  or g2978 (n_1864, A[35], wc45);
  not gc45 (wc45, n_687);
  xnor g2979 (n_1918, n_687, A[35]);
  xnor g2980 (n_2034, n_760, A[35]);
  or g2981 (n_2035, A[35], wc46);
  not gc46 (wc46, n_760);
  or g2982 (n_2037, A[35], wc47);
  not gc47 (wc47, n_776);
  xnor g2983 (n_48, n_1734, n_795);
  or g2984 (n_2072, A[39], wc48);
  not gc48 (wc48, n_795);
  and g2985 (n_2257, A[41], wc49);
  not gc49 (wc49, n_108);
  or g2986 (n_2258, A[41], wc50);
  not gc50 (wc50, n_108);
  or g2987 (n_2830, wc51, n_2099);
  not gc51 (wc51, n_2094);
  or g2988 (n_2975, wc52, n_2265);
  not gc52 (wc52, n_2262);
  and g2989 (n_2272, wc53, n_2096);
  not gc53 (wc53, n_2097);
  or g2990 (n_2416, wc54, n_2105);
  not gc54 (wc54, n_2275);
  not g2991 (Z[2], n_2826);
  or g2992 (n_2833, wc55, n_2095);
  not gc55 (wc55, n_2096);
  or g2993 (n_2835, wc56, n_2105);
  not gc56 (wc56, n_2100);
  and g2994 (n_2279, wc57, n_2102);
  not gc57 (wc57, n_2103);
  or g2997 (n_2838, wc58, n_2101);
  not gc58 (wc58, n_2102);
  or g2998 (n_2972, wc59, n_2257);
  not gc59 (wc59, n_2258);
  and g2999 (n_2282, wc60, n_2108);
  not gc60 (wc60, n_2109);
  and g3000 (n_2418, wc61, n_2100);
  not gc61 (wc61, n_2273);
  and g3001 (n_2280, wc62, n_2277);
  not gc62 (wc62, n_2272);
  or g3002 (n_2414, n_2099, n_2270);
  or g3003 (n_2415, n_2270, wc63);
  not gc63 (wc63, n_2275);
  or g3004 (n_2419, n_2270, n_2416);
  xor g3005 (Z[3], n_803, n_2829);
  xor g3006 (Z[4], n_2270, n_2830);
  or g3007 (n_2839, wc64, n_2111);
  not gc64 (wc64, n_2106);
  or g3008 (n_2842, wc65, n_2107);
  not gc65 (wc65, n_2108);
  and g3009 (n_2409, n_2258, wc66);
  not gc66 (wc66, n_2259);
  and g3010 (n_2422, wc67, n_2279);
  not gc67 (wc67, n_2280);
  or g3011 (n_2522, wc68, n_2117);
  not gc68 (wc68, n_2285);
  or g3012 (n_2423, n_2420, n_2270);
  or g3013 (n_2844, wc69, n_2117);
  not gc69 (wc69, n_2112);
  or g3014 (n_2967, wc70, n_2251);
  not gc70 (wc70, n_2252);
  or g3015 (n_2969, wc71, n_2261);
  not gc71 (wc71, n_2256);
  and g3016 (n_2289, wc72, n_2114);
  not gc72 (wc72, n_2115);
  and g3017 (n_2292, wc73, n_2120);
  not gc73 (wc73, n_2121);
  and g3018 (n_2524, wc74, n_2112);
  not gc74 (wc74, n_2283);
  or g3019 (n_2847, wc75, n_2113);
  not gc75 (wc75, n_2114);
  or g3020 (n_2850, wc76, n_2123);
  not gc76 (wc76, n_2118);
  or g3021 (n_2853, wc77, n_2119);
  not gc77 (wc77, n_2120);
  and g3022 (n_2299, wc78, n_2126);
  not gc78 (wc78, n_2127);
  and g3023 (n_2399, wc79, n_2246);
  not gc79 (wc79, n_2247);
  and g3024 (n_2402, wc80, n_2252);
  not gc80 (wc80, n_2253);
  and g3025 (n_2290, wc81, n_2287);
  not gc81 (wc81, n_2282);
  or g3026 (n_2431, wc82, n_2129);
  not gc82 (wc82, n_2295);
  or g3027 (n_2620, wc83, n_2261);
  not gc83 (wc83, n_2405);
  and g3028 (n_2531, wc84, n_2295);
  not gc84 (wc84, n_2427);
  or g3029 (n_2520, wc85, n_2111);
  not gc85 (wc85, n_2518);
  or g3030 (n_2525, n_2522, wc86);
  not gc86 (wc86, n_2518);
  or g3031 (n_2855, wc87, n_2129);
  not gc87 (wc87, n_2124);
  or g3032 (n_2858, wc88, n_2125);
  not gc88 (wc88, n_2126);
  or g3033 (n_2959, wc89, n_2249);
  not gc89 (wc89, n_2244);
  or g3034 (n_2962, wc90, n_2245);
  not gc90 (wc90, n_2246);
  or g3035 (n_2964, wc91, n_2255);
  not gc91 (wc91, n_2250);
  and g3036 (n_2302, wc92, n_2132);
  not gc92 (wc92, n_2133);
  and g3037 (n_2309, wc93, n_2138);
  not gc93 (wc93, n_2139);
  and g3038 (n_2424, wc94, n_2289);
  not gc94 (wc94, n_2290);
  and g3039 (n_2432, wc95, n_2124);
  not gc95 (wc95, n_2293);
  and g3040 (n_2300, wc96, n_2297);
  not gc96 (wc96, n_2292);
  or g3041 (n_2637, wc97, n_2141);
  not gc97 (wc97, n_2305);
  and g3042 (n_2410, wc98, n_2407);
  not gc98 (wc98, n_2402);
  or g3043 (n_2527, wc99, n_2427);
  not gc99 (wc99, n_2518);
  or g3044 (n_2859, wc100, n_2135);
  not gc100 (wc100, n_2130);
  or g3045 (n_2862, wc101, n_2131);
  not gc101 (wc101, n_2132);
  or g3046 (n_2864, wc102, n_2141);
  not gc102 (wc102, n_2136);
  or g3047 (n_2867, wc103, n_2137);
  not gc103 (wc103, n_2138);
  or g3048 (n_2870, wc104, n_2147);
  not gc104 (wc104, n_2142);
  or g3049 (n_2954, wc105, n_2243);
  not gc105 (wc105, n_2238);
  and g3050 (n_2312, wc106, n_2144);
  not gc106 (wc106, n_2145);
  and g3051 (n_2389, wc107, n_2234);
  not gc107 (wc107, n_2235);
  and g3052 (n_2392, wc108, n_2240);
  not gc108 (wc108, n_2241);
  and g3053 (n_2436, wc109, n_2299);
  not gc109 (wc109, n_2300);
  and g3054 (n_2310, wc110, n_2307);
  not gc110 (wc110, n_2302);
  or g3055 (n_2446, wc111, n_2153);
  not gc111 (wc111, n_2315);
  or g3056 (n_2506, wc112, n_2249);
  not gc112 (wc112, n_2395);
  and g3057 (n_2621, wc113, n_2256);
  not gc113 (wc113, n_2403);
  and g3058 (n_2514, wc114, n_2409);
  not gc114 (wc114, n_2410);
  and g3059 (n_2429, wc115, n_2295);
  not gc115 (wc115, n_2424);
  or g3060 (n_2873, wc116, n_2143);
  not gc116 (wc116, n_2144);
  or g3061 (n_2875, wc117, n_2153);
  not gc117 (wc117, n_2148);
  or g3062 (n_2948, wc118, n_2237);
  not gc118 (wc118, n_2232);
  or g3063 (n_2951, wc119, n_2233);
  not gc119 (wc119, n_2234);
  or g3064 (n_2957, wc120, n_2239);
  not gc120 (wc120, n_2240);
  and g3065 (n_2319, wc121, n_2150);
  not gc121 (wc121, n_2151);
  and g3066 (n_2322, wc122, n_2156);
  not gc122 (wc122, n_2157);
  and g3067 (n_2329, wc123, n_2162);
  not gc123 (wc123, n_2163);
  and g3068 (n_2332, wc124, n_2168);
  not gc124 (wc124, n_2169);
  and g3069 (n_2339, wc125, n_2174);
  not gc125 (wc125, n_2175);
  and g3070 (n_2342, wc126, n_2180);
  not gc126 (wc126, n_2181);
  and g3071 (n_2349, wc127, n_2186);
  not gc127 (wc127, n_2187);
  and g3072 (n_2352, wc128, n_2192);
  not gc128 (wc128, n_2193);
  and g3073 (n_2359, wc129, n_2198);
  not gc129 (wc129, n_2199);
  and g3074 (n_2362, wc130, n_2204);
  not gc130 (wc130, n_2205);
  and g3075 (n_2369, wc131, n_2210);
  not gc131 (wc131, n_2211);
  and g3076 (n_2639, wc132, n_2136);
  not gc132 (wc132, n_2303);
  and g3077 (n_2439, wc133, n_2309);
  not gc133 (wc133, n_2310);
  or g3078 (n_2548, wc134, n_2165);
  not gc134 (wc134, n_2325);
  or g3079 (n_2461, wc135, n_2177);
  not gc135 (wc135, n_2335);
  or g3080 (n_2740, wc136, n_2189);
  not gc136 (wc136, n_2345);
  or g3081 (n_2476, wc137, n_2201);
  not gc137 (wc137, n_2355);
  or g3082 (n_2584, wc138, n_2213);
  not gc138 (wc138, n_2365);
  and g3083 (n_2400, wc139, n_2397);
  not gc139 (wc139, n_2392);
  and g3084 (n_2529, wc140, n_2118);
  not gc140 (wc140, n_2425);
  and g3085 (n_2532, wc141, n_2292);
  not gc141 (wc141, n_2429);
  and g3086 (n_2535, n_2432, wc142);
  not gc142 (wc142, n_2433);
  and g3087 (n_2646, wc143, n_2315);
  not gc143 (wc143, n_2442);
  or g3088 (n_2878, wc144, n_2149);
  not gc144 (wc144, n_2150);
  or g3089 (n_2880, wc145, n_2159);
  not gc145 (wc145, n_2154);
  or g3090 (n_2883, wc146, n_2155);
  not gc146 (wc146, n_2156);
  or g3091 (n_2885, wc147, n_2165);
  not gc147 (wc147, n_2160);
  or g3092 (n_2888, wc148, n_2161);
  not gc148 (wc148, n_2162);
  or g3093 (n_2891, wc149, n_2171);
  not gc149 (wc149, n_2166);
  or g3094 (n_2894, wc150, n_2167);
  not gc150 (wc150, n_2168);
  or g3095 (n_2896, wc151, n_2177);
  not gc151 (wc151, n_2172);
  or g3096 (n_2899, wc152, n_2173);
  not gc152 (wc152, n_2174);
  or g3097 (n_2900, wc153, n_2183);
  not gc153 (wc153, n_2178);
  or g3098 (n_2903, wc154, n_2179);
  not gc154 (wc154, n_2180);
  or g3099 (n_2905, wc155, n_2189);
  not gc155 (wc155, n_2184);
  or g3100 (n_2908, wc156, n_2185);
  not gc156 (wc156, n_2186);
  or g3101 (n_2911, wc157, n_2195);
  not gc157 (wc157, n_2190);
  or g3102 (n_2914, wc158, n_2191);
  not gc158 (wc158, n_2192);
  or g3103 (n_2916, wc159, n_2201);
  not gc159 (wc159, n_2196);
  or g3104 (n_2919, wc160, n_2197);
  not gc160 (wc160, n_2198);
  or g3105 (n_2921, wc161, n_2207);
  not gc161 (wc161, n_2202);
  or g3106 (n_2924, wc162, n_2203);
  not gc162 (wc162, n_2204);
  or g3107 (n_2926, wc163, n_2213);
  not gc163 (wc163, n_2208);
  or g3108 (n_2929, wc164, n_2209);
  not gc164 (wc164, n_2210);
  and g3109 (n_2372, wc165, n_2216);
  not gc165 (wc165, n_2217);
  and g3110 (n_2382, wc166, n_2228);
  not gc166 (wc166, n_2229);
  and g3111 (n_2447, wc167, n_2148);
  not gc167 (wc167, n_2313);
  and g3112 (n_2320, wc168, n_2317);
  not gc168 (wc168, n_2312);
  and g3113 (n_2330, wc169, n_2327);
  not gc169 (wc169, n_2322);
  and g3114 (n_2340, wc170, n_2337);
  not gc170 (wc170, n_2332);
  and g3115 (n_2350, wc171, n_2347);
  not gc171 (wc171, n_2342);
  and g3116 (n_2360, wc172, n_2357);
  not gc172 (wc172, n_2352);
  and g3117 (n_2370, wc173, n_2367);
  not gc173 (wc173, n_2362);
  or g3118 (n_2692, wc174, n_2237);
  not gc174 (wc174, n_2385);
  and g3119 (n_2507, wc175, n_2244);
  not gc175 (wc175, n_2393);
  and g3120 (n_2511, wc176, n_2399);
  not gc176 (wc176, n_2400);
  and g3121 (n_2538, n_2436, wc177);
  not gc177 (wc177, n_2437);
  and g3122 (n_2444, wc178, n_2315);
  not gc178 (wc178, n_2439);
  and g3123 (n_2561, wc179, n_2335);
  not gc179 (wc179, n_2457);
  and g3124 (n_2749, wc180, n_2355);
  not gc180 (wc180, n_2472);
  and g3125 (n_2630, n_2262, wc181);
  not gc181 (wc181, n_2515);
  or g3126 (n_2932, wc182, n_2219);
  not gc182 (wc182, n_2214);
  or g3127 (n_2935, wc183, n_2215);
  not gc183 (wc183, n_2216);
  or g3128 (n_2943, wc184, n_2231);
  not gc184 (wc184, n_2226);
  or g3129 (n_2946, wc185, n_2227);
  not gc185 (wc185, n_2228);
  and g3130 (n_2379, wc186, n_2222);
  not gc186 (wc186, n_2223);
  and g3131 (n_2451, wc187, n_2319);
  not gc187 (wc187, n_2320);
  and g3132 (n_2549, wc188, n_2160);
  not gc188 (wc188, n_2323);
  and g3133 (n_2454, wc189, n_2329);
  not gc189 (wc189, n_2330);
  and g3134 (n_2462, wc190, n_2172);
  not gc190 (wc190, n_2333);
  and g3135 (n_2466, wc191, n_2339);
  not gc191 (wc191, n_2340);
  and g3136 (n_2742, wc192, n_2184);
  not gc192 (wc192, n_2343);
  and g3137 (n_2469, wc193, n_2349);
  not gc193 (wc193, n_2350);
  and g3138 (n_2477, wc194, n_2196);
  not gc194 (wc194, n_2353);
  and g3139 (n_2481, wc195, n_2359);
  not gc195 (wc195, n_2360);
  and g3140 (n_2585, wc196, n_2208);
  not gc196 (wc196, n_2363);
  and g3141 (n_2484, wc197, n_2369);
  not gc197 (wc197, n_2370);
  or g3142 (n_2491, wc198, n_2225);
  not gc198 (wc198, n_2375);
  and g3143 (n_2390, wc199, n_2387);
  not gc199 (wc199, n_2382);
  and g3144 (n_2644, wc200, n_2142);
  not gc200 (wc200, n_2440);
  and g3145 (n_2647, wc201, n_2312);
  not gc201 (wc201, n_2444);
  and g3146 (n_2597, wc202, n_2375);
  not gc202 (wc202, n_2487);
  and g3147 (n_2703, wc203, n_2395);
  not gc203 (wc203, n_2502);
  or g3148 (n_2653, wc204, n_2159);
  not gc204 (wc204, n_2543);
  or g3149 (n_2661, n_2548, wc205);
  not gc205 (wc205, n_2543);
  or g3150 (n_2665, wc206, n_2457);
  not gc206 (wc206, n_2543);
  or g3151 (n_2756, wc207, n_2207);
  not gc207 (wc207, n_2579);
  or g3152 (n_2764, n_2584, wc208);
  not gc208 (wc208, n_2579);
  or g3153 (n_2768, wc209, n_2487);
  not gc209 (wc209, n_2579);
  or g3154 (n_2937, wc210, n_2225);
  not gc210 (wc210, n_2220);
  or g3155 (n_2940, wc211, n_2221);
  not gc211 (wc211, n_2222);
  and g3156 (n_2492, wc212, n_2220);
  not gc212 (wc212, n_2373);
  and g3157 (n_2380, wc213, n_2377);
  not gc213 (wc213, n_2372);
  and g3158 (n_2693, wc214, n_2232);
  not gc214 (wc214, n_2383);
  and g3159 (n_2499, wc215, n_2389);
  not gc215 (wc215, n_2390);
  and g3160 (n_2650, n_2447, wc216);
  not gc216 (wc216, n_2448);
  and g3161 (n_2459, wc217, n_2335);
  not gc217 (wc217, n_2454);
  and g3162 (n_2474, wc218, n_2355);
  not gc218 (wc218, n_2469);
  and g3163 (n_2489, wc219, n_2375);
  not gc219 (wc219, n_2484);
  or g3164 (n_2716, wc220, n_2255);
  not gc220 (wc220, n_2615);
  or g3165 (n_2724, n_2620, wc221);
  not gc221 (wc221, n_2615);
  or g3166 (n_2728, wc222, n_2517);
  not gc222 (wc222, n_2615);
  or g3167 (n_2635, wc223, n_2135);
  not gc223 (wc223, n_2633);
  or g3168 (n_2640, n_2637, wc224);
  not gc224 (wc224, n_2633);
  or g3169 (n_2642, wc225, n_2442);
  not gc225 (wc225, n_2633);
  and g3170 (n_2496, wc226, n_2379);
  not gc226 (wc226, n_2380);
  and g3171 (n_2540, n_2451, wc227);
  not gc227 (wc227, n_2452);
  and g3172 (n_2558, wc228, n_2166);
  not gc228 (wc228, n_2455);
  and g3173 (n_2563, wc229, n_2332);
  not gc229 (wc229, n_2459);
  and g3174 (n_2568, n_2462, wc230);
  not gc230 (wc230, n_2463);
  and g3175 (n_2573, n_2466, wc231);
  not gc231 (wc231, n_2467);
  and g3176 (n_2747, wc232, n_2190);
  not gc232 (wc232, n_2470);
  and g3177 (n_2750, wc233, n_2352);
  not gc233 (wc233, n_2474);
  and g3178 (n_2753, n_2477, wc234);
  not gc234 (wc234, n_2478);
  and g3179 (n_2576, n_2481, wc235);
  not gc235 (wc235, n_2482);
  and g3180 (n_2594, wc236, n_2214);
  not gc236 (wc236, n_2485);
  and g3181 (n_2599, wc237, n_2372);
  not gc237 (wc237, n_2489);
  and g3182 (n_2504, wc238, n_2395);
  not gc238 (wc238, n_2499);
  or g3183 (n_2656, n_2653, wc239);
  not gc239 (wc239, n_2633);
  or g3184 (n_2660, n_2657, wc240);
  not gc240 (wc240, n_2633);
  or g3185 (n_2664, n_2661, wc241);
  not gc241 (wc241, n_2633);
  or g3186 (n_2668, n_2665, wc242);
  not gc242 (wc242, n_2633);
  or g3187 (n_2672, n_2669, wc243);
  not gc243 (wc243, n_2633);
  or g3188 (n_2676, n_2673, wc244);
  not gc244 (wc244, n_2633);
  or g3189 (n_2680, n_2677, wc245);
  not gc245 (wc245, n_2633);
  or g3190 (n_2684, n_2681, wc246);
  not gc246 (wc246, n_2633);
  and g3191 (n_2604, n_2492, wc247);
  not gc247 (wc247, n_2493);
  and g3192 (n_2700, wc248, n_2238);
  not gc248 (wc248, n_2500);
  and g3193 (n_2705, wc249, n_2392);
  not gc249 (wc249, n_2504);
  and g3194 (n_2710, n_2507, wc250);
  not gc250 (wc250, n_2508);
  and g3195 (n_2612, n_2511, wc251);
  not gc251 (wc251, n_2512);
  and g3196 (n_2546, wc252, n_2325);
  not gc252 (wc252, n_2540);
  and g3197 (n_2559, wc253, n_2556);
  not gc253 (wc253, n_2540);
  and g3198 (n_2564, wc254, n_2561);
  not gc254 (wc254, n_2540);
  and g3199 (n_2569, wc255, n_2566);
  not gc255 (wc255, n_2540);
  and g3200 (n_2574, wc256, n_2571);
  not gc256 (wc256, n_2540);
  and g3201 (n_2582, wc257, n_2365);
  not gc257 (wc257, n_2576);
  and g3202 (n_2595, wc258, n_2592);
  not gc258 (wc258, n_2576);
  and g3203 (n_2600, wc259, n_2597);
  not gc259 (wc259, n_2576);
  and g3204 (n_2605, wc260, n_2602);
  not gc260 (wc260, n_2576);
  and g3205 (n_2610, wc261, n_2607);
  not gc261 (wc261, n_2576);
  and g3206 (n_2789, wc262, n_2385);
  not gc262 (wc262, n_2688);
  and g3207 (n_2798, wc263, n_2698);
  not gc263 (wc263, n_2688);
  and g3208 (n_2801, n_2703, wc264);
  not gc264 (wc264, n_2688);
  and g3209 (n_2804, wc265, n_2708);
  not gc265 (wc265, n_2688);
  and g3210 (n_2807, wc266, n_2615);
  not gc266 (wc266, n_2688);
  and g3211 (n_2609, n_2496, wc267);
  not gc267 (wc267, n_2497);
  and g3212 (n_2655, wc268, n_2154);
  not gc268 (wc268, n_2541);
  and g3213 (n_2659, wc269, n_2322);
  not gc269 (wc269, n_2546);
  and g3214 (n_2663, n_2549, wc270);
  not gc270 (wc270, n_2550);
  and g3215 (n_2667, n_2454, wc271);
  not gc271 (wc271, n_2553);
  and g3216 (n_2671, wc272, n_2558);
  not gc272 (wc272, n_2559);
  and g3217 (n_2675, wc273, n_2563);
  not gc273 (wc273, n_2564);
  and g3218 (n_2679, wc274, n_2568);
  not gc274 (wc274, n_2569);
  and g3219 (n_2683, wc275, n_2573);
  not gc275 (wc275, n_2574);
  and g3220 (n_2758, wc276, n_2202);
  not gc276 (wc276, n_2577);
  and g3221 (n_2762, wc277, n_2362);
  not gc277 (wc277, n_2582);
  and g3222 (n_2766, n_2585, wc278);
  not gc278 (wc278, n_2586);
  and g3223 (n_2770, n_2484, wc279);
  not gc279 (wc279, n_2589);
  and g3224 (n_2774, wc280, n_2594);
  not gc280 (wc280, n_2595);
  and g3225 (n_2778, wc281, n_2599);
  not gc281 (wc281, n_2600);
  and g3226 (n_2618, wc282, n_2405);
  not gc282 (wc282, n_2612);
  and g3227 (n_2631, wc283, n_2628);
  not gc283 (wc283, n_2612);
  and g3228 (n_2782, wc284, n_2604);
  not gc284 (wc284, n_2605);
  and g3229 (n_2717, wc285, n_2250);
  not gc285 (wc285, n_2613);
  and g3230 (n_2721, wc286, n_2402);
  not gc286 (wc286, n_2618);
  and g3231 (n_2725, n_2621, wc287);
  not gc287 (wc287, n_2622);
  and g3232 (n_2729, n_2514, wc288);
  not gc288 (wc288, n_2625);
  and g3233 (n_2733, wc289, n_2630);
  not gc289 (wc289, n_2631);
  and g3234 (n_2685, n_2609, wc290);
  not gc290 (wc290, n_2610);
  or g3235 (n_2738, wc291, n_2183);
  not gc291 (wc291, n_2736);
  or g3236 (n_2743, n_2740, wc292);
  not gc292 (wc292, n_2736);
  or g3237 (n_2745, wc293, n_2472);
  not gc293 (wc293, n_2736);
  or g3238 (n_2759, n_2756, wc294);
  not gc294 (wc294, n_2736);
  or g3239 (n_2763, wc295, n_2760);
  not gc295 (wc295, n_2736);
  or g3240 (n_2767, n_2764, wc296);
  not gc296 (wc296, n_2736);
  or g3241 (n_2771, n_2768, wc297);
  not gc297 (wc297, n_2736);
  or g3242 (n_2775, wc298, n_2772);
  not gc298 (wc298, n_2736);
  or g3243 (n_2779, wc299, n_2776);
  not gc299 (wc299, n_2736);
  or g3244 (n_2783, wc300, n_2780);
  not gc300 (wc300, n_2736);
  or g3245 (n_2785, wc301, n_2688);
  not gc301 (wc301, n_2736);
  and g3246 (n_2690, wc302, n_2385);
  not gc302 (wc302, n_2685);
  and g3247 (n_2701, wc303, n_2698);
  not gc303 (wc303, n_2685);
  and g3248 (n_2706, wc304, n_2703);
  not gc304 (wc304, n_2685);
  and g3249 (n_2711, wc305, n_2708);
  not gc305 (wc305, n_2685);
  and g3250 (n_2714, wc306, n_2615);
  not gc306 (wc306, n_2685);
  and g3251 (n_2787, wc307, n_2226);
  not gc307 (wc307, n_2686);
  and g3252 (n_2790, wc308, n_2382);
  not gc308 (wc308, n_2690);
  and g3253 (n_2793, n_2693, wc309);
  not gc309 (wc309, n_2694);
  and g3254 (n_2796, n_2499, wc310);
  not gc310 (wc310, n_2696);
  and g3255 (n_2799, wc311, n_2700);
  not gc311 (wc311, n_2701);
  and g3256 (n_2802, wc312, n_2705);
  not gc312 (wc312, n_2706);
  and g3257 (n_2805, wc313, n_2710);
  not gc313 (wc313, n_2711);
  and g3258 (n_2808, wc314, n_2612);
  not gc314 (wc314, n_2714);
  and g3259 (n_2811, n_2717, wc315);
  not gc315 (wc315, n_2718);
  and g3260 (n_2814, n_2721, wc316);
  not gc316 (wc316, n_2722);
  and g3261 (n_2817, n_2725, wc317);
  not gc317 (wc317, n_2726);
  and g3262 (n_2820, n_2729, wc318);
  not gc318 (wc318, n_2730);
  and g3263 (n_2823, n_2733, wc319);
  not gc319 (wc319, n_2734);
  not g3264 (Z[61], n_2977);
endmodule

module mult_signed_const_GENERIC(A, Z);
  input [42:0] A;
  output [61:0] Z;
  wire [42:0] A;
  wire [61:0] Z;
  mult_signed_const_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_10350_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [46:0] A;
  output [65:0] Z;
  wire [46:0] A;
  wire [65:0] Z;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_113, n_116, n_117;
  wire n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125;
  wire n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133;
  wire n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_263, n_264, n_265, n_266;
  wire n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395;
  wire n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403;
  wire n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411;
  wire n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419;
  wire n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451;
  wire n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459;
  wire n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467;
  wire n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475;
  wire n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483;
  wire n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491;
  wire n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499;
  wire n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507;
  wire n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515;
  wire n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523;
  wire n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531;
  wire n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539;
  wire n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555;
  wire n_556, n_557, n_558, n_559, n_560, n_561, n_562, n_563;
  wire n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571;
  wire n_572, n_573, n_574, n_575, n_576, n_577, n_578, n_579;
  wire n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587;
  wire n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595;
  wire n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603;
  wire n_604, n_605, n_606, n_607, n_608, n_609, n_610, n_611;
  wire n_612, n_613, n_614, n_615, n_616, n_617, n_618, n_619;
  wire n_620, n_621, n_622, n_623, n_624, n_625, n_626, n_627;
  wire n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635;
  wire n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643;
  wire n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651;
  wire n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_660;
  wire n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668;
  wire n_669, n_670, n_671, n_674, n_675, n_676, n_677, n_678;
  wire n_679, n_680, n_681, n_682, n_683, n_684, n_686, n_687;
  wire n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_695;
  wire n_696, n_697, n_698, n_699, n_700, n_701, n_702, n_703;
  wire n_704, n_705, n_706, n_707, n_708, n_709, n_712, n_713;
  wire n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721;
  wire n_722, n_723, n_724, n_725, n_729, n_730, n_731, n_732;
  wire n_733, n_735, n_736, n_737, n_738, n_739, n_740, n_741;
  wire n_742, n_745, n_746, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_755, n_756, n_757, n_760, n_761, n_762;
  wire n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771;
  wire n_772, n_775, n_776, n_777, n_778, n_779, n_780, n_781;
  wire n_782, n_783, n_784, n_785, n_788, n_789, n_790, n_791;
  wire n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_800;
  wire n_801, n_803, n_804, n_805, n_806, n_807, n_808, n_809;
  wire n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820;
  wire n_822, n_825, n_826, n_827, n_828, n_829, n_835, n_836;
  wire n_837, n_838, n_842, n_843, n_844, n_845, n_849, n_850;
  wire n_851, n_852, n_854, n_856, n_857, n_861, n_862, n_864;
  wire n_865, n_868, n_871, n_872, n_873, n_874, n_875, n_876;
  wire n_877, n_878, n_879, n_880, n_881, n_883, n_884, n_885;
  wire n_886, n_890, n_891, n_892, n_893, n_894, n_895, n_896;
  wire n_897, n_899, n_901, n_902, n_903, n_904, n_905, n_906;
  wire n_907, n_909, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_921, n_923, n_924, n_925, n_926, n_927;
  wire n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_937;
  wire n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948;
  wire n_949, n_950, n_951, n_952, n_955, n_956, n_957, n_959;
  wire n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967;
  wire n_968, n_969, n_970, n_971, n_972, n_973, n_975, n_976;
  wire n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985;
  wire n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993;
  wire n_994, n_995, n_996, n_998, n_999, n_1001, n_1002, n_1003;
  wire n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011;
  wire n_1012, n_1013, n_1014, n_1015, n_1018, n_1019, n_1020, n_1021;
  wire n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030;
  wire n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038;
  wire n_1039, n_1040, n_1041, n_1047, n_1048, n_1051, n_1052, n_1053;
  wire n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061;
  wire n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1070;
  wire n_1071, n_1073, n_1074, n_1077, n_1078, n_1079, n_1080, n_1081;
  wire n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089;
  wire n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097;
  wire n_1101, n_1102, n_1103, n_1104, n_1105, n_1107, n_1108, n_1109;
  wire n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117;
  wire n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125;
  wire n_1126, n_1127, n_1128, n_1129, n_1130, n_1135, n_1136, n_1137;
  wire n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146;
  wire n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154;
  wire n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162;
  wire n_1167, n_1169, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176;
  wire n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184;
  wire n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192;
  wire n_1193, n_1194, n_1197, n_1198, n_1199, n_1200, n_1201, n_1203;
  wire n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211;
  wire n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219;
  wire n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1229;
  wire n_1231, n_1232, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240;
  wire n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248;
  wire n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1257, n_1258, n_1261, n_1263, n_1264, n_1267, n_1268, n_1269;
  wire n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
  wire n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285;
  wire n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1293, n_1295;
  wire n_1296, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305;
  wire n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313;
  wire n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321;
  wire n_1322, n_1325, n_1327, n_1328, n_1331, n_1332, n_1333, n_1334;
  wire n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342;
  wire n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350;
  wire n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1359;
  wire n_1360, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369;
  wire n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377;
  wire n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385;
  wire n_1386, n_1389, n_1391, n_1392, n_1395, n_1396, n_1397, n_1398;
  wire n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406;
  wire n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414;
  wire n_1415, n_1416, n_1417, n_1418, n_1419, n_1421, n_1423, n_1424;
  wire n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434;
  wire n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442;
  wire n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450;
  wire n_1453, n_1455, n_1456, n_1459, n_1460, n_1461, n_1462, n_1463;
  wire n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471;
  wire n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479;
  wire n_1480, n_1481, n_1482, n_1483, n_1485, n_1487, n_1488, n_1491;
  wire n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499;
  wire n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507;
  wire n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1517;
  wire n_1519, n_1520, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528;
  wire n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536;
  wire n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544;
  wire n_1545, n_1546, n_1547, n_1548, n_1549, n_1551, n_1552, n_1555;
  wire n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563;
  wire n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571;
  wire n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579;
  wire n_1580, n_1581, n_1583, n_1586, n_1587, n_1588, n_1589, n_1590;
  wire n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598;
  wire n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606;
  wire n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1615;
  wire n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625;
  wire n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633;
  wire n_1634, n_1635, n_1636, n_1637, n_1638, n_1642, n_1643, n_1645;
  wire n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656;
  wire n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664;
  wire n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1674, n_1675;
  wire n_1677, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687;
  wire n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695;
  wire n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1706;
  wire n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718;
  wire n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726;
  wire n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734;
  wire n_1738, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749;
  wire n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757;
  wire n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765;
  wire n_1766, n_1767, n_1771, n_1775, n_1776, n_1777, n_1778, n_1779;
  wire n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787;
  wire n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795;
  wire n_1796, n_1797, n_1798, n_1799, n_1803, n_1807, n_1808, n_1809;
  wire n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817;
  wire n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825;
  wire n_1826, n_1827, n_1828, n_1829, n_1830, n_1837, n_1838, n_1843;
  wire n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851;
  wire n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859;
  wire n_1860, n_1861, n_1862, n_1869, n_1870, n_1875, n_1876, n_1877;
  wire n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885;
  wire n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893;
  wire n_1894, n_1899, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906;
  wire n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914;
  wire n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922;
  wire n_1923, n_1924, n_1925, n_1926, n_1931, n_1933, n_1934, n_1935;
  wire n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943;
  wire n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951;
  wire n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959;
  wire n_1960, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1969;
  wire n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978;
  wire n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986;
  wire n_1987, n_1988, n_1989, n_1990, n_1995, n_1997, n_1998, n_2003;
  wire n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011;
  wire n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019;
  wire n_2020, n_2021, n_2022, n_2023, n_2024, n_2026, n_2027, n_2029;
  wire n_2031, n_2032, n_2034, n_2037, n_2038, n_2039, n_2040, n_2041;
  wire n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049;
  wire n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2058;
  wire n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070;
  wire n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078;
  wire n_2079, n_2080, n_2081, n_2082, n_2085, n_2086, n_2087, n_2090;
  wire n_2091, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099;
  wire n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107;
  wire n_2108, n_2109, n_2110, n_2114, n_2115, n_2118, n_2119, n_2120;
  wire n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128;
  wire n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2138;
  wire n_2143, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151;
  wire n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159;
  wire n_2162, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171;
  wire n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2187;
  wire n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195;
  wire n_2196, n_2197, n_2198, n_2205, n_2207, n_2209, n_2210, n_2211;
  wire n_2212, n_2213, n_2214, n_2221, n_2222, n_2223, n_2224, n_2225;
  wire n_2226, n_2227, n_2228, n_2229, n_2230, n_2233, n_2235, n_2236;
  wire n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2247, n_2248;
  wire n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2257;
  wire n_2258, n_2259, n_2260, n_2261, n_2262, n_2265, n_2267, n_2268;
  wire n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2277, n_2278;
  wire n_2290, n_2292, n_2294, n_2295, n_2296, n_2297, n_2298, n_2300;
  wire n_2301, n_2302, n_2303, n_2304, n_2306, n_2307, n_2308, n_2309;
  wire n_2310, n_2312, n_2313, n_2314, n_2315, n_2316, n_2318, n_2319;
  wire n_2320, n_2321, n_2322, n_2324, n_2325, n_2326, n_2327, n_2328;
  wire n_2330, n_2331, n_2332, n_2333, n_2334, n_2336, n_2337, n_2338;
  wire n_2339, n_2340, n_2342, n_2343, n_2344, n_2345, n_2346, n_2348;
  wire n_2349, n_2350, n_2351, n_2352, n_2354, n_2355, n_2356, n_2357;
  wire n_2358, n_2360, n_2361, n_2362, n_2363, n_2364, n_2366, n_2367;
  wire n_2368, n_2369, n_2370, n_2372, n_2373, n_2374, n_2375, n_2376;
  wire n_2378, n_2379, n_2380, n_2381, n_2382, n_2384, n_2385, n_2386;
  wire n_2387, n_2388, n_2390, n_2391, n_2392, n_2393, n_2394, n_2396;
  wire n_2397, n_2398, n_2399, n_2400, n_2402, n_2403, n_2404, n_2405;
  wire n_2406, n_2408, n_2409, n_2410, n_2411, n_2412, n_2414, n_2415;
  wire n_2416, n_2417, n_2418, n_2420, n_2421, n_2422, n_2423, n_2424;
  wire n_2426, n_2427, n_2428, n_2429, n_2430, n_2432, n_2433, n_2434;
  wire n_2435, n_2436, n_2438, n_2439, n_2440, n_2441, n_2442, n_2444;
  wire n_2445, n_2446, n_2447, n_2448, n_2450, n_2451, n_2452, n_2453;
  wire n_2454, n_2456, n_2457, n_2458, n_2459, n_2460, n_2462, n_2463;
  wire n_2464, n_2465, n_2466, n_2468, n_2469, n_2470, n_2471, n_2472;
  wire n_2474, n_2475, n_2478, n_2483, n_2485, n_2486, n_2488, n_2490;
  wire n_2492, n_2493, n_2495, n_2496, n_2498, n_2500, n_2502, n_2503;
  wire n_2505, n_2506, n_2508, n_2510, n_2512, n_2513, n_2515, n_2516;
  wire n_2518, n_2520, n_2522, n_2523, n_2525, n_2526, n_2528, n_2530;
  wire n_2532, n_2533, n_2535, n_2536, n_2538, n_2540, n_2542, n_2543;
  wire n_2545, n_2546, n_2548, n_2550, n_2552, n_2553, n_2555, n_2556;
  wire n_2558, n_2560, n_2562, n_2563, n_2565, n_2566, n_2568, n_2570;
  wire n_2572, n_2573, n_2575, n_2576, n_2578, n_2580, n_2582, n_2583;
  wire n_2585, n_2586, n_2588, n_2590, n_2592, n_2593, n_2595, n_2596;
  wire n_2598, n_2600, n_2602, n_2603, n_2605, n_2606, n_2608, n_2610;
  wire n_2612, n_2613, n_2615, n_2616, n_2618, n_2620, n_2622, n_2623;
  wire n_2625, n_2626, n_2628, n_2630, n_2632, n_2633, n_2637, n_2638;
  wire n_2639, n_2641, n_2642, n_2643, n_2645, n_2646, n_2647, n_2648;
  wire n_2650, n_2652, n_2654, n_2655, n_2656, n_2658, n_2659, n_2660;
  wire n_2662, n_2663, n_2665, n_2667, n_2669, n_2670, n_2671, n_2673;
  wire n_2674, n_2675, n_2677, n_2678, n_2680, n_2682, n_2684, n_2685;
  wire n_2686, n_2688, n_2689, n_2690, n_2692, n_2693, n_2695, n_2697;
  wire n_2699, n_2700, n_2701, n_2703, n_2704, n_2705, n_2707, n_2708;
  wire n_2710, n_2712, n_2714, n_2715, n_2716, n_2718, n_2719, n_2720;
  wire n_2722, n_2723, n_2725, n_2727, n_2729, n_2730, n_2731, n_2733;
  wire n_2734, n_2735, n_2737, n_2738, n_2740, n_2742, n_2744, n_2745;
  wire n_2746, n_2748, n_2749, n_2750, n_2752, n_2754, n_2755, n_2756;
  wire n_2758, n_2759, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766;
  wire n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774;
  wire n_2775, n_2777, n_2780, n_2782, n_2783, n_2784, n_2787, n_2790;
  wire n_2792, n_2793, n_2795, n_2797, n_2798, n_2800, n_2802, n_2803;
  wire n_2805, n_2807, n_2808, n_2810, n_2811, n_2813, n_2816, n_2818;
  wire n_2819, n_2820, n_2823, n_2826, n_2828, n_2829, n_2831, n_2833;
  wire n_2834, n_2836, n_2838, n_2839, n_2841, n_2843, n_2844, n_2846;
  wire n_2847, n_2849, n_2852, n_2854, n_2855, n_2856, n_2859, n_2862;
  wire n_2864, n_2865, n_2867, n_2869, n_2870, n_2872, n_2874, n_2875;
  wire n_2877, n_2879, n_2880, n_2882, n_2884, n_2885, n_2886, n_2888;
  wire n_2889, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897;
  wire n_2898, n_2899, n_2900, n_2901, n_2902, n_2904, n_2905, n_2906;
  wire n_2908, n_2909, n_2910, n_2912, n_2913, n_2914, n_2916, n_2917;
  wire n_2918, n_2920, n_2921, n_2922, n_2924, n_2925, n_2926, n_2928;
  wire n_2929, n_2930, n_2932, n_2933, n_2934, n_2935, n_2937, n_2939;
  wire n_2941, n_2942, n_2943, n_2945, n_2947, n_2949, n_2950, n_2952;
  wire n_2954, n_2955, n_2957, n_2959, n_2960, n_2963, n_2965, n_2966;
  wire n_2967, n_2969, n_2970, n_2971, n_2973, n_2974, n_2975, n_2977;
  wire n_2978, n_2979, n_2981, n_2982, n_2983, n_2985, n_2986, n_2987;
  wire n_2989, n_2990, n_2991, n_2993, n_2994, n_2995, n_2997, n_2999;
  wire n_3000, n_3001, n_3003, n_3004, n_3006, n_3007, n_3008, n_3009;
  wire n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017;
  wire n_3019, n_3020, n_3021, n_3023, n_3024, n_3025, n_3027, n_3028;
  wire n_3029, n_3031, n_3032, n_3033, n_3035, n_3036, n_3037, n_3039;
  wire n_3040, n_3041, n_3043, n_3044, n_3046, n_3047, n_3048, n_3049;
  wire n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057;
  wire n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065;
  wire n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073;
  wire n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081;
  wire n_3082, n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089;
  wire n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3097, n_3099;
  wire n_3102, n_3103, n_3105, n_3106, n_3107, n_3108, n_3110, n_3111;
  wire n_3112, n_3114, n_3115, n_3116, n_3117, n_3119, n_3120, n_3122;
  wire n_3123, n_3125, n_3126, n_3127, n_3128, n_3130, n_3131, n_3132;
  wire n_3134, n_3135, n_3136, n_3137, n_3139, n_3140, n_3142, n_3143;
  wire n_3145, n_3146, n_3147, n_3148, n_3150, n_3151, n_3152, n_3153;
  wire n_3155, n_3156, n_3157, n_3158, n_3160, n_3161, n_3163, n_3164;
  wire n_3166, n_3167, n_3168, n_3169, n_3171, n_3172, n_3173, n_3175;
  wire n_3176, n_3177, n_3178, n_3180, n_3181, n_3183, n_3184, n_3186;
  wire n_3187, n_3188, n_3189, n_3191, n_3192, n_3193, n_3194, n_3196;
  wire n_3197, n_3198, n_3199, n_3201, n_3202, n_3204, n_3205, n_3207;
  wire n_3208, n_3209, n_3210, n_3212, n_3213, n_3215, n_3216, n_3218;
  wire n_3219, n_3220, n_3221, n_3223, n_3224, n_3226, n_3227, n_3229;
  wire n_3230, n_3231, n_3232, n_3234, n_3235, n_3236, n_3237, n_3239;
  wire n_3240, n_3241, n_3242, n_3244, n_3245, n_3247, n_3248, n_3250;
  wire n_3251, n_3252, n_3253, n_3255, n_3256, n_3257, n_3259;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g372 (n_175, A[4], A[0]);
  and g2 (n_108, A[4], A[0]);
  xor g373 (n_871, A[1], A[3]);
  xor g374 (n_174, n_871, A[5]);
  nand g3 (n_872, A[1], A[3]);
  nand g375 (n_873, A[5], A[3]);
  nand g376 (n_874, A[1], A[5]);
  nand g377 (n_107, n_872, n_873, n_874);
  xor g378 (n_247, A[6], A[4]);
  and g379 (n_248, A[6], A[4]);
  xor g380 (n_875, A[0], A[2]);
  xor g381 (n_173, n_875, n_247);
  nand g382 (n_876, A[0], A[2]);
  nand g4 (n_877, n_247, A[2]);
  nand g5 (n_878, A[0], n_247);
  nand g383 (n_106, n_876, n_877, n_878);
  xor g384 (n_879, A[1], A[7]);
  xor g385 (n_249, n_879, A[5]);
  nand g386 (n_880, A[1], A[7]);
  nand g387 (n_881, A[5], A[7]);
  nand g6 (n_251, n_880, n_881, n_874);
  xor g389 (n_883, A[3], n_248);
  xor g390 (n_172, n_883, n_249);
  nand g391 (n_884, A[3], n_248);
  nand g392 (n_885, n_249, n_248);
  nand g393 (n_886, A[3], n_249);
  nand g394 (n_105, n_884, n_885, n_886);
  xor g395 (n_250, A[8], A[6]);
  and g396 (n_253, A[8], A[6]);
  xor g398 (n_252, n_875, A[4]);
  nand g401 (n_890, A[2], A[4]);
  xor g403 (n_891, n_250, n_251);
  xor g404 (n_171, n_891, n_252);
  nand g405 (n_892, n_250, n_251);
  nand g406 (n_893, n_252, n_251);
  nand g407 (n_894, n_250, n_252);
  nand g408 (n_104, n_892, n_893, n_894);
  xor g409 (n_895, A[1], A[9]);
  xor g410 (n_255, n_895, A[3]);
  nand g411 (n_896, A[1], A[9]);
  nand g412 (n_897, A[3], A[9]);
  nand g414 (n_258, n_896, n_897, n_872);
  xor g415 (n_899, A[7], A[5]);
  xor g416 (n_256, n_899, n_253);
  nand g418 (n_901, n_253, A[5]);
  nand g419 (n_902, A[7], n_253);
  nand g420 (n_260, n_881, n_901, n_902);
  xor g421 (n_903, n_254, n_255);
  xor g422 (n_170, n_903, n_256);
  nand g423 (n_904, n_254, n_255);
  nand g424 (n_905, n_256, n_255);
  nand g425 (n_906, n_254, n_256);
  nand g426 (n_103, n_904, n_905, n_906);
  xor g427 (n_257, A[10], A[8]);
  and g428 (n_262, A[10], A[8]);
  xor g429 (n_907, A[4], A[2]);
  xor g430 (n_259, n_907, A[6]);
  nand g432 (n_909, A[6], A[2]);
  xor g435 (n_911, A[0], n_257);
  xor g436 (n_261, n_911, n_258);
  nand g437 (n_912, A[0], n_257);
  nand g438 (n_913, n_258, n_257);
  nand g439 (n_914, A[0], n_258);
  nand g440 (n_266, n_912, n_913, n_914);
  xor g441 (n_915, n_259, n_260);
  xor g442 (n_169, n_915, n_261);
  nand g443 (n_916, n_259, n_260);
  nand g444 (n_917, n_261, n_260);
  nand g445 (n_918, n_259, n_261);
  nand g446 (n_102, n_916, n_917, n_918);
  xor g448 (n_264, n_895, A[5]);
  nand g450 (n_921, A[5], A[9]);
  nand g452 (n_269, n_896, n_921, n_874);
  xor g453 (n_923, A[3], A[11]);
  xor g454 (n_265, n_923, A[7]);
  nand g455 (n_924, A[3], A[11]);
  nand g456 (n_925, A[7], A[11]);
  nand g457 (n_926, A[3], A[7]);
  nand g458 (n_270, n_924, n_925, n_926);
  xor g459 (n_927, n_262, n_263);
  xor g460 (n_267, n_927, n_264);
  nand g461 (n_928, n_262, n_263);
  nand g462 (n_929, n_264, n_263);
  nand g463 (n_930, n_262, n_264);
  nand g464 (n_274, n_928, n_929, n_930);
  xor g465 (n_931, n_265, n_266);
  xor g466 (n_168, n_931, n_267);
  nand g467 (n_932, n_265, n_266);
  nand g468 (n_933, n_267, n_266);
  nand g469 (n_934, n_265, n_267);
  nand g470 (n_101, n_932, n_933, n_934);
  xor g471 (n_268, A[12], A[10]);
  and g472 (n_275, A[12], A[10]);
  xor g474 (n_271, n_247, A[8]);
  nand g476 (n_937, A[8], A[4]);
  xor g480 (n_272, n_875, n_268);
  nand g482 (n_941, n_268, A[0]);
  nand g483 (n_942, A[2], n_268);
  nand g484 (n_279, n_876, n_941, n_942);
  xor g485 (n_943, n_269, n_270);
  xor g486 (n_273, n_943, n_271);
  nand g487 (n_944, n_269, n_270);
  nand g488 (n_945, n_271, n_270);
  nand g489 (n_946, n_269, n_271);
  nand g490 (n_281, n_944, n_945, n_946);
  xor g491 (n_947, n_272, n_273);
  xor g492 (n_167, n_947, n_274);
  nand g493 (n_948, n_272, n_273);
  nand g494 (n_949, n_274, n_273);
  nand g495 (n_950, n_272, n_274);
  nand g496 (n_100, n_948, n_949, n_950);
  xor g497 (n_951, A[1], A[11]);
  xor g498 (n_278, n_951, A[7]);
  nand g499 (n_952, A[1], A[11]);
  nand g502 (n_284, n_952, n_925, n_880);
  xor g503 (n_955, A[5], A[13]);
  xor g504 (n_277, n_955, A[3]);
  nand g505 (n_956, A[5], A[13]);
  nand g506 (n_957, A[3], A[13]);
  nand g508 (n_285, n_956, n_957, n_873);
  xor g509 (n_959, A[9], n_275);
  xor g510 (n_280, n_959, n_276);
  nand g511 (n_960, A[9], n_275);
  nand g512 (n_961, n_276, n_275);
  nand g513 (n_962, A[9], n_276);
  nand g514 (n_288, n_960, n_961, n_962);
  xor g515 (n_963, n_277, n_278);
  xor g516 (n_282, n_963, n_279);
  nand g517 (n_964, n_277, n_278);
  nand g518 (n_965, n_279, n_278);
  nand g519 (n_966, n_277, n_279);
  nand g520 (n_290, n_964, n_965, n_966);
  xor g521 (n_967, n_280, n_281);
  xor g522 (n_166, n_967, n_282);
  nand g523 (n_968, n_280, n_281);
  nand g524 (n_969, n_282, n_281);
  nand g525 (n_970, n_280, n_282);
  nand g526 (n_99, n_968, n_969, n_970);
  xor g527 (n_283, A[14], A[12]);
  and g528 (n_292, A[14], A[12]);
  xor g529 (n_971, A[8], A[0]);
  xor g530 (n_287, n_971, A[6]);
  nand g531 (n_972, A[8], A[0]);
  nand g532 (n_973, A[6], A[0]);
  xor g535 (n_975, A[10], A[4]);
  xor g536 (n_286, n_975, A[2]);
  nand g537 (n_976, A[10], A[4]);
  nand g539 (n_978, A[10], A[2]);
  nand g540 (n_294, n_976, n_890, n_978);
  xor g541 (n_979, n_283, n_284);
  xor g542 (n_289, n_979, n_285);
  nand g543 (n_980, n_283, n_284);
  nand g544 (n_981, n_285, n_284);
  nand g545 (n_982, n_283, n_285);
  nand g546 (n_298, n_980, n_981, n_982);
  xor g547 (n_983, n_286, n_287);
  xor g548 (n_291, n_983, n_288);
  nand g549 (n_984, n_286, n_287);
  nand g550 (n_985, n_288, n_287);
  nand g551 (n_986, n_286, n_288);
  nand g552 (n_301, n_984, n_985, n_986);
  xor g553 (n_987, n_289, n_290);
  xor g554 (n_165, n_987, n_291);
  nand g555 (n_988, n_289, n_290);
  nand g556 (n_989, n_291, n_290);
  nand g557 (n_990, n_289, n_291);
  nand g558 (n_98, n_988, n_989, n_990);
  xor g559 (n_991, A[1], A[15]);
  xor g560 (n_295, n_991, A[13]);
  nand g561 (n_992, A[1], A[15]);
  nand g562 (n_993, A[13], A[15]);
  nand g563 (n_994, A[1], A[13]);
  nand g564 (n_303, n_992, n_993, n_994);
  xor g565 (n_995, A[9], A[7]);
  xor g566 (n_296, n_995, A[11]);
  nand g567 (n_996, A[9], A[7]);
  nand g569 (n_998, A[9], A[11]);
  nand g570 (n_304, n_996, n_925, n_998);
  xor g571 (n_999, A[5], A[3]);
  xor g572 (n_297, n_999, n_292);
  nand g574 (n_1001, n_292, A[3]);
  nand g575 (n_1002, A[5], n_292);
  nand g576 (n_307, n_873, n_1001, n_1002);
  xor g577 (n_1003, n_293, n_294);
  xor g578 (n_299, n_1003, n_295);
  nand g579 (n_1004, n_293, n_294);
  nand g580 (n_1005, n_295, n_294);
  nand g581 (n_1006, n_293, n_295);
  nand g582 (n_309, n_1004, n_1005, n_1006);
  xor g583 (n_1007, n_296, n_297);
  xor g584 (n_300, n_1007, n_298);
  nand g585 (n_1008, n_296, n_297);
  nand g586 (n_1009, n_298, n_297);
  nand g587 (n_1010, n_296, n_298);
  nand g588 (n_311, n_1008, n_1009, n_1010);
  xor g589 (n_1011, n_299, n_300);
  xor g590 (n_164, n_1011, n_301);
  nand g591 (n_1012, n_299, n_300);
  nand g592 (n_1013, n_301, n_300);
  nand g593 (n_1014, n_299, n_301);
  nand g594 (n_97, n_1012, n_1013, n_1014);
  xor g595 (n_302, A[16], A[14]);
  and g596 (n_313, A[16], A[14]);
  xor g597 (n_1015, A[10], A[2]);
  xor g598 (n_306, n_1015, A[0]);
  nand g601 (n_1018, A[10], A[0]);
  nand g602 (n_314, n_978, n_876, n_1018);
  xor g603 (n_1019, A[8], A[12]);
  xor g604 (n_305, n_1019, A[6]);
  nand g605 (n_1020, A[8], A[12]);
  nand g606 (n_1021, A[6], A[12]);
  xor g609 (n_1023, A[4], n_302);
  xor g610 (n_308, n_1023, n_303);
  nand g611 (n_1024, A[4], n_302);
  nand g612 (n_1025, n_303, n_302);
  nand g613 (n_1026, A[4], n_303);
  nand g614 (n_319, n_1024, n_1025, n_1026);
  xor g615 (n_1027, n_304, n_305);
  xor g616 (n_310, n_1027, n_306);
  nand g617 (n_1028, n_304, n_305);
  nand g618 (n_1029, n_306, n_305);
  nand g619 (n_1030, n_304, n_306);
  nand g620 (n_321, n_1028, n_1029, n_1030);
  xor g621 (n_1031, n_307, n_308);
  xor g622 (n_312, n_1031, n_309);
  nand g623 (n_1032, n_307, n_308);
  nand g624 (n_1033, n_309, n_308);
  nand g625 (n_1034, n_307, n_309);
  nand g626 (n_323, n_1032, n_1033, n_1034);
  xor g627 (n_1035, n_310, n_311);
  xor g628 (n_163, n_1035, n_312);
  nand g629 (n_1036, n_310, n_311);
  nand g630 (n_1037, n_312, n_311);
  nand g631 (n_1038, n_310, n_312);
  nand g632 (n_96, n_1036, n_1037, n_1038);
  xor g633 (n_1039, A[1], A[17]);
  xor g634 (n_317, n_1039, A[15]);
  nand g635 (n_1040, A[1], A[17]);
  nand g636 (n_1041, A[15], A[17]);
  nand g638 (n_326, n_1040, n_1041, n_992);
  xor g640 (n_318, n_923, A[9]);
  nand g644 (n_328, n_924, n_998, n_897);
  xor g645 (n_1047, A[13], A[7]);
  xor g646 (n_316, n_1047, A[5]);
  nand g647 (n_1048, A[13], A[7]);
  nand g650 (n_327, n_1048, n_881, n_956);
  xor g651 (n_1051, n_313, n_314);
  xor g652 (n_320, n_1051, n_315);
  nand g653 (n_1052, n_313, n_314);
  nand g654 (n_1053, n_315, n_314);
  nand g655 (n_1054, n_313, n_315);
  nand g656 (n_332, n_1052, n_1053, n_1054);
  xor g657 (n_1055, n_316, n_317);
  xor g658 (n_322, n_1055, n_318);
  nand g659 (n_1056, n_316, n_317);
  nand g660 (n_1057, n_318, n_317);
  nand g661 (n_1058, n_316, n_318);
  nand g662 (n_334, n_1056, n_1057, n_1058);
  xor g663 (n_1059, n_319, n_320);
  xor g664 (n_324, n_1059, n_321);
  nand g665 (n_1060, n_319, n_320);
  nand g666 (n_1061, n_321, n_320);
  nand g667 (n_1062, n_319, n_321);
  nand g668 (n_110, n_1060, n_1061, n_1062);
  xor g669 (n_1063, n_322, n_323);
  xor g670 (n_162, n_1063, n_324);
  nand g671 (n_1064, n_322, n_323);
  nand g672 (n_1065, n_324, n_323);
  nand g673 (n_1066, n_322, n_324);
  nand g674 (n_95, n_1064, n_1065, n_1066);
  xor g675 (n_325, A[18], A[16]);
  and g676 (n_113, A[18], A[16]);
  xor g677 (n_1067, A[12], A[4]);
  xor g678 (n_329, n_1067, A[2]);
  nand g679 (n_1068, A[12], A[4]);
  nand g681 (n_1070, A[12], A[2]);
  nand g682 (n_335, n_1068, n_890, n_1070);
  xor g683 (n_1071, A[10], A[0]);
  xor g684 (n_330, n_1071, A[14]);
  nand g686 (n_1073, A[14], A[0]);
  nand g687 (n_1074, A[10], A[14]);
  nand g688 (n_336, n_1018, n_1073, n_1074);
  xor g690 (n_331, n_250, n_325);
  nand g692 (n_1077, n_325, A[6]);
  nand g693 (n_1078, A[8], n_325);
  xor g695 (n_1079, n_326, n_327);
  xor g696 (n_333, n_1079, n_328);
  nand g697 (n_1080, n_326, n_327);
  nand g698 (n_1081, n_328, n_327);
  nand g699 (n_1082, n_326, n_328);
  nand g700 (n_342, n_1080, n_1081, n_1082);
  xor g701 (n_1083, n_329, n_330);
  xor g702 (n_109, n_1083, n_331);
  nand g703 (n_1084, n_329, n_330);
  nand g704 (n_1085, n_331, n_330);
  nand g705 (n_1086, n_329, n_331);
  nand g706 (n_343, n_1084, n_1085, n_1086);
  xor g707 (n_1087, n_332, n_333);
  xor g708 (n_111, n_1087, n_334);
  nand g709 (n_1088, n_332, n_333);
  nand g710 (n_1089, n_334, n_333);
  nand g711 (n_1090, n_332, n_334);
  nand g712 (n_346, n_1088, n_1089, n_1090);
  xor g713 (n_1091, n_109, n_110);
  xor g714 (n_161, n_1091, n_111);
  nand g715 (n_1092, n_109, n_110);
  nand g716 (n_1093, n_111, n_110);
  nand g717 (n_1094, n_109, n_111);
  nand g718 (n_94, n_1092, n_1093, n_1094);
  xor g719 (n_1095, A[1], A[19]);
  xor g720 (n_338, n_1095, A[13]);
  nand g721 (n_1096, A[1], A[19]);
  nand g722 (n_1097, A[13], A[19]);
  nand g724 (n_348, n_1096, n_1097, n_994);
  xor g726 (n_339, n_999, A[17]);
  nand g728 (n_1101, A[17], A[3]);
  nand g729 (n_1102, A[5], A[17]);
  nand g730 (n_349, n_873, n_1101, n_1102);
  xor g731 (n_1103, A[11], A[15]);
  xor g732 (n_337, n_1103, A[9]);
  nand g733 (n_1104, A[11], A[15]);
  nand g734 (n_1105, A[9], A[15]);
  nand g736 (n_350, n_1104, n_1105, n_998);
  xor g737 (n_1107, A[7], n_113);
  xor g738 (n_341, n_1107, n_335);
  nand g739 (n_1108, A[7], n_113);
  nand g740 (n_1109, n_335, n_113);
  nand g741 (n_1110, A[7], n_335);
  nand g742 (n_354, n_1108, n_1109, n_1110);
  xor g743 (n_1111, n_336, n_337);
  xor g744 (n_344, n_1111, n_338);
  nand g745 (n_1112, n_336, n_337);
  nand g746 (n_1113, n_338, n_337);
  nand g747 (n_1114, n_336, n_338);
  nand g748 (n_356, n_1112, n_1113, n_1114);
  xor g749 (n_1115, n_339, n_340);
  xor g750 (n_345, n_1115, n_341);
  nand g751 (n_1116, n_339, n_340);
  nand g752 (n_1117, n_341, n_340);
  nand g753 (n_1118, n_339, n_341);
  nand g754 (n_358, n_1116, n_1117, n_1118);
  xor g755 (n_1119, n_342, n_343);
  xor g756 (n_347, n_1119, n_344);
  nand g757 (n_1120, n_342, n_343);
  nand g758 (n_1121, n_344, n_343);
  nand g759 (n_1122, n_342, n_344);
  nand g760 (n_360, n_1120, n_1121, n_1122);
  xor g761 (n_1123, n_345, n_346);
  xor g762 (n_160, n_1123, n_347);
  nand g763 (n_1124, n_345, n_346);
  nand g764 (n_1125, n_347, n_346);
  nand g765 (n_1126, n_345, n_347);
  nand g766 (n_93, n_1124, n_1125, n_1126);
  xor g767 (n_1127, A[20], A[18]);
  xor g768 (n_352, n_1127, A[14]);
  nand g769 (n_1128, A[20], A[18]);
  nand g770 (n_1129, A[14], A[18]);
  nand g771 (n_1130, A[20], A[14]);
  nand g772 (n_362, n_1128, n_1129, n_1130);
  xor g774 (n_353, n_247, A[12]);
  xor g779 (n_1135, A[2], A[16]);
  xor g780 (n_351, n_1135, A[10]);
  nand g781 (n_1136, A[2], A[16]);
  nand g782 (n_1137, A[10], A[16]);
  nand g784 (n_364, n_1136, n_1137, n_978);
  xor g785 (n_1139, A[8], n_348);
  xor g786 (n_355, n_1139, n_349);
  nand g787 (n_1140, A[8], n_348);
  nand g788 (n_1141, n_349, n_348);
  nand g789 (n_1142, A[8], n_349);
  nand g790 (n_368, n_1140, n_1141, n_1142);
  xor g791 (n_1143, n_350, n_351);
  xor g792 (n_357, n_1143, n_352);
  nand g793 (n_1144, n_350, n_351);
  nand g794 (n_1145, n_352, n_351);
  nand g795 (n_1146, n_350, n_352);
  nand g796 (n_370, n_1144, n_1145, n_1146);
  xor g797 (n_1147, n_353, n_354);
  xor g798 (n_359, n_1147, n_355);
  nand g799 (n_1148, n_353, n_354);
  nand g800 (n_1149, n_355, n_354);
  nand g801 (n_1150, n_353, n_355);
  nand g802 (n_372, n_1148, n_1149, n_1150);
  xor g803 (n_1151, n_356, n_357);
  xor g804 (n_361, n_1151, n_358);
  nand g805 (n_1152, n_356, n_357);
  nand g806 (n_1153, n_358, n_357);
  nand g807 (n_1154, n_356, n_358);
  nand g808 (n_374, n_1152, n_1153, n_1154);
  xor g809 (n_1155, n_359, n_360);
  xor g810 (n_159, n_1155, n_361);
  nand g811 (n_1156, n_359, n_360);
  nand g812 (n_1157, n_361, n_360);
  nand g813 (n_1158, n_359, n_361);
  nand g814 (n_92, n_1156, n_1157, n_1158);
  xor g815 (n_1159, A[21], A[19]);
  xor g816 (n_366, n_1159, A[15]);
  nand g817 (n_1160, A[21], A[19]);
  nand g818 (n_1161, A[15], A[19]);
  nand g819 (n_1162, A[21], A[15]);
  nand g820 (n_376, n_1160, n_1161, n_1162);
  xor g822 (n_367, n_899, A[13]);
  xor g827 (n_1167, A[3], A[17]);
  xor g828 (n_365, n_1167, A[11]);
  nand g830 (n_1169, A[11], A[17]);
  nand g832 (n_378, n_1101, n_1169, n_924);
  xor g833 (n_1171, A[9], n_362);
  xor g834 (n_369, n_1171, n_363);
  nand g835 (n_1172, A[9], n_362);
  nand g836 (n_1173, n_363, n_362);
  nand g837 (n_1174, A[9], n_363);
  nand g838 (n_382, n_1172, n_1173, n_1174);
  xor g839 (n_1175, n_364, n_365);
  xor g840 (n_371, n_1175, n_366);
  nand g841 (n_1176, n_364, n_365);
  nand g842 (n_1177, n_366, n_365);
  nand g843 (n_1178, n_364, n_366);
  nand g844 (n_384, n_1176, n_1177, n_1178);
  xor g845 (n_1179, n_367, n_368);
  xor g846 (n_373, n_1179, n_369);
  nand g847 (n_1180, n_367, n_368);
  nand g848 (n_1181, n_369, n_368);
  nand g849 (n_1182, n_367, n_369);
  nand g850 (n_386, n_1180, n_1181, n_1182);
  xor g851 (n_1183, n_370, n_371);
  xor g852 (n_375, n_1183, n_372);
  nand g853 (n_1184, n_370, n_371);
  nand g854 (n_1185, n_372, n_371);
  nand g855 (n_1186, n_370, n_372);
  nand g856 (n_389, n_1184, n_1185, n_1186);
  xor g857 (n_1187, n_373, n_374);
  xor g858 (n_158, n_1187, n_375);
  nand g859 (n_1188, n_373, n_374);
  nand g860 (n_1189, n_375, n_374);
  nand g861 (n_1190, n_373, n_375);
  nand g862 (n_91, n_1188, n_1189, n_1190);
  xor g863 (n_1191, A[22], A[20]);
  xor g864 (n_380, n_1191, A[16]);
  nand g865 (n_1192, A[22], A[20]);
  nand g866 (n_1193, A[16], A[20]);
  nand g867 (n_1194, A[22], A[16]);
  nand g868 (n_390, n_1192, n_1193, n_1194);
  xor g870 (n_381, n_250, A[14]);
  nand g872 (n_1197, A[14], A[6]);
  nand g873 (n_1198, A[8], A[14]);
  xor g875 (n_1199, A[4], A[18]);
  xor g876 (n_379, n_1199, A[12]);
  nand g877 (n_1200, A[4], A[18]);
  nand g878 (n_1201, A[12], A[18]);
  nand g880 (n_392, n_1200, n_1201, n_1068);
  xor g881 (n_1203, A[10], n_376);
  xor g882 (n_383, n_1203, n_327);
  nand g883 (n_1204, A[10], n_376);
  nand g884 (n_1205, n_327, n_376);
  nand g885 (n_1206, A[10], n_327);
  nand g886 (n_394, n_1204, n_1205, n_1206);
  xor g887 (n_1207, n_378, n_379);
  xor g888 (n_385, n_1207, n_380);
  nand g889 (n_1208, n_378, n_379);
  nand g890 (n_1209, n_380, n_379);
  nand g891 (n_1210, n_378, n_380);
  nand g892 (n_396, n_1208, n_1209, n_1210);
  xor g893 (n_1211, n_381, n_382);
  xor g894 (n_387, n_1211, n_383);
  nand g895 (n_1212, n_381, n_382);
  nand g896 (n_1213, n_383, n_382);
  nand g897 (n_1214, n_381, n_383);
  nand g898 (n_398, n_1212, n_1213, n_1214);
  xor g899 (n_1215, n_384, n_385);
  xor g900 (n_388, n_1215, n_386);
  nand g901 (n_1216, n_384, n_385);
  nand g902 (n_1217, n_386, n_385);
  nand g903 (n_1218, n_384, n_386);
  nand g904 (n_401, n_1216, n_1217, n_1218);
  xor g905 (n_1219, n_387, n_388);
  xor g906 (n_157, n_1219, n_389);
  nand g907 (n_1220, n_387, n_388);
  nand g908 (n_1221, n_389, n_388);
  nand g909 (n_1222, n_387, n_389);
  nand g910 (n_90, n_1220, n_1221, n_1222);
  xor g911 (n_1223, A[23], A[21]);
  xor g912 (n_177, n_1223, A[17]);
  nand g913 (n_1224, A[23], A[21]);
  nand g914 (n_1225, A[17], A[21]);
  nand g915 (n_1226, A[23], A[17]);
  nand g916 (n_402, n_1224, n_1225, n_1226);
  xor g918 (n_393, n_995, A[15]);
  nand g920 (n_1229, A[15], A[7]);
  nand g922 (n_403, n_996, n_1229, n_1105);
  xor g923 (n_1231, A[5], A[19]);
  xor g924 (n_176, n_1231, A[13]);
  nand g925 (n_1232, A[5], A[19]);
  nand g928 (n_404, n_1232, n_1097, n_956);
  xor g929 (n_1235, A[11], n_390);
  xor g930 (n_395, n_1235, n_391);
  nand g931 (n_1236, A[11], n_390);
  nand g932 (n_1237, n_391, n_390);
  nand g933 (n_1238, A[11], n_391);
  nand g934 (n_408, n_1236, n_1237, n_1238);
  xor g935 (n_1239, n_392, n_176);
  xor g936 (n_397, n_1239, n_177);
  nand g937 (n_1240, n_392, n_176);
  nand g938 (n_1241, n_177, n_176);
  nand g939 (n_1242, n_392, n_177);
  nand g940 (n_410, n_1240, n_1241, n_1242);
  xor g941 (n_1243, n_393, n_394);
  xor g942 (n_399, n_1243, n_395);
  nand g943 (n_1244, n_393, n_394);
  nand g944 (n_1245, n_395, n_394);
  nand g945 (n_1246, n_393, n_395);
  nand g946 (n_412, n_1244, n_1245, n_1246);
  xor g947 (n_1247, n_396, n_397);
  xor g948 (n_400, n_1247, n_398);
  nand g949 (n_1248, n_396, n_397);
  nand g950 (n_1249, n_398, n_397);
  nand g951 (n_1250, n_396, n_398);
  nand g952 (n_415, n_1248, n_1249, n_1250);
  xor g953 (n_1251, n_399, n_400);
  xor g954 (n_156, n_1251, n_401);
  nand g955 (n_1252, n_399, n_400);
  nand g956 (n_1253, n_401, n_400);
  nand g957 (n_1254, n_399, n_401);
  nand g958 (n_89, n_1252, n_1253, n_1254);
  xor g959 (n_1255, A[24], A[22]);
  xor g960 (n_406, n_1255, A[18]);
  nand g961 (n_1256, A[24], A[22]);
  nand g962 (n_1257, A[18], A[22]);
  nand g963 (n_1258, A[24], A[18]);
  nand g964 (n_416, n_1256, n_1257, n_1258);
  xor g966 (n_407, n_257, A[16]);
  nand g968 (n_1261, A[16], A[8]);
  xor g971 (n_1263, A[6], A[20]);
  xor g972 (n_405, n_1263, A[14]);
  nand g973 (n_1264, A[6], A[20]);
  nand g976 (n_418, n_1264, n_1130, n_1197);
  xor g977 (n_1267, A[12], n_402);
  xor g978 (n_409, n_1267, n_403);
  nand g979 (n_1268, A[12], n_402);
  nand g980 (n_1269, n_403, n_402);
  nand g981 (n_1270, A[12], n_403);
  nand g982 (n_422, n_1268, n_1269, n_1270);
  xor g983 (n_1271, n_404, n_405);
  xor g984 (n_411, n_1271, n_406);
  nand g985 (n_1272, n_404, n_405);
  nand g986 (n_1273, n_406, n_405);
  nand g987 (n_1274, n_404, n_406);
  nand g988 (n_424, n_1272, n_1273, n_1274);
  xor g989 (n_1275, n_407, n_408);
  xor g990 (n_413, n_1275, n_409);
  nand g991 (n_1276, n_407, n_408);
  nand g992 (n_1277, n_409, n_408);
  nand g993 (n_1278, n_407, n_409);
  nand g994 (n_426, n_1276, n_1277, n_1278);
  xor g995 (n_1279, n_410, n_411);
  xor g996 (n_414, n_1279, n_412);
  nand g997 (n_1280, n_410, n_411);
  nand g998 (n_1281, n_412, n_411);
  nand g999 (n_1282, n_410, n_412);
  nand g1000 (n_429, n_1280, n_1281, n_1282);
  xor g1001 (n_1283, n_413, n_414);
  xor g1002 (n_155, n_1283, n_415);
  nand g1003 (n_1284, n_413, n_414);
  nand g1004 (n_1285, n_415, n_414);
  nand g1005 (n_1286, n_413, n_415);
  nand g1006 (n_88, n_1284, n_1285, n_1286);
  xor g1007 (n_1287, A[25], A[23]);
  xor g1008 (n_420, n_1287, A[19]);
  nand g1009 (n_1288, A[25], A[23]);
  nand g1010 (n_1289, A[19], A[23]);
  nand g1011 (n_1290, A[25], A[19]);
  nand g1012 (n_430, n_1288, n_1289, n_1290);
  xor g1013 (n_1291, A[11], A[9]);
  xor g1014 (n_421, n_1291, A[17]);
  nand g1016 (n_1293, A[17], A[9]);
  nand g1018 (n_431, n_998, n_1293, n_1169);
  xor g1019 (n_1295, A[7], A[21]);
  xor g1020 (n_419, n_1295, A[15]);
  nand g1021 (n_1296, A[7], A[21]);
  nand g1024 (n_432, n_1296, n_1162, n_1229);
  xor g1025 (n_1299, A[13], n_416);
  xor g1026 (n_423, n_1299, n_417);
  nand g1027 (n_1300, A[13], n_416);
  nand g1028 (n_1301, n_417, n_416);
  nand g1029 (n_1302, A[13], n_417);
  nand g1030 (n_436, n_1300, n_1301, n_1302);
  xor g1031 (n_1303, n_418, n_419);
  xor g1032 (n_425, n_1303, n_420);
  nand g1033 (n_1304, n_418, n_419);
  nand g1034 (n_1305, n_420, n_419);
  nand g1035 (n_1306, n_418, n_420);
  nand g1036 (n_438, n_1304, n_1305, n_1306);
  xor g1037 (n_1307, n_421, n_422);
  xor g1038 (n_427, n_1307, n_423);
  nand g1039 (n_1308, n_421, n_422);
  nand g1040 (n_1309, n_423, n_422);
  nand g1041 (n_1310, n_421, n_423);
  nand g1042 (n_440, n_1308, n_1309, n_1310);
  xor g1043 (n_1311, n_424, n_425);
  xor g1044 (n_428, n_1311, n_426);
  nand g1045 (n_1312, n_424, n_425);
  nand g1046 (n_1313, n_426, n_425);
  nand g1047 (n_1314, n_424, n_426);
  nand g1048 (n_443, n_1312, n_1313, n_1314);
  xor g1049 (n_1315, n_427, n_428);
  xor g1050 (n_154, n_1315, n_429);
  nand g1051 (n_1316, n_427, n_428);
  nand g1052 (n_1317, n_429, n_428);
  nand g1053 (n_1318, n_427, n_429);
  nand g1054 (n_87, n_1316, n_1317, n_1318);
  xor g1055 (n_1319, A[26], A[24]);
  xor g1056 (n_434, n_1319, A[20]);
  nand g1057 (n_1320, A[26], A[24]);
  nand g1058 (n_1321, A[20], A[24]);
  nand g1059 (n_1322, A[26], A[20]);
  nand g1060 (n_444, n_1320, n_1321, n_1322);
  xor g1062 (n_435, n_268, A[18]);
  nand g1064 (n_1325, A[18], A[10]);
  xor g1067 (n_1327, A[8], A[22]);
  xor g1068 (n_433, n_1327, A[16]);
  nand g1069 (n_1328, A[8], A[22]);
  nand g1072 (n_446, n_1328, n_1194, n_1261);
  xor g1073 (n_1331, A[14], n_430);
  xor g1074 (n_437, n_1331, n_431);
  nand g1075 (n_1332, A[14], n_430);
  nand g1076 (n_1333, n_431, n_430);
  nand g1077 (n_1334, A[14], n_431);
  nand g1078 (n_450, n_1332, n_1333, n_1334);
  xor g1079 (n_1335, n_432, n_433);
  xor g1080 (n_439, n_1335, n_434);
  nand g1081 (n_1336, n_432, n_433);
  nand g1082 (n_1337, n_434, n_433);
  nand g1083 (n_1338, n_432, n_434);
  nand g1084 (n_452, n_1336, n_1337, n_1338);
  xor g1085 (n_1339, n_435, n_436);
  xor g1086 (n_441, n_1339, n_437);
  nand g1087 (n_1340, n_435, n_436);
  nand g1088 (n_1341, n_437, n_436);
  nand g1089 (n_1342, n_435, n_437);
  nand g1090 (n_454, n_1340, n_1341, n_1342);
  xor g1091 (n_1343, n_438, n_439);
  xor g1092 (n_442, n_1343, n_440);
  nand g1093 (n_1344, n_438, n_439);
  nand g1094 (n_1345, n_440, n_439);
  nand g1095 (n_1346, n_438, n_440);
  nand g1096 (n_457, n_1344, n_1345, n_1346);
  xor g1097 (n_1347, n_441, n_442);
  xor g1098 (n_153, n_1347, n_443);
  nand g1099 (n_1348, n_441, n_442);
  nand g1100 (n_1349, n_443, n_442);
  nand g1101 (n_1350, n_441, n_443);
  nand g1102 (n_86, n_1348, n_1349, n_1350);
  xor g1103 (n_1351, A[27], A[25]);
  xor g1104 (n_448, n_1351, A[21]);
  nand g1105 (n_1352, A[27], A[25]);
  nand g1106 (n_1353, A[21], A[25]);
  nand g1107 (n_1354, A[27], A[21]);
  nand g1108 (n_458, n_1352, n_1353, n_1354);
  xor g1109 (n_1355, A[13], A[11]);
  xor g1110 (n_449, n_1355, A[19]);
  nand g1111 (n_1356, A[13], A[11]);
  nand g1112 (n_1357, A[19], A[11]);
  nand g1114 (n_459, n_1356, n_1357, n_1097);
  xor g1115 (n_1359, A[9], A[23]);
  xor g1116 (n_447, n_1359, A[17]);
  nand g1117 (n_1360, A[9], A[23]);
  nand g1120 (n_460, n_1360, n_1226, n_1293);
  xor g1121 (n_1363, A[15], n_444);
  xor g1122 (n_451, n_1363, n_445);
  nand g1123 (n_1364, A[15], n_444);
  nand g1124 (n_1365, n_445, n_444);
  nand g1125 (n_1366, A[15], n_445);
  nand g1126 (n_464, n_1364, n_1365, n_1366);
  xor g1127 (n_1367, n_446, n_447);
  xor g1128 (n_453, n_1367, n_448);
  nand g1129 (n_1368, n_446, n_447);
  nand g1130 (n_1369, n_448, n_447);
  nand g1131 (n_1370, n_446, n_448);
  nand g1132 (n_466, n_1368, n_1369, n_1370);
  xor g1133 (n_1371, n_449, n_450);
  xor g1134 (n_455, n_1371, n_451);
  nand g1135 (n_1372, n_449, n_450);
  nand g1136 (n_1373, n_451, n_450);
  nand g1137 (n_1374, n_449, n_451);
  nand g1138 (n_468, n_1372, n_1373, n_1374);
  xor g1139 (n_1375, n_452, n_453);
  xor g1140 (n_456, n_1375, n_454);
  nand g1141 (n_1376, n_452, n_453);
  nand g1142 (n_1377, n_454, n_453);
  nand g1143 (n_1378, n_452, n_454);
  nand g1144 (n_471, n_1376, n_1377, n_1378);
  xor g1145 (n_1379, n_455, n_456);
  xor g1146 (n_152, n_1379, n_457);
  nand g1147 (n_1380, n_455, n_456);
  nand g1148 (n_1381, n_457, n_456);
  nand g1149 (n_1382, n_455, n_457);
  nand g1150 (n_85, n_1380, n_1381, n_1382);
  xor g1151 (n_1383, A[28], A[26]);
  xor g1152 (n_462, n_1383, A[22]);
  nand g1153 (n_1384, A[28], A[26]);
  nand g1154 (n_1385, A[22], A[26]);
  nand g1155 (n_1386, A[28], A[22]);
  nand g1156 (n_472, n_1384, n_1385, n_1386);
  xor g1158 (n_463, n_283, A[20]);
  nand g1160 (n_1389, A[20], A[12]);
  xor g1163 (n_1391, A[10], A[24]);
  xor g1164 (n_461, n_1391, A[18]);
  nand g1165 (n_1392, A[10], A[24]);
  nand g1168 (n_474, n_1392, n_1258, n_1325);
  xor g1169 (n_1395, A[16], n_458);
  xor g1170 (n_465, n_1395, n_459);
  nand g1171 (n_1396, A[16], n_458);
  nand g1172 (n_1397, n_459, n_458);
  nand g1173 (n_1398, A[16], n_459);
  nand g1174 (n_478, n_1396, n_1397, n_1398);
  xor g1175 (n_1399, n_460, n_461);
  xor g1176 (n_467, n_1399, n_462);
  nand g1177 (n_1400, n_460, n_461);
  nand g1178 (n_1401, n_462, n_461);
  nand g1179 (n_1402, n_460, n_462);
  nand g1180 (n_480, n_1400, n_1401, n_1402);
  xor g1181 (n_1403, n_463, n_464);
  xor g1182 (n_469, n_1403, n_465);
  nand g1183 (n_1404, n_463, n_464);
  nand g1184 (n_1405, n_465, n_464);
  nand g1185 (n_1406, n_463, n_465);
  nand g1186 (n_482, n_1404, n_1405, n_1406);
  xor g1187 (n_1407, n_466, n_467);
  xor g1188 (n_470, n_1407, n_468);
  nand g1189 (n_1408, n_466, n_467);
  nand g1190 (n_1409, n_468, n_467);
  nand g1191 (n_1410, n_466, n_468);
  nand g1192 (n_485, n_1408, n_1409, n_1410);
  xor g1193 (n_1411, n_469, n_470);
  xor g1194 (n_151, n_1411, n_471);
  nand g1195 (n_1412, n_469, n_470);
  nand g1196 (n_1413, n_471, n_470);
  nand g1197 (n_1414, n_469, n_471);
  nand g1198 (n_84, n_1412, n_1413, n_1414);
  xor g1199 (n_1415, A[29], A[27]);
  xor g1200 (n_476, n_1415, A[23]);
  nand g1201 (n_1416, A[29], A[27]);
  nand g1202 (n_1417, A[23], A[27]);
  nand g1203 (n_1418, A[29], A[23]);
  nand g1204 (n_486, n_1416, n_1417, n_1418);
  xor g1205 (n_1419, A[15], A[13]);
  xor g1206 (n_477, n_1419, A[21]);
  nand g1208 (n_1421, A[21], A[13]);
  nand g1210 (n_487, n_993, n_1421, n_1162);
  xor g1211 (n_1423, A[11], A[25]);
  xor g1212 (n_475, n_1423, A[19]);
  nand g1213 (n_1424, A[11], A[25]);
  nand g1216 (n_488, n_1424, n_1290, n_1357);
  xor g1217 (n_1427, A[17], n_472);
  xor g1218 (n_479, n_1427, n_473);
  nand g1219 (n_1428, A[17], n_472);
  nand g1220 (n_1429, n_473, n_472);
  nand g1221 (n_1430, A[17], n_473);
  nand g1222 (n_492, n_1428, n_1429, n_1430);
  xor g1223 (n_1431, n_474, n_475);
  xor g1224 (n_481, n_1431, n_476);
  nand g1225 (n_1432, n_474, n_475);
  nand g1226 (n_1433, n_476, n_475);
  nand g1227 (n_1434, n_474, n_476);
  nand g1228 (n_494, n_1432, n_1433, n_1434);
  xor g1229 (n_1435, n_477, n_478);
  xor g1230 (n_483, n_1435, n_479);
  nand g1231 (n_1436, n_477, n_478);
  nand g1232 (n_1437, n_479, n_478);
  nand g1233 (n_1438, n_477, n_479);
  nand g1234 (n_496, n_1436, n_1437, n_1438);
  xor g1235 (n_1439, n_480, n_481);
  xor g1236 (n_484, n_1439, n_482);
  nand g1237 (n_1440, n_480, n_481);
  nand g1238 (n_1441, n_482, n_481);
  nand g1239 (n_1442, n_480, n_482);
  nand g1240 (n_499, n_1440, n_1441, n_1442);
  xor g1241 (n_1443, n_483, n_484);
  xor g1242 (n_150, n_1443, n_485);
  nand g1243 (n_1444, n_483, n_484);
  nand g1244 (n_1445, n_485, n_484);
  nand g1245 (n_1446, n_483, n_485);
  nand g1246 (n_83, n_1444, n_1445, n_1446);
  xor g1247 (n_1447, A[30], A[28]);
  xor g1248 (n_490, n_1447, A[24]);
  nand g1249 (n_1448, A[30], A[28]);
  nand g1250 (n_1449, A[24], A[28]);
  nand g1251 (n_1450, A[30], A[24]);
  nand g1252 (n_500, n_1448, n_1449, n_1450);
  xor g1254 (n_491, n_302, A[22]);
  nand g1256 (n_1453, A[22], A[14]);
  xor g1259 (n_1455, A[12], A[26]);
  xor g1260 (n_489, n_1455, A[20]);
  nand g1261 (n_1456, A[12], A[26]);
  nand g1264 (n_502, n_1456, n_1322, n_1389);
  xor g1265 (n_1459, A[18], n_486);
  xor g1266 (n_493, n_1459, n_487);
  nand g1267 (n_1460, A[18], n_486);
  nand g1268 (n_1461, n_487, n_486);
  nand g1269 (n_1462, A[18], n_487);
  nand g1270 (n_506, n_1460, n_1461, n_1462);
  xor g1271 (n_1463, n_488, n_489);
  xor g1272 (n_495, n_1463, n_490);
  nand g1273 (n_1464, n_488, n_489);
  nand g1274 (n_1465, n_490, n_489);
  nand g1275 (n_1466, n_488, n_490);
  nand g1276 (n_508, n_1464, n_1465, n_1466);
  xor g1277 (n_1467, n_491, n_492);
  xor g1278 (n_497, n_1467, n_493);
  nand g1279 (n_1468, n_491, n_492);
  nand g1280 (n_1469, n_493, n_492);
  nand g1281 (n_1470, n_491, n_493);
  nand g1282 (n_510, n_1468, n_1469, n_1470);
  xor g1283 (n_1471, n_494, n_495);
  xor g1284 (n_498, n_1471, n_496);
  nand g1285 (n_1472, n_494, n_495);
  nand g1286 (n_1473, n_496, n_495);
  nand g1287 (n_1474, n_494, n_496);
  nand g1288 (n_513, n_1472, n_1473, n_1474);
  xor g1289 (n_1475, n_497, n_498);
  xor g1290 (n_149, n_1475, n_499);
  nand g1291 (n_1476, n_497, n_498);
  nand g1292 (n_1477, n_499, n_498);
  nand g1293 (n_1478, n_497, n_499);
  nand g1294 (n_82, n_1476, n_1477, n_1478);
  xor g1295 (n_1479, A[31], A[29]);
  xor g1296 (n_504, n_1479, A[25]);
  nand g1297 (n_1480, A[31], A[29]);
  nand g1298 (n_1481, A[25], A[29]);
  nand g1299 (n_1482, A[31], A[25]);
  nand g1300 (n_514, n_1480, n_1481, n_1482);
  xor g1301 (n_1483, A[17], A[15]);
  xor g1302 (n_505, n_1483, A[23]);
  nand g1304 (n_1485, A[23], A[15]);
  nand g1306 (n_515, n_1041, n_1485, n_1226);
  xor g1307 (n_1487, A[13], A[27]);
  xor g1308 (n_503, n_1487, A[21]);
  nand g1309 (n_1488, A[13], A[27]);
  nand g1312 (n_516, n_1488, n_1354, n_1421);
  xor g1313 (n_1491, A[19], n_500);
  xor g1314 (n_507, n_1491, n_501);
  nand g1315 (n_1492, A[19], n_500);
  nand g1316 (n_1493, n_501, n_500);
  nand g1317 (n_1494, A[19], n_501);
  nand g1318 (n_520, n_1492, n_1493, n_1494);
  xor g1319 (n_1495, n_502, n_503);
  xor g1320 (n_509, n_1495, n_504);
  nand g1321 (n_1496, n_502, n_503);
  nand g1322 (n_1497, n_504, n_503);
  nand g1323 (n_1498, n_502, n_504);
  nand g1324 (n_522, n_1496, n_1497, n_1498);
  xor g1325 (n_1499, n_505, n_506);
  xor g1326 (n_511, n_1499, n_507);
  nand g1327 (n_1500, n_505, n_506);
  nand g1328 (n_1501, n_507, n_506);
  nand g1329 (n_1502, n_505, n_507);
  nand g1330 (n_524, n_1500, n_1501, n_1502);
  xor g1331 (n_1503, n_508, n_509);
  xor g1332 (n_512, n_1503, n_510);
  nand g1333 (n_1504, n_508, n_509);
  nand g1334 (n_1505, n_510, n_509);
  nand g1335 (n_1506, n_508, n_510);
  nand g1336 (n_527, n_1504, n_1505, n_1506);
  xor g1337 (n_1507, n_511, n_512);
  xor g1338 (n_148, n_1507, n_513);
  nand g1339 (n_1508, n_511, n_512);
  nand g1340 (n_1509, n_513, n_512);
  nand g1341 (n_1510, n_511, n_513);
  nand g1342 (n_81, n_1508, n_1509, n_1510);
  xor g1343 (n_1511, A[32], A[30]);
  xor g1344 (n_518, n_1511, A[26]);
  nand g1345 (n_1512, A[32], A[30]);
  nand g1346 (n_1513, A[26], A[30]);
  nand g1347 (n_1514, A[32], A[26]);
  nand g1348 (n_528, n_1512, n_1513, n_1514);
  xor g1350 (n_519, n_325, A[24]);
  nand g1352 (n_1517, A[24], A[16]);
  xor g1355 (n_1519, A[14], A[28]);
  xor g1356 (n_517, n_1519, A[22]);
  nand g1357 (n_1520, A[14], A[28]);
  nand g1360 (n_530, n_1520, n_1386, n_1453);
  xor g1361 (n_1523, A[20], n_514);
  xor g1362 (n_521, n_1523, n_515);
  nand g1363 (n_1524, A[20], n_514);
  nand g1364 (n_1525, n_515, n_514);
  nand g1365 (n_1526, A[20], n_515);
  nand g1366 (n_534, n_1524, n_1525, n_1526);
  xor g1367 (n_1527, n_516, n_517);
  xor g1368 (n_523, n_1527, n_518);
  nand g1369 (n_1528, n_516, n_517);
  nand g1370 (n_1529, n_518, n_517);
  nand g1371 (n_1530, n_516, n_518);
  nand g1372 (n_536, n_1528, n_1529, n_1530);
  xor g1373 (n_1531, n_519, n_520);
  xor g1374 (n_525, n_1531, n_521);
  nand g1375 (n_1532, n_519, n_520);
  nand g1376 (n_1533, n_521, n_520);
  nand g1377 (n_1534, n_519, n_521);
  nand g1378 (n_538, n_1532, n_1533, n_1534);
  xor g1379 (n_1535, n_522, n_523);
  xor g1380 (n_526, n_1535, n_524);
  nand g1381 (n_1536, n_522, n_523);
  nand g1382 (n_1537, n_524, n_523);
  nand g1383 (n_1538, n_522, n_524);
  nand g1384 (n_541, n_1536, n_1537, n_1538);
  xor g1385 (n_1539, n_525, n_526);
  xor g1386 (n_147, n_1539, n_527);
  nand g1387 (n_1540, n_525, n_526);
  nand g1388 (n_1541, n_527, n_526);
  nand g1389 (n_1542, n_525, n_527);
  nand g1390 (n_80, n_1540, n_1541, n_1542);
  xor g1391 (n_1543, A[33], A[31]);
  xor g1392 (n_532, n_1543, A[27]);
  nand g1393 (n_1544, A[33], A[31]);
  nand g1394 (n_1545, A[27], A[31]);
  nand g1395 (n_1546, A[33], A[27]);
  nand g1396 (n_542, n_1544, n_1545, n_1546);
  xor g1397 (n_1547, A[19], A[17]);
  xor g1398 (n_533, n_1547, A[25]);
  nand g1399 (n_1548, A[19], A[17]);
  nand g1400 (n_1549, A[25], A[17]);
  nand g1402 (n_544, n_1548, n_1549, n_1290);
  xor g1403 (n_1551, A[15], A[29]);
  xor g1404 (n_531, n_1551, A[23]);
  nand g1405 (n_1552, A[15], A[29]);
  nand g1408 (n_543, n_1552, n_1418, n_1485);
  xor g1409 (n_1555, A[21], n_528);
  xor g1410 (n_535, n_1555, n_529);
  nand g1411 (n_1556, A[21], n_528);
  nand g1412 (n_1557, n_529, n_528);
  nand g1413 (n_1558, A[21], n_529);
  nand g1414 (n_548, n_1556, n_1557, n_1558);
  xor g1415 (n_1559, n_530, n_531);
  xor g1416 (n_537, n_1559, n_532);
  nand g1417 (n_1560, n_530, n_531);
  nand g1418 (n_1561, n_532, n_531);
  nand g1419 (n_1562, n_530, n_532);
  nand g1420 (n_550, n_1560, n_1561, n_1562);
  xor g1421 (n_1563, n_533, n_534);
  xor g1422 (n_539, n_1563, n_535);
  nand g1423 (n_1564, n_533, n_534);
  nand g1424 (n_1565, n_535, n_534);
  nand g1425 (n_1566, n_533, n_535);
  nand g1426 (n_553, n_1564, n_1565, n_1566);
  xor g1427 (n_1567, n_536, n_537);
  xor g1428 (n_540, n_1567, n_538);
  nand g1429 (n_1568, n_536, n_537);
  nand g1430 (n_1569, n_538, n_537);
  nand g1431 (n_1570, n_536, n_538);
  nand g1432 (n_555, n_1568, n_1569, n_1570);
  xor g1433 (n_1571, n_539, n_540);
  xor g1434 (n_146, n_1571, n_541);
  nand g1435 (n_1572, n_539, n_540);
  nand g1436 (n_1573, n_541, n_540);
  nand g1437 (n_1574, n_539, n_541);
  nand g1438 (n_79, n_1572, n_1573, n_1574);
  xor g1439 (n_1575, A[32], A[28]);
  xor g1440 (n_546, n_1575, A[20]);
  nand g1441 (n_1576, A[32], A[28]);
  nand g1442 (n_1577, A[20], A[28]);
  nand g1443 (n_1578, A[32], A[20]);
  nand g1444 (n_556, n_1576, n_1577, n_1578);
  xor g1445 (n_1579, A[18], A[26]);
  xor g1446 (n_547, n_1579, A[16]);
  nand g1447 (n_1580, A[18], A[26]);
  nand g1448 (n_1581, A[16], A[26]);
  xor g1451 (n_1583, A[30], A[24]);
  xor g1452 (n_545, n_1583, A[22]);
  nand g1455 (n_1586, A[30], A[22]);
  nand g1456 (n_557, n_1450, n_1256, n_1586);
  xor g1457 (n_1587, A[34], n_542);
  xor g1458 (n_549, n_1587, n_543);
  nand g1459 (n_1588, A[34], n_542);
  nand g1460 (n_1589, n_543, n_542);
  nand g1461 (n_1590, A[34], n_543);
  nand g1462 (n_562, n_1588, n_1589, n_1590);
  xor g1463 (n_1591, n_544, n_545);
  xor g1464 (n_551, n_1591, n_546);
  nand g1465 (n_1592, n_544, n_545);
  nand g1466 (n_1593, n_546, n_545);
  nand g1467 (n_1594, n_544, n_546);
  nand g1468 (n_564, n_1592, n_1593, n_1594);
  xor g1469 (n_1595, n_547, n_548);
  xor g1470 (n_552, n_1595, n_549);
  nand g1471 (n_1596, n_547, n_548);
  nand g1472 (n_1597, n_549, n_548);
  nand g1473 (n_1598, n_547, n_549);
  nand g1474 (n_567, n_1596, n_1597, n_1598);
  xor g1475 (n_1599, n_550, n_551);
  xor g1476 (n_554, n_1599, n_552);
  nand g1477 (n_1600, n_550, n_551);
  nand g1478 (n_1601, n_552, n_551);
  nand g1479 (n_1602, n_550, n_552);
  nand g1480 (n_569, n_1600, n_1601, n_1602);
  xor g1481 (n_1603, n_553, n_554);
  xor g1482 (n_145, n_1603, n_555);
  nand g1483 (n_1604, n_553, n_554);
  nand g1484 (n_1605, n_555, n_554);
  nand g1485 (n_1606, n_553, n_555);
  nand g1486 (n_78, n_1604, n_1605, n_1606);
  xor g1487 (n_1607, A[33], A[29]);
  xor g1488 (n_560, n_1607, A[21]);
  nand g1489 (n_1608, A[33], A[29]);
  nand g1490 (n_1609, A[21], A[29]);
  nand g1491 (n_1610, A[33], A[21]);
  nand g1492 (n_571, n_1608, n_1609, n_1610);
  xor g1493 (n_1611, A[19], A[27]);
  xor g1494 (n_561, n_1611, A[17]);
  nand g1495 (n_1612, A[19], A[27]);
  nand g1496 (n_1613, A[17], A[27]);
  nand g1498 (n_572, n_1612, n_1613, n_1548);
  xor g1499 (n_1615, A[31], A[25]);
  xor g1500 (n_559, n_1615, A[23]);
  nand g1503 (n_1618, A[31], A[23]);
  nand g1504 (n_570, n_1482, n_1288, n_1618);
  xor g1505 (n_1619, A[35], n_556);
  xor g1506 (n_563, n_1619, n_557);
  nand g1507 (n_1620, A[35], n_556);
  nand g1508 (n_1621, n_557, n_556);
  nand g1509 (n_1622, A[35], n_557);
  nand g1510 (n_576, n_1620, n_1621, n_1622);
  xor g1511 (n_1623, n_558, n_559);
  xor g1512 (n_565, n_1623, n_560);
  nand g1513 (n_1624, n_558, n_559);
  nand g1514 (n_1625, n_560, n_559);
  nand g1515 (n_1626, n_558, n_560);
  nand g1516 (n_577, n_1624, n_1625, n_1626);
  xor g1517 (n_1627, n_561, n_562);
  xor g1518 (n_566, n_1627, n_563);
  nand g1519 (n_1628, n_561, n_562);
  nand g1520 (n_1629, n_563, n_562);
  nand g1521 (n_1630, n_561, n_563);
  nand g1522 (n_581, n_1628, n_1629, n_1630);
  xor g1523 (n_1631, n_564, n_565);
  xor g1524 (n_568, n_1631, n_566);
  nand g1525 (n_1632, n_564, n_565);
  nand g1526 (n_1633, n_566, n_565);
  nand g1527 (n_1634, n_564, n_566);
  nand g1528 (n_583, n_1632, n_1633, n_1634);
  xor g1529 (n_1635, n_567, n_568);
  xor g1530 (n_144, n_1635, n_569);
  nand g1531 (n_1636, n_567, n_568);
  nand g1532 (n_1637, n_569, n_568);
  nand g1533 (n_1638, n_567, n_569);
  nand g1534 (n_77, n_1636, n_1637, n_1638);
  xor g1536 (n_573, n_1511, A[22]);
  nand g1539 (n_1642, A[32], A[22]);
  nand g1540 (n_584, n_1512, n_1586, n_1642);
  xor g1541 (n_1643, A[20], A[28]);
  xor g1542 (n_575, n_1643, A[18]);
  nand g1544 (n_1645, A[18], A[28]);
  nand g1546 (n_585, n_1577, n_1645, n_1128);
  xor g1548 (n_574, n_1319, A[34]);
  nand g1550 (n_1649, A[34], A[24]);
  nand g1551 (n_1650, A[26], A[34]);
  nand g1552 (n_587, n_1320, n_1649, n_1650);
  xor g1553 (n_1651, A[36], n_570);
  xor g1554 (n_578, n_1651, n_571);
  nand g1555 (n_1652, A[36], n_570);
  nand g1556 (n_1653, n_571, n_570);
  nand g1557 (n_1654, A[36], n_571);
  nand g1558 (n_590, n_1652, n_1653, n_1654);
  xor g1559 (n_1655, n_572, n_573);
  xor g1560 (n_579, n_1655, n_574);
  nand g1561 (n_1656, n_572, n_573);
  nand g1562 (n_1657, n_574, n_573);
  nand g1563 (n_1658, n_572, n_574);
  nand g1564 (n_591, n_1656, n_1657, n_1658);
  xor g1565 (n_1659, n_575, n_576);
  xor g1566 (n_580, n_1659, n_577);
  nand g1567 (n_1660, n_575, n_576);
  nand g1568 (n_1661, n_577, n_576);
  nand g1569 (n_1662, n_575, n_577);
  nand g1570 (n_595, n_1660, n_1661, n_1662);
  xor g1571 (n_1663, n_578, n_579);
  xor g1572 (n_582, n_1663, n_580);
  nand g1573 (n_1664, n_578, n_579);
  nand g1574 (n_1665, n_580, n_579);
  nand g1575 (n_1666, n_578, n_580);
  nand g1576 (n_597, n_1664, n_1665, n_1666);
  xor g1577 (n_1667, n_581, n_582);
  xor g1578 (n_143, n_1667, n_583);
  nand g1579 (n_1668, n_581, n_582);
  nand g1580 (n_1669, n_583, n_582);
  nand g1581 (n_1670, n_581, n_583);
  nand g1582 (n_76, n_1668, n_1669, n_1670);
  xor g1584 (n_586, n_1543, A[23]);
  nand g1587 (n_1674, A[33], A[23]);
  nand g1588 (n_598, n_1544, n_1618, n_1674);
  xor g1589 (n_1675, A[21], A[29]);
  xor g1590 (n_589, n_1675, A[19]);
  nand g1592 (n_1677, A[19], A[29]);
  nand g1594 (n_599, n_1609, n_1677, n_1160);
  xor g1596 (n_588, n_1351, A[35]);
  nand g1598 (n_1681, A[35], A[25]);
  nand g1599 (n_1682, A[27], A[35]);
  nand g1600 (n_601, n_1352, n_1681, n_1682);
  xor g1601 (n_1683, A[37], n_584);
  xor g1602 (n_592, n_1683, n_585);
  nand g1603 (n_1684, A[37], n_584);
  nand g1604 (n_1685, n_585, n_584);
  nand g1605 (n_1686, A[37], n_585);
  nand g1606 (n_604, n_1684, n_1685, n_1686);
  xor g1607 (n_1687, n_586, n_587);
  xor g1608 (n_593, n_1687, n_588);
  nand g1609 (n_1688, n_586, n_587);
  nand g1610 (n_1689, n_588, n_587);
  nand g1611 (n_1690, n_586, n_588);
  nand g1612 (n_605, n_1688, n_1689, n_1690);
  xor g1613 (n_1691, n_589, n_590);
  xor g1614 (n_594, n_1691, n_591);
  nand g1615 (n_1692, n_589, n_590);
  nand g1616 (n_1693, n_591, n_590);
  nand g1617 (n_1694, n_589, n_591);
  nand g1618 (n_609, n_1692, n_1693, n_1694);
  xor g1619 (n_1695, n_592, n_593);
  xor g1620 (n_596, n_1695, n_594);
  nand g1621 (n_1696, n_592, n_593);
  nand g1622 (n_1697, n_594, n_593);
  nand g1623 (n_1698, n_592, n_594);
  nand g1624 (n_611, n_1696, n_1697, n_1698);
  xor g1625 (n_1699, n_595, n_596);
  xor g1626 (n_142, n_1699, n_597);
  nand g1627 (n_1700, n_595, n_596);
  nand g1628 (n_1701, n_597, n_596);
  nand g1629 (n_1702, n_595, n_597);
  nand g1630 (n_75, n_1700, n_1701, n_1702);
  xor g1632 (n_600, n_1511, A[24]);
  nand g1635 (n_1706, A[32], A[24]);
  nand g1636 (n_612, n_1512, n_1450, n_1706);
  xor g1638 (n_602, n_1191, A[28]);
  nand g1642 (n_613, n_1192, n_1577, n_1386);
  xor g1643 (n_1711, A[26], A[36]);
  xor g1644 (n_603, n_1711, A[38]);
  nand g1645 (n_1712, A[26], A[36]);
  nand g1646 (n_1713, A[38], A[36]);
  nand g1647 (n_1714, A[26], A[38]);
  nand g1648 (n_615, n_1712, n_1713, n_1714);
  xor g1649 (n_1715, A[34], n_598);
  xor g1650 (n_606, n_1715, n_599);
  nand g1651 (n_1716, A[34], n_598);
  nand g1652 (n_1717, n_599, n_598);
  nand g1653 (n_1718, A[34], n_599);
  nand g1654 (n_618, n_1716, n_1717, n_1718);
  xor g1655 (n_1719, n_600, n_601);
  xor g1656 (n_607, n_1719, n_602);
  nand g1657 (n_1720, n_600, n_601);
  nand g1658 (n_1721, n_602, n_601);
  nand g1659 (n_1722, n_600, n_602);
  nand g1660 (n_619, n_1720, n_1721, n_1722);
  xor g1661 (n_1723, n_603, n_604);
  xor g1662 (n_608, n_1723, n_605);
  nand g1663 (n_1724, n_603, n_604);
  nand g1664 (n_1725, n_605, n_604);
  nand g1665 (n_1726, n_603, n_605);
  nand g1666 (n_623, n_1724, n_1725, n_1726);
  xor g1667 (n_1727, n_606, n_607);
  xor g1668 (n_610, n_1727, n_608);
  nand g1669 (n_1728, n_606, n_607);
  nand g1670 (n_1729, n_608, n_607);
  nand g1671 (n_1730, n_606, n_608);
  nand g1672 (n_625, n_1728, n_1729, n_1730);
  xor g1673 (n_1731, n_609, n_610);
  xor g1674 (n_141, n_1731, n_611);
  nand g1675 (n_1732, n_609, n_610);
  nand g1676 (n_1733, n_611, n_610);
  nand g1677 (n_1734, n_609, n_611);
  nand g1678 (n_74, n_1732, n_1733, n_1734);
  xor g1680 (n_614, n_1543, A[25]);
  nand g1683 (n_1738, A[33], A[25]);
  nand g1684 (n_626, n_1544, n_1482, n_1738);
  xor g1686 (n_616, n_1223, A[29]);
  nand g1690 (n_627, n_1224, n_1609, n_1418);
  xor g1691 (n_1743, A[27], A[37]);
  xor g1692 (n_617, n_1743, A[39]);
  nand g1693 (n_1744, A[27], A[37]);
  nand g1694 (n_1745, A[39], A[37]);
  nand g1695 (n_1746, A[27], A[39]);
  nand g1696 (n_629, n_1744, n_1745, n_1746);
  xor g1697 (n_1747, A[35], n_612);
  xor g1698 (n_620, n_1747, n_613);
  nand g1699 (n_1748, A[35], n_612);
  nand g1700 (n_1749, n_613, n_612);
  nand g1701 (n_1750, A[35], n_613);
  nand g1702 (n_632, n_1748, n_1749, n_1750);
  xor g1703 (n_1751, n_614, n_615);
  xor g1704 (n_621, n_1751, n_616);
  nand g1705 (n_1752, n_614, n_615);
  nand g1706 (n_1753, n_616, n_615);
  nand g1707 (n_1754, n_614, n_616);
  nand g1708 (n_633, n_1752, n_1753, n_1754);
  xor g1709 (n_1755, n_617, n_618);
  xor g1710 (n_622, n_1755, n_619);
  nand g1711 (n_1756, n_617, n_618);
  nand g1712 (n_1757, n_619, n_618);
  nand g1713 (n_1758, n_617, n_619);
  nand g1714 (n_637, n_1756, n_1757, n_1758);
  xor g1715 (n_1759, n_620, n_621);
  xor g1716 (n_624, n_1759, n_622);
  nand g1717 (n_1760, n_620, n_621);
  nand g1718 (n_1761, n_622, n_621);
  nand g1719 (n_1762, n_620, n_622);
  nand g1720 (n_639, n_1760, n_1761, n_1762);
  xor g1721 (n_1763, n_623, n_624);
  xor g1722 (n_140, n_1763, n_625);
  nand g1723 (n_1764, n_623, n_624);
  nand g1724 (n_1765, n_625, n_624);
  nand g1725 (n_1766, n_623, n_625);
  nand g1726 (n_73, n_1764, n_1765, n_1766);
  xor g1727 (n_1767, A[32], A[26]);
  xor g1728 (n_628, n_1767, A[24]);
  nand g1732 (n_640, n_1514, n_1320, n_1706);
  xor g1733 (n_1771, A[22], A[30]);
  xor g1734 (n_630, n_1771, A[28]);
  nand g1738 (n_641, n_1586, n_1448, n_1386);
  xor g1739 (n_1775, A[34], A[40]);
  xor g1740 (n_631, n_1775, A[38]);
  nand g1741 (n_1776, A[34], A[40]);
  nand g1742 (n_1777, A[38], A[40]);
  nand g1743 (n_1778, A[34], A[38]);
  nand g1744 (n_643, n_1776, n_1777, n_1778);
  xor g1745 (n_1779, A[36], n_626);
  xor g1746 (n_634, n_1779, n_627);
  nand g1747 (n_1780, A[36], n_626);
  nand g1748 (n_1781, n_627, n_626);
  nand g1749 (n_1782, A[36], n_627);
  nand g1750 (n_646, n_1780, n_1781, n_1782);
  xor g1751 (n_1783, n_628, n_629);
  xor g1752 (n_635, n_1783, n_630);
  nand g1753 (n_1784, n_628, n_629);
  nand g1754 (n_1785, n_630, n_629);
  nand g1755 (n_1786, n_628, n_630);
  nand g1756 (n_647, n_1784, n_1785, n_1786);
  xor g1757 (n_1787, n_631, n_632);
  xor g1758 (n_636, n_1787, n_633);
  nand g1759 (n_1788, n_631, n_632);
  nand g1760 (n_1789, n_633, n_632);
  nand g1761 (n_1790, n_631, n_633);
  nand g1762 (n_651, n_1788, n_1789, n_1790);
  xor g1763 (n_1791, n_634, n_635);
  xor g1764 (n_638, n_1791, n_636);
  nand g1765 (n_1792, n_634, n_635);
  nand g1766 (n_1793, n_636, n_635);
  nand g1767 (n_1794, n_634, n_636);
  nand g1768 (n_653, n_1792, n_1793, n_1794);
  xor g1769 (n_1795, n_637, n_638);
  xor g1770 (n_139, n_1795, n_639);
  nand g1771 (n_1796, n_637, n_638);
  nand g1772 (n_1797, n_639, n_638);
  nand g1773 (n_1798, n_637, n_639);
  nand g1774 (n_72, n_1796, n_1797, n_1798);
  xor g1775 (n_1799, A[33], A[27]);
  xor g1776 (n_642, n_1799, A[25]);
  nand g1780 (n_654, n_1546, n_1352, n_1738);
  xor g1781 (n_1803, A[23], A[31]);
  xor g1782 (n_644, n_1803, A[29]);
  nand g1786 (n_655, n_1618, n_1480, n_1418);
  xor g1787 (n_1807, A[35], A[41]);
  xor g1788 (n_645, n_1807, A[39]);
  nand g1789 (n_1808, A[35], A[41]);
  nand g1790 (n_1809, A[39], A[41]);
  nand g1791 (n_1810, A[35], A[39]);
  nand g1792 (n_658, n_1808, n_1809, n_1810);
  xor g1793 (n_1811, A[37], n_640);
  xor g1794 (n_648, n_1811, n_641);
  nand g1795 (n_1812, A[37], n_640);
  nand g1796 (n_1813, n_641, n_640);
  nand g1797 (n_1814, A[37], n_641);
  nand g1798 (n_660, n_1812, n_1813, n_1814);
  xor g1799 (n_1815, n_642, n_643);
  xor g1800 (n_649, n_1815, n_644);
  nand g1801 (n_1816, n_642, n_643);
  nand g1802 (n_1817, n_644, n_643);
  nand g1803 (n_1818, n_642, n_644);
  nand g1804 (n_661, n_1816, n_1817, n_1818);
  xor g1805 (n_1819, n_645, n_646);
  xor g1806 (n_650, n_1819, n_647);
  nand g1807 (n_1820, n_645, n_646);
  nand g1808 (n_1821, n_647, n_646);
  nand g1809 (n_1822, n_645, n_647);
  nand g1810 (n_665, n_1820, n_1821, n_1822);
  xor g1811 (n_1823, n_648, n_649);
  xor g1812 (n_652, n_1823, n_650);
  nand g1813 (n_1824, n_648, n_649);
  nand g1814 (n_1825, n_650, n_649);
  nand g1815 (n_1826, n_648, n_650);
  nand g1816 (n_667, n_1824, n_1825, n_1826);
  xor g1817 (n_1827, n_651, n_652);
  xor g1818 (n_138, n_1827, n_653);
  nand g1819 (n_1828, n_651, n_652);
  nand g1820 (n_1829, n_653, n_652);
  nand g1821 (n_1830, n_651, n_653);
  nand g1822 (n_71, n_1828, n_1829, n_1830);
  xor g1824 (n_656, n_1575, A[26]);
  nand g1828 (n_668, n_1576, n_1384, n_1514);
  xor g1830 (n_657, n_1583, A[36]);
  nand g1832 (n_1837, A[36], A[30]);
  nand g1833 (n_1838, A[24], A[36]);
  nand g1834 (n_671, n_1450, n_1837, n_1838);
  xor g1841 (n_1843, A[42], n_654);
  xor g1842 (n_662, n_1843, n_655);
  nand g1843 (n_1844, A[42], n_654);
  nand g1844 (n_1845, n_655, n_654);
  nand g1845 (n_1846, A[42], n_655);
  nand g1846 (n_674, n_1844, n_1845, n_1846);
  xor g1847 (n_1847, n_656, n_657);
  xor g1848 (n_663, n_1847, n_658);
  nand g1849 (n_1848, n_656, n_657);
  nand g1850 (n_1849, n_658, n_657);
  nand g1851 (n_1850, n_656, n_658);
  nand g1852 (n_675, n_1848, n_1849, n_1850);
  xor g1853 (n_1851, n_631, n_660);
  xor g1854 (n_664, n_1851, n_661);
  nand g1855 (n_1852, n_631, n_660);
  nand g1856 (n_1853, n_661, n_660);
  nand g1857 (n_1854, n_631, n_661);
  nand g1858 (n_679, n_1852, n_1853, n_1854);
  xor g1859 (n_1855, n_662, n_663);
  xor g1860 (n_666, n_1855, n_664);
  nand g1861 (n_1856, n_662, n_663);
  nand g1862 (n_1857, n_664, n_663);
  nand g1863 (n_1858, n_662, n_664);
  nand g1864 (n_681, n_1856, n_1857, n_1858);
  xor g1865 (n_1859, n_665, n_666);
  xor g1866 (n_137, n_1859, n_667);
  nand g1867 (n_1860, n_665, n_666);
  nand g1868 (n_1861, n_667, n_666);
  nand g1869 (n_1862, n_665, n_667);
  nand g1870 (n_70, n_1860, n_1861, n_1862);
  xor g1872 (n_669, n_1607, A[27]);
  nand g1876 (n_682, n_1608, n_1416, n_1546);
  xor g1878 (n_670, n_1615, A[37]);
  nand g1880 (n_1869, A[37], A[31]);
  nand g1881 (n_1870, A[25], A[37]);
  nand g1882 (n_684, n_1482, n_1869, n_1870);
  xor g1889 (n_1875, A[43], n_668);
  xor g1890 (n_676, n_1875, n_669);
  nand g1891 (n_1876, A[43], n_668);
  nand g1892 (n_1877, n_669, n_668);
  nand g1893 (n_1878, A[43], n_669);
  nand g1894 (n_689, n_1876, n_1877, n_1878);
  xor g1895 (n_1879, n_670, n_671);
  xor g1896 (n_677, n_1879, n_643);
  nand g1897 (n_1880, n_670, n_671);
  nand g1898 (n_1881, n_643, n_671);
  nand g1899 (n_1882, n_670, n_643);
  nand g1900 (n_688, n_1880, n_1881, n_1882);
  xor g1901 (n_1883, n_645, n_674);
  xor g1902 (n_678, n_1883, n_675);
  nand g1903 (n_1884, n_645, n_674);
  nand g1904 (n_1885, n_675, n_674);
  nand g1905 (n_1886, n_645, n_675);
  nand g1906 (n_692, n_1884, n_1885, n_1886);
  xor g1907 (n_1887, n_676, n_677);
  xor g1908 (n_680, n_1887, n_678);
  nand g1909 (n_1888, n_676, n_677);
  nand g1910 (n_1889, n_678, n_677);
  nand g1911 (n_1890, n_676, n_678);
  nand g1912 (n_695, n_1888, n_1889, n_1890);
  xor g1913 (n_1891, n_679, n_680);
  xor g1914 (n_136, n_1891, n_681);
  nand g1915 (n_1892, n_679, n_680);
  nand g1916 (n_1893, n_681, n_680);
  nand g1917 (n_1894, n_679, n_681);
  nand g1918 (n_69, n_1892, n_1893, n_1894);
  xor g1920 (n_683, n_1511, A[28]);
  nand g1924 (n_696, n_1512, n_1448, n_1576);
  xor g1925 (n_1899, A[26], A[38]);
  xor g1926 (n_687, n_1899, A[42]);
  nand g1928 (n_1901, A[42], A[38]);
  nand g1929 (n_1902, A[26], A[42]);
  nand g1930 (n_698, n_1714, n_1901, n_1902);
  xor g1931 (n_1903, A[36], A[44]);
  xor g1932 (n_686, n_1903, A[34]);
  nand g1933 (n_1904, A[36], A[44]);
  nand g1934 (n_1905, A[34], A[44]);
  nand g1935 (n_1906, A[36], A[34]);
  nand g1936 (n_699, n_1904, n_1905, n_1906);
  xor g1937 (n_1907, A[40], n_682);
  xor g1938 (n_690, n_1907, n_683);
  nand g1939 (n_1908, A[40], n_682);
  nand g1940 (n_1909, n_683, n_682);
  nand g1941 (n_1910, A[40], n_683);
  nand g1942 (n_702, n_1908, n_1909, n_1910);
  xor g1943 (n_1911, n_684, n_658);
  xor g1944 (n_691, n_1911, n_686);
  nand g1945 (n_1912, n_684, n_658);
  nand g1946 (n_1913, n_686, n_658);
  nand g1947 (n_1914, n_684, n_686);
  nand g1948 (n_705, n_1912, n_1913, n_1914);
  xor g1949 (n_1915, n_687, n_688);
  xor g1950 (n_693, n_1915, n_689);
  nand g1951 (n_1916, n_687, n_688);
  nand g1952 (n_1917, n_689, n_688);
  nand g1953 (n_1918, n_687, n_689);
  nand g1954 (n_706, n_1916, n_1917, n_1918);
  xor g1955 (n_1919, n_690, n_691);
  xor g1956 (n_694, n_1919, n_692);
  nand g1957 (n_1920, n_690, n_691);
  nand g1958 (n_1921, n_692, n_691);
  nand g1959 (n_1922, n_690, n_692);
  nand g1960 (n_709, n_1920, n_1921, n_1922);
  xor g1961 (n_1923, n_693, n_694);
  xor g1962 (n_135, n_1923, n_695);
  nand g1963 (n_1924, n_693, n_694);
  nand g1964 (n_1925, n_695, n_694);
  nand g1965 (n_1926, n_693, n_695);
  nand g1966 (n_68, n_1924, n_1925, n_1926);
  xor g1968 (n_697, n_1543, A[29]);
  nand g1972 (n_712, n_1544, n_1480, n_1608);
  xor g1973 (n_1931, A[27], A[39]);
  xor g1974 (n_701, n_1931, A[43]);
  nand g1976 (n_1933, A[43], A[39]);
  nand g1977 (n_1934, A[27], A[43]);
  nand g1978 (n_715, n_1746, n_1933, n_1934);
  xor g1979 (n_1935, A[37], A[45]);
  xor g1980 (n_700, n_1935, A[35]);
  nand g1981 (n_1936, A[37], A[45]);
  nand g1982 (n_1937, A[35], A[45]);
  nand g1983 (n_1938, A[37], A[35]);
  nand g1984 (n_713, n_1936, n_1937, n_1938);
  xor g1985 (n_1939, A[41], n_696);
  xor g1986 (n_703, n_1939, n_697);
  nand g1987 (n_1940, A[41], n_696);
  nand g1988 (n_1941, n_697, n_696);
  nand g1989 (n_1942, A[41], n_697);
  nand g1990 (n_718, n_1940, n_1941, n_1942);
  xor g1991 (n_1943, n_698, n_699);
  xor g1992 (n_704, n_1943, n_700);
  nand g1993 (n_1944, n_698, n_699);
  nand g1994 (n_1945, n_700, n_699);
  nand g1995 (n_1946, n_698, n_700);
  nand g1996 (n_720, n_1944, n_1945, n_1946);
  xor g1997 (n_1947, n_701, n_702);
  xor g1998 (n_707, n_1947, n_703);
  nand g1999 (n_1948, n_701, n_702);
  nand g2000 (n_1949, n_703, n_702);
  nand g2001 (n_1950, n_701, n_703);
  nand g2002 (n_722, n_1948, n_1949, n_1950);
  xor g2003 (n_1951, n_704, n_705);
  xor g2004 (n_708, n_1951, n_706);
  nand g2005 (n_1952, n_704, n_705);
  nand g2006 (n_1953, n_706, n_705);
  nand g2007 (n_1954, n_704, n_706);
  nand g2008 (n_725, n_1952, n_1953, n_1954);
  xor g2009 (n_1955, n_707, n_708);
  xor g2010 (n_134, n_1955, n_709);
  nand g2011 (n_1956, n_707, n_708);
  nand g2012 (n_1957, n_709, n_708);
  nand g2013 (n_1958, n_707, n_709);
  nand g2014 (n_67, n_1956, n_1957, n_1958);
  xor g2017 (n_1959, A[46], A[30]);
  xor g2018 (n_714, n_1959, A[32]);
  nand g2019 (n_1960, A[46], A[30]);
  nand g2021 (n_1962, A[46], A[32]);
  nand g2022 (n_729, n_1960, n_1512, n_1962);
  xor g2023 (n_1963, A[28], A[44]);
  xor g2024 (n_716, n_1963, A[40]);
  nand g2025 (n_1964, A[28], A[44]);
  nand g2026 (n_1965, A[40], A[44]);
  nand g2027 (n_1966, A[28], A[40]);
  nand g2028 (n_732, n_1964, n_1965, n_1966);
  xor g2029 (n_1967, A[38], A[42]);
  xor g2030 (n_717, n_1967, A[36]);
  nand g2032 (n_1969, A[36], A[42]);
  nand g2034 (n_730, n_1901, n_1969, n_1713);
  xor g2035 (n_1971, A[34], n_712);
  xor g2036 (n_719, n_1971, n_713);
  nand g2037 (n_1972, A[34], n_712);
  nand g2038 (n_1973, n_713, n_712);
  nand g2039 (n_1974, A[34], n_713);
  nand g2040 (n_735, n_1972, n_1973, n_1974);
  xor g2041 (n_1975, n_714, n_715);
  xor g2042 (n_721, n_1975, n_716);
  nand g2043 (n_1976, n_714, n_715);
  nand g2044 (n_1977, n_716, n_715);
  nand g2045 (n_1978, n_714, n_716);
  nand g2046 (n_737, n_1976, n_1977, n_1978);
  xor g2047 (n_1979, n_717, n_718);
  xor g2048 (n_723, n_1979, n_719);
  nand g2049 (n_1980, n_717, n_718);
  nand g2050 (n_1981, n_719, n_718);
  nand g2051 (n_1982, n_717, n_719);
  nand g2052 (n_739, n_1980, n_1981, n_1982);
  xor g2053 (n_1983, n_720, n_721);
  xor g2054 (n_724, n_1983, n_722);
  nand g2055 (n_1984, n_720, n_721);
  nand g2056 (n_1985, n_722, n_721);
  nand g2057 (n_1986, n_720, n_722);
  nand g2058 (n_742, n_1984, n_1985, n_1986);
  xor g2059 (n_1987, n_723, n_724);
  xor g2060 (n_133, n_1987, n_725);
  nand g2061 (n_1988, n_723, n_724);
  nand g2062 (n_1989, n_725, n_724);
  nand g2063 (n_1990, n_723, n_725);
  nand g2064 (n_66, n_1988, n_1989, n_1990);
  xor g2068 (n_731, n_1607, A[31]);
  xor g2073 (n_1995, A[39], A[43]);
  xor g2074 (n_733, n_1995, A[46]);
  nand g2076 (n_1997, A[46], A[43]);
  nand g2077 (n_1998, A[39], A[46]);
  nand g2078 (n_746, n_1933, n_1997, n_1998);
  xor g2085 (n_2003, A[41], n_729);
  xor g2086 (n_736, n_2003, n_730);
  nand g2087 (n_2004, A[41], n_729);
  nand g2088 (n_2005, n_730, n_729);
  nand g2089 (n_2006, A[41], n_730);
  nand g2090 (n_750, n_2004, n_2005, n_2006);
  xor g2091 (n_2007, n_731, n_732);
  xor g2092 (n_738, n_2007, n_733);
  nand g2093 (n_2008, n_731, n_732);
  nand g2094 (n_2009, n_733, n_732);
  nand g2095 (n_2010, n_731, n_733);
  nand g2096 (n_753, n_2008, n_2009, n_2010);
  xor g2097 (n_2011, n_700, n_735);
  xor g2098 (n_740, n_2011, n_736);
  nand g2099 (n_2012, n_700, n_735);
  nand g2100 (n_2013, n_736, n_735);
  nand g2101 (n_2014, n_700, n_736);
  nand g2102 (n_754, n_2012, n_2013, n_2014);
  xor g2103 (n_2015, n_737, n_738);
  xor g2104 (n_741, n_2015, n_739);
  nand g2105 (n_2016, n_737, n_738);
  nand g2106 (n_2017, n_739, n_738);
  nand g2107 (n_2018, n_737, n_739);
  nand g2108 (n_757, n_2016, n_2017, n_2018);
  xor g2109 (n_2019, n_740, n_741);
  xor g2110 (n_132, n_2019, n_742);
  nand g2111 (n_2020, n_740, n_741);
  nand g2112 (n_2021, n_742, n_741);
  nand g2113 (n_2022, n_740, n_742);
  nand g2114 (n_65, n_2020, n_2021, n_2022);
  xor g2116 (n_745, n_2023, A[30]);
  nand g2120 (n_760, n_2024, n_1512, n_2026);
  xor g2121 (n_2027, A[40], A[44]);
  xor g2122 (n_749, n_2027, A[38]);
  nand g2124 (n_2029, A[38], A[44]);
  nand g2126 (n_761, n_1965, n_2029, n_1777);
  xor g2128 (n_748, n_2031, A[36]);
  nand g2132 (n_762, n_2032, n_1969, n_2034);
  xor g2134 (n_751, n_1971, n_745);
  nand g2136 (n_2037, n_745, n_712);
  nand g2137 (n_2038, A[34], n_745);
  nand g2138 (n_766, n_1972, n_2037, n_2038);
  xor g2139 (n_2039, n_746, n_713);
  xor g2140 (n_752, n_2039, n_748);
  nand g2141 (n_2040, n_746, n_713);
  nand g2142 (n_2041, n_748, n_713);
  nand g2143 (n_2042, n_746, n_748);
  nand g2144 (n_768, n_2040, n_2041, n_2042);
  xor g2145 (n_2043, n_749, n_750);
  xor g2146 (n_755, n_2043, n_751);
  nand g2147 (n_2044, n_749, n_750);
  nand g2148 (n_2045, n_751, n_750);
  nand g2149 (n_2046, n_749, n_751);
  nand g2150 (n_770, n_2044, n_2045, n_2046);
  xor g2151 (n_2047, n_752, n_753);
  xor g2152 (n_756, n_2047, n_754);
  nand g2153 (n_2048, n_752, n_753);
  nand g2154 (n_2049, n_754, n_753);
  nand g2155 (n_2050, n_752, n_754);
  nand g2156 (n_772, n_2048, n_2049, n_2050);
  xor g2157 (n_2051, n_755, n_756);
  xor g2158 (n_131, n_2051, n_757);
  nand g2159 (n_2052, n_755, n_756);
  nand g2160 (n_2053, n_757, n_756);
  nand g2161 (n_2054, n_755, n_757);
  nand g2162 (n_64, n_2052, n_2053, n_2054);
  xor g2165 (n_2055, A[31], A[39]);
  xor g2166 (n_764, n_2055, A[43]);
  nand g2167 (n_2056, A[31], A[39]);
  nand g2169 (n_2058, A[31], A[43]);
  nand g2170 (n_776, n_2056, n_1933, n_2058);
  xor g2178 (n_765, n_2063, n_760);
  nand g2181 (n_2066, A[41], n_760);
  nand g2182 (n_779, n_2064, n_2065, n_2066);
  xor g2183 (n_2067, n_761, n_762);
  xor g2184 (n_767, n_2067, n_700);
  nand g2185 (n_2068, n_761, n_762);
  nand g2186 (n_2069, n_700, n_762);
  nand g2187 (n_2070, n_761, n_700);
  nand g2188 (n_781, n_2068, n_2069, n_2070);
  xor g2189 (n_2071, n_764, n_765);
  xor g2190 (n_769, n_2071, n_766);
  nand g2191 (n_2072, n_764, n_765);
  nand g2192 (n_2073, n_766, n_765);
  nand g2193 (n_2074, n_764, n_766);
  nand g2194 (n_783, n_2072, n_2073, n_2074);
  xor g2195 (n_2075, n_767, n_768);
  xor g2196 (n_771, n_2075, n_769);
  nand g2197 (n_2076, n_767, n_768);
  nand g2198 (n_2077, n_769, n_768);
  nand g2199 (n_2078, n_767, n_769);
  nand g2200 (n_785, n_2076, n_2077, n_2078);
  xor g2201 (n_2079, n_770, n_771);
  xor g2202 (n_130, n_2079, n_772);
  nand g2203 (n_2080, n_770, n_771);
  nand g2204 (n_2081, n_772, n_771);
  nand g2205 (n_2082, n_770, n_772);
  nand g2206 (n_63, n_2080, n_2081, n_2082);
  xor g2208 (n_775, n_2023, A[44]);
  nand g2210 (n_2085, A[44], A[32]);
  nand g2212 (n_788, n_2024, n_2085, n_2086);
  xor g2213 (n_2087, A[40], A[38]);
  xor g2214 (n_778, n_2087, A[42]);
  nand g2217 (n_2090, A[40], A[42]);
  nand g2218 (n_789, n_1777, n_1901, n_2090);
  xor g2219 (n_2091, A[36], A[34]);
  xor g2220 (n_777, n_2091, A[33]);
  nand g2222 (n_2093, A[33], A[34]);
  nand g2223 (n_2094, A[36], A[33]);
  nand g2224 (n_791, n_1906, n_2093, n_2094);
  xor g2225 (n_2095, n_713, n_775);
  xor g2226 (n_780, n_2095, n_776);
  nand g2227 (n_2096, n_713, n_775);
  nand g2228 (n_2097, n_776, n_775);
  nand g2229 (n_2098, n_713, n_776);
  nand g2230 (n_793, n_2096, n_2097, n_2098);
  xor g2231 (n_2099, n_777, n_778);
  xor g2232 (n_782, n_2099, n_779);
  nand g2233 (n_2100, n_777, n_778);
  nand g2234 (n_2101, n_779, n_778);
  nand g2235 (n_2102, n_777, n_779);
  nand g2236 (n_795, n_2100, n_2101, n_2102);
  xor g2237 (n_2103, n_780, n_781);
  xor g2238 (n_784, n_2103, n_782);
  nand g2239 (n_2104, n_780, n_781);
  nand g2240 (n_2105, n_782, n_781);
  nand g2241 (n_2106, n_780, n_782);
  nand g2242 (n_798, n_2104, n_2105, n_2106);
  xor g2243 (n_2107, n_783, n_784);
  xor g2244 (n_129, n_2107, n_785);
  nand g2245 (n_2108, n_783, n_784);
  nand g2246 (n_2109, n_785, n_784);
  nand g2247 (n_2110, n_783, n_785);
  nand g2248 (n_62, n_2108, n_2109, n_2110);
  xor g2252 (n_792, n_1995, A[37]);
  nand g2255 (n_2114, A[43], A[37]);
  nand g2256 (n_800, n_1933, n_1745, n_2114);
  xor g2257 (n_2115, A[45], A[35]);
  xor g2258 (n_790, n_2115, A[41]);
  nand g2261 (n_2118, A[45], A[41]);
  nand g2262 (n_801, n_1937, n_1808, n_2118);
  xor g2264 (n_794, n_2119, n_789);
  nand g2266 (n_2121, n_789, n_788);
  nand g2268 (n_805, n_2120, n_2121, n_2122);
  xor g2269 (n_2123, n_790, n_791);
  xor g2270 (n_796, n_2123, n_792);
  nand g2271 (n_2124, n_790, n_791);
  nand g2272 (n_2125, n_792, n_791);
  nand g2273 (n_2126, n_790, n_792);
  nand g2274 (n_806, n_2124, n_2125, n_2126);
  xor g2275 (n_2127, n_793, n_794);
  xor g2276 (n_797, n_2127, n_795);
  nand g2277 (n_2128, n_793, n_794);
  nand g2278 (n_2129, n_795, n_794);
  nand g2279 (n_2130, n_793, n_795);
  nand g2280 (n_809, n_2128, n_2129, n_2130);
  xor g2281 (n_2131, n_796, n_797);
  xor g2282 (n_128, n_2131, n_798);
  nand g2283 (n_2132, n_796, n_797);
  nand g2284 (n_2133, n_798, n_797);
  nand g2285 (n_2134, n_796, n_798);
  nand g2286 (n_61, n_2132, n_2133, n_2134);
  xor g2288 (n_803, n_2135, A[40]);
  nand g2292 (n_813, n_2086, n_1965, n_2138);
  xor g2299 (n_2143, A[34], A[33]);
  xor g2300 (n_804, n_2143, n_800);
  nand g2302 (n_2145, n_800, A[33]);
  nand g2303 (n_2146, A[34], n_800);
  nand g2304 (n_816, n_2093, n_2145, n_2146);
  xor g2305 (n_2147, n_801, n_717);
  xor g2306 (n_807, n_2147, n_803);
  nand g2307 (n_2148, n_801, n_717);
  nand g2308 (n_2149, n_803, n_717);
  nand g2309 (n_2150, n_801, n_803);
  nand g2310 (n_817, n_2148, n_2149, n_2150);
  xor g2311 (n_2151, n_804, n_805);
  xor g2312 (n_808, n_2151, n_806);
  nand g2313 (n_2152, n_804, n_805);
  nand g2314 (n_2153, n_806, n_805);
  nand g2315 (n_2154, n_804, n_806);
  nand g2316 (n_820, n_2152, n_2153, n_2154);
  xor g2317 (n_2155, n_807, n_808);
  xor g2318 (n_127, n_2155, n_809);
  nand g2319 (n_2156, n_807, n_808);
  nand g2320 (n_2157, n_809, n_808);
  nand g2321 (n_2158, n_807, n_809);
  nand g2322 (n_60, n_2156, n_2157, n_2158);
  xor g2325 (n_2159, A[39], A[37]);
  xor g2326 (n_814, n_2159, A[45]);
  nand g2329 (n_2162, A[39], A[45]);
  nand g2330 (n_822, n_1745, n_1936, n_2162);
  nand g2336 (n_825, n_1808, n_2165, n_2166);
  xor g2337 (n_2167, n_730, n_813);
  xor g2338 (n_818, n_2167, n_814);
  nand g2339 (n_2168, n_730, n_813);
  nand g2340 (n_2169, n_814, n_813);
  nand g2341 (n_2170, n_730, n_814);
  nand g2342 (n_827, n_2168, n_2169, n_2170);
  xor g2343 (n_2171, n_815, n_816);
  xor g2344 (n_819, n_2171, n_817);
  nand g2345 (n_2172, n_815, n_816);
  nand g2346 (n_2173, n_817, n_816);
  nand g2347 (n_2174, n_815, n_817);
  nand g2348 (n_829, n_2172, n_2173, n_2174);
  xor g2349 (n_2175, n_818, n_819);
  xor g2350 (n_126, n_2175, n_820);
  nand g2351 (n_2176, n_818, n_819);
  nand g2352 (n_2177, n_820, n_819);
  nand g2353 (n_2178, n_818, n_820);
  nand g2354 (n_59, n_2176, n_2177, n_2178);
  xor g2367 (n_2187, A[43], n_822);
  xor g2368 (n_826, n_2187, n_717);
  nand g2369 (n_2188, A[43], n_822);
  nand g2370 (n_2189, n_717, n_822);
  nand g2371 (n_2190, A[43], n_717);
  nand g2372 (n_836, n_2188, n_2189, n_2190);
  xor g2373 (n_2191, n_803, n_825);
  xor g2374 (n_828, n_2191, n_826);
  nand g2375 (n_2192, n_803, n_825);
  nand g2376 (n_2193, n_826, n_825);
  nand g2377 (n_2194, n_803, n_826);
  nand g2378 (n_838, n_2192, n_2193, n_2194);
  xor g2379 (n_2195, n_827, n_828);
  xor g2380 (n_125, n_2195, n_829);
  nand g2381 (n_2196, n_827, n_828);
  nand g2382 (n_2197, n_829, n_828);
  nand g2383 (n_2198, n_827, n_829);
  nand g2384 (n_58, n_2196, n_2197, n_2198);
  nand g2398 (n_843, n_2165, n_2205, n_2006);
  xor g2399 (n_2207, n_813, n_814);
  xor g2400 (n_837, n_2207, n_835);
  nand g2402 (n_2209, n_835, n_814);
  nand g2403 (n_2210, n_813, n_835);
  nand g2404 (n_845, n_2169, n_2209, n_2210);
  xor g2405 (n_2211, n_836, n_837);
  xor g2406 (n_124, n_2211, n_838);
  nand g2407 (n_2212, n_836, n_837);
  nand g2408 (n_2213, n_838, n_837);
  nand g2409 (n_2214, n_836, n_838);
  nand g2410 (n_123, n_2212, n_2213, n_2214);
  xor g2418 (n_842, n_1967, A[43]);
  nand g2420 (n_2221, A[43], A[42]);
  nand g2421 (n_2222, A[38], A[43]);
  nand g2422 (n_850, n_1901, n_2221, n_2222);
  xor g2423 (n_2223, n_822, n_803);
  xor g2424 (n_844, n_2223, n_842);
  nand g2425 (n_2224, n_822, n_803);
  nand g2426 (n_2225, n_842, n_803);
  nand g2427 (n_2226, n_822, n_842);
  nand g2428 (n_852, n_2224, n_2225, n_2226);
  xor g2429 (n_2227, n_843, n_844);
  xor g2430 (n_57, n_2227, n_845);
  nand g2431 (n_2228, n_843, n_844);
  nand g2432 (n_2229, n_845, n_844);
  nand g2433 (n_2230, n_843, n_845);
  nand g2434 (n_122, n_2228, n_2229, n_2230);
  xor g2438 (n_849, n_1995, A[41]);
  nand g2440 (n_2233, A[41], A[43]);
  nand g2442 (n_854, n_1933, n_2233, n_1809);
  xor g2444 (n_851, n_2235, n_849);
  nand g2446 (n_2237, n_849, n_813);
  nand g2448 (n_857, n_2236, n_2237, n_2238);
  xor g2449 (n_2239, n_850, n_851);
  xor g2450 (n_56, n_2239, n_852);
  nand g2451 (n_2240, n_850, n_851);
  nand g2452 (n_2241, n_852, n_851);
  nand g2453 (n_2242, n_850, n_852);
  nand g2454 (n_121, n_2240, n_2241, n_2242);
  xor g2461 (n_2247, A[42], A[45]);
  xor g2462 (n_856, n_2247, n_854);
  nand g2463 (n_2248, A[42], A[45]);
  nand g2464 (n_2249, n_854, A[45]);
  nand g2465 (n_2250, A[42], n_854);
  nand g2466 (n_862, n_2248, n_2249, n_2250);
  xor g2467 (n_2251, n_803, n_856);
  xor g2468 (n_55, n_2251, n_857);
  nand g2469 (n_2252, n_803, n_856);
  nand g2470 (n_2253, n_857, n_856);
  nand g2471 (n_2254, n_803, n_857);
  nand g2472 (n_120, n_2252, n_2253, n_2254);
  xor g2475 (n_2255, A[43], A[41]);
  nand g2480 (n_865, n_2233, n_2257, n_2258);
  xor g2481 (n_2259, n_813, n_861);
  xor g2482 (n_54, n_2259, n_862);
  nand g2483 (n_2260, n_813, n_861);
  nand g2484 (n_2261, n_862, n_861);
  nand g2485 (n_2262, n_813, n_862);
  nand g2486 (n_119, n_2260, n_2261, n_2262);
  xor g2488 (n_864, n_2135, A[42]);
  nand g2490 (n_2265, A[42], A[44]);
  nand g2492 (n_868, n_2086, n_2265, n_2032);
  xor g2493 (n_2267, A[45], n_864);
  xor g2494 (n_53, n_2267, n_865);
  nand g2495 (n_2268, A[45], n_864);
  nand g2496 (n_2269, n_865, n_864);
  nand g2497 (n_2270, A[45], n_865);
  nand g2498 (n_118, n_2268, n_2269, n_2270);
  xor g2502 (n_52, n_2271, n_868);
  nand g2505 (n_2274, A[45], n_868);
  nand g2506 (n_117, n_2272, n_2273, n_2274);
  xor g2508 (n_51, n_2135, A[43]);
  nand g2510 (n_2277, A[43], A[44]);
  nand g2512 (n_116, n_2086, n_2277, n_2278);
  nor g11 (n_2294, A[2], A[0]);
  nor g13 (n_2290, A[1], A[3]);
  nor g15 (n_2300, A[2], n_175);
  nand g16 (n_2295, A[2], n_175);
  nor g17 (n_2296, n_108, n_174);
  nand g18 (n_2297, n_108, n_174);
  nor g19 (n_2306, n_107, n_173);
  nand g20 (n_2301, n_107, n_173);
  nor g21 (n_2302, n_106, n_172);
  nand g22 (n_2303, n_106, n_172);
  nor g23 (n_2312, n_105, n_171);
  nand g24 (n_2307, n_105, n_171);
  nor g25 (n_2308, n_104, n_170);
  nand g26 (n_2309, n_104, n_170);
  nor g27 (n_2318, n_103, n_169);
  nand g28 (n_2313, n_103, n_169);
  nor g29 (n_2314, n_102, n_168);
  nand g30 (n_2315, n_102, n_168);
  nor g31 (n_2324, n_101, n_167);
  nand g32 (n_2319, n_101, n_167);
  nor g33 (n_2320, n_100, n_166);
  nand g34 (n_2321, n_100, n_166);
  nor g35 (n_2330, n_99, n_165);
  nand g36 (n_2325, n_99, n_165);
  nor g37 (n_2326, n_98, n_164);
  nand g38 (n_2327, n_98, n_164);
  nor g39 (n_2336, n_97, n_163);
  nand g40 (n_2331, n_97, n_163);
  nor g41 (n_2332, n_96, n_162);
  nand g42 (n_2333, n_96, n_162);
  nor g43 (n_2342, n_95, n_161);
  nand g44 (n_2337, n_95, n_161);
  nor g45 (n_2338, n_94, n_160);
  nand g46 (n_2339, n_94, n_160);
  nor g47 (n_2348, n_93, n_159);
  nand g48 (n_2343, n_93, n_159);
  nor g49 (n_2344, n_92, n_158);
  nand g50 (n_2345, n_92, n_158);
  nor g51 (n_2354, n_91, n_157);
  nand g52 (n_2349, n_91, n_157);
  nor g53 (n_2350, n_90, n_156);
  nand g54 (n_2351, n_90, n_156);
  nor g55 (n_2360, n_89, n_155);
  nand g56 (n_2355, n_89, n_155);
  nor g57 (n_2356, n_88, n_154);
  nand g58 (n_2357, n_88, n_154);
  nor g59 (n_2366, n_87, n_153);
  nand g60 (n_2361, n_87, n_153);
  nor g61 (n_2362, n_86, n_152);
  nand g62 (n_2363, n_86, n_152);
  nor g63 (n_2372, n_85, n_151);
  nand g64 (n_2367, n_85, n_151);
  nor g65 (n_2368, n_84, n_150);
  nand g66 (n_2369, n_84, n_150);
  nor g67 (n_2378, n_83, n_149);
  nand g68 (n_2373, n_83, n_149);
  nor g69 (n_2374, n_82, n_148);
  nand g70 (n_2375, n_82, n_148);
  nor g71 (n_2384, n_81, n_147);
  nand g72 (n_2379, n_81, n_147);
  nor g73 (n_2380, n_80, n_146);
  nand g74 (n_2381, n_80, n_146);
  nor g75 (n_2390, n_79, n_145);
  nand g76 (n_2385, n_79, n_145);
  nor g77 (n_2386, n_78, n_144);
  nand g78 (n_2387, n_78, n_144);
  nor g79 (n_2396, n_77, n_143);
  nand g80 (n_2391, n_77, n_143);
  nor g81 (n_2392, n_76, n_142);
  nand g82 (n_2393, n_76, n_142);
  nor g83 (n_2402, n_75, n_141);
  nand g84 (n_2397, n_75, n_141);
  nor g85 (n_2398, n_74, n_140);
  nand g86 (n_2399, n_74, n_140);
  nor g87 (n_2408, n_73, n_139);
  nand g88 (n_2403, n_73, n_139);
  nor g89 (n_2404, n_72, n_138);
  nand g90 (n_2405, n_72, n_138);
  nor g91 (n_2414, n_71, n_137);
  nand g92 (n_2409, n_71, n_137);
  nor g93 (n_2410, n_70, n_136);
  nand g94 (n_2411, n_70, n_136);
  nor g95 (n_2420, n_69, n_135);
  nand g96 (n_2415, n_69, n_135);
  nor g97 (n_2416, n_68, n_134);
  nand g98 (n_2417, n_68, n_134);
  nor g99 (n_2426, n_67, n_133);
  nand g100 (n_2421, n_67, n_133);
  nor g101 (n_2422, n_66, n_132);
  nand g102 (n_2423, n_66, n_132);
  nor g103 (n_2432, n_65, n_131);
  nand g104 (n_2427, n_65, n_131);
  nor g105 (n_2428, n_64, n_130);
  nand g106 (n_2429, n_64, n_130);
  nor g107 (n_2438, n_63, n_129);
  nand g108 (n_2433, n_63, n_129);
  nor g109 (n_2434, n_62, n_128);
  nand g110 (n_2435, n_62, n_128);
  nor g111 (n_2444, n_61, n_127);
  nand g112 (n_2439, n_61, n_127);
  nor g113 (n_2440, n_60, n_126);
  nand g114 (n_2441, n_60, n_126);
  nor g115 (n_2450, n_59, n_125);
  nand g116 (n_2445, n_59, n_125);
  nor g117 (n_2446, n_58, n_124);
  nand g118 (n_2447, n_58, n_124);
  nor g119 (n_2456, n_57, n_123);
  nand g120 (n_2451, n_57, n_123);
  nor g121 (n_2452, n_56, n_122);
  nand g122 (n_2453, n_56, n_122);
  nor g123 (n_2462, n_55, n_121);
  nand g124 (n_2457, n_55, n_121);
  nor g125 (n_2458, n_54, n_120);
  nand g126 (n_2459, n_54, n_120);
  nor g127 (n_2468, n_53, n_119);
  nand g128 (n_2463, n_53, n_119);
  nor g129 (n_2464, n_52, n_118);
  nand g130 (n_2465, n_52, n_118);
  nor g131 (n_2474, n_51, n_117);
  nand g132 (n_2469, n_51, n_117);
  nor g142 (n_2292, n_876, n_2290);
  nor g146 (n_2298, n_2295, n_2296);
  nor g149 (n_2488, n_2300, n_2296);
  nor g150 (n_2304, n_2301, n_2302);
  nor g153 (n_2490, n_2306, n_2302);
  nor g154 (n_2310, n_2307, n_2308);
  nor g157 (n_2498, n_2312, n_2308);
  nor g158 (n_2316, n_2313, n_2314);
  nor g161 (n_2500, n_2318, n_2314);
  nor g162 (n_2322, n_2319, n_2320);
  nor g165 (n_2508, n_2324, n_2320);
  nor g166 (n_2328, n_2325, n_2326);
  nor g169 (n_2510, n_2330, n_2326);
  nor g170 (n_2334, n_2331, n_2332);
  nor g173 (n_2518, n_2336, n_2332);
  nor g174 (n_2340, n_2337, n_2338);
  nor g177 (n_2520, n_2342, n_2338);
  nor g178 (n_2346, n_2343, n_2344);
  nor g181 (n_2528, n_2348, n_2344);
  nor g182 (n_2352, n_2349, n_2350);
  nor g185 (n_2530, n_2354, n_2350);
  nor g186 (n_2358, n_2355, n_2356);
  nor g189 (n_2538, n_2360, n_2356);
  nor g190 (n_2364, n_2361, n_2362);
  nor g193 (n_2540, n_2366, n_2362);
  nor g194 (n_2370, n_2367, n_2368);
  nor g197 (n_2548, n_2372, n_2368);
  nor g198 (n_2376, n_2373, n_2374);
  nor g201 (n_2550, n_2378, n_2374);
  nor g202 (n_2382, n_2379, n_2380);
  nor g205 (n_2558, n_2384, n_2380);
  nor g206 (n_2388, n_2385, n_2386);
  nor g209 (n_2560, n_2390, n_2386);
  nor g210 (n_2394, n_2391, n_2392);
  nor g213 (n_2568, n_2396, n_2392);
  nor g214 (n_2400, n_2397, n_2398);
  nor g217 (n_2570, n_2402, n_2398);
  nor g218 (n_2406, n_2403, n_2404);
  nor g221 (n_2578, n_2408, n_2404);
  nor g222 (n_2412, n_2409, n_2410);
  nor g225 (n_2580, n_2414, n_2410);
  nor g226 (n_2418, n_2415, n_2416);
  nor g229 (n_2588, n_2420, n_2416);
  nor g230 (n_2424, n_2421, n_2422);
  nor g233 (n_2590, n_2426, n_2422);
  nor g234 (n_2430, n_2427, n_2428);
  nor g237 (n_2598, n_2432, n_2428);
  nor g238 (n_2436, n_2433, n_2434);
  nor g241 (n_2600, n_2438, n_2434);
  nor g242 (n_2442, n_2439, n_2440);
  nor g245 (n_2608, n_2444, n_2440);
  nor g246 (n_2448, n_2445, n_2446);
  nor g249 (n_2610, n_2450, n_2446);
  nor g250 (n_2454, n_2451, n_2452);
  nor g253 (n_2618, n_2456, n_2452);
  nor g254 (n_2460, n_2457, n_2458);
  nor g257 (n_2620, n_2462, n_2458);
  nor g258 (n_2466, n_2463, n_2464);
  nor g261 (n_2628, n_2468, n_2464);
  nor g262 (n_2472, n_2469, n_2470);
  nor g265 (n_2630, n_2474, n_2470);
  nor g275 (n_2486, n_2306, n_2485);
  nand g284 (n_2643, n_2488, n_2490);
  nor g285 (n_2496, n_2318, n_2495);
  nand g294 (n_2650, n_2498, n_2500);
  nor g295 (n_2506, n_2330, n_2505);
  nand g304 (n_2658, n_2508, n_2510);
  nor g305 (n_2516, n_2342, n_2515);
  nand g314 (n_2665, n_2518, n_2520);
  nor g315 (n_2526, n_2354, n_2525);
  nand g324 (n_2673, n_2528, n_2530);
  nor g325 (n_2536, n_2366, n_2535);
  nand g334 (n_2680, n_2538, n_2540);
  nor g335 (n_2546, n_2378, n_2545);
  nand g344 (n_2688, n_2548, n_2550);
  nor g345 (n_2556, n_2390, n_2555);
  nand g354 (n_2695, n_2558, n_2560);
  nor g355 (n_2566, n_2402, n_2565);
  nand g364 (n_2703, n_2568, n_2570);
  nor g365 (n_2576, n_2414, n_2575);
  nand g2522 (n_2710, n_2578, n_2580);
  nor g2523 (n_2586, n_2426, n_2585);
  nand g2532 (n_2718, n_2588, n_2590);
  nor g2533 (n_2596, n_2438, n_2595);
  nand g2542 (n_2725, n_2598, n_2600);
  nor g2543 (n_2606, n_2450, n_2605);
  nand g2552 (n_2733, n_2608, n_2610);
  nor g2553 (n_2616, n_2462, n_2615);
  nand g2562 (n_2740, n_2618, n_2620);
  nor g2563 (n_2626, n_2474, n_2625);
  nand g2572 (n_2748, n_2628, n_2630);
  nand g2575 (n_3105, n_2295, n_2637);
  nand g2577 (n_3107, n_2485, n_2638);
  nand g2580 (n_3110, n_2641, n_2642);
  nand g2583 (n_2752, n_2645, n_2646);
  nor g2584 (n_2648, n_2324, n_2647);
  nor g2587 (n_2762, n_2324, n_2650);
  nor g2593 (n_2656, n_2654, n_2647);
  nor g2596 (n_2768, n_2650, n_2654);
  nor g2597 (n_2660, n_2658, n_2647);
  nor g2600 (n_2771, n_2650, n_2658);
  nor g2601 (n_2663, n_2348, n_2662);
  nor g2604 (n_2892, n_2348, n_2665);
  nor g2610 (n_2671, n_2669, n_2662);
  nor g2613 (n_2898, n_2665, n_2669);
  nor g2614 (n_2675, n_2673, n_2662);
  nor g2617 (n_2777, n_2665, n_2673);
  nor g2618 (n_2678, n_2372, n_2677);
  nor g2621 (n_2790, n_2372, n_2680);
  nor g2627 (n_2686, n_2684, n_2677);
  nor g2630 (n_2800, n_2680, n_2684);
  nor g2631 (n_2690, n_2688, n_2677);
  nor g2634 (n_2805, n_2680, n_2688);
  nor g2635 (n_2693, n_2396, n_2692);
  nor g2638 (n_3007, n_2396, n_2695);
  nor g2644 (n_2701, n_2699, n_2692);
  nor g2647 (n_3013, n_2695, n_2699);
  nor g2648 (n_2705, n_2703, n_2692);
  nor g2651 (n_2813, n_2695, n_2703);
  nor g2652 (n_2708, n_2420, n_2707);
  nor g2655 (n_2826, n_2420, n_2710);
  nor g2661 (n_2716, n_2714, n_2707);
  nor g2664 (n_2836, n_2710, n_2714);
  nor g2665 (n_2720, n_2718, n_2707);
  nor g2668 (n_2841, n_2710, n_2718);
  nor g2669 (n_2723, n_2444, n_2722);
  nor g2672 (n_2947, n_2444, n_2725);
  nor g2678 (n_2731, n_2729, n_2722);
  nor g2681 (n_2957, n_2725, n_2729);
  nor g2682 (n_2735, n_2733, n_2722);
  nor g2685 (n_2849, n_2725, n_2733);
  nor g2686 (n_2738, n_2468, n_2737);
  nor g2689 (n_2862, n_2468, n_2740);
  nor g2695 (n_2746, n_2744, n_2737);
  nor g2698 (n_2872, n_2740, n_2744);
  nor g2699 (n_2750, n_2748, n_2737);
  nor g2702 (n_2877, n_2740, n_2748);
  nand g2705 (n_3114, n_2307, n_2754);
  nand g2706 (n_2755, n_2498, n_2752);
  nand g2707 (n_3116, n_2495, n_2755);
  nand g2710 (n_3119, n_2758, n_2759);
  nand g2713 (n_3122, n_2647, n_2761);
  nand g2714 (n_2764, n_2762, n_2752);
  nand g2715 (n_3125, n_2763, n_2764);
  nand g2716 (n_2767, n_2765, n_2752);
  nand g2717 (n_3127, n_2766, n_2767);
  nand g2718 (n_2770, n_2768, n_2752);
  nand g2719 (n_3130, n_2769, n_2770);
  nand g2720 (n_2773, n_2771, n_2752);
  nand g2721 (n_2882, n_2772, n_2773);
  nor g2722 (n_2775, n_2360, n_2774);
  nand g2731 (n_2906, n_2538, n_2777);
  nor g2732 (n_2784, n_2782, n_2774);
  nor g2737 (n_2787, n_2680, n_2774);
  nand g2746 (n_2918, n_2777, n_2790);
  nand g2751 (n_2922, n_2777, n_2795);
  nand g2756 (n_2926, n_2777, n_2800);
  nand g2761 (n_2930, n_2777, n_2805);
  nor g2762 (n_2811, n_2408, n_2810);
  nand g2771 (n_3021, n_2578, n_2813);
  nor g2772 (n_2820, n_2818, n_2810);
  nor g2777 (n_2823, n_2710, n_2810);
  nand g2786 (n_3033, n_2813, n_2826);
  nand g2791 (n_3037, n_2813, n_2831);
  nand g2796 (n_3041, n_2813, n_2836);
  nand g2801 (n_2937, n_2813, n_2841);
  nor g2802 (n_2847, n_2456, n_2846);
  nand g2811 (n_2969, n_2618, n_2849);
  nor g2812 (n_2856, n_2854, n_2846);
  nor g2817 (n_2859, n_2740, n_2846);
  nand g2826 (n_2981, n_2849, n_2862);
  nand g2831 (n_2985, n_2849, n_2867);
  nand g2836 (n_2989, n_2849, n_2872);
  nand g2841 (n_2993, n_2849, n_2877);
  nand g2844 (n_3134, n_2331, n_2884);
  nand g2845 (n_2885, n_2518, n_2882);
  nand g2846 (n_3136, n_2515, n_2885);
  nand g2849 (n_3139, n_2888, n_2889);
  nand g2852 (n_3142, n_2662, n_2891);
  nand g2853 (n_2894, n_2892, n_2882);
  nand g2854 (n_3145, n_2893, n_2894);
  nand g2855 (n_2897, n_2895, n_2882);
  nand g2856 (n_3147, n_2896, n_2897);
  nand g2857 (n_2900, n_2898, n_2882);
  nand g2858 (n_3150, n_2899, n_2900);
  nand g2859 (n_2901, n_2777, n_2882);
  nand g2860 (n_3152, n_2774, n_2901);
  nand g2863 (n_3155, n_2904, n_2905);
  nand g2866 (n_3157, n_2908, n_2909);
  nand g2869 (n_3160, n_2912, n_2913);
  nand g2872 (n_3163, n_2916, n_2917);
  nand g2875 (n_3166, n_2920, n_2921);
  nand g2878 (n_3168, n_2924, n_2925);
  nand g2881 (n_3171, n_2928, n_2929);
  nand g2884 (n_2997, n_2932, n_2933);
  nor g2885 (n_2935, n_2432, n_2934);
  nor g2888 (n_3047, n_2432, n_2937);
  nor g2894 (n_2943, n_2941, n_2934);
  nor g2897 (n_3053, n_2941, n_2937);
  nor g2898 (n_2945, n_2725, n_2934);
  nor g2901 (n_3056, n_2725, n_2937);
  nor g2922 (n_2967, n_2965, n_2934);
  nor g2925 (n_3071, n_2937, n_2965);
  nor g2926 (n_2971, n_2969, n_2934);
  nor g2929 (n_3074, n_2937, n_2969);
  nor g2930 (n_2975, n_2973, n_2934);
  nor g2933 (n_3077, n_2937, n_2973);
  nor g2934 (n_2979, n_2977, n_2934);
  nor g2937 (n_3080, n_2937, n_2977);
  nor g2938 (n_2983, n_2981, n_2934);
  nor g2941 (n_3083, n_2937, n_2981);
  nor g2942 (n_2987, n_2985, n_2934);
  nor g2945 (n_3086, n_2937, n_2985);
  nor g2946 (n_2991, n_2989, n_2934);
  nor g2949 (n_3089, n_2937, n_2989);
  nor g2950 (n_2995, n_2993, n_2934);
  nor g2953 (n_3092, n_2937, n_2993);
  nand g2956 (n_3175, n_2379, n_2999);
  nand g2957 (n_3000, n_2558, n_2997);
  nand g2958 (n_3177, n_2555, n_3000);
  nand g2961 (n_3180, n_3003, n_3004);
  nand g2964 (n_3183, n_2692, n_3006);
  nand g2965 (n_3009, n_3007, n_2997);
  nand g2966 (n_3186, n_3008, n_3009);
  nand g2967 (n_3012, n_3010, n_2997);
  nand g2968 (n_3188, n_3011, n_3012);
  nand g2969 (n_3015, n_3013, n_2997);
  nand g2970 (n_3191, n_3014, n_3015);
  nand g2971 (n_3016, n_2813, n_2997);
  nand g2972 (n_3193, n_2810, n_3016);
  nand g2975 (n_3196, n_3019, n_3020);
  nand g2978 (n_3198, n_3023, n_3024);
  nand g2981 (n_3201, n_3027, n_3028);
  nand g2984 (n_3204, n_3031, n_3032);
  nand g2987 (n_3207, n_3035, n_3036);
  nand g2990 (n_3209, n_3039, n_3040);
  nand g2993 (n_3212, n_3043, n_3044);
  nand g2996 (n_3215, n_2934, n_3046);
  nand g2997 (n_3049, n_3047, n_2997);
  nand g2998 (n_3218, n_3048, n_3049);
  nand g2999 (n_3052, n_3050, n_2997);
  nand g3000 (n_3220, n_3051, n_3052);
  nand g3001 (n_3055, n_3053, n_2997);
  nand g3002 (n_3223, n_3054, n_3055);
  nand g3003 (n_3058, n_3056, n_2997);
  nand g3004 (n_3226, n_3057, n_3058);
  nand g3005 (n_3061, n_3059, n_2997);
  nand g3006 (n_3229, n_3060, n_3061);
  nand g3007 (n_3064, n_3062, n_2997);
  nand g3008 (n_3231, n_3063, n_3064);
  nand g3009 (n_3067, n_3065, n_2997);
  nand g3010 (n_3234, n_3066, n_3067);
  nand g3011 (n_3070, n_3068, n_2997);
  nand g3012 (n_3236, n_3069, n_3070);
  nand g3013 (n_3073, n_3071, n_2997);
  nand g3014 (n_3239, n_3072, n_3073);
  nand g3015 (n_3076, n_3074, n_2997);
  nand g3016 (n_3241, n_3075, n_3076);
  nand g3017 (n_3079, n_3077, n_2997);
  nand g3018 (n_3244, n_3078, n_3079);
  nand g3019 (n_3082, n_3080, n_2997);
  nand g3020 (n_3247, n_3081, n_3082);
  nand g3021 (n_3085, n_3083, n_2997);
  nand g3022 (n_3250, n_3084, n_3085);
  nand g3023 (n_3088, n_3086, n_2997);
  nand g3024 (n_3252, n_3087, n_3088);
  nand g3025 (n_3091, n_3089, n_2997);
  nand g3026 (n_3255, n_3090, n_3091);
  nand g3027 (n_3094, n_3092, n_2997);
  nand g3028 (n_3095, n_3093, n_3094);
  nand g3031 (n_3259, n_2475, n_3097);
  xnor g3043 (Z[5], n_3105, n_3106);
  xnor g3045 (Z[6], n_3107, n_3108);
  xnor g3048 (Z[7], n_3110, n_3111);
  xnor g3050 (Z[8], n_2752, n_3112);
  xnor g3053 (Z[9], n_3114, n_3115);
  xnor g3055 (Z[10], n_3116, n_3117);
  xnor g3058 (Z[11], n_3119, n_3120);
  xnor g3061 (Z[12], n_3122, n_3123);
  xnor g3064 (Z[13], n_3125, n_3126);
  xnor g3066 (Z[14], n_3127, n_3128);
  xnor g3069 (Z[15], n_3130, n_3131);
  xnor g3071 (Z[16], n_2882, n_3132);
  xnor g3074 (Z[17], n_3134, n_3135);
  xnor g3076 (Z[18], n_3136, n_3137);
  xnor g3079 (Z[19], n_3139, n_3140);
  xnor g3082 (Z[20], n_3142, n_3143);
  xnor g3085 (Z[21], n_3145, n_3146);
  xnor g3087 (Z[22], n_3147, n_3148);
  xnor g3090 (Z[23], n_3150, n_3151);
  xnor g3092 (Z[24], n_3152, n_3153);
  xnor g3095 (Z[25], n_3155, n_3156);
  xnor g3097 (Z[26], n_3157, n_3158);
  xnor g3100 (Z[27], n_3160, n_3161);
  xnor g3103 (Z[28], n_3163, n_3164);
  xnor g3106 (Z[29], n_3166, n_3167);
  xnor g3108 (Z[30], n_3168, n_3169);
  xnor g3111 (Z[31], n_3171, n_3172);
  xnor g3113 (Z[32], n_2997, n_3173);
  xnor g3116 (Z[33], n_3175, n_3176);
  xnor g3118 (Z[34], n_3177, n_3178);
  xnor g3121 (Z[35], n_3180, n_3181);
  xnor g3124 (Z[36], n_3183, n_3184);
  xnor g3127 (Z[37], n_3186, n_3187);
  xnor g3129 (Z[38], n_3188, n_3189);
  xnor g3132 (Z[39], n_3191, n_3192);
  xnor g3134 (Z[40], n_3193, n_3194);
  xnor g3137 (Z[41], n_3196, n_3197);
  xnor g3139 (Z[42], n_3198, n_3199);
  xnor g3142 (Z[43], n_3201, n_3202);
  xnor g3145 (Z[44], n_3204, n_3205);
  xnor g3148 (Z[45], n_3207, n_3208);
  xnor g3150 (Z[46], n_3209, n_3210);
  xnor g3153 (Z[47], n_3212, n_3213);
  xnor g3156 (Z[48], n_3215, n_3216);
  xnor g3159 (Z[49], n_3218, n_3219);
  xnor g3161 (Z[50], n_3220, n_3221);
  xnor g3164 (Z[51], n_3223, n_3224);
  xnor g3167 (Z[52], n_3226, n_3227);
  xnor g3170 (Z[53], n_3229, n_3230);
  xnor g3172 (Z[54], n_3231, n_3232);
  xnor g3175 (Z[55], n_3234, n_3235);
  xnor g3177 (Z[56], n_3236, n_3237);
  xnor g3180 (Z[57], n_3239, n_3240);
  xnor g3182 (Z[58], n_3241, n_3242);
  xnor g3185 (Z[59], n_3244, n_3245);
  xnor g3188 (Z[60], n_3247, n_3248);
  xnor g3191 (Z[61], n_3250, n_3251);
  xnor g3193 (Z[62], n_3252, n_3253);
  xnor g3196 (Z[63], n_3255, n_3256);
  xnor g3198 (Z[64], n_3095, n_3257);
  or g3215 (n_254, wc, wc0, n_108);
  not gc0 (wc0, n_876);
  not gc (wc, n_890);
  or g3216 (n_263, wc1, wc2, n_248);
  not gc2 (wc2, n_890);
  not gc1 (wc1, n_909);
  or g3217 (n_276, wc3, n_253, n_248);
  not gc3 (wc3, n_937);
  or g3218 (n_293, wc4, wc5, n_253);
  not gc5 (wc5, n_972);
  not gc4 (wc4, n_973);
  or g3219 (n_315, wc6, wc7, n_253);
  not gc7 (wc7, n_1020);
  not gc6 (wc6, n_1021);
  or g3220 (n_363, wc8, wc9, n_248);
  not gc9 (wc9, n_1021);
  not gc8 (wc8, n_1068);
  or g3221 (n_391, wc10, wc11, n_253);
  not gc11 (wc11, n_1197);
  not gc10 (wc10, n_1198);
  or g3222 (n_417, wc12, wc13, n_262);
  not gc13 (wc13, n_1137);
  not gc12 (wc12, n_1261);
  or g3223 (n_445, wc14, wc15, n_275);
  not gc15 (wc15, n_1201);
  not gc14 (wc14, n_1325);
  or g3224 (n_473, wc16, wc17, n_292);
  not gc17 (wc17, n_1130);
  not gc16 (wc16, n_1389);
  or g3225 (n_501, wc18, wc19, n_313);
  not gc19 (wc19, n_1194);
  not gc18 (wc18, n_1453);
  or g3226 (n_529, wc20, wc21, n_113);
  not gc21 (wc21, n_1258);
  not gc20 (wc20, n_1517);
  or g3227 (n_558, wc22, wc23, n_113);
  not gc23 (wc23, n_1580);
  not gc22 (wc22, n_1581);
  xnor g3228 (n_2023, A[46], A[32]);
  or g3229 (n_2024, wc24, A[46]);
  not gc24 (wc24, A[32]);
  or g3230 (n_2026, wc25, A[46]);
  not gc25 (wc25, A[30]);
  xnor g3231 (n_2063, A[41], A[33]);
  or g3232 (n_2064, A[33], wc26);
  not gc26 (wc26, A[41]);
  or g3233 (n_2086, wc27, A[46]);
  not gc27 (wc27, A[44]);
  xnor g3234 (n_2135, A[46], A[44]);
  or g3235 (n_2138, wc28, A[46]);
  not gc28 (wc28, A[40]);
  xnor g3236 (n_815, n_1807, A[43]);
  or g3237 (n_2165, wc29, A[43]);
  not gc29 (wc29, A[41]);
  or g3238 (n_2166, wc30, A[43]);
  not gc30 (wc30, A[35]);
  xnor g3240 (n_861, n_2255, A[45]);
  or g3241 (n_2257, wc31, A[45]);
  not gc31 (wc31, A[41]);
  or g3242 (n_2258, wc32, A[45]);
  not gc32 (wc32, A[43]);
  or g3243 (n_2032, wc33, A[46]);
  not gc33 (wc33, A[42]);
  xnor g3244 (n_2271, A[45], A[43]);
  or g3245 (n_2272, A[43], wc34);
  not gc34 (wc34, A[45]);
  or g3246 (n_2278, wc35, A[46]);
  not gc35 (wc35, A[43]);
  and g3247 (n_2478, wc36, A[46]);
  not gc36 (wc36, A[45]);
  or g3248 (n_2475, wc37, A[46]);
  not gc37 (wc37, A[45]);
  or g3249 (n_340, wc38, wc39, n_253);
  not gc39 (wc39, n_1077);
  not gc38 (wc38, n_1078);
  or g3250 (n_2122, A[33], wc40);
  not gc40 (wc40, n_789);
  xnor g3251 (n_835, n_730, n_2255);
  or g3252 (n_2205, A[43], wc41);
  not gc41 (wc41, n_730);
  or g3253 (n_2238, A[45], wc42);
  not gc42 (wc42, n_849);
  and g3254 (n_2483, wc43, n_872);
  not gc43 (wc43, n_2292);
  or g3256 (n_3099, n_2294, wc44);
  not gc44 (wc44, n_876);
  or g3257 (n_3102, n_2290, wc45);
  not gc45 (wc45, n_872);
  xnor g3258 (n_2031, A[46], A[42]);
  or g3259 (n_2034, wc46, A[46]);
  not gc46 (wc46, A[36]);
  or g3260 (n_2065, A[33], wc47);
  not gc47 (wc47, n_760);
  xnor g3261 (n_2119, n_788, A[33]);
  or g3262 (n_2120, A[33], wc48);
  not gc48 (wc48, n_788);
  xnor g3263 (n_2235, n_813, A[45]);
  or g3264 (n_2236, A[45], wc49);
  not gc49 (wc49, n_813);
  or g3265 (n_2273, A[43], wc50);
  not gc50 (wc50, n_868);
  and g3266 (n_2470, A[45], wc51);
  not gc51 (wc51, n_116);
  or g3267 (n_2471, A[45], wc52);
  not gc52 (wc52, n_116);
  or g3268 (n_3103, wc53, n_2300);
  not gc53 (wc53, n_2295);
  or g3269 (n_3257, wc54, n_2478);
  not gc54 (wc54, n_2475);
  and g3270 (n_2485, wc55, n_2297);
  not gc55 (wc55, n_2298);
  or g3271 (n_2639, wc56, n_2306);
  not gc56 (wc56, n_2488);
  not g3272 (Z[2], n_3099);
  or g3273 (n_3106, wc57, n_2296);
  not gc57 (wc57, n_2297);
  or g3274 (n_3108, wc58, n_2306);
  not gc58 (wc58, n_2301);
  and g3275 (n_2492, wc59, n_2303);
  not gc59 (wc59, n_2304);
  or g3278 (n_3111, wc60, n_2302);
  not gc60 (wc60, n_2303);
  or g3279 (n_3256, wc61, n_2470);
  not gc61 (wc61, n_2471);
  and g3280 (n_2495, wc62, n_2309);
  not gc62 (wc62, n_2310);
  and g3281 (n_2641, wc63, n_2301);
  not gc63 (wc63, n_2486);
  and g3282 (n_2493, wc64, n_2490);
  not gc64 (wc64, n_2485);
  or g3283 (n_2637, n_2300, n_2483);
  or g3284 (n_2638, n_2483, wc65);
  not gc65 (wc65, n_2488);
  or g3285 (n_2642, n_2483, n_2639);
  xor g3286 (Z[3], n_876, n_3102);
  xor g3287 (Z[4], n_2483, n_3103);
  or g3288 (n_3112, wc66, n_2312);
  not gc66 (wc66, n_2307);
  or g3289 (n_3115, wc67, n_2308);
  not gc67 (wc67, n_2309);
  and g3290 (n_2632, n_2471, wc68);
  not gc68 (wc68, n_2472);
  and g3291 (n_2645, wc69, n_2492);
  not gc69 (wc69, n_2493);
  or g3292 (n_2756, wc70, n_2318);
  not gc70 (wc70, n_2498);
  or g3293 (n_2646, n_2643, n_2483);
  or g3294 (n_3117, wc71, n_2318);
  not gc71 (wc71, n_2313);
  or g3295 (n_3251, wc72, n_2464);
  not gc72 (wc72, n_2465);
  or g3296 (n_3253, wc73, n_2474);
  not gc73 (wc73, n_2469);
  and g3297 (n_2502, wc74, n_2315);
  not gc74 (wc74, n_2316);
  and g3298 (n_2505, wc75, n_2321);
  not gc75 (wc75, n_2322);
  and g3299 (n_2625, wc76, n_2465);
  not gc76 (wc76, n_2466);
  and g3300 (n_2758, wc77, n_2313);
  not gc77 (wc77, n_2496);
  or g3301 (n_2744, wc78, n_2474);
  not gc78 (wc78, n_2628);
  or g3302 (n_3120, wc79, n_2314);
  not gc79 (wc79, n_2315);
  or g3303 (n_3123, wc80, n_2324);
  not gc80 (wc80, n_2319);
  or g3304 (n_3126, wc81, n_2320);
  not gc81 (wc81, n_2321);
  or g3305 (n_3248, wc82, n_2468);
  not gc82 (wc82, n_2463);
  and g3306 (n_2512, wc83, n_2327);
  not gc83 (wc83, n_2328);
  and g3307 (n_2622, wc84, n_2459);
  not gc84 (wc84, n_2460);
  and g3308 (n_2503, wc85, n_2500);
  not gc85 (wc85, n_2495);
  or g3309 (n_2654, wc86, n_2330);
  not gc86 (wc86, n_2508);
  and g3310 (n_2633, wc87, n_2630);
  not gc87 (wc87, n_2625);
  and g3311 (n_2765, wc88, n_2508);
  not gc88 (wc88, n_2650);
  or g3312 (n_2754, wc89, n_2312);
  not gc89 (wc89, n_2752);
  or g3313 (n_2759, n_2756, wc90);
  not gc90 (wc90, n_2752);
  or g3314 (n_3128, wc91, n_2330);
  not gc91 (wc91, n_2325);
  or g3315 (n_3131, wc92, n_2326);
  not gc92 (wc92, n_2327);
  or g3316 (n_3240, wc93, n_2452);
  not gc93 (wc93, n_2453);
  or g3317 (n_3242, wc94, n_2462);
  not gc94 (wc94, n_2457);
  or g3318 (n_3245, wc95, n_2458);
  not gc95 (wc95, n_2459);
  and g3319 (n_2515, wc96, n_2333);
  not gc96 (wc96, n_2334);
  and g3320 (n_2522, wc97, n_2339);
  not gc97 (wc97, n_2340);
  and g3321 (n_2615, wc98, n_2453);
  not gc98 (wc98, n_2454);
  and g3322 (n_2647, wc99, n_2502);
  not gc99 (wc99, n_2503);
  and g3323 (n_2655, wc100, n_2325);
  not gc100 (wc100, n_2506);
  and g3324 (n_2513, wc101, n_2510);
  not gc101 (wc101, n_2505);
  or g3325 (n_2886, wc102, n_2342);
  not gc102 (wc102, n_2518);
  or g3326 (n_2854, wc103, n_2462);
  not gc103 (wc103, n_2618);
  and g3327 (n_2745, wc104, n_2469);
  not gc104 (wc104, n_2626);
  and g3328 (n_2749, wc105, n_2632);
  not gc105 (wc105, n_2633);
  or g3329 (n_2761, wc106, n_2650);
  not gc106 (wc106, n_2752);
  or g3330 (n_3132, wc107, n_2336);
  not gc107 (wc107, n_2331);
  or g3331 (n_3135, wc108, n_2332);
  not gc108 (wc108, n_2333);
  or g3332 (n_3137, wc109, n_2342);
  not gc109 (wc109, n_2337);
  or g3333 (n_3140, wc110, n_2338);
  not gc110 (wc110, n_2339);
  or g3334 (n_3143, wc111, n_2348);
  not gc111 (wc111, n_2343);
  or g3335 (n_3237, wc112, n_2456);
  not gc112 (wc112, n_2451);
  and g3336 (n_2525, wc113, n_2345);
  not gc113 (wc113, n_2346);
  and g3337 (n_2612, wc114, n_2447);
  not gc114 (wc114, n_2448);
  and g3338 (n_2659, wc115, n_2512);
  not gc115 (wc115, n_2513);
  and g3339 (n_2523, wc116, n_2520);
  not gc116 (wc116, n_2515);
  or g3340 (n_2669, wc117, n_2354);
  not gc117 (wc117, n_2528);
  and g3341 (n_2623, wc118, n_2620);
  not gc118 (wc118, n_2615);
  and g3342 (n_2652, wc119, n_2508);
  not gc119 (wc119, n_2647);
  and g3343 (n_2867, wc120, n_2628);
  not gc120 (wc120, n_2740);
  or g3344 (n_3146, wc121, n_2344);
  not gc121 (wc121, n_2345);
  or g3345 (n_3148, wc122, n_2354);
  not gc122 (wc122, n_2349);
  or g3346 (n_3232, wc123, n_2450);
  not gc123 (wc123, n_2445);
  or g3347 (n_3235, wc124, n_2446);
  not gc124 (wc124, n_2447);
  and g3348 (n_2532, wc125, n_2351);
  not gc125 (wc125, n_2352);
  and g3349 (n_2535, wc126, n_2357);
  not gc126 (wc126, n_2358);
  and g3350 (n_2542, wc127, n_2363);
  not gc127 (wc127, n_2364);
  and g3351 (n_2545, wc128, n_2369);
  not gc128 (wc128, n_2370);
  and g3352 (n_2552, wc129, n_2375);
  not gc129 (wc129, n_2376);
  and g3353 (n_2555, wc130, n_2381);
  not gc130 (wc130, n_2382);
  and g3354 (n_2562, wc131, n_2387);
  not gc131 (wc131, n_2388);
  and g3355 (n_2565, wc132, n_2393);
  not gc132 (wc132, n_2394);
  and g3356 (n_2572, wc133, n_2399);
  not gc133 (wc133, n_2400);
  and g3357 (n_2575, wc134, n_2405);
  not gc134 (wc134, n_2406);
  and g3358 (n_2582, wc135, n_2411);
  not gc135 (wc135, n_2412);
  and g3359 (n_2585, wc136, n_2417);
  not gc136 (wc136, n_2418);
  and g3360 (n_2592, wc137, n_2423);
  not gc137 (wc137, n_2424);
  and g3361 (n_2888, wc138, n_2337);
  not gc138 (wc138, n_2516);
  and g3362 (n_2662, wc139, n_2522);
  not gc139 (wc139, n_2523);
  or g3363 (n_2782, wc140, n_2366);
  not gc140 (wc140, n_2538);
  or g3364 (n_2684, wc141, n_2378);
  not gc141 (wc141, n_2548);
  or g3365 (n_3001, wc142, n_2390);
  not gc142 (wc142, n_2558);
  or g3366 (n_2699, wc143, n_2402);
  not gc143 (wc143, n_2568);
  or g3367 (n_2818, wc144, n_2414);
  not gc144 (wc144, n_2578);
  or g3368 (n_2714, wc145, n_2426);
  not gc145 (wc145, n_2588);
  and g3369 (n_2855, wc146, n_2457);
  not gc146 (wc146, n_2616);
  and g3370 (n_2737, wc147, n_2622);
  not gc147 (wc147, n_2623);
  and g3371 (n_2763, wc148, n_2319);
  not gc148 (wc148, n_2648);
  and g3372 (n_2766, wc149, n_2505);
  not gc149 (wc149, n_2652);
  and g3373 (n_2769, n_2655, wc150);
  not gc150 (wc150, n_2656);
  and g3374 (n_2895, wc151, n_2528);
  not gc151 (wc151, n_2665);
  or g3375 (n_3151, wc152, n_2350);
  not gc152 (wc152, n_2351);
  or g3376 (n_3153, wc153, n_2360);
  not gc153 (wc153, n_2355);
  or g3377 (n_3156, wc154, n_2356);
  not gc154 (wc154, n_2357);
  or g3378 (n_3158, wc155, n_2366);
  not gc155 (wc155, n_2361);
  or g3379 (n_3161, wc156, n_2362);
  not gc156 (wc156, n_2363);
  or g3380 (n_3164, wc157, n_2372);
  not gc157 (wc157, n_2367);
  or g3381 (n_3167, wc158, n_2368);
  not gc158 (wc158, n_2369);
  or g3382 (n_3169, wc159, n_2378);
  not gc159 (wc159, n_2373);
  or g3383 (n_3172, wc160, n_2374);
  not gc160 (wc160, n_2375);
  or g3384 (n_3173, wc161, n_2384);
  not gc161 (wc161, n_2379);
  or g3385 (n_3176, wc162, n_2380);
  not gc162 (wc162, n_2381);
  or g3386 (n_3178, wc163, n_2390);
  not gc163 (wc163, n_2385);
  or g3387 (n_3181, wc164, n_2386);
  not gc164 (wc164, n_2387);
  or g3388 (n_3184, wc165, n_2396);
  not gc165 (wc165, n_2391);
  or g3389 (n_3187, wc166, n_2392);
  not gc166 (wc166, n_2393);
  or g3390 (n_3189, wc167, n_2402);
  not gc167 (wc167, n_2397);
  or g3391 (n_3192, wc168, n_2398);
  not gc168 (wc168, n_2399);
  or g3392 (n_3194, wc169, n_2408);
  not gc169 (wc169, n_2403);
  or g3393 (n_3197, wc170, n_2404);
  not gc170 (wc170, n_2405);
  or g3394 (n_3199, wc171, n_2414);
  not gc171 (wc171, n_2409);
  or g3395 (n_3202, wc172, n_2410);
  not gc172 (wc172, n_2411);
  or g3396 (n_3205, wc173, n_2420);
  not gc173 (wc173, n_2415);
  or g3397 (n_3208, wc174, n_2416);
  not gc174 (wc174, n_2417);
  or g3398 (n_3210, wc175, n_2426);
  not gc175 (wc175, n_2421);
  or g3399 (n_3213, wc176, n_2422);
  not gc176 (wc176, n_2423);
  and g3400 (n_2595, wc177, n_2429);
  not gc177 (wc177, n_2430);
  and g3401 (n_2605, wc178, n_2441);
  not gc178 (wc178, n_2442);
  and g3402 (n_2670, wc179, n_2349);
  not gc179 (wc179, n_2526);
  and g3403 (n_2533, wc180, n_2530);
  not gc180 (wc180, n_2525);
  and g3404 (n_2543, wc181, n_2540);
  not gc181 (wc181, n_2535);
  and g3405 (n_2553, wc182, n_2550);
  not gc182 (wc182, n_2545);
  and g3406 (n_2563, wc183, n_2560);
  not gc183 (wc183, n_2555);
  and g3407 (n_2573, wc184, n_2570);
  not gc184 (wc184, n_2565);
  and g3408 (n_2583, wc185, n_2580);
  not gc185 (wc185, n_2575);
  and g3409 (n_2593, wc186, n_2590);
  not gc186 (wc186, n_2585);
  or g3410 (n_2729, wc187, n_2450);
  not gc187 (wc187, n_2608);
  and g3411 (n_2772, n_2659, wc188);
  not gc188 (wc188, n_2660);
  and g3412 (n_2667, wc189, n_2528);
  not gc189 (wc189, n_2662);
  and g3413 (n_2795, wc190, n_2548);
  not gc190 (wc190, n_2680);
  and g3414 (n_3010, wc191, n_2568);
  not gc191 (wc191, n_2695);
  and g3415 (n_2831, wc192, n_2588);
  not gc192 (wc192, n_2710);
  and g3416 (n_2742, wc193, n_2628);
  not gc193 (wc193, n_2737);
  or g3417 (n_3216, wc194, n_2432);
  not gc194 (wc194, n_2427);
  or g3418 (n_3219, wc195, n_2428);
  not gc195 (wc195, n_2429);
  or g3419 (n_3224, wc196, n_2434);
  not gc196 (wc196, n_2435);
  or g3420 (n_3227, wc197, n_2444);
  not gc197 (wc197, n_2439);
  or g3421 (n_3230, wc198, n_2440);
  not gc198 (wc198, n_2441);
  and g3422 (n_2602, wc199, n_2435);
  not gc199 (wc199, n_2436);
  and g3423 (n_2674, wc200, n_2532);
  not gc200 (wc200, n_2533);
  and g3424 (n_2783, wc201, n_2361);
  not gc201 (wc201, n_2536);
  and g3425 (n_2677, wc202, n_2542);
  not gc202 (wc202, n_2543);
  and g3426 (n_2685, wc203, n_2373);
  not gc203 (wc203, n_2546);
  and g3427 (n_2689, wc204, n_2552);
  not gc204 (wc204, n_2553);
  and g3428 (n_3003, wc205, n_2385);
  not gc205 (wc205, n_2556);
  and g3429 (n_2692, wc206, n_2562);
  not gc206 (wc206, n_2563);
  and g3430 (n_2700, wc207, n_2397);
  not gc207 (wc207, n_2566);
  and g3431 (n_2704, wc208, n_2572);
  not gc208 (wc208, n_2573);
  and g3432 (n_2819, wc209, n_2409);
  not gc209 (wc209, n_2576);
  and g3433 (n_2707, wc210, n_2582);
  not gc210 (wc210, n_2583);
  and g3434 (n_2715, wc211, n_2421);
  not gc211 (wc211, n_2586);
  and g3435 (n_2719, wc212, n_2592);
  not gc212 (wc212, n_2593);
  or g3436 (n_2941, wc213, n_2438);
  not gc213 (wc213, n_2598);
  and g3437 (n_2613, wc214, n_2610);
  not gc214 (wc214, n_2605);
  and g3438 (n_2893, wc215, n_2343);
  not gc215 (wc215, n_2663);
  and g3439 (n_2896, wc216, n_2525);
  not gc216 (wc216, n_2667);
  and g3440 (n_2864, wc217, n_2463);
  not gc217 (wc217, n_2738);
  and g3441 (n_2869, wc218, n_2625);
  not gc218 (wc218, n_2742);
  and g3442 (n_2874, n_2745, wc219);
  not gc219 (wc219, n_2746);
  and g3443 (n_2879, n_2749, wc220);
  not gc220 (wc220, n_2750);
  or g3444 (n_2902, wc221, n_2360);
  not gc221 (wc221, n_2777);
  or g3445 (n_2910, n_2782, wc222);
  not gc222 (wc222, n_2777);
  or g3446 (n_2914, wc223, n_2680);
  not gc223 (wc223, n_2777);
  or g3447 (n_3017, wc224, n_2408);
  not gc224 (wc224, n_2813);
  or g3448 (n_3025, n_2818, wc225);
  not gc225 (wc225, n_2813);
  or g3449 (n_3029, wc226, n_2710);
  not gc226 (wc226, n_2813);
  or g3450 (n_3221, wc227, n_2438);
  not gc227 (wc227, n_2433);
  and g3451 (n_2942, wc228, n_2433);
  not gc228 (wc228, n_2596);
  and g3452 (n_2603, wc229, n_2600);
  not gc229 (wc229, n_2595);
  and g3453 (n_2730, wc230, n_2445);
  not gc230 (wc230, n_2606);
  and g3454 (n_2734, wc231, n_2612);
  not gc231 (wc231, n_2613);
  and g3455 (n_2899, n_2670, wc232);
  not gc232 (wc232, n_2671);
  and g3456 (n_2682, wc233, n_2548);
  not gc233 (wc233, n_2677);
  and g3457 (n_2697, wc234, n_2568);
  not gc234 (wc234, n_2692);
  and g3458 (n_2712, wc235, n_2588);
  not gc235 (wc235, n_2707);
  and g3459 (n_2952, wc236, n_2608);
  not gc236 (wc236, n_2725);
  or g3460 (n_2884, wc237, n_2336);
  not gc237 (wc237, n_2882);
  or g3461 (n_2889, n_2886, wc238);
  not gc238 (wc238, n_2882);
  or g3462 (n_2891, wc239, n_2665);
  not gc239 (wc239, n_2882);
  and g3463 (n_3050, wc240, n_2598);
  not gc240 (wc240, n_2937);
  and g3464 (n_2722, wc241, n_2602);
  not gc241 (wc241, n_2603);
  and g3465 (n_2774, n_2674, wc242);
  not gc242 (wc242, n_2675);
  and g3466 (n_2792, wc243, n_2367);
  not gc243 (wc243, n_2678);
  and g3467 (n_2797, wc244, n_2545);
  not gc244 (wc244, n_2682);
  and g3468 (n_2802, n_2685, wc245);
  not gc245 (wc245, n_2686);
  and g3469 (n_2807, n_2689, wc246);
  not gc246 (wc246, n_2690);
  and g3470 (n_3008, wc247, n_2391);
  not gc247 (wc247, n_2693);
  and g3471 (n_3011, wc248, n_2565);
  not gc248 (wc248, n_2697);
  and g3472 (n_3014, n_2700, wc249);
  not gc249 (wc249, n_2701);
  and g3473 (n_2810, n_2704, wc250);
  not gc250 (wc250, n_2705);
  and g3474 (n_2828, wc251, n_2415);
  not gc251 (wc251, n_2708);
  and g3475 (n_2833, wc252, n_2585);
  not gc252 (wc252, n_2712);
  and g3476 (n_2838, n_2715, wc253);
  not gc253 (wc253, n_2716);
  and g3477 (n_2843, n_2719, wc254);
  not gc254 (wc254, n_2720);
  or g3478 (n_2965, wc255, n_2456);
  not gc255 (wc255, n_2849);
  or g3479 (n_2973, n_2854, wc256);
  not gc256 (wc256, n_2849);
  or g3480 (n_2977, wc257, n_2740);
  not gc257 (wc257, n_2849);
  or g3481 (n_2905, n_2902, wc258);
  not gc258 (wc258, n_2882);
  or g3482 (n_2909, n_2906, wc259);
  not gc259 (wc259, n_2882);
  or g3483 (n_2913, n_2910, wc260);
  not gc260 (wc260, n_2882);
  or g3484 (n_2917, n_2914, wc261);
  not gc261 (wc261, n_2882);
  or g3485 (n_2921, n_2918, wc262);
  not gc262 (wc262, n_2882);
  or g3486 (n_2925, n_2922, wc263);
  not gc263 (wc263, n_2882);
  or g3487 (n_2929, n_2926, wc264);
  not gc264 (wc264, n_2882);
  or g3488 (n_2933, n_2930, wc265);
  not gc265 (wc265, n_2882);
  and g3489 (n_2727, wc266, n_2608);
  not gc266 (wc266, n_2722);
  and g3490 (n_2780, wc267, n_2538);
  not gc267 (wc267, n_2774);
  and g3491 (n_2793, wc268, n_2790);
  not gc268 (wc268, n_2774);
  and g3492 (n_2798, wc269, n_2795);
  not gc269 (wc269, n_2774);
  and g3493 (n_2803, wc270, n_2800);
  not gc270 (wc270, n_2774);
  and g3494 (n_2808, wc271, n_2805);
  not gc271 (wc271, n_2774);
  and g3495 (n_2816, wc272, n_2578);
  not gc272 (wc272, n_2810);
  and g3496 (n_2829, wc273, n_2826);
  not gc273 (wc273, n_2810);
  and g3497 (n_2834, wc274, n_2831);
  not gc274 (wc274, n_2810);
  and g3498 (n_2839, wc275, n_2836);
  not gc275 (wc275, n_2810);
  and g3499 (n_2844, wc276, n_2841);
  not gc276 (wc276, n_2810);
  and g3500 (n_3059, wc277, n_2947);
  not gc277 (wc277, n_2937);
  and g3501 (n_3062, n_2952, wc278);
  not gc278 (wc278, n_2937);
  and g3502 (n_3065, wc279, n_2957);
  not gc279 (wc279, n_2937);
  and g3503 (n_3068, wc280, n_2849);
  not gc280 (wc280, n_2937);
  and g3504 (n_2949, wc281, n_2439);
  not gc281 (wc281, n_2723);
  and g3505 (n_2954, wc282, n_2605);
  not gc282 (wc282, n_2727);
  and g3506 (n_2959, n_2730, wc283);
  not gc283 (wc283, n_2731);
  and g3507 (n_2846, n_2734, wc284);
  not gc284 (wc284, n_2735);
  and g3508 (n_2904, wc285, n_2355);
  not gc285 (wc285, n_2775);
  and g3509 (n_2908, wc286, n_2535);
  not gc286 (wc286, n_2780);
  and g3510 (n_2912, n_2783, wc287);
  not gc287 (wc287, n_2784);
  and g3511 (n_2916, n_2677, wc288);
  not gc288 (wc288, n_2787);
  and g3512 (n_2920, wc289, n_2792);
  not gc289 (wc289, n_2793);
  and g3513 (n_2924, wc290, n_2797);
  not gc290 (wc290, n_2798);
  and g3514 (n_2928, wc291, n_2802);
  not gc291 (wc291, n_2803);
  and g3515 (n_2932, wc292, n_2807);
  not gc292 (wc292, n_2808);
  and g3516 (n_3019, wc293, n_2403);
  not gc293 (wc293, n_2811);
  and g3517 (n_3023, wc294, n_2575);
  not gc294 (wc294, n_2816);
  and g3518 (n_3027, n_2819, wc295);
  not gc295 (wc295, n_2820);
  and g3519 (n_3031, n_2707, wc296);
  not gc296 (wc296, n_2823);
  and g3520 (n_3035, wc297, n_2828);
  not gc297 (wc297, n_2829);
  and g3521 (n_3039, wc298, n_2833);
  not gc298 (wc298, n_2834);
  and g3522 (n_3043, wc299, n_2838);
  not gc299 (wc299, n_2839);
  and g3523 (n_2934, wc300, n_2843);
  not gc300 (wc300, n_2844);
  and g3524 (n_2852, wc301, n_2618);
  not gc301 (wc301, n_2846);
  and g3525 (n_2865, wc302, n_2862);
  not gc302 (wc302, n_2846);
  and g3526 (n_2870, wc303, n_2867);
  not gc303 (wc303, n_2846);
  and g3527 (n_2875, wc304, n_2872);
  not gc304 (wc304, n_2846);
  and g3528 (n_2880, wc305, n_2877);
  not gc305 (wc305, n_2846);
  and g3529 (n_2939, wc306, n_2598);
  not gc306 (wc306, n_2934);
  and g3530 (n_2950, wc307, n_2947);
  not gc307 (wc307, n_2934);
  and g3531 (n_2955, wc308, n_2952);
  not gc308 (wc308, n_2934);
  and g3532 (n_2960, wc309, n_2957);
  not gc309 (wc309, n_2934);
  and g3533 (n_2963, wc310, n_2849);
  not gc310 (wc310, n_2934);
  and g3534 (n_2966, wc311, n_2451);
  not gc311 (wc311, n_2847);
  and g3535 (n_2970, wc312, n_2615);
  not gc312 (wc312, n_2852);
  and g3536 (n_2974, n_2855, wc313);
  not gc313 (wc313, n_2856);
  and g3537 (n_2978, n_2737, wc314);
  not gc314 (wc314, n_2859);
  and g3538 (n_2982, wc315, n_2864);
  not gc315 (wc315, n_2865);
  and g3539 (n_2986, wc316, n_2869);
  not gc316 (wc316, n_2870);
  and g3540 (n_2990, wc317, n_2874);
  not gc317 (wc317, n_2875);
  and g3541 (n_2994, wc318, n_2879);
  not gc318 (wc318, n_2880);
  and g3542 (n_3048, wc319, n_2427);
  not gc319 (wc319, n_2935);
  and g3543 (n_3051, wc320, n_2595);
  not gc320 (wc320, n_2939);
  and g3544 (n_3054, n_2942, wc321);
  not gc321 (wc321, n_2943);
  and g3545 (n_3057, n_2722, wc322);
  not gc322 (wc322, n_2945);
  and g3546 (n_3060, wc323, n_2949);
  not gc323 (wc323, n_2950);
  and g3547 (n_3063, wc324, n_2954);
  not gc324 (wc324, n_2955);
  and g3548 (n_3066, wc325, n_2959);
  not gc325 (wc325, n_2960);
  and g3549 (n_3069, wc326, n_2846);
  not gc326 (wc326, n_2963);
  or g3550 (n_2999, wc327, n_2384);
  not gc327 (wc327, n_2997);
  or g3551 (n_3004, n_3001, wc328);
  not gc328 (wc328, n_2997);
  or g3552 (n_3006, wc329, n_2695);
  not gc329 (wc329, n_2997);
  or g3553 (n_3020, n_3017, wc330);
  not gc330 (wc330, n_2997);
  or g3554 (n_3024, wc331, n_3021);
  not gc331 (wc331, n_2997);
  or g3555 (n_3028, n_3025, wc332);
  not gc332 (wc332, n_2997);
  or g3556 (n_3032, n_3029, wc333);
  not gc333 (wc333, n_2997);
  or g3557 (n_3036, wc334, n_3033);
  not gc334 (wc334, n_2997);
  or g3558 (n_3040, wc335, n_3037);
  not gc335 (wc335, n_2997);
  or g3559 (n_3044, wc336, n_3041);
  not gc336 (wc336, n_2997);
  or g3560 (n_3046, wc337, n_2937);
  not gc337 (wc337, n_2997);
  and g3561 (n_3072, n_2966, wc338);
  not gc338 (wc338, n_2967);
  and g3562 (n_3075, n_2970, wc339);
  not gc339 (wc339, n_2971);
  and g3563 (n_3078, n_2974, wc340);
  not gc340 (wc340, n_2975);
  and g3564 (n_3081, n_2978, wc341);
  not gc341 (wc341, n_2979);
  and g3565 (n_3084, n_2982, wc342);
  not gc342 (wc342, n_2983);
  and g3566 (n_3087, n_2986, wc343);
  not gc343 (wc343, n_2987);
  and g3567 (n_3090, n_2990, wc344);
  not gc344 (wc344, n_2991);
  and g3568 (n_3093, n_2994, wc345);
  not gc345 (wc345, n_2995);
  or g3569 (n_3097, n_2478, wc346);
  not gc346 (wc346, n_3095);
  not g3570 (Z[65], n_3259);
endmodule

module mult_signed_const_10350_GENERIC(A, Z);
  input [46:0] A;
  output [65:0] Z;
  wire [46:0] A;
  wire [65:0] Z;
  mult_signed_const_10350_GENERIC_REAL g1(.A ({A[46:2], A[0], A[0]}),
       .Z (Z));
endmodule

module mult_signed_const_10729_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [47:0] A;
  output [66:0] Z;
  wire [47:0] A;
  wire [66:0] Z;
  wire n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59;
  wire n_60, n_61, n_62, n_63, n_64, n_65, n_66, n_67;
  wire n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_113, n_114, n_115, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_251, n_252;
  wire n_253, n_254, n_255, n_256, n_257, n_258, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_265, n_266, n_267, n_268;
  wire n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276;
  wire n_277, n_278, n_279, n_280, n_281, n_282, n_283, n_284;
  wire n_285, n_286, n_287, n_288, n_289, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_328, n_329, n_330, n_331, n_332, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560;
  wire n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584;
  wire n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592;
  wire n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600;
  wire n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608;
  wire n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616;
  wire n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648;
  wire n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656;
  wire n_657, n_658, n_659, n_660, n_661, n_662, n_664, n_665;
  wire n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_678, n_679, n_680, n_681, n_682, n_683;
  wire n_684, n_685, n_686, n_687, n_688, n_690, n_691, n_692;
  wire n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700;
  wire n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708;
  wire n_709, n_710, n_711, n_712, n_713, n_714, n_716, n_717;
  wire n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725;
  wire n_726, n_727, n_731, n_732, n_733, n_734, n_735, n_736;
  wire n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_747;
  wire n_748, n_749, n_750, n_753, n_754, n_755, n_756, n_757;
  wire n_758, n_759, n_760, n_762, n_763, n_766, n_767, n_768;
  wire n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_778;
  wire n_779, n_780, n_783, n_784, n_785, n_786, n_787, n_788;
  wire n_789, n_790, n_793, n_795, n_796, n_797, n_798, n_799;
  wire n_800, n_801, n_802, n_803, n_806, n_807, n_808, n_809;
  wire n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_818;
  wire n_819, n_821, n_822, n_823, n_824, n_825, n_826, n_827;
  wire n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838;
  wire n_840, n_843, n_844, n_845, n_846, n_847, n_853, n_854;
  wire n_855, n_856, n_860, n_861, n_862, n_863, n_867, n_868;
  wire n_869, n_870, n_872, n_874, n_875, n_879, n_880, n_882;
  wire n_883, n_886, n_889, n_890, n_891, n_892, n_893, n_894;
  wire n_895, n_896, n_897, n_898, n_900, n_901, n_902, n_903;
  wire n_904, n_907, n_909, n_910, n_911, n_912, n_913, n_914;
  wire n_915, n_916, n_917, n_919, n_920, n_921, n_922, n_923;
  wire n_924, n_927, n_929, n_930, n_931, n_932, n_933, n_934;
  wire n_935, n_936, n_937, n_938, n_939, n_940, n_941, n_945;
  wire n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_955;
  wire n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966;
  wire n_967, n_968, n_969, n_970, n_971, n_972, n_973, n_977;
  wire n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985;
  wire n_986, n_987, n_988, n_991, n_997, n_998, n_999, n_1000;
  wire n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008;
  wire n_1009, n_1010, n_1011, n_1012, n_1013, n_1016, n_1019, n_1020;
  wire n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028;
  wire n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1037;
  wire n_1038, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046;
  wire n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054;
  wire n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1063;
  wire n_1065, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074;
  wire n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082;
  wire n_1083, n_1084, n_1085, n_1088, n_1089, n_1090, n_1091, n_1093;
  wire n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101;
  wire n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109;
  wire n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1119;
  wire n_1121, n_1122, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130;
  wire n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138;
  wire n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146;
  wire n_1147, n_1148, n_1153, n_1154, n_1155, n_1157, n_1158, n_1159;
  wire n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167;
  wire n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175;
  wire n_1176, n_1177, n_1178, n_1179, n_1180, n_1185, n_1186, n_1189;
  wire n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197;
  wire n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205;
  wire n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1215;
  wire n_1217, n_1218, n_1219, n_1221, n_1222, n_1223, n_1224, n_1225;
  wire n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233;
  wire n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241;
  wire n_1242, n_1243, n_1244, n_1247, n_1249, n_1250, n_1253, n_1254;
  wire n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262;
  wire n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270;
  wire n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1279, n_1281;
  wire n_1282, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291;
  wire n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299;
  wire n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307;
  wire n_1308, n_1311, n_1313, n_1314, n_1317, n_1318, n_1319, n_1320;
  wire n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328;
  wire n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336;
  wire n_1337, n_1338, n_1339, n_1340, n_1343, n_1345, n_1346, n_1349;
  wire n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1375;
  wire n_1377, n_1378, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386;
  wire n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394;
  wire n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402;
  wire n_1403, n_1404, n_1407, n_1409, n_1410, n_1413, n_1414, n_1415;
  wire n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423;
  wire n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431;
  wire n_1432, n_1433, n_1434, n_1435, n_1436, n_1439, n_1441, n_1442;
  wire n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452;
  wire n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460;
  wire n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468;
  wire n_1471, n_1473, n_1474, n_1477, n_1478, n_1479, n_1480, n_1481;
  wire n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489;
  wire n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
  wire n_1498, n_1499, n_1500, n_1503, n_1505, n_1506, n_1509, n_1510;
  wire n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518;
  wire n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526;
  wire n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1535, n_1537;
  wire n_1538, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547;
  wire n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555;
  wire n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563;
  wire n_1564, n_1567, n_1569, n_1570, n_1573, n_1574, n_1575, n_1576;
  wire n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584;
  wire n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592;
  wire n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1601;
  wire n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611;
  wire n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619;
  wire n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627;
  wire n_1628, n_1629, n_1630, n_1631, n_1633, n_1636, n_1637, n_1638;
  wire n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646;
  wire n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654;
  wire n_1655, n_1656, n_1660, n_1661, n_1663, n_1667, n_1668, n_1669;
  wire n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677;
  wire n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685;
  wire n_1686, n_1687, n_1688, n_1692, n_1693, n_1695, n_1699, n_1700;
  wire n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708;
  wire n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716;
  wire n_1717, n_1718, n_1719, n_1720, n_1724, n_1729, n_1730, n_1731;
  wire n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739;
  wire n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747;
  wire n_1748, n_1749, n_1750, n_1751, n_1752, n_1756, n_1761, n_1762;
  wire n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770;
  wire n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778;
  wire n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1789;
  wire n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800;
  wire n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1821, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830;
  wire n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838;
  wire n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846;
  wire n_1847, n_1848, n_1855, n_1856, n_1861, n_1862, n_1863, n_1864;
  wire n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872;
  wire n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880;
  wire n_1887, n_1888, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898;
  wire n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906;
  wire n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1917, n_1919;
  wire n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927;
  wire n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935;
  wire n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943;
  wire n_1944, n_1949, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956;
  wire n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964;
  wire n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972;
  wire n_1973, n_1974, n_1975, n_1976, n_1981, n_1982, n_1983, n_1984;
  wire n_1985, n_1987, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994;
  wire n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002;
  wire n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010;
  wire n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2019, n_2021;
  wire n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029;
  wire n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037;
  wire n_2038, n_2039, n_2040, n_2043, n_2044, n_2053, n_2054, n_2055;
  wire n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063;
  wire n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071;
  wire n_2072, n_2073, n_2074, n_2076, n_2077, n_2079, n_2081, n_2082;
  wire n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091;
  wire n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099;
  wire n_2100, n_2101, n_2102, n_2103, n_2104, n_2113, n_2114, n_2115;
  wire n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123;
  wire n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131;
  wire n_2132, n_2135, n_2136, n_2137, n_2140, n_2141, n_2143, n_2144;
  wire n_2145, n_2146, n_2147, n_2149, n_2150, n_2151, n_2152, n_2153;
  wire n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161;
  wire n_2164, n_2165, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173;
  wire n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181;
  wire n_2182, n_2183, n_2184, n_2185, n_2188, n_2193, n_2194, n_2195;
  wire n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203;
  wire n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2211, n_2215;
  wire n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223;
  wire n_2224, n_2225, n_2226, n_2227, n_2228, n_2237, n_2238, n_2239;
  wire n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247;
  wire n_2248, n_2255, n_2256, n_2257, n_2259, n_2260, n_2261, n_2262;
  wire n_2263, n_2264, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276;
  wire n_2277, n_2278, n_2279, n_2280, n_2283, n_2284, n_2285, n_2286;
  wire n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2297, n_2298;
  wire n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2307;
  wire n_2308, n_2309, n_2310, n_2311, n_2312, n_2315, n_2317, n_2318;
  wire n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2327, n_2328;
  wire n_2340, n_2342, n_2344, n_2345, n_2346, n_2347, n_2348, n_2350;
  wire n_2351, n_2352, n_2353, n_2354, n_2356, n_2357, n_2358, n_2359;
  wire n_2360, n_2362, n_2363, n_2364, n_2365, n_2366, n_2368, n_2369;
  wire n_2370, n_2371, n_2372, n_2374, n_2375, n_2376, n_2377, n_2378;
  wire n_2380, n_2381, n_2382, n_2383, n_2384, n_2386, n_2387, n_2388;
  wire n_2389, n_2390, n_2392, n_2393, n_2394, n_2395, n_2396, n_2398;
  wire n_2399, n_2400, n_2401, n_2402, n_2404, n_2405, n_2406, n_2407;
  wire n_2408, n_2410, n_2411, n_2412, n_2413, n_2414, n_2416, n_2417;
  wire n_2418, n_2419, n_2420, n_2422, n_2423, n_2424, n_2425, n_2426;
  wire n_2428, n_2429, n_2430, n_2431, n_2432, n_2434, n_2435, n_2436;
  wire n_2437, n_2438, n_2440, n_2441, n_2442, n_2443, n_2444, n_2446;
  wire n_2447, n_2448, n_2449, n_2450, n_2452, n_2453, n_2454, n_2455;
  wire n_2456, n_2458, n_2459, n_2460, n_2461, n_2462, n_2464, n_2465;
  wire n_2466, n_2467, n_2468, n_2470, n_2471, n_2472, n_2473, n_2474;
  wire n_2476, n_2477, n_2478, n_2479, n_2480, n_2482, n_2483, n_2484;
  wire n_2485, n_2486, n_2488, n_2489, n_2490, n_2491, n_2492, n_2494;
  wire n_2495, n_2496, n_2497, n_2498, n_2500, n_2501, n_2502, n_2503;
  wire n_2504, n_2506, n_2507, n_2508, n_2509, n_2510, n_2512, n_2513;
  wire n_2514, n_2515, n_2516, n_2518, n_2519, n_2520, n_2521, n_2522;
  wire n_2524, n_2525, n_2526, n_2527, n_2528, n_2530, n_2533, n_2535;
  wire n_2536, n_2538, n_2539, n_2541, n_2542, n_2543, n_2545, n_2546;
  wire n_2548, n_2549, n_2550, n_2552, n_2553, n_2555, n_2556, n_2557;
  wire n_2559, n_2560, n_2562, n_2563, n_2564, n_2566, n_2567, n_2569;
  wire n_2570, n_2571, n_2573, n_2574, n_2576, n_2577, n_2578, n_2580;
  wire n_2581, n_2583, n_2584, n_2585, n_2587, n_2588, n_2590, n_2591;
  wire n_2592, n_2594, n_2595, n_2597, n_2598, n_2599, n_2601, n_2602;
  wire n_2604, n_2605, n_2606, n_2608, n_2609, n_2611, n_2612, n_2613;
  wire n_2615, n_2616, n_2618, n_2619, n_2620, n_2622, n_2623, n_2625;
  wire n_2626, n_2627, n_2629, n_2630, n_2632, n_2633, n_2634, n_2636;
  wire n_2637, n_2639, n_2640, n_2643, n_2644, n_2645, n_2646, n_2647;
  wire n_2648, n_2650, n_2651, n_2652, n_2653, n_2654, n_2656, n_2657;
  wire n_2658, n_2659, n_2660, n_2662, n_2663, n_2664, n_2665, n_2666;
  wire n_2668, n_2669, n_2670, n_2671, n_2672, n_2674, n_2675, n_2676;
  wire n_2677, n_2678, n_2680, n_2681, n_2682, n_2683, n_2684, n_2686;
  wire n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2694, n_2695;
  wire n_2697, n_2698, n_2699, n_2701, n_2702, n_2704, n_2705, n_2706;
  wire n_2708, n_2709, n_2711, n_2712, n_2713, n_2715, n_2716, n_2717;
  wire n_2718, n_2719, n_2720, n_2722, n_2723, n_2724, n_2725, n_2726;
  wire n_2728, n_2729, n_2730, n_2731, n_2732, n_2734, n_2736, n_2737;
  wire n_2739, n_2741, n_2742, n_2744, n_2746, n_2747, n_2749, n_2750;
  wire n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758;
  wire n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766;
  wire n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774;
  wire n_2775, n_2779, n_2780, n_2782, n_2784, n_2785, n_2787, n_2789;
  wire n_2790, n_2792, n_2794, n_2795, n_2797, n_2799, n_2800, n_2802;
  wire n_2804, n_2805, n_2807, n_2809, n_2810, n_2812, n_2814, n_2815;
  wire n_2817, n_2819, n_2820, n_2822, n_2824, n_2825, n_2827, n_2829;
  wire n_2830, n_2832, n_2834, n_2835, n_2837, n_2839, n_2840, n_2842;
  wire n_2844, n_2845, n_2847, n_2849, n_2850, n_2852, n_2854, n_2856;
  wire n_2860, n_2863, n_2864, n_2866, n_2867, n_2868, n_2870, n_2871;
  wire n_2872, n_2874, n_2875, n_2876, n_2878, n_2879, n_2880, n_2882;
  wire n_2883, n_2884, n_2886, n_2887, n_2888, n_2890, n_2891, n_2892;
  wire n_2894, n_2895, n_2896, n_2898, n_2899, n_2900, n_2902, n_2903;
  wire n_2904, n_2906, n_2907, n_2908, n_2910, n_2911, n_2912, n_2914;
  wire n_2915, n_2916, n_2918, n_2919, n_2920, n_2922, n_2923, n_2924;
  wire n_2926, n_2927, n_2928, n_2930, n_2931, n_2932, n_2934, n_2935;
  wire n_2936, n_2938, n_2939, n_2940, n_2942, n_2943, n_2944, n_2946;
  wire n_2947, n_2948, n_2950, n_2951, n_2952, n_2954, n_2955, n_2956;
  wire n_2958, n_2959, n_2960, n_2962, n_2963, n_2964, n_2966, n_2967;
  wire n_2968, n_2970, n_2971, n_2972, n_2974, n_2975, n_2976, n_2978;
  wire n_2979, n_2980, n_2982, n_2983, n_2984, n_2986, n_2987;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g380 (n_178, A[4], A[2]);
  and g2 (n_110, A[4], A[2]);
  xor g381 (n_889, A[5], A[3]);
  xor g382 (n_177, n_889, A[1]);
  nand g3 (n_890, A[5], A[3]);
  nand g383 (n_891, A[1], A[3]);
  nand g384 (n_892, A[5], A[1]);
  nand g385 (n_109, n_890, n_891, n_892);
  xor g386 (n_251, A[6], A[4]);
  and g387 (n_252, A[6], A[4]);
  xor g388 (n_893, A[2], A[0]);
  xor g389 (n_176, n_893, n_251);
  nand g390 (n_894, A[2], A[0]);
  nand g4 (n_895, n_251, A[0]);
  nand g5 (n_896, A[2], n_251);
  nand g391 (n_108, n_894, n_895, n_896);
  xor g392 (n_897, A[7], A[5]);
  xor g393 (n_253, n_897, A[1]);
  nand g394 (n_898, A[7], A[5]);
  nand g396 (n_900, A[7], A[1]);
  nand g6 (n_255, n_898, n_892, n_900);
  xor g397 (n_901, A[3], n_252);
  xor g398 (n_175, n_901, n_253);
  nand g399 (n_902, A[3], n_252);
  nand g400 (n_903, n_253, n_252);
  nand g401 (n_904, A[3], n_253);
  nand g402 (n_107, n_902, n_903, n_904);
  xor g403 (n_254, A[8], A[6]);
  and g404 (n_257, A[8], A[6]);
  xor g406 (n_256, n_178, A[0]);
  nand g408 (n_907, A[0], A[4]);
  xor g411 (n_909, n_254, n_255);
  xor g412 (n_174, n_909, n_256);
  nand g413 (n_910, n_254, n_255);
  nand g414 (n_911, n_256, n_255);
  nand g415 (n_912, n_254, n_256);
  nand g416 (n_106, n_910, n_911, n_912);
  xor g417 (n_913, A[9], A[7]);
  xor g418 (n_259, n_913, A[3]);
  nand g419 (n_914, A[9], A[7]);
  nand g420 (n_915, A[3], A[7]);
  nand g421 (n_916, A[9], A[3]);
  nand g422 (n_262, n_914, n_915, n_916);
  xor g423 (n_917, A[1], A[5]);
  xor g424 (n_260, n_917, n_257);
  nand g426 (n_919, n_257, A[5]);
  nand g427 (n_920, A[1], n_257);
  nand g428 (n_264, n_892, n_919, n_920);
  xor g429 (n_921, n_258, n_259);
  xor g430 (n_173, n_921, n_260);
  nand g431 (n_922, n_258, n_259);
  nand g432 (n_923, n_260, n_259);
  nand g433 (n_924, n_258, n_260);
  nand g434 (n_105, n_922, n_923, n_924);
  xor g435 (n_261, A[10], A[8]);
  and g436 (n_266, A[10], A[8]);
  xor g438 (n_263, n_178, A[6]);
  nand g440 (n_927, A[6], A[2]);
  xor g443 (n_929, A[0], n_261);
  xor g444 (n_265, n_929, n_262);
  nand g445 (n_930, A[0], n_261);
  nand g446 (n_931, n_262, n_261);
  nand g447 (n_932, A[0], n_262);
  nand g448 (n_270, n_930, n_931, n_932);
  xor g449 (n_933, n_263, n_264);
  xor g450 (n_172, n_933, n_265);
  nand g451 (n_934, n_263, n_264);
  nand g452 (n_935, n_265, n_264);
  nand g453 (n_936, n_263, n_265);
  nand g454 (n_104, n_934, n_935, n_936);
  xor g455 (n_937, A[11], A[9]);
  xor g456 (n_268, n_937, A[5]);
  nand g457 (n_938, A[11], A[9]);
  nand g458 (n_939, A[5], A[9]);
  nand g459 (n_940, A[11], A[5]);
  nand g460 (n_273, n_938, n_939, n_940);
  xor g461 (n_941, A[3], A[7]);
  xor g462 (n_269, n_941, A[1]);
  nand g466 (n_274, n_915, n_900, n_891);
  xor g467 (n_945, n_266, n_267);
  xor g468 (n_271, n_945, n_268);
  nand g469 (n_946, n_266, n_267);
  nand g470 (n_947, n_268, n_267);
  nand g471 (n_948, n_266, n_268);
  nand g472 (n_278, n_946, n_947, n_948);
  xor g473 (n_949, n_269, n_270);
  xor g474 (n_171, n_949, n_271);
  nand g475 (n_950, n_269, n_270);
  nand g476 (n_951, n_271, n_270);
  nand g477 (n_952, n_269, n_271);
  nand g478 (n_103, n_950, n_951, n_952);
  xor g479 (n_272, A[12], A[10]);
  and g480 (n_279, A[12], A[10]);
  xor g482 (n_275, n_251, A[8]);
  nand g484 (n_955, A[8], A[4]);
  xor g488 (n_276, n_893, n_272);
  nand g490 (n_959, n_272, A[0]);
  nand g491 (n_960, A[2], n_272);
  nand g492 (n_283, n_894, n_959, n_960);
  xor g493 (n_961, n_273, n_274);
  xor g494 (n_277, n_961, n_275);
  nand g495 (n_962, n_273, n_274);
  nand g496 (n_963, n_275, n_274);
  nand g497 (n_964, n_273, n_275);
  nand g498 (n_285, n_962, n_963, n_964);
  xor g499 (n_965, n_276, n_277);
  xor g500 (n_170, n_965, n_278);
  nand g501 (n_966, n_276, n_277);
  nand g502 (n_967, n_278, n_277);
  nand g503 (n_968, n_276, n_278);
  nand g504 (n_102, n_966, n_967, n_968);
  xor g505 (n_969, A[13], A[11]);
  xor g506 (n_282, n_969, A[7]);
  nand g507 (n_970, A[13], A[11]);
  nand g508 (n_971, A[7], A[11]);
  nand g509 (n_972, A[13], A[7]);
  nand g510 (n_288, n_970, n_971, n_972);
  xor g511 (n_973, A[5], A[9]);
  xor g512 (n_281, n_973, A[3]);
  nand g516 (n_289, n_939, n_916, n_890);
  xor g517 (n_977, A[1], n_279);
  xor g518 (n_284, n_977, n_280);
  nand g519 (n_978, A[1], n_279);
  nand g520 (n_979, n_280, n_279);
  nand g521 (n_980, A[1], n_280);
  nand g522 (n_292, n_978, n_979, n_980);
  xor g523 (n_981, n_281, n_282);
  xor g524 (n_286, n_981, n_283);
  nand g525 (n_982, n_281, n_282);
  nand g526 (n_983, n_283, n_282);
  nand g527 (n_984, n_281, n_283);
  nand g528 (n_294, n_982, n_983, n_984);
  xor g529 (n_985, n_284, n_285);
  xor g530 (n_169, n_985, n_286);
  nand g531 (n_986, n_284, n_285);
  nand g532 (n_987, n_286, n_285);
  nand g533 (n_988, n_284, n_286);
  nand g534 (n_101, n_986, n_987, n_988);
  xor g535 (n_287, A[14], A[12]);
  and g536 (n_296, A[14], A[12]);
  xor g538 (n_291, n_254, A[10]);
  nand g540 (n_991, A[10], A[6]);
  xor g549 (n_997, n_287, n_288);
  xor g550 (n_293, n_997, n_289);
  nand g551 (n_998, n_287, n_288);
  nand g552 (n_999, n_289, n_288);
  nand g553 (n_1000, n_287, n_289);
  nand g554 (n_302, n_998, n_999, n_1000);
  xor g555 (n_1001, n_256, n_291);
  xor g556 (n_295, n_1001, n_292);
  nand g557 (n_1002, n_256, n_291);
  nand g558 (n_1003, n_292, n_291);
  nand g559 (n_1004, n_256, n_292);
  nand g560 (n_305, n_1002, n_1003, n_1004);
  xor g561 (n_1005, n_293, n_294);
  xor g562 (n_168, n_1005, n_295);
  nand g563 (n_1006, n_293, n_294);
  nand g564 (n_1007, n_295, n_294);
  nand g565 (n_1008, n_293, n_295);
  nand g566 (n_100, n_1006, n_1007, n_1008);
  xor g567 (n_1009, A[15], A[13]);
  xor g568 (n_298, n_1009, A[9]);
  nand g569 (n_1010, A[15], A[13]);
  nand g570 (n_1011, A[9], A[13]);
  nand g571 (n_1012, A[15], A[9]);
  nand g572 (n_307, n_1010, n_1011, n_1012);
  xor g573 (n_1013, A[1], A[7]);
  xor g574 (n_299, n_1013, A[11]);
  nand g577 (n_1016, A[1], A[11]);
  nand g578 (n_308, n_900, n_971, n_1016);
  xor g580 (n_301, n_889, n_296);
  nand g582 (n_1019, n_296, A[3]);
  nand g583 (n_1020, A[5], n_296);
  nand g584 (n_311, n_890, n_1019, n_1020);
  xor g585 (n_1021, n_297, n_298);
  xor g586 (n_303, n_1021, n_299);
  nand g587 (n_1022, n_297, n_298);
  nand g588 (n_1023, n_299, n_298);
  nand g589 (n_1024, n_297, n_299);
  nand g590 (n_313, n_1022, n_1023, n_1024);
  xor g591 (n_1025, n_258, n_301);
  xor g592 (n_304, n_1025, n_302);
  nand g593 (n_1026, n_258, n_301);
  nand g594 (n_1027, n_302, n_301);
  nand g595 (n_1028, n_258, n_302);
  nand g596 (n_315, n_1026, n_1027, n_1028);
  xor g597 (n_1029, n_303, n_304);
  xor g598 (n_167, n_1029, n_305);
  nand g599 (n_1030, n_303, n_304);
  nand g600 (n_1031, n_305, n_304);
  nand g601 (n_1032, n_303, n_305);
  nand g602 (n_99, n_1030, n_1031, n_1032);
  xor g603 (n_306, A[16], A[14]);
  and g604 (n_317, A[16], A[14]);
  xor g605 (n_1033, A[10], A[2]);
  xor g606 (n_310, n_1033, A[8]);
  nand g607 (n_1034, A[10], A[2]);
  nand g608 (n_1035, A[8], A[2]);
  xor g611 (n_1037, A[12], A[6]);
  xor g612 (n_309, n_1037, A[4]);
  nand g613 (n_1038, A[12], A[6]);
  nand g615 (n_1040, A[12], A[4]);
  xor g617 (n_1041, A[0], n_306);
  xor g618 (n_312, n_1041, n_307);
  nand g619 (n_1042, A[0], n_306);
  nand g620 (n_1043, n_307, n_306);
  nand g621 (n_1044, A[0], n_307);
  nand g622 (n_323, n_1042, n_1043, n_1044);
  xor g623 (n_1045, n_308, n_309);
  xor g624 (n_314, n_1045, n_310);
  nand g625 (n_1046, n_308, n_309);
  nand g626 (n_1047, n_310, n_309);
  nand g627 (n_1048, n_308, n_310);
  nand g628 (n_325, n_1046, n_1047, n_1048);
  xor g629 (n_1049, n_311, n_312);
  xor g630 (n_316, n_1049, n_313);
  nand g631 (n_1050, n_311, n_312);
  nand g632 (n_1051, n_313, n_312);
  nand g633 (n_1052, n_311, n_313);
  nand g634 (n_327, n_1050, n_1051, n_1052);
  xor g635 (n_1053, n_314, n_315);
  xor g636 (n_166, n_1053, n_316);
  nand g637 (n_1054, n_314, n_315);
  nand g638 (n_1055, n_316, n_315);
  nand g639 (n_1056, n_314, n_316);
  nand g640 (n_98, n_1054, n_1055, n_1056);
  xor g641 (n_1057, A[17], A[15]);
  xor g642 (n_321, n_1057, A[11]);
  nand g643 (n_1058, A[17], A[15]);
  nand g644 (n_1059, A[11], A[15]);
  nand g645 (n_1060, A[17], A[11]);
  nand g646 (n_330, n_1058, n_1059, n_1060);
  xor g647 (n_1061, A[3], A[1]);
  xor g648 (n_322, n_1061, A[9]);
  nand g650 (n_1063, A[9], A[1]);
  nand g652 (n_331, n_891, n_1063, n_916);
  xor g653 (n_1065, A[13], A[7]);
  xor g654 (n_320, n_1065, A[5]);
  nand g657 (n_1068, A[13], A[5]);
  nand g658 (n_332, n_972, n_898, n_1068);
  xor g659 (n_1069, n_317, n_318);
  xor g660 (n_324, n_1069, n_319);
  nand g661 (n_1070, n_317, n_318);
  nand g662 (n_1071, n_319, n_318);
  nand g663 (n_1072, n_317, n_319);
  nand g664 (n_336, n_1070, n_1071, n_1072);
  xor g665 (n_1073, n_320, n_321);
  xor g666 (n_326, n_1073, n_322);
  nand g667 (n_1074, n_320, n_321);
  nand g668 (n_1075, n_322, n_321);
  nand g669 (n_1076, n_320, n_322);
  nand g670 (n_338, n_1074, n_1075, n_1076);
  xor g671 (n_1077, n_323, n_324);
  xor g672 (n_328, n_1077, n_325);
  nand g673 (n_1078, n_323, n_324);
  nand g674 (n_1079, n_325, n_324);
  nand g675 (n_1080, n_323, n_325);
  nand g676 (n_340, n_1078, n_1079, n_1080);
  xor g677 (n_1081, n_326, n_327);
  xor g678 (n_165, n_1081, n_328);
  nand g679 (n_1082, n_326, n_327);
  nand g680 (n_1083, n_328, n_327);
  nand g681 (n_1084, n_326, n_328);
  nand g682 (n_97, n_1082, n_1083, n_1084);
  xor g683 (n_329, A[18], A[16]);
  and g684 (n_113, A[18], A[16]);
  xor g685 (n_1085, A[12], A[4]);
  xor g686 (n_334, n_1085, A[2]);
  nand g689 (n_1088, A[12], A[2]);
  xor g691 (n_1089, A[10], A[14]);
  xor g692 (n_333, n_1089, A[8]);
  nand g693 (n_1090, A[10], A[14]);
  nand g694 (n_1091, A[8], A[14]);
  xor g697 (n_1093, A[6], A[0]);
  xor g698 (n_335, n_1093, n_329);
  nand g699 (n_1094, A[6], A[0]);
  nand g700 (n_1095, n_329, A[0]);
  nand g701 (n_1096, A[6], n_329);
  nand g702 (n_344, n_1094, n_1095, n_1096);
  xor g703 (n_1097, n_330, n_331);
  xor g704 (n_337, n_1097, n_332);
  nand g705 (n_1098, n_330, n_331);
  nand g706 (n_1099, n_332, n_331);
  nand g707 (n_1100, n_330, n_332);
  nand g708 (n_346, n_1098, n_1099, n_1100);
  xor g709 (n_1101, n_333, n_334);
  xor g710 (n_339, n_1101, n_335);
  nand g711 (n_1102, n_333, n_334);
  nand g712 (n_1103, n_335, n_334);
  nand g713 (n_1104, n_333, n_335);
  nand g714 (n_347, n_1102, n_1103, n_1104);
  xor g715 (n_1105, n_336, n_337);
  xor g716 (n_111, n_1105, n_338);
  nand g717 (n_1106, n_336, n_337);
  nand g718 (n_1107, n_338, n_337);
  nand g719 (n_1108, n_336, n_338);
  nand g720 (n_350, n_1106, n_1107, n_1108);
  xor g721 (n_1109, n_339, n_340);
  xor g722 (n_164, n_1109, n_111);
  nand g723 (n_1110, n_339, n_340);
  nand g724 (n_1111, n_111, n_340);
  nand g725 (n_1112, n_339, n_111);
  nand g726 (n_96, n_1110, n_1111, n_1112);
  xor g727 (n_1113, A[19], A[17]);
  xor g728 (n_342, n_1113, A[13]);
  nand g729 (n_1114, A[19], A[17]);
  nand g730 (n_1115, A[13], A[17]);
  nand g731 (n_1116, A[19], A[13]);
  nand g732 (n_352, n_1114, n_1115, n_1116);
  xor g734 (n_343, n_889, A[11]);
  nand g736 (n_1119, A[11], A[3]);
  nand g738 (n_353, n_890, n_1119, n_940);
  xor g739 (n_1121, A[1], A[15]);
  xor g740 (n_341, n_1121, A[9]);
  nand g741 (n_1122, A[1], A[15]);
  nand g744 (n_354, n_1122, n_1012, n_1063);
  xor g745 (n_1125, A[7], n_113);
  xor g746 (n_345, n_1125, n_114);
  nand g747 (n_1126, A[7], n_113);
  nand g748 (n_1127, n_114, n_113);
  nand g749 (n_1128, A[7], n_114);
  nand g750 (n_358, n_1126, n_1127, n_1128);
  xor g751 (n_1129, n_115, n_341);
  xor g752 (n_348, n_1129, n_342);
  nand g753 (n_1130, n_115, n_341);
  nand g754 (n_1131, n_342, n_341);
  nand g755 (n_1132, n_115, n_342);
  nand g756 (n_360, n_1130, n_1131, n_1132);
  xor g757 (n_1133, n_343, n_344);
  xor g758 (n_349, n_1133, n_345);
  nand g759 (n_1134, n_343, n_344);
  nand g760 (n_1135, n_345, n_344);
  nand g761 (n_1136, n_343, n_345);
  nand g762 (n_362, n_1134, n_1135, n_1136);
  xor g763 (n_1137, n_346, n_347);
  xor g764 (n_351, n_1137, n_348);
  nand g765 (n_1138, n_346, n_347);
  nand g766 (n_1139, n_348, n_347);
  nand g767 (n_1140, n_346, n_348);
  nand g768 (n_364, n_1138, n_1139, n_1140);
  xor g769 (n_1141, n_349, n_350);
  xor g770 (n_163, n_1141, n_351);
  nand g771 (n_1142, n_349, n_350);
  nand g772 (n_1143, n_351, n_350);
  nand g773 (n_1144, n_349, n_351);
  nand g774 (n_95, n_1142, n_1143, n_1144);
  xor g775 (n_1145, A[20], A[18]);
  xor g776 (n_356, n_1145, A[14]);
  nand g777 (n_1146, A[20], A[18]);
  nand g778 (n_1147, A[14], A[18]);
  nand g779 (n_1148, A[20], A[14]);
  nand g780 (n_366, n_1146, n_1147, n_1148);
  xor g782 (n_357, n_251, A[12]);
  xor g787 (n_1153, A[2], A[16]);
  xor g788 (n_355, n_1153, A[10]);
  nand g789 (n_1154, A[2], A[16]);
  nand g790 (n_1155, A[10], A[16]);
  nand g792 (n_368, n_1154, n_1155, n_1034);
  xor g793 (n_1157, A[8], n_352);
  xor g794 (n_359, n_1157, n_353);
  nand g795 (n_1158, A[8], n_352);
  nand g796 (n_1159, n_353, n_352);
  nand g797 (n_1160, A[8], n_353);
  nand g798 (n_372, n_1158, n_1159, n_1160);
  xor g799 (n_1161, n_354, n_355);
  xor g800 (n_361, n_1161, n_356);
  nand g801 (n_1162, n_354, n_355);
  nand g802 (n_1163, n_356, n_355);
  nand g803 (n_1164, n_354, n_356);
  nand g804 (n_374, n_1162, n_1163, n_1164);
  xor g805 (n_1165, n_357, n_358);
  xor g806 (n_363, n_1165, n_359);
  nand g807 (n_1166, n_357, n_358);
  nand g808 (n_1167, n_359, n_358);
  nand g809 (n_1168, n_357, n_359);
  nand g810 (n_376, n_1166, n_1167, n_1168);
  xor g811 (n_1169, n_360, n_361);
  xor g812 (n_365, n_1169, n_362);
  nand g813 (n_1170, n_360, n_361);
  nand g814 (n_1171, n_362, n_361);
  nand g815 (n_1172, n_360, n_362);
  nand g816 (n_378, n_1170, n_1171, n_1172);
  xor g817 (n_1173, n_363, n_364);
  xor g818 (n_162, n_1173, n_365);
  nand g819 (n_1174, n_363, n_364);
  nand g820 (n_1175, n_365, n_364);
  nand g821 (n_1176, n_363, n_365);
  nand g822 (n_94, n_1174, n_1175, n_1176);
  xor g823 (n_1177, A[21], A[19]);
  xor g824 (n_370, n_1177, A[15]);
  nand g825 (n_1178, A[21], A[19]);
  nand g826 (n_1179, A[15], A[19]);
  nand g827 (n_1180, A[21], A[15]);
  nand g828 (n_380, n_1178, n_1179, n_1180);
  xor g830 (n_371, n_897, A[13]);
  xor g835 (n_1185, A[3], A[17]);
  xor g836 (n_369, n_1185, A[11]);
  nand g837 (n_1186, A[3], A[17]);
  nand g840 (n_382, n_1186, n_1060, n_1119);
  xor g841 (n_1189, A[9], n_366);
  xor g842 (n_373, n_1189, n_319);
  nand g843 (n_1190, A[9], n_366);
  nand g844 (n_1191, n_319, n_366);
  nand g845 (n_1192, A[9], n_319);
  nand g846 (n_386, n_1190, n_1191, n_1192);
  xor g847 (n_1193, n_368, n_369);
  xor g848 (n_375, n_1193, n_370);
  nand g849 (n_1194, n_368, n_369);
  nand g850 (n_1195, n_370, n_369);
  nand g851 (n_1196, n_368, n_370);
  nand g852 (n_388, n_1194, n_1195, n_1196);
  xor g853 (n_1197, n_371, n_372);
  xor g854 (n_377, n_1197, n_373);
  nand g855 (n_1198, n_371, n_372);
  nand g856 (n_1199, n_373, n_372);
  nand g857 (n_1200, n_371, n_373);
  nand g858 (n_390, n_1198, n_1199, n_1200);
  xor g859 (n_1201, n_374, n_375);
  xor g860 (n_379, n_1201, n_376);
  nand g861 (n_1202, n_374, n_375);
  nand g862 (n_1203, n_376, n_375);
  nand g863 (n_1204, n_374, n_376);
  nand g864 (n_393, n_1202, n_1203, n_1204);
  xor g865 (n_1205, n_377, n_378);
  xor g866 (n_161, n_1205, n_379);
  nand g867 (n_1206, n_377, n_378);
  nand g868 (n_1207, n_379, n_378);
  nand g869 (n_1208, n_377, n_379);
  nand g870 (n_93, n_1206, n_1207, n_1208);
  xor g871 (n_1209, A[22], A[20]);
  xor g872 (n_384, n_1209, A[16]);
  nand g873 (n_1210, A[22], A[20]);
  nand g874 (n_1211, A[16], A[20]);
  nand g875 (n_1212, A[22], A[16]);
  nand g876 (n_394, n_1210, n_1211, n_1212);
  xor g878 (n_385, n_254, A[14]);
  nand g880 (n_1215, A[14], A[6]);
  xor g883 (n_1217, A[4], A[18]);
  xor g884 (n_383, n_1217, A[12]);
  nand g885 (n_1218, A[4], A[18]);
  nand g886 (n_1219, A[12], A[18]);
  nand g888 (n_396, n_1218, n_1219, n_1040);
  xor g889 (n_1221, A[10], n_380);
  xor g890 (n_387, n_1221, n_332);
  nand g891 (n_1222, A[10], n_380);
  nand g892 (n_1223, n_332, n_380);
  nand g893 (n_1224, A[10], n_332);
  nand g894 (n_179, n_1222, n_1223, n_1224);
  xor g895 (n_1225, n_382, n_383);
  xor g896 (n_389, n_1225, n_384);
  nand g897 (n_1226, n_382, n_383);
  nand g898 (n_1227, n_384, n_383);
  nand g899 (n_1228, n_382, n_384);
  nand g900 (n_400, n_1226, n_1227, n_1228);
  xor g901 (n_1229, n_385, n_386);
  xor g902 (n_391, n_1229, n_387);
  nand g903 (n_1230, n_385, n_386);
  nand g904 (n_1231, n_387, n_386);
  nand g905 (n_1232, n_385, n_387);
  nand g906 (n_402, n_1230, n_1231, n_1232);
  xor g907 (n_1233, n_388, n_389);
  xor g908 (n_392, n_1233, n_390);
  nand g909 (n_1234, n_388, n_389);
  nand g910 (n_1235, n_390, n_389);
  nand g911 (n_1236, n_388, n_390);
  nand g912 (n_405, n_1234, n_1235, n_1236);
  xor g913 (n_1237, n_391, n_392);
  xor g914 (n_160, n_1237, n_393);
  nand g915 (n_1238, n_391, n_392);
  nand g916 (n_1239, n_393, n_392);
  nand g917 (n_1240, n_391, n_393);
  nand g918 (n_92, n_1238, n_1239, n_1240);
  xor g919 (n_1241, A[23], A[21]);
  xor g920 (n_398, n_1241, A[17]);
  nand g921 (n_1242, A[23], A[21]);
  nand g922 (n_1243, A[17], A[21]);
  nand g923 (n_1244, A[23], A[17]);
  nand g924 (n_406, n_1242, n_1243, n_1244);
  xor g926 (n_399, n_913, A[15]);
  nand g928 (n_1247, A[15], A[7]);
  nand g930 (n_407, n_914, n_1247, n_1012);
  xor g931 (n_1249, A[5], A[19]);
  xor g932 (n_397, n_1249, A[13]);
  nand g933 (n_1250, A[5], A[19]);
  nand g936 (n_408, n_1250, n_1116, n_1068);
  xor g937 (n_1253, A[11], n_394);
  xor g938 (n_180, n_1253, n_395);
  nand g939 (n_1254, A[11], n_394);
  nand g940 (n_1255, n_395, n_394);
  nand g941 (n_1256, A[11], n_395);
  nand g942 (n_412, n_1254, n_1255, n_1256);
  xor g943 (n_1257, n_396, n_397);
  xor g944 (n_401, n_1257, n_398);
  nand g945 (n_1258, n_396, n_397);
  nand g946 (n_1259, n_398, n_397);
  nand g947 (n_1260, n_396, n_398);
  nand g948 (n_414, n_1258, n_1259, n_1260);
  xor g949 (n_1261, n_399, n_179);
  xor g950 (n_403, n_1261, n_180);
  nand g951 (n_1262, n_399, n_179);
  nand g952 (n_1263, n_180, n_179);
  nand g953 (n_1264, n_399, n_180);
  nand g954 (n_416, n_1262, n_1263, n_1264);
  xor g955 (n_1265, n_400, n_401);
  xor g956 (n_404, n_1265, n_402);
  nand g957 (n_1266, n_400, n_401);
  nand g958 (n_1267, n_402, n_401);
  nand g959 (n_1268, n_400, n_402);
  nand g960 (n_419, n_1266, n_1267, n_1268);
  xor g961 (n_1269, n_403, n_404);
  xor g962 (n_159, n_1269, n_405);
  nand g963 (n_1270, n_403, n_404);
  nand g964 (n_1271, n_405, n_404);
  nand g965 (n_1272, n_403, n_405);
  nand g966 (n_91, n_1270, n_1271, n_1272);
  xor g967 (n_1273, A[24], A[22]);
  xor g968 (n_410, n_1273, A[18]);
  nand g969 (n_1274, A[24], A[22]);
  nand g970 (n_1275, A[18], A[22]);
  nand g971 (n_1276, A[24], A[18]);
  nand g972 (n_420, n_1274, n_1275, n_1276);
  xor g974 (n_411, n_261, A[16]);
  nand g976 (n_1279, A[16], A[8]);
  xor g979 (n_1281, A[6], A[20]);
  xor g980 (n_409, n_1281, A[14]);
  nand g981 (n_1282, A[6], A[20]);
  nand g984 (n_422, n_1282, n_1148, n_1215);
  xor g985 (n_1285, A[12], n_406);
  xor g986 (n_413, n_1285, n_407);
  nand g987 (n_1286, A[12], n_406);
  nand g988 (n_1287, n_407, n_406);
  nand g989 (n_1288, A[12], n_407);
  nand g990 (n_426, n_1286, n_1287, n_1288);
  xor g991 (n_1289, n_408, n_409);
  xor g992 (n_415, n_1289, n_410);
  nand g993 (n_1290, n_408, n_409);
  nand g994 (n_1291, n_410, n_409);
  nand g995 (n_1292, n_408, n_410);
  nand g996 (n_428, n_1290, n_1291, n_1292);
  xor g997 (n_1293, n_411, n_412);
  xor g998 (n_417, n_1293, n_413);
  nand g999 (n_1294, n_411, n_412);
  nand g1000 (n_1295, n_413, n_412);
  nand g1001 (n_1296, n_411, n_413);
  nand g1002 (n_430, n_1294, n_1295, n_1296);
  xor g1003 (n_1297, n_414, n_415);
  xor g1004 (n_418, n_1297, n_416);
  nand g1005 (n_1298, n_414, n_415);
  nand g1006 (n_1299, n_416, n_415);
  nand g1007 (n_1300, n_414, n_416);
  nand g1008 (n_433, n_1298, n_1299, n_1300);
  xor g1009 (n_1301, n_417, n_418);
  xor g1010 (n_158, n_1301, n_419);
  nand g1011 (n_1302, n_417, n_418);
  nand g1012 (n_1303, n_419, n_418);
  nand g1013 (n_1304, n_417, n_419);
  nand g1014 (n_90, n_1302, n_1303, n_1304);
  xor g1015 (n_1305, A[25], A[23]);
  xor g1016 (n_424, n_1305, A[19]);
  nand g1017 (n_1306, A[25], A[23]);
  nand g1018 (n_1307, A[19], A[23]);
  nand g1019 (n_1308, A[25], A[19]);
  nand g1020 (n_434, n_1306, n_1307, n_1308);
  xor g1022 (n_425, n_937, A[17]);
  nand g1024 (n_1311, A[17], A[9]);
  nand g1026 (n_435, n_938, n_1311, n_1060);
  xor g1027 (n_1313, A[7], A[21]);
  xor g1028 (n_423, n_1313, A[15]);
  nand g1029 (n_1314, A[7], A[21]);
  nand g1032 (n_436, n_1314, n_1180, n_1247);
  xor g1033 (n_1317, A[13], n_420);
  xor g1034 (n_427, n_1317, n_421);
  nand g1035 (n_1318, A[13], n_420);
  nand g1036 (n_1319, n_421, n_420);
  nand g1037 (n_1320, A[13], n_421);
  nand g1038 (n_440, n_1318, n_1319, n_1320);
  xor g1039 (n_1321, n_422, n_423);
  xor g1040 (n_429, n_1321, n_424);
  nand g1041 (n_1322, n_422, n_423);
  nand g1042 (n_1323, n_424, n_423);
  nand g1043 (n_1324, n_422, n_424);
  nand g1044 (n_442, n_1322, n_1323, n_1324);
  xor g1045 (n_1325, n_425, n_426);
  xor g1046 (n_431, n_1325, n_427);
  nand g1047 (n_1326, n_425, n_426);
  nand g1048 (n_1327, n_427, n_426);
  nand g1049 (n_1328, n_425, n_427);
  nand g1050 (n_444, n_1326, n_1327, n_1328);
  xor g1051 (n_1329, n_428, n_429);
  xor g1052 (n_432, n_1329, n_430);
  nand g1053 (n_1330, n_428, n_429);
  nand g1054 (n_1331, n_430, n_429);
  nand g1055 (n_1332, n_428, n_430);
  nand g1056 (n_447, n_1330, n_1331, n_1332);
  xor g1057 (n_1333, n_431, n_432);
  xor g1058 (n_157, n_1333, n_433);
  nand g1059 (n_1334, n_431, n_432);
  nand g1060 (n_1335, n_433, n_432);
  nand g1061 (n_1336, n_431, n_433);
  nand g1062 (n_89, n_1334, n_1335, n_1336);
  xor g1063 (n_1337, A[26], A[24]);
  xor g1064 (n_438, n_1337, A[20]);
  nand g1065 (n_1338, A[26], A[24]);
  nand g1066 (n_1339, A[20], A[24]);
  nand g1067 (n_1340, A[26], A[20]);
  nand g1068 (n_448, n_1338, n_1339, n_1340);
  xor g1070 (n_439, n_272, A[18]);
  nand g1072 (n_1343, A[18], A[10]);
  xor g1075 (n_1345, A[8], A[22]);
  xor g1076 (n_437, n_1345, A[16]);
  nand g1077 (n_1346, A[8], A[22]);
  nand g1080 (n_450, n_1346, n_1212, n_1279);
  xor g1081 (n_1349, A[14], n_434);
  xor g1082 (n_441, n_1349, n_435);
  nand g1083 (n_1350, A[14], n_434);
  nand g1084 (n_1351, n_435, n_434);
  nand g1085 (n_1352, A[14], n_435);
  nand g1086 (n_454, n_1350, n_1351, n_1352);
  xor g1087 (n_1353, n_436, n_437);
  xor g1088 (n_443, n_1353, n_438);
  nand g1089 (n_1354, n_436, n_437);
  nand g1090 (n_1355, n_438, n_437);
  nand g1091 (n_1356, n_436, n_438);
  nand g1092 (n_456, n_1354, n_1355, n_1356);
  xor g1093 (n_1357, n_439, n_440);
  xor g1094 (n_445, n_1357, n_441);
  nand g1095 (n_1358, n_439, n_440);
  nand g1096 (n_1359, n_441, n_440);
  nand g1097 (n_1360, n_439, n_441);
  nand g1098 (n_458, n_1358, n_1359, n_1360);
  xor g1099 (n_1361, n_442, n_443);
  xor g1100 (n_446, n_1361, n_444);
  nand g1101 (n_1362, n_442, n_443);
  nand g1102 (n_1363, n_444, n_443);
  nand g1103 (n_1364, n_442, n_444);
  nand g1104 (n_461, n_1362, n_1363, n_1364);
  xor g1105 (n_1365, n_445, n_446);
  xor g1106 (n_156, n_1365, n_447);
  nand g1107 (n_1366, n_445, n_446);
  nand g1108 (n_1367, n_447, n_446);
  nand g1109 (n_1368, n_445, n_447);
  nand g1110 (n_88, n_1366, n_1367, n_1368);
  xor g1111 (n_1369, A[27], A[25]);
  xor g1112 (n_452, n_1369, A[21]);
  nand g1113 (n_1370, A[27], A[25]);
  nand g1114 (n_1371, A[21], A[25]);
  nand g1115 (n_1372, A[27], A[21]);
  nand g1116 (n_462, n_1370, n_1371, n_1372);
  xor g1118 (n_453, n_969, A[19]);
  nand g1120 (n_1375, A[19], A[11]);
  nand g1122 (n_463, n_970, n_1375, n_1116);
  xor g1123 (n_1377, A[9], A[23]);
  xor g1124 (n_451, n_1377, A[17]);
  nand g1125 (n_1378, A[9], A[23]);
  nand g1128 (n_464, n_1378, n_1244, n_1311);
  xor g1129 (n_1381, A[15], n_448);
  xor g1130 (n_455, n_1381, n_449);
  nand g1131 (n_1382, A[15], n_448);
  nand g1132 (n_1383, n_449, n_448);
  nand g1133 (n_1384, A[15], n_449);
  nand g1134 (n_468, n_1382, n_1383, n_1384);
  xor g1135 (n_1385, n_450, n_451);
  xor g1136 (n_457, n_1385, n_452);
  nand g1137 (n_1386, n_450, n_451);
  nand g1138 (n_1387, n_452, n_451);
  nand g1139 (n_1388, n_450, n_452);
  nand g1140 (n_470, n_1386, n_1387, n_1388);
  xor g1141 (n_1389, n_453, n_454);
  xor g1142 (n_459, n_1389, n_455);
  nand g1143 (n_1390, n_453, n_454);
  nand g1144 (n_1391, n_455, n_454);
  nand g1145 (n_1392, n_453, n_455);
  nand g1146 (n_472, n_1390, n_1391, n_1392);
  xor g1147 (n_1393, n_456, n_457);
  xor g1148 (n_460, n_1393, n_458);
  nand g1149 (n_1394, n_456, n_457);
  nand g1150 (n_1395, n_458, n_457);
  nand g1151 (n_1396, n_456, n_458);
  nand g1152 (n_475, n_1394, n_1395, n_1396);
  xor g1153 (n_1397, n_459, n_460);
  xor g1154 (n_155, n_1397, n_461);
  nand g1155 (n_1398, n_459, n_460);
  nand g1156 (n_1399, n_461, n_460);
  nand g1157 (n_1400, n_459, n_461);
  nand g1158 (n_87, n_1398, n_1399, n_1400);
  xor g1159 (n_1401, A[28], A[26]);
  xor g1160 (n_466, n_1401, A[22]);
  nand g1161 (n_1402, A[28], A[26]);
  nand g1162 (n_1403, A[22], A[26]);
  nand g1163 (n_1404, A[28], A[22]);
  nand g1164 (n_476, n_1402, n_1403, n_1404);
  xor g1166 (n_467, n_287, A[20]);
  nand g1168 (n_1407, A[20], A[12]);
  xor g1171 (n_1409, A[10], A[24]);
  xor g1172 (n_465, n_1409, A[18]);
  nand g1173 (n_1410, A[10], A[24]);
  nand g1176 (n_478, n_1410, n_1276, n_1343);
  xor g1177 (n_1413, A[16], n_462);
  xor g1178 (n_469, n_1413, n_463);
  nand g1179 (n_1414, A[16], n_462);
  nand g1180 (n_1415, n_463, n_462);
  nand g1181 (n_1416, A[16], n_463);
  nand g1182 (n_482, n_1414, n_1415, n_1416);
  xor g1183 (n_1417, n_464, n_465);
  xor g1184 (n_471, n_1417, n_466);
  nand g1185 (n_1418, n_464, n_465);
  nand g1186 (n_1419, n_466, n_465);
  nand g1187 (n_1420, n_464, n_466);
  nand g1188 (n_484, n_1418, n_1419, n_1420);
  xor g1189 (n_1421, n_467, n_468);
  xor g1190 (n_473, n_1421, n_469);
  nand g1191 (n_1422, n_467, n_468);
  nand g1192 (n_1423, n_469, n_468);
  nand g1193 (n_1424, n_467, n_469);
  nand g1194 (n_486, n_1422, n_1423, n_1424);
  xor g1195 (n_1425, n_470, n_471);
  xor g1196 (n_474, n_1425, n_472);
  nand g1197 (n_1426, n_470, n_471);
  nand g1198 (n_1427, n_472, n_471);
  nand g1199 (n_1428, n_470, n_472);
  nand g1200 (n_489, n_1426, n_1427, n_1428);
  xor g1201 (n_1429, n_473, n_474);
  xor g1202 (n_154, n_1429, n_475);
  nand g1203 (n_1430, n_473, n_474);
  nand g1204 (n_1431, n_475, n_474);
  nand g1205 (n_1432, n_473, n_475);
  nand g1206 (n_86, n_1430, n_1431, n_1432);
  xor g1207 (n_1433, A[29], A[27]);
  xor g1208 (n_480, n_1433, A[23]);
  nand g1209 (n_1434, A[29], A[27]);
  nand g1210 (n_1435, A[23], A[27]);
  nand g1211 (n_1436, A[29], A[23]);
  nand g1212 (n_490, n_1434, n_1435, n_1436);
  xor g1214 (n_481, n_1009, A[21]);
  nand g1216 (n_1439, A[21], A[13]);
  nand g1218 (n_491, n_1010, n_1439, n_1180);
  xor g1219 (n_1441, A[11], A[25]);
  xor g1220 (n_479, n_1441, A[19]);
  nand g1221 (n_1442, A[11], A[25]);
  nand g1224 (n_492, n_1442, n_1308, n_1375);
  xor g1225 (n_1445, A[17], n_476);
  xor g1226 (n_483, n_1445, n_477);
  nand g1227 (n_1446, A[17], n_476);
  nand g1228 (n_1447, n_477, n_476);
  nand g1229 (n_1448, A[17], n_477);
  nand g1230 (n_496, n_1446, n_1447, n_1448);
  xor g1231 (n_1449, n_478, n_479);
  xor g1232 (n_485, n_1449, n_480);
  nand g1233 (n_1450, n_478, n_479);
  nand g1234 (n_1451, n_480, n_479);
  nand g1235 (n_1452, n_478, n_480);
  nand g1236 (n_498, n_1450, n_1451, n_1452);
  xor g1237 (n_1453, n_481, n_482);
  xor g1238 (n_487, n_1453, n_483);
  nand g1239 (n_1454, n_481, n_482);
  nand g1240 (n_1455, n_483, n_482);
  nand g1241 (n_1456, n_481, n_483);
  nand g1242 (n_500, n_1454, n_1455, n_1456);
  xor g1243 (n_1457, n_484, n_485);
  xor g1244 (n_488, n_1457, n_486);
  nand g1245 (n_1458, n_484, n_485);
  nand g1246 (n_1459, n_486, n_485);
  nand g1247 (n_1460, n_484, n_486);
  nand g1248 (n_503, n_1458, n_1459, n_1460);
  xor g1249 (n_1461, n_487, n_488);
  xor g1250 (n_153, n_1461, n_489);
  nand g1251 (n_1462, n_487, n_488);
  nand g1252 (n_1463, n_489, n_488);
  nand g1253 (n_1464, n_487, n_489);
  nand g1254 (n_85, n_1462, n_1463, n_1464);
  xor g1255 (n_1465, A[30], A[28]);
  xor g1256 (n_494, n_1465, A[24]);
  nand g1257 (n_1466, A[30], A[28]);
  nand g1258 (n_1467, A[24], A[28]);
  nand g1259 (n_1468, A[30], A[24]);
  nand g1260 (n_504, n_1466, n_1467, n_1468);
  xor g1262 (n_495, n_306, A[22]);
  nand g1264 (n_1471, A[22], A[14]);
  xor g1267 (n_1473, A[12], A[26]);
  xor g1268 (n_493, n_1473, A[20]);
  nand g1269 (n_1474, A[12], A[26]);
  nand g1272 (n_506, n_1474, n_1340, n_1407);
  xor g1273 (n_1477, A[18], n_490);
  xor g1274 (n_497, n_1477, n_491);
  nand g1275 (n_1478, A[18], n_490);
  nand g1276 (n_1479, n_491, n_490);
  nand g1277 (n_1480, A[18], n_491);
  nand g1278 (n_510, n_1478, n_1479, n_1480);
  xor g1279 (n_1481, n_492, n_493);
  xor g1280 (n_499, n_1481, n_494);
  nand g1281 (n_1482, n_492, n_493);
  nand g1282 (n_1483, n_494, n_493);
  nand g1283 (n_1484, n_492, n_494);
  nand g1284 (n_512, n_1482, n_1483, n_1484);
  xor g1285 (n_1485, n_495, n_496);
  xor g1286 (n_501, n_1485, n_497);
  nand g1287 (n_1486, n_495, n_496);
  nand g1288 (n_1487, n_497, n_496);
  nand g1289 (n_1488, n_495, n_497);
  nand g1290 (n_514, n_1486, n_1487, n_1488);
  xor g1291 (n_1489, n_498, n_499);
  xor g1292 (n_502, n_1489, n_500);
  nand g1293 (n_1490, n_498, n_499);
  nand g1294 (n_1491, n_500, n_499);
  nand g1295 (n_1492, n_498, n_500);
  nand g1296 (n_517, n_1490, n_1491, n_1492);
  xor g1297 (n_1493, n_501, n_502);
  xor g1298 (n_152, n_1493, n_503);
  nand g1299 (n_1494, n_501, n_502);
  nand g1300 (n_1495, n_503, n_502);
  nand g1301 (n_1496, n_501, n_503);
  nand g1302 (n_84, n_1494, n_1495, n_1496);
  xor g1303 (n_1497, A[31], A[29]);
  xor g1304 (n_508, n_1497, A[25]);
  nand g1305 (n_1498, A[31], A[29]);
  nand g1306 (n_1499, A[25], A[29]);
  nand g1307 (n_1500, A[31], A[25]);
  nand g1308 (n_518, n_1498, n_1499, n_1500);
  xor g1310 (n_509, n_1057, A[23]);
  nand g1312 (n_1503, A[23], A[15]);
  nand g1314 (n_519, n_1058, n_1503, n_1244);
  xor g1315 (n_1505, A[13], A[27]);
  xor g1316 (n_507, n_1505, A[21]);
  nand g1317 (n_1506, A[13], A[27]);
  nand g1320 (n_520, n_1506, n_1372, n_1439);
  xor g1321 (n_1509, A[19], n_504);
  xor g1322 (n_511, n_1509, n_505);
  nand g1323 (n_1510, A[19], n_504);
  nand g1324 (n_1511, n_505, n_504);
  nand g1325 (n_1512, A[19], n_505);
  nand g1326 (n_524, n_1510, n_1511, n_1512);
  xor g1327 (n_1513, n_506, n_507);
  xor g1328 (n_513, n_1513, n_508);
  nand g1329 (n_1514, n_506, n_507);
  nand g1330 (n_1515, n_508, n_507);
  nand g1331 (n_1516, n_506, n_508);
  nand g1332 (n_526, n_1514, n_1515, n_1516);
  xor g1333 (n_1517, n_509, n_510);
  xor g1334 (n_515, n_1517, n_511);
  nand g1335 (n_1518, n_509, n_510);
  nand g1336 (n_1519, n_511, n_510);
  nand g1337 (n_1520, n_509, n_511);
  nand g1338 (n_528, n_1518, n_1519, n_1520);
  xor g1339 (n_1521, n_512, n_513);
  xor g1340 (n_516, n_1521, n_514);
  nand g1341 (n_1522, n_512, n_513);
  nand g1342 (n_1523, n_514, n_513);
  nand g1343 (n_1524, n_512, n_514);
  nand g1344 (n_531, n_1522, n_1523, n_1524);
  xor g1345 (n_1525, n_515, n_516);
  xor g1346 (n_151, n_1525, n_517);
  nand g1347 (n_1526, n_515, n_516);
  nand g1348 (n_1527, n_517, n_516);
  nand g1349 (n_1528, n_515, n_517);
  nand g1350 (n_83, n_1526, n_1527, n_1528);
  xor g1351 (n_1529, A[32], A[30]);
  xor g1352 (n_522, n_1529, A[26]);
  nand g1353 (n_1530, A[32], A[30]);
  nand g1354 (n_1531, A[26], A[30]);
  nand g1355 (n_1532, A[32], A[26]);
  nand g1356 (n_532, n_1530, n_1531, n_1532);
  xor g1358 (n_523, n_329, A[24]);
  nand g1360 (n_1535, A[24], A[16]);
  xor g1363 (n_1537, A[14], A[28]);
  xor g1364 (n_521, n_1537, A[22]);
  nand g1365 (n_1538, A[14], A[28]);
  nand g1368 (n_534, n_1538, n_1404, n_1471);
  xor g1369 (n_1541, A[20], n_518);
  xor g1370 (n_525, n_1541, n_519);
  nand g1371 (n_1542, A[20], n_518);
  nand g1372 (n_1543, n_519, n_518);
  nand g1373 (n_1544, A[20], n_519);
  nand g1374 (n_538, n_1542, n_1543, n_1544);
  xor g1375 (n_1545, n_520, n_521);
  xor g1376 (n_527, n_1545, n_522);
  nand g1377 (n_1546, n_520, n_521);
  nand g1378 (n_1547, n_522, n_521);
  nand g1379 (n_1548, n_520, n_522);
  nand g1380 (n_540, n_1546, n_1547, n_1548);
  xor g1381 (n_1549, n_523, n_524);
  xor g1382 (n_529, n_1549, n_525);
  nand g1383 (n_1550, n_523, n_524);
  nand g1384 (n_1551, n_525, n_524);
  nand g1385 (n_1552, n_523, n_525);
  nand g1386 (n_542, n_1550, n_1551, n_1552);
  xor g1387 (n_1553, n_526, n_527);
  xor g1388 (n_530, n_1553, n_528);
  nand g1389 (n_1554, n_526, n_527);
  nand g1390 (n_1555, n_528, n_527);
  nand g1391 (n_1556, n_526, n_528);
  nand g1392 (n_545, n_1554, n_1555, n_1556);
  xor g1393 (n_1557, n_529, n_530);
  xor g1394 (n_150, n_1557, n_531);
  nand g1395 (n_1558, n_529, n_530);
  nand g1396 (n_1559, n_531, n_530);
  nand g1397 (n_1560, n_529, n_531);
  nand g1398 (n_82, n_1558, n_1559, n_1560);
  xor g1399 (n_1561, A[33], A[31]);
  xor g1400 (n_536, n_1561, A[27]);
  nand g1401 (n_1562, A[33], A[31]);
  nand g1402 (n_1563, A[27], A[31]);
  nand g1403 (n_1564, A[33], A[27]);
  nand g1404 (n_546, n_1562, n_1563, n_1564);
  xor g1406 (n_537, n_1113, A[25]);
  nand g1408 (n_1567, A[25], A[17]);
  nand g1410 (n_548, n_1114, n_1567, n_1308);
  xor g1411 (n_1569, A[15], A[29]);
  xor g1412 (n_535, n_1569, A[23]);
  nand g1413 (n_1570, A[15], A[29]);
  nand g1416 (n_547, n_1570, n_1436, n_1503);
  xor g1417 (n_1573, A[21], n_532);
  xor g1418 (n_539, n_1573, n_533);
  nand g1419 (n_1574, A[21], n_532);
  nand g1420 (n_1575, n_533, n_532);
  nand g1421 (n_1576, A[21], n_533);
  nand g1422 (n_552, n_1574, n_1575, n_1576);
  xor g1423 (n_1577, n_534, n_535);
  xor g1424 (n_541, n_1577, n_536);
  nand g1425 (n_1578, n_534, n_535);
  nand g1426 (n_1579, n_536, n_535);
  nand g1427 (n_1580, n_534, n_536);
  nand g1428 (n_554, n_1578, n_1579, n_1580);
  xor g1429 (n_1581, n_537, n_538);
  xor g1430 (n_543, n_1581, n_539);
  nand g1431 (n_1582, n_537, n_538);
  nand g1432 (n_1583, n_539, n_538);
  nand g1433 (n_1584, n_537, n_539);
  nand g1434 (n_557, n_1582, n_1583, n_1584);
  xor g1435 (n_1585, n_540, n_541);
  xor g1436 (n_544, n_1585, n_542);
  nand g1437 (n_1586, n_540, n_541);
  nand g1438 (n_1587, n_542, n_541);
  nand g1439 (n_1588, n_540, n_542);
  nand g1440 (n_559, n_1586, n_1587, n_1588);
  xor g1441 (n_1589, n_543, n_544);
  xor g1442 (n_149, n_1589, n_545);
  nand g1443 (n_1590, n_543, n_544);
  nand g1444 (n_1591, n_545, n_544);
  nand g1445 (n_1592, n_543, n_545);
  nand g1446 (n_81, n_1590, n_1591, n_1592);
  xor g1447 (n_1593, A[32], A[28]);
  xor g1448 (n_550, n_1593, A[20]);
  nand g1449 (n_1594, A[32], A[28]);
  nand g1450 (n_1595, A[20], A[28]);
  nand g1451 (n_1596, A[32], A[20]);
  nand g1452 (n_560, n_1594, n_1595, n_1596);
  xor g1453 (n_1597, A[18], A[26]);
  xor g1454 (n_551, n_1597, A[16]);
  nand g1455 (n_1598, A[18], A[26]);
  nand g1456 (n_1599, A[16], A[26]);
  xor g1459 (n_1601, A[30], A[24]);
  xor g1460 (n_549, n_1601, A[22]);
  nand g1463 (n_1604, A[30], A[22]);
  nand g1464 (n_561, n_1468, n_1274, n_1604);
  xor g1465 (n_1605, A[34], n_546);
  xor g1466 (n_553, n_1605, n_547);
  nand g1467 (n_1606, A[34], n_546);
  nand g1468 (n_1607, n_547, n_546);
  nand g1469 (n_1608, A[34], n_547);
  nand g1470 (n_566, n_1606, n_1607, n_1608);
  xor g1471 (n_1609, n_548, n_549);
  xor g1472 (n_555, n_1609, n_550);
  nand g1473 (n_1610, n_548, n_549);
  nand g1474 (n_1611, n_550, n_549);
  nand g1475 (n_1612, n_548, n_550);
  nand g1476 (n_568, n_1610, n_1611, n_1612);
  xor g1477 (n_1613, n_551, n_552);
  xor g1478 (n_556, n_1613, n_553);
  nand g1479 (n_1614, n_551, n_552);
  nand g1480 (n_1615, n_553, n_552);
  nand g1481 (n_1616, n_551, n_553);
  nand g1482 (n_571, n_1614, n_1615, n_1616);
  xor g1483 (n_1617, n_554, n_555);
  xor g1484 (n_558, n_1617, n_556);
  nand g1485 (n_1618, n_554, n_555);
  nand g1486 (n_1619, n_556, n_555);
  nand g1487 (n_1620, n_554, n_556);
  nand g1488 (n_573, n_1618, n_1619, n_1620);
  xor g1489 (n_1621, n_557, n_558);
  xor g1490 (n_148, n_1621, n_559);
  nand g1491 (n_1622, n_557, n_558);
  nand g1492 (n_1623, n_559, n_558);
  nand g1493 (n_1624, n_557, n_559);
  nand g1494 (n_80, n_1622, n_1623, n_1624);
  xor g1495 (n_1625, A[33], A[29]);
  xor g1496 (n_564, n_1625, A[21]);
  nand g1497 (n_1626, A[33], A[29]);
  nand g1498 (n_1627, A[21], A[29]);
  nand g1499 (n_1628, A[33], A[21]);
  nand g1500 (n_575, n_1626, n_1627, n_1628);
  xor g1501 (n_1629, A[19], A[27]);
  xor g1502 (n_565, n_1629, A[17]);
  nand g1503 (n_1630, A[19], A[27]);
  nand g1504 (n_1631, A[17], A[27]);
  nand g1506 (n_576, n_1630, n_1631, n_1114);
  xor g1507 (n_1633, A[31], A[25]);
  xor g1508 (n_563, n_1633, A[23]);
  nand g1511 (n_1636, A[31], A[23]);
  nand g1512 (n_574, n_1500, n_1306, n_1636);
  xor g1513 (n_1637, A[35], n_560);
  xor g1514 (n_567, n_1637, n_561);
  nand g1515 (n_1638, A[35], n_560);
  nand g1516 (n_1639, n_561, n_560);
  nand g1517 (n_1640, A[35], n_561);
  nand g1518 (n_580, n_1638, n_1639, n_1640);
  xor g1519 (n_1641, n_562, n_563);
  xor g1520 (n_569, n_1641, n_564);
  nand g1521 (n_1642, n_562, n_563);
  nand g1522 (n_1643, n_564, n_563);
  nand g1523 (n_1644, n_562, n_564);
  nand g1524 (n_581, n_1642, n_1643, n_1644);
  xor g1525 (n_1645, n_565, n_566);
  xor g1526 (n_570, n_1645, n_567);
  nand g1527 (n_1646, n_565, n_566);
  nand g1528 (n_1647, n_567, n_566);
  nand g1529 (n_1648, n_565, n_567);
  nand g1530 (n_585, n_1646, n_1647, n_1648);
  xor g1531 (n_1649, n_568, n_569);
  xor g1532 (n_572, n_1649, n_570);
  nand g1533 (n_1650, n_568, n_569);
  nand g1534 (n_1651, n_570, n_569);
  nand g1535 (n_1652, n_568, n_570);
  nand g1536 (n_587, n_1650, n_1651, n_1652);
  xor g1537 (n_1653, n_571, n_572);
  xor g1538 (n_147, n_1653, n_573);
  nand g1539 (n_1654, n_571, n_572);
  nand g1540 (n_1655, n_573, n_572);
  nand g1541 (n_1656, n_571, n_573);
  nand g1542 (n_79, n_1654, n_1655, n_1656);
  xor g1544 (n_577, n_1529, A[22]);
  nand g1547 (n_1660, A[32], A[22]);
  nand g1548 (n_588, n_1530, n_1604, n_1660);
  xor g1549 (n_1661, A[20], A[28]);
  xor g1550 (n_579, n_1661, A[18]);
  nand g1552 (n_1663, A[18], A[28]);
  nand g1554 (n_589, n_1595, n_1663, n_1146);
  xor g1556 (n_578, n_1337, A[34]);
  nand g1558 (n_1667, A[34], A[24]);
  nand g1559 (n_1668, A[26], A[34]);
  nand g1560 (n_591, n_1338, n_1667, n_1668);
  xor g1561 (n_1669, A[36], n_574);
  xor g1562 (n_582, n_1669, n_575);
  nand g1563 (n_1670, A[36], n_574);
  nand g1564 (n_1671, n_575, n_574);
  nand g1565 (n_1672, A[36], n_575);
  nand g1566 (n_594, n_1670, n_1671, n_1672);
  xor g1567 (n_1673, n_576, n_577);
  xor g1568 (n_583, n_1673, n_578);
  nand g1569 (n_1674, n_576, n_577);
  nand g1570 (n_1675, n_578, n_577);
  nand g1571 (n_1676, n_576, n_578);
  nand g1572 (n_595, n_1674, n_1675, n_1676);
  xor g1573 (n_1677, n_579, n_580);
  xor g1574 (n_584, n_1677, n_581);
  nand g1575 (n_1678, n_579, n_580);
  nand g1576 (n_1679, n_581, n_580);
  nand g1577 (n_1680, n_579, n_581);
  nand g1578 (n_599, n_1678, n_1679, n_1680);
  xor g1579 (n_1681, n_582, n_583);
  xor g1580 (n_586, n_1681, n_584);
  nand g1581 (n_1682, n_582, n_583);
  nand g1582 (n_1683, n_584, n_583);
  nand g1583 (n_1684, n_582, n_584);
  nand g1584 (n_601, n_1682, n_1683, n_1684);
  xor g1585 (n_1685, n_585, n_586);
  xor g1586 (n_146, n_1685, n_587);
  nand g1587 (n_1686, n_585, n_586);
  nand g1588 (n_1687, n_587, n_586);
  nand g1589 (n_1688, n_585, n_587);
  nand g1590 (n_78, n_1686, n_1687, n_1688);
  xor g1592 (n_590, n_1561, A[23]);
  nand g1595 (n_1692, A[33], A[23]);
  nand g1596 (n_602, n_1562, n_1636, n_1692);
  xor g1597 (n_1693, A[21], A[29]);
  xor g1598 (n_593, n_1693, A[19]);
  nand g1600 (n_1695, A[19], A[29]);
  nand g1602 (n_603, n_1627, n_1695, n_1178);
  xor g1604 (n_592, n_1369, A[35]);
  nand g1606 (n_1699, A[35], A[25]);
  nand g1607 (n_1700, A[27], A[35]);
  nand g1608 (n_605, n_1370, n_1699, n_1700);
  xor g1609 (n_1701, A[37], n_588);
  xor g1610 (n_596, n_1701, n_589);
  nand g1611 (n_1702, A[37], n_588);
  nand g1612 (n_1703, n_589, n_588);
  nand g1613 (n_1704, A[37], n_589);
  nand g1614 (n_608, n_1702, n_1703, n_1704);
  xor g1615 (n_1705, n_590, n_591);
  xor g1616 (n_597, n_1705, n_592);
  nand g1617 (n_1706, n_590, n_591);
  nand g1618 (n_1707, n_592, n_591);
  nand g1619 (n_1708, n_590, n_592);
  nand g1620 (n_609, n_1706, n_1707, n_1708);
  xor g1621 (n_1709, n_593, n_594);
  xor g1622 (n_598, n_1709, n_595);
  nand g1623 (n_1710, n_593, n_594);
  nand g1624 (n_1711, n_595, n_594);
  nand g1625 (n_1712, n_593, n_595);
  nand g1626 (n_613, n_1710, n_1711, n_1712);
  xor g1627 (n_1713, n_596, n_597);
  xor g1628 (n_600, n_1713, n_598);
  nand g1629 (n_1714, n_596, n_597);
  nand g1630 (n_1715, n_598, n_597);
  nand g1631 (n_1716, n_596, n_598);
  nand g1632 (n_615, n_1714, n_1715, n_1716);
  xor g1633 (n_1717, n_599, n_600);
  xor g1634 (n_145, n_1717, n_601);
  nand g1635 (n_1718, n_599, n_600);
  nand g1636 (n_1719, n_601, n_600);
  nand g1637 (n_1720, n_599, n_601);
  nand g1638 (n_77, n_1718, n_1719, n_1720);
  xor g1640 (n_604, n_1529, A[24]);
  nand g1643 (n_1724, A[32], A[24]);
  nand g1644 (n_616, n_1530, n_1468, n_1724);
  xor g1646 (n_606, n_1209, A[28]);
  nand g1650 (n_617, n_1210, n_1595, n_1404);
  xor g1651 (n_1729, A[26], A[36]);
  xor g1652 (n_607, n_1729, A[38]);
  nand g1653 (n_1730, A[26], A[36]);
  nand g1654 (n_1731, A[38], A[36]);
  nand g1655 (n_1732, A[26], A[38]);
  nand g1656 (n_619, n_1730, n_1731, n_1732);
  xor g1657 (n_1733, A[34], n_602);
  xor g1658 (n_610, n_1733, n_603);
  nand g1659 (n_1734, A[34], n_602);
  nand g1660 (n_1735, n_603, n_602);
  nand g1661 (n_1736, A[34], n_603);
  nand g1662 (n_622, n_1734, n_1735, n_1736);
  xor g1663 (n_1737, n_604, n_605);
  xor g1664 (n_611, n_1737, n_606);
  nand g1665 (n_1738, n_604, n_605);
  nand g1666 (n_1739, n_606, n_605);
  nand g1667 (n_1740, n_604, n_606);
  nand g1668 (n_623, n_1738, n_1739, n_1740);
  xor g1669 (n_1741, n_607, n_608);
  xor g1670 (n_612, n_1741, n_609);
  nand g1671 (n_1742, n_607, n_608);
  nand g1672 (n_1743, n_609, n_608);
  nand g1673 (n_1744, n_607, n_609);
  nand g1674 (n_627, n_1742, n_1743, n_1744);
  xor g1675 (n_1745, n_610, n_611);
  xor g1676 (n_614, n_1745, n_612);
  nand g1677 (n_1746, n_610, n_611);
  nand g1678 (n_1747, n_612, n_611);
  nand g1679 (n_1748, n_610, n_612);
  nand g1680 (n_629, n_1746, n_1747, n_1748);
  xor g1681 (n_1749, n_613, n_614);
  xor g1682 (n_144, n_1749, n_615);
  nand g1683 (n_1750, n_613, n_614);
  nand g1684 (n_1751, n_615, n_614);
  nand g1685 (n_1752, n_613, n_615);
  nand g1686 (n_76, n_1750, n_1751, n_1752);
  xor g1688 (n_618, n_1561, A[25]);
  nand g1691 (n_1756, A[33], A[25]);
  nand g1692 (n_630, n_1562, n_1500, n_1756);
  xor g1694 (n_620, n_1241, A[29]);
  nand g1698 (n_631, n_1242, n_1627, n_1436);
  xor g1699 (n_1761, A[27], A[37]);
  xor g1700 (n_621, n_1761, A[39]);
  nand g1701 (n_1762, A[27], A[37]);
  nand g1702 (n_1763, A[39], A[37]);
  nand g1703 (n_1764, A[27], A[39]);
  nand g1704 (n_633, n_1762, n_1763, n_1764);
  xor g1705 (n_1765, A[35], n_616);
  xor g1706 (n_624, n_1765, n_617);
  nand g1707 (n_1766, A[35], n_616);
  nand g1708 (n_1767, n_617, n_616);
  nand g1709 (n_1768, A[35], n_617);
  nand g1710 (n_636, n_1766, n_1767, n_1768);
  xor g1711 (n_1769, n_618, n_619);
  xor g1712 (n_625, n_1769, n_620);
  nand g1713 (n_1770, n_618, n_619);
  nand g1714 (n_1771, n_620, n_619);
  nand g1715 (n_1772, n_618, n_620);
  nand g1716 (n_637, n_1770, n_1771, n_1772);
  xor g1717 (n_1773, n_621, n_622);
  xor g1718 (n_626, n_1773, n_623);
  nand g1719 (n_1774, n_621, n_622);
  nand g1720 (n_1775, n_623, n_622);
  nand g1721 (n_1776, n_621, n_623);
  nand g1722 (n_641, n_1774, n_1775, n_1776);
  xor g1723 (n_1777, n_624, n_625);
  xor g1724 (n_628, n_1777, n_626);
  nand g1725 (n_1778, n_624, n_625);
  nand g1726 (n_1779, n_626, n_625);
  nand g1727 (n_1780, n_624, n_626);
  nand g1728 (n_643, n_1778, n_1779, n_1780);
  xor g1729 (n_1781, n_627, n_628);
  xor g1730 (n_143, n_1781, n_629);
  nand g1731 (n_1782, n_627, n_628);
  nand g1732 (n_1783, n_629, n_628);
  nand g1733 (n_1784, n_627, n_629);
  nand g1734 (n_75, n_1782, n_1783, n_1784);
  xor g1735 (n_1785, A[32], A[26]);
  xor g1736 (n_632, n_1785, A[24]);
  nand g1740 (n_644, n_1532, n_1338, n_1724);
  xor g1741 (n_1789, A[22], A[30]);
  xor g1742 (n_634, n_1789, A[28]);
  nand g1746 (n_645, n_1604, n_1466, n_1404);
  xor g1747 (n_1793, A[34], A[40]);
  xor g1748 (n_635, n_1793, A[38]);
  nand g1749 (n_1794, A[34], A[40]);
  nand g1750 (n_1795, A[38], A[40]);
  nand g1751 (n_1796, A[34], A[38]);
  nand g1752 (n_647, n_1794, n_1795, n_1796);
  xor g1753 (n_1797, A[36], n_630);
  xor g1754 (n_638, n_1797, n_631);
  nand g1755 (n_1798, A[36], n_630);
  nand g1756 (n_1799, n_631, n_630);
  nand g1757 (n_1800, A[36], n_631);
  nand g1758 (n_650, n_1798, n_1799, n_1800);
  xor g1759 (n_1801, n_632, n_633);
  xor g1760 (n_639, n_1801, n_634);
  nand g1761 (n_1802, n_632, n_633);
  nand g1762 (n_1803, n_634, n_633);
  nand g1763 (n_1804, n_632, n_634);
  nand g1764 (n_651, n_1802, n_1803, n_1804);
  xor g1765 (n_1805, n_635, n_636);
  xor g1766 (n_640, n_1805, n_637);
  nand g1767 (n_1806, n_635, n_636);
  nand g1768 (n_1807, n_637, n_636);
  nand g1769 (n_1808, n_635, n_637);
  nand g1770 (n_655, n_1806, n_1807, n_1808);
  xor g1771 (n_1809, n_638, n_639);
  xor g1772 (n_642, n_1809, n_640);
  nand g1773 (n_1810, n_638, n_639);
  nand g1774 (n_1811, n_640, n_639);
  nand g1775 (n_1812, n_638, n_640);
  nand g1776 (n_657, n_1810, n_1811, n_1812);
  xor g1777 (n_1813, n_641, n_642);
  xor g1778 (n_142, n_1813, n_643);
  nand g1779 (n_1814, n_641, n_642);
  nand g1780 (n_1815, n_643, n_642);
  nand g1781 (n_1816, n_641, n_643);
  nand g1782 (n_74, n_1814, n_1815, n_1816);
  xor g1783 (n_1817, A[33], A[27]);
  xor g1784 (n_646, n_1817, A[25]);
  nand g1788 (n_658, n_1564, n_1370, n_1756);
  xor g1789 (n_1821, A[23], A[31]);
  xor g1790 (n_648, n_1821, A[29]);
  nand g1794 (n_659, n_1636, n_1498, n_1436);
  xor g1795 (n_1825, A[35], A[41]);
  xor g1796 (n_649, n_1825, A[39]);
  nand g1797 (n_1826, A[35], A[41]);
  nand g1798 (n_1827, A[39], A[41]);
  nand g1799 (n_1828, A[35], A[39]);
  nand g1800 (n_662, n_1826, n_1827, n_1828);
  xor g1801 (n_1829, A[37], n_644);
  xor g1802 (n_652, n_1829, n_645);
  nand g1803 (n_1830, A[37], n_644);
  nand g1804 (n_1831, n_645, n_644);
  nand g1805 (n_1832, A[37], n_645);
  nand g1806 (n_664, n_1830, n_1831, n_1832);
  xor g1807 (n_1833, n_646, n_647);
  xor g1808 (n_653, n_1833, n_648);
  nand g1809 (n_1834, n_646, n_647);
  nand g1810 (n_1835, n_648, n_647);
  nand g1811 (n_1836, n_646, n_648);
  nand g1812 (n_665, n_1834, n_1835, n_1836);
  xor g1813 (n_1837, n_649, n_650);
  xor g1814 (n_654, n_1837, n_651);
  nand g1815 (n_1838, n_649, n_650);
  nand g1816 (n_1839, n_651, n_650);
  nand g1817 (n_1840, n_649, n_651);
  nand g1818 (n_669, n_1838, n_1839, n_1840);
  xor g1819 (n_1841, n_652, n_653);
  xor g1820 (n_656, n_1841, n_654);
  nand g1821 (n_1842, n_652, n_653);
  nand g1822 (n_1843, n_654, n_653);
  nand g1823 (n_1844, n_652, n_654);
  nand g1824 (n_671, n_1842, n_1843, n_1844);
  xor g1825 (n_1845, n_655, n_656);
  xor g1826 (n_141, n_1845, n_657);
  nand g1827 (n_1846, n_655, n_656);
  nand g1828 (n_1847, n_657, n_656);
  nand g1829 (n_1848, n_655, n_657);
  nand g1830 (n_73, n_1846, n_1847, n_1848);
  xor g1832 (n_660, n_1593, A[26]);
  nand g1836 (n_672, n_1594, n_1402, n_1532);
  xor g1838 (n_661, n_1601, A[36]);
  nand g1840 (n_1855, A[36], A[30]);
  nand g1841 (n_1856, A[24], A[36]);
  nand g1842 (n_675, n_1468, n_1855, n_1856);
  xor g1849 (n_1861, A[42], n_658);
  xor g1850 (n_666, n_1861, n_659);
  nand g1851 (n_1862, A[42], n_658);
  nand g1852 (n_1863, n_659, n_658);
  nand g1853 (n_1864, A[42], n_659);
  nand g1854 (n_678, n_1862, n_1863, n_1864);
  xor g1855 (n_1865, n_660, n_661);
  xor g1856 (n_667, n_1865, n_662);
  nand g1857 (n_1866, n_660, n_661);
  nand g1858 (n_1867, n_662, n_661);
  nand g1859 (n_1868, n_660, n_662);
  nand g1860 (n_679, n_1866, n_1867, n_1868);
  xor g1861 (n_1869, n_635, n_664);
  xor g1862 (n_668, n_1869, n_665);
  nand g1863 (n_1870, n_635, n_664);
  nand g1864 (n_1871, n_665, n_664);
  nand g1865 (n_1872, n_635, n_665);
  nand g1866 (n_683, n_1870, n_1871, n_1872);
  xor g1867 (n_1873, n_666, n_667);
  xor g1868 (n_670, n_1873, n_668);
  nand g1869 (n_1874, n_666, n_667);
  nand g1870 (n_1875, n_668, n_667);
  nand g1871 (n_1876, n_666, n_668);
  nand g1872 (n_685, n_1874, n_1875, n_1876);
  xor g1873 (n_1877, n_669, n_670);
  xor g1874 (n_140, n_1877, n_671);
  nand g1875 (n_1878, n_669, n_670);
  nand g1876 (n_1879, n_671, n_670);
  nand g1877 (n_1880, n_669, n_671);
  nand g1878 (n_72, n_1878, n_1879, n_1880);
  xor g1880 (n_673, n_1625, A[27]);
  nand g1884 (n_686, n_1626, n_1434, n_1564);
  xor g1886 (n_674, n_1633, A[37]);
  nand g1888 (n_1887, A[37], A[31]);
  nand g1889 (n_1888, A[25], A[37]);
  nand g1890 (n_688, n_1500, n_1887, n_1888);
  xor g1897 (n_1893, A[43], n_672);
  xor g1898 (n_680, n_1893, n_673);
  nand g1899 (n_1894, A[43], n_672);
  nand g1900 (n_1895, n_673, n_672);
  nand g1901 (n_1896, A[43], n_673);
  nand g1902 (n_693, n_1894, n_1895, n_1896);
  xor g1903 (n_1897, n_674, n_675);
  xor g1904 (n_681, n_1897, n_647);
  nand g1905 (n_1898, n_674, n_675);
  nand g1906 (n_1899, n_647, n_675);
  nand g1907 (n_1900, n_674, n_647);
  nand g1908 (n_692, n_1898, n_1899, n_1900);
  xor g1909 (n_1901, n_649, n_678);
  xor g1910 (n_682, n_1901, n_679);
  nand g1911 (n_1902, n_649, n_678);
  nand g1912 (n_1903, n_679, n_678);
  nand g1913 (n_1904, n_649, n_679);
  nand g1914 (n_696, n_1902, n_1903, n_1904);
  xor g1915 (n_1905, n_680, n_681);
  xor g1916 (n_684, n_1905, n_682);
  nand g1917 (n_1906, n_680, n_681);
  nand g1918 (n_1907, n_682, n_681);
  nand g1919 (n_1908, n_680, n_682);
  nand g1920 (n_699, n_1906, n_1907, n_1908);
  xor g1921 (n_1909, n_683, n_684);
  xor g1922 (n_139, n_1909, n_685);
  nand g1923 (n_1910, n_683, n_684);
  nand g1924 (n_1911, n_685, n_684);
  nand g1925 (n_1912, n_683, n_685);
  nand g1926 (n_71, n_1910, n_1911, n_1912);
  xor g1928 (n_687, n_1529, A[28]);
  nand g1932 (n_700, n_1530, n_1466, n_1594);
  xor g1933 (n_1917, A[26], A[38]);
  xor g1934 (n_691, n_1917, A[42]);
  nand g1936 (n_1919, A[42], A[38]);
  nand g1937 (n_1920, A[26], A[42]);
  nand g1938 (n_702, n_1732, n_1919, n_1920);
  xor g1939 (n_1921, A[36], A[44]);
  xor g1940 (n_690, n_1921, A[34]);
  nand g1941 (n_1922, A[36], A[44]);
  nand g1942 (n_1923, A[34], A[44]);
  nand g1943 (n_1924, A[36], A[34]);
  nand g1944 (n_703, n_1922, n_1923, n_1924);
  xor g1945 (n_1925, A[40], n_686);
  xor g1946 (n_694, n_1925, n_687);
  nand g1947 (n_1926, A[40], n_686);
  nand g1948 (n_1927, n_687, n_686);
  nand g1949 (n_1928, A[40], n_687);
  nand g1950 (n_706, n_1926, n_1927, n_1928);
  xor g1951 (n_1929, n_688, n_662);
  xor g1952 (n_695, n_1929, n_690);
  nand g1953 (n_1930, n_688, n_662);
  nand g1954 (n_1931, n_690, n_662);
  nand g1955 (n_1932, n_688, n_690);
  nand g1956 (n_709, n_1930, n_1931, n_1932);
  xor g1957 (n_1933, n_691, n_692);
  xor g1958 (n_697, n_1933, n_693);
  nand g1959 (n_1934, n_691, n_692);
  nand g1960 (n_1935, n_693, n_692);
  nand g1961 (n_1936, n_691, n_693);
  nand g1962 (n_710, n_1934, n_1935, n_1936);
  xor g1963 (n_1937, n_694, n_695);
  xor g1964 (n_698, n_1937, n_696);
  nand g1965 (n_1938, n_694, n_695);
  nand g1966 (n_1939, n_696, n_695);
  nand g1967 (n_1940, n_694, n_696);
  nand g1968 (n_713, n_1938, n_1939, n_1940);
  xor g1969 (n_1941, n_697, n_698);
  xor g1970 (n_138, n_1941, n_699);
  nand g1971 (n_1942, n_697, n_698);
  nand g1972 (n_1943, n_699, n_698);
  nand g1973 (n_1944, n_697, n_699);
  nand g1974 (n_70, n_1942, n_1943, n_1944);
  xor g1976 (n_701, n_1561, A[29]);
  nand g1980 (n_714, n_1562, n_1498, n_1626);
  xor g1981 (n_1949, A[27], A[39]);
  xor g1982 (n_705, n_1949, A[43]);
  nand g1984 (n_1951, A[43], A[39]);
  nand g1985 (n_1952, A[27], A[43]);
  nand g1986 (n_716, n_1764, n_1951, n_1952);
  xor g1987 (n_1953, A[37], A[45]);
  xor g1988 (n_704, n_1953, A[35]);
  nand g1989 (n_1954, A[37], A[45]);
  nand g1990 (n_1955, A[35], A[45]);
  nand g1991 (n_1956, A[37], A[35]);
  nand g1992 (n_717, n_1954, n_1955, n_1956);
  xor g1993 (n_1957, A[41], n_700);
  xor g1994 (n_707, n_1957, n_701);
  nand g1995 (n_1958, A[41], n_700);
  nand g1996 (n_1959, n_701, n_700);
  nand g1997 (n_1960, A[41], n_701);
  nand g1998 (n_720, n_1958, n_1959, n_1960);
  xor g1999 (n_1961, n_702, n_703);
  xor g2000 (n_708, n_1961, n_704);
  nand g2001 (n_1962, n_702, n_703);
  nand g2002 (n_1963, n_704, n_703);
  nand g2003 (n_1964, n_702, n_704);
  nand g2004 (n_723, n_1962, n_1963, n_1964);
  xor g2005 (n_1965, n_705, n_706);
  xor g2006 (n_711, n_1965, n_707);
  nand g2007 (n_1966, n_705, n_706);
  nand g2008 (n_1967, n_707, n_706);
  nand g2009 (n_1968, n_705, n_707);
  nand g2010 (n_724, n_1966, n_1967, n_1968);
  xor g2011 (n_1969, n_708, n_709);
  xor g2012 (n_712, n_1969, n_710);
  nand g2013 (n_1970, n_708, n_709);
  nand g2014 (n_1971, n_710, n_709);
  nand g2015 (n_1972, n_708, n_710);
  nand g2016 (n_727, n_1970, n_1971, n_1972);
  xor g2017 (n_1973, n_711, n_712);
  xor g2018 (n_137, n_1973, n_713);
  nand g2019 (n_1974, n_711, n_712);
  nand g2020 (n_1975, n_713, n_712);
  nand g2021 (n_1976, n_711, n_713);
  nand g2022 (n_69, n_1974, n_1975, n_1976);
  xor g2029 (n_1981, A[46], A[40]);
  xor g2030 (n_719, n_1981, A[44]);
  nand g2031 (n_1982, A[46], A[40]);
  nand g2032 (n_1983, A[44], A[40]);
  nand g2033 (n_1984, A[46], A[44]);
  nand g2034 (n_733, n_1982, n_1983, n_1984);
  xor g2035 (n_1985, A[38], A[42]);
  xor g2036 (n_718, n_1985, A[36]);
  nand g2038 (n_1987, A[36], A[42]);
  nand g2040 (n_731, n_1919, n_1987, n_1731);
  xor g2041 (n_1989, A[34], n_714);
  xor g2042 (n_721, n_1989, n_687);
  nand g2043 (n_1990, A[34], n_714);
  nand g2044 (n_1991, n_687, n_714);
  nand g2045 (n_1992, A[34], n_687);
  nand g2046 (n_736, n_1990, n_1991, n_1992);
  xor g2047 (n_1993, n_716, n_717);
  xor g2048 (n_722, n_1993, n_718);
  nand g2049 (n_1994, n_716, n_717);
  nand g2050 (n_1995, n_718, n_717);
  nand g2051 (n_1996, n_716, n_718);
  nand g2052 (n_738, n_1994, n_1995, n_1996);
  xor g2053 (n_1997, n_719, n_720);
  xor g2054 (n_725, n_1997, n_721);
  nand g2055 (n_1998, n_719, n_720);
  nand g2056 (n_1999, n_721, n_720);
  nand g2057 (n_2000, n_719, n_721);
  nand g2058 (n_740, n_1998, n_1999, n_2000);
  xor g2059 (n_2001, n_722, n_723);
  xor g2060 (n_726, n_2001, n_724);
  nand g2061 (n_2002, n_722, n_723);
  nand g2062 (n_2003, n_724, n_723);
  nand g2063 (n_2004, n_722, n_724);
  nand g2064 (n_743, n_2002, n_2003, n_2004);
  xor g2065 (n_2005, n_725, n_726);
  xor g2066 (n_136, n_2005, n_727);
  nand g2067 (n_2006, n_725, n_726);
  nand g2068 (n_2007, n_727, n_726);
  nand g2069 (n_2008, n_725, n_727);
  nand g2070 (n_68, n_2006, n_2007, n_2008);
  xor g2073 (n_2009, A[47], A[31]);
  xor g2074 (n_732, n_2009, A[33]);
  nand g2075 (n_2010, A[47], A[31]);
  nand g2077 (n_2012, A[47], A[33]);
  nand g2078 (n_747, n_2010, n_1562, n_2012);
  xor g2079 (n_2013, A[29], A[45]);
  xor g2080 (n_734, n_2013, A[41]);
  nand g2081 (n_2014, A[29], A[45]);
  nand g2082 (n_2015, A[41], A[45]);
  nand g2083 (n_2016, A[29], A[41]);
  nand g2084 (n_750, n_2014, n_2015, n_2016);
  xor g2085 (n_2017, A[39], A[43]);
  xor g2086 (n_735, n_2017, A[37]);
  nand g2088 (n_2019, A[37], A[43]);
  nand g2090 (n_748, n_1951, n_2019, n_1763);
  xor g2091 (n_2021, A[35], n_700);
  xor g2092 (n_737, n_2021, n_731);
  nand g2093 (n_2022, A[35], n_700);
  nand g2094 (n_2023, n_731, n_700);
  nand g2095 (n_2024, A[35], n_731);
  nand g2096 (n_753, n_2022, n_2023, n_2024);
  xor g2097 (n_2025, n_732, n_733);
  xor g2098 (n_739, n_2025, n_734);
  nand g2099 (n_2026, n_732, n_733);
  nand g2100 (n_2027, n_734, n_733);
  nand g2101 (n_2028, n_732, n_734);
  nand g2102 (n_755, n_2026, n_2027, n_2028);
  xor g2103 (n_2029, n_735, n_736);
  xor g2104 (n_741, n_2029, n_737);
  nand g2105 (n_2030, n_735, n_736);
  nand g2106 (n_2031, n_737, n_736);
  nand g2107 (n_2032, n_735, n_737);
  nand g2108 (n_757, n_2030, n_2031, n_2032);
  xor g2109 (n_2033, n_738, n_739);
  xor g2110 (n_742, n_2033, n_740);
  nand g2111 (n_2034, n_738, n_739);
  nand g2112 (n_2035, n_740, n_739);
  nand g2113 (n_2036, n_738, n_740);
  nand g2114 (n_760, n_2034, n_2035, n_2036);
  xor g2115 (n_2037, n_741, n_742);
  xor g2116 (n_135, n_2037, n_743);
  nand g2117 (n_2038, n_741, n_742);
  nand g2118 (n_2039, n_743, n_742);
  nand g2119 (n_2040, n_741, n_743);
  nand g2120 (n_67, n_2038, n_2039, n_2040);
  xor g2124 (n_749, n_1529, A[47]);
  nand g2126 (n_2043, A[47], A[30]);
  nand g2127 (n_2044, A[32], A[47]);
  nand g2128 (n_763, n_1530, n_2043, n_2044);
  xor g2141 (n_2053, A[34], n_747);
  xor g2142 (n_754, n_2053, n_748);
  nand g2143 (n_2054, A[34], n_747);
  nand g2144 (n_2055, n_748, n_747);
  nand g2145 (n_2056, A[34], n_748);
  nand g2146 (n_768, n_2054, n_2055, n_2056);
  xor g2147 (n_2057, n_749, n_750);
  xor g2148 (n_756, n_2057, n_719);
  nand g2149 (n_2058, n_749, n_750);
  nand g2150 (n_2059, n_719, n_750);
  nand g2151 (n_2060, n_749, n_719);
  nand g2152 (n_770, n_2058, n_2059, n_2060);
  xor g2153 (n_2061, n_718, n_753);
  xor g2154 (n_758, n_2061, n_754);
  nand g2155 (n_2062, n_718, n_753);
  nand g2156 (n_2063, n_754, n_753);
  nand g2157 (n_2064, n_718, n_754);
  nand g2158 (n_772, n_2062, n_2063, n_2064);
  xor g2159 (n_2065, n_755, n_756);
  xor g2160 (n_759, n_2065, n_757);
  nand g2161 (n_2066, n_755, n_756);
  nand g2162 (n_2067, n_757, n_756);
  nand g2163 (n_2068, n_755, n_757);
  nand g2164 (n_775, n_2066, n_2067, n_2068);
  xor g2165 (n_2069, n_758, n_759);
  xor g2166 (n_134, n_2069, n_760);
  nand g2167 (n_2070, n_758, n_759);
  nand g2168 (n_2071, n_760, n_759);
  nand g2169 (n_2072, n_758, n_760);
  nand g2170 (n_66, n_2070, n_2071, n_2072);
  xor g2172 (n_762, n_2073, A[31]);
  nand g2176 (n_778, n_2074, n_1562, n_2076);
  xor g2177 (n_2077, A[41], A[45]);
  xor g2178 (n_767, n_2077, A[39]);
  nand g2180 (n_2079, A[39], A[45]);
  nand g2182 (n_779, n_2015, n_2079, n_1827);
  xor g2184 (n_766, n_2081, A[37]);
  nand g2188 (n_780, n_2082, n_2019, n_2084);
  xor g2189 (n_2085, A[35], n_762);
  xor g2190 (n_771, n_2085, n_763);
  nand g2191 (n_2086, A[35], n_762);
  nand g2192 (n_2087, n_763, n_762);
  nand g2193 (n_2088, A[35], n_763);
  nand g2194 (n_784, n_2086, n_2087, n_2088);
  xor g2195 (n_2089, n_733, n_731);
  xor g2196 (n_769, n_2089, n_766);
  nand g2197 (n_2090, n_733, n_731);
  nand g2198 (n_2091, n_766, n_731);
  nand g2199 (n_2092, n_733, n_766);
  nand g2200 (n_786, n_2090, n_2091, n_2092);
  xor g2201 (n_2093, n_767, n_768);
  xor g2202 (n_773, n_2093, n_769);
  nand g2203 (n_2094, n_767, n_768);
  nand g2204 (n_2095, n_769, n_768);
  nand g2205 (n_2096, n_767, n_769);
  nand g2206 (n_788, n_2094, n_2095, n_2096);
  xor g2207 (n_2097, n_770, n_771);
  xor g2208 (n_774, n_2097, n_772);
  nand g2209 (n_2098, n_770, n_771);
  nand g2210 (n_2099, n_772, n_771);
  nand g2211 (n_2100, n_770, n_772);
  nand g2212 (n_790, n_2098, n_2099, n_2100);
  xor g2213 (n_2101, n_773, n_774);
  xor g2214 (n_133, n_2101, n_775);
  nand g2215 (n_2102, n_773, n_774);
  nand g2216 (n_2103, n_775, n_774);
  nand g2217 (n_2104, n_773, n_775);
  nand g2218 (n_65, n_2102, n_2103, n_2104);
  xor g2234 (n_783, n_2113, n_778);
  nand g2237 (n_2116, A[34], n_778);
  nand g2238 (n_797, n_2114, n_2115, n_2116);
  xor g2239 (n_2117, n_779, n_780);
  xor g2240 (n_785, n_2117, n_718);
  nand g2241 (n_2118, n_779, n_780);
  nand g2242 (n_2119, n_718, n_780);
  nand g2243 (n_2120, n_779, n_718);
  nand g2244 (n_799, n_2118, n_2119, n_2120);
  xor g2245 (n_2121, n_719, n_783);
  xor g2246 (n_787, n_2121, n_784);
  nand g2247 (n_2122, n_719, n_783);
  nand g2248 (n_2123, n_784, n_783);
  nand g2249 (n_2124, n_719, n_784);
  nand g2250 (n_801, n_2122, n_2123, n_2124);
  xor g2251 (n_2125, n_785, n_786);
  xor g2252 (n_789, n_2125, n_787);
  nand g2253 (n_2126, n_785, n_786);
  nand g2254 (n_2127, n_787, n_786);
  nand g2255 (n_2128, n_785, n_787);
  nand g2256 (n_803, n_2126, n_2127, n_2128);
  xor g2257 (n_2129, n_788, n_789);
  xor g2258 (n_132, n_2129, n_790);
  nand g2259 (n_2130, n_788, n_789);
  nand g2260 (n_2131, n_790, n_789);
  nand g2261 (n_2132, n_788, n_790);
  nand g2262 (n_64, n_2130, n_2131, n_2132);
  xor g2264 (n_793, n_2073, A[45]);
  nand g2266 (n_2135, A[45], A[33]);
  nand g2268 (n_806, n_2074, n_2135, n_2136);
  xor g2269 (n_2137, A[41], A[39]);
  xor g2270 (n_796, n_2137, A[43]);
  nand g2273 (n_2140, A[41], A[43]);
  nand g2274 (n_807, n_1827, n_1951, n_2140);
  xor g2275 (n_2141, A[37], A[35]);
  xor g2276 (n_795, n_2141, A[32]);
  nand g2278 (n_2143, A[32], A[35]);
  nand g2279 (n_2144, A[37], A[32]);
  nand g2280 (n_809, n_1956, n_2143, n_2144);
  xor g2281 (n_2145, n_731, n_793);
  xor g2282 (n_798, n_2145, n_733);
  nand g2283 (n_2146, n_731, n_793);
  nand g2284 (n_2147, n_733, n_793);
  nand g2286 (n_811, n_2146, n_2147, n_2090);
  xor g2287 (n_2149, n_795, n_796);
  xor g2288 (n_800, n_2149, n_797);
  nand g2289 (n_2150, n_795, n_796);
  nand g2290 (n_2151, n_797, n_796);
  nand g2291 (n_2152, n_795, n_797);
  nand g2292 (n_813, n_2150, n_2151, n_2152);
  xor g2293 (n_2153, n_798, n_799);
  xor g2294 (n_802, n_2153, n_800);
  nand g2295 (n_2154, n_798, n_799);
  nand g2296 (n_2155, n_800, n_799);
  nand g2297 (n_2156, n_798, n_800);
  nand g2298 (n_816, n_2154, n_2155, n_2156);
  xor g2299 (n_2157, n_801, n_802);
  xor g2300 (n_131, n_2157, n_803);
  nand g2301 (n_2158, n_801, n_802);
  nand g2302 (n_2159, n_803, n_802);
  nand g2303 (n_2160, n_801, n_803);
  nand g2304 (n_63, n_2158, n_2159, n_2160);
  xor g2307 (n_2161, A[44], A[40]);
  xor g2308 (n_810, n_2161, A[38]);
  nand g2311 (n_2164, A[44], A[38]);
  nand g2312 (n_818, n_1983, n_1795, n_2164);
  xor g2313 (n_2165, A[42], A[36]);
  xor g2314 (n_808, n_2165, A[34]);
  nand g2317 (n_2168, A[42], A[34]);
  nand g2318 (n_819, n_1987, n_1924, n_2168);
  xor g2320 (n_812, n_2169, n_807);
  nand g2322 (n_2171, n_807, n_806);
  nand g2324 (n_823, n_2170, n_2171, n_2172);
  xor g2325 (n_2173, n_808, n_809);
  xor g2326 (n_814, n_2173, n_810);
  nand g2327 (n_2174, n_808, n_809);
  nand g2328 (n_2175, n_810, n_809);
  nand g2329 (n_2176, n_808, n_810);
  nand g2330 (n_824, n_2174, n_2175, n_2176);
  xor g2331 (n_2177, n_811, n_812);
  xor g2332 (n_815, n_2177, n_813);
  nand g2333 (n_2178, n_811, n_812);
  nand g2334 (n_2179, n_813, n_812);
  nand g2335 (n_2180, n_811, n_813);
  nand g2336 (n_827, n_2178, n_2179, n_2180);
  xor g2337 (n_2181, n_814, n_815);
  xor g2338 (n_130, n_2181, n_816);
  nand g2339 (n_2182, n_814, n_815);
  nand g2340 (n_2183, n_816, n_815);
  nand g2341 (n_2184, n_814, n_816);
  nand g2342 (n_62, n_2182, n_2183, n_2184);
  xor g2344 (n_821, n_2185, A[41]);
  nand g2348 (n_831, n_2136, n_2015, n_2188);
  xor g2355 (n_2193, A[35], A[46]);
  xor g2356 (n_822, n_2193, n_818);
  nand g2357 (n_2194, A[35], A[46]);
  nand g2358 (n_2195, n_818, A[46]);
  nand g2359 (n_2196, A[35], n_818);
  nand g2360 (n_834, n_2194, n_2195, n_2196);
  xor g2361 (n_2197, n_819, n_735);
  xor g2362 (n_825, n_2197, n_821);
  nand g2363 (n_2198, n_819, n_735);
  nand g2364 (n_2199, n_821, n_735);
  nand g2365 (n_2200, n_819, n_821);
  nand g2366 (n_835, n_2198, n_2199, n_2200);
  xor g2367 (n_2201, n_822, n_823);
  xor g2368 (n_826, n_2201, n_824);
  nand g2369 (n_2202, n_822, n_823);
  nand g2370 (n_2203, n_824, n_823);
  nand g2371 (n_2204, n_822, n_824);
  nand g2372 (n_838, n_2202, n_2203, n_2204);
  xor g2373 (n_2205, n_825, n_826);
  xor g2374 (n_129, n_2205, n_827);
  nand g2375 (n_2206, n_825, n_826);
  nand g2376 (n_2207, n_827, n_826);
  nand g2377 (n_2208, n_825, n_827);
  nand g2378 (n_61, n_2206, n_2207, n_2208);
  xor g2381 (n_2209, A[40], A[38]);
  xor g2382 (n_832, n_2209, A[46]);
  nand g2384 (n_2211, A[46], A[38]);
  nand g2386 (n_840, n_1795, n_2211, n_1982);
  nand g2392 (n_843, n_1987, n_2215, n_2216);
  xor g2393 (n_2217, n_748, n_831);
  xor g2394 (n_836, n_2217, n_832);
  nand g2395 (n_2218, n_748, n_831);
  nand g2396 (n_2219, n_832, n_831);
  nand g2397 (n_2220, n_748, n_832);
  nand g2398 (n_845, n_2218, n_2219, n_2220);
  xor g2399 (n_2221, n_833, n_834);
  xor g2400 (n_837, n_2221, n_835);
  nand g2401 (n_2222, n_833, n_834);
  nand g2402 (n_2223, n_835, n_834);
  nand g2403 (n_2224, n_833, n_835);
  nand g2404 (n_847, n_2222, n_2223, n_2224);
  xor g2405 (n_2225, n_836, n_837);
  xor g2406 (n_128, n_2225, n_838);
  nand g2407 (n_2226, n_836, n_837);
  nand g2408 (n_2227, n_838, n_837);
  nand g2409 (n_2228, n_836, n_838);
  nand g2410 (n_60, n_2226, n_2227, n_2228);
  xor g2423 (n_2237, A[44], n_840);
  xor g2424 (n_844, n_2237, n_735);
  nand g2425 (n_2238, A[44], n_840);
  nand g2426 (n_2239, n_735, n_840);
  nand g2427 (n_2240, A[44], n_735);
  nand g2428 (n_854, n_2238, n_2239, n_2240);
  xor g2429 (n_2241, n_821, n_843);
  xor g2430 (n_846, n_2241, n_844);
  nand g2431 (n_2242, n_821, n_843);
  nand g2432 (n_2243, n_844, n_843);
  nand g2433 (n_2244, n_821, n_844);
  nand g2434 (n_856, n_2242, n_2243, n_2244);
  xor g2435 (n_2245, n_845, n_846);
  xor g2436 (n_127, n_2245, n_847);
  nand g2437 (n_2246, n_845, n_846);
  nand g2438 (n_2247, n_847, n_846);
  nand g2439 (n_2248, n_845, n_847);
  nand g2440 (n_59, n_2246, n_2247, n_2248);
  nand g2453 (n_2256, A[42], n_748);
  nand g2454 (n_861, n_2215, n_2255, n_2256);
  xor g2455 (n_2257, n_831, n_832);
  xor g2456 (n_855, n_2257, n_853);
  nand g2458 (n_2259, n_853, n_832);
  nand g2459 (n_2260, n_831, n_853);
  nand g2460 (n_863, n_2219, n_2259, n_2260);
  xor g2461 (n_2261, n_854, n_855);
  xor g2462 (n_126, n_2261, n_856);
  nand g2463 (n_2262, n_854, n_855);
  nand g2464 (n_2263, n_856, n_855);
  nand g2465 (n_2264, n_854, n_856);
  nand g2466 (n_125, n_2262, n_2263, n_2264);
  xor g2474 (n_860, n_2017, A[44]);
  nand g2476 (n_2271, A[44], A[43]);
  nand g2477 (n_2272, A[39], A[44]);
  nand g2478 (n_868, n_1951, n_2271, n_2272);
  xor g2479 (n_2273, n_840, n_821);
  xor g2480 (n_862, n_2273, n_860);
  nand g2481 (n_2274, n_840, n_821);
  nand g2482 (n_2275, n_860, n_821);
  nand g2483 (n_2276, n_840, n_860);
  nand g2484 (n_870, n_2274, n_2275, n_2276);
  xor g2485 (n_2277, n_861, n_862);
  xor g2486 (n_58, n_2277, n_863);
  nand g2487 (n_2278, n_861, n_862);
  nand g2488 (n_2279, n_863, n_862);
  nand g2489 (n_2280, n_861, n_863);
  nand g2490 (n_124, n_2278, n_2279, n_2280);
  xor g2494 (n_867, n_2161, A[42]);
  nand g2496 (n_2283, A[42], A[44]);
  nand g2497 (n_2284, A[40], A[42]);
  nand g2498 (n_872, n_1983, n_2283, n_2284);
  xor g2500 (n_869, n_2285, n_867);
  nand g2502 (n_2287, n_867, n_831);
  nand g2504 (n_875, n_2286, n_2287, n_2288);
  xor g2505 (n_2289, n_868, n_869);
  xor g2506 (n_57, n_2289, n_870);
  nand g2507 (n_2290, n_868, n_869);
  nand g2508 (n_2291, n_870, n_869);
  nand g2509 (n_2292, n_868, n_870);
  nand g2510 (n_123, n_2290, n_2291, n_2292);
  xor g2517 (n_2297, A[43], A[46]);
  xor g2518 (n_874, n_2297, n_872);
  nand g2519 (n_2298, A[43], A[46]);
  nand g2520 (n_2299, n_872, A[46]);
  nand g2521 (n_2300, A[43], n_872);
  nand g2522 (n_880, n_2298, n_2299, n_2300);
  xor g2523 (n_2301, n_821, n_874);
  xor g2524 (n_56, n_2301, n_875);
  nand g2525 (n_2302, n_821, n_874);
  nand g2526 (n_2303, n_875, n_874);
  nand g2527 (n_2304, n_821, n_875);
  nand g2528 (n_122, n_2302, n_2303, n_2304);
  xor g2531 (n_2305, A[44], A[42]);
  nand g2536 (n_883, n_2283, n_2307, n_2308);
  xor g2537 (n_2309, n_831, n_879);
  xor g2538 (n_55, n_2309, n_880);
  nand g2539 (n_2310, n_831, n_879);
  nand g2540 (n_2311, n_880, n_879);
  nand g2541 (n_2312, n_831, n_880);
  nand g2542 (n_121, n_2310, n_2311, n_2312);
  xor g2544 (n_882, n_2185, A[43]);
  nand g2546 (n_2315, A[43], A[45]);
  nand g2548 (n_886, n_2136, n_2315, n_2082);
  xor g2549 (n_2317, A[46], n_882);
  xor g2550 (n_54, n_2317, n_883);
  nand g2551 (n_2318, A[46], n_882);
  nand g2552 (n_2319, n_883, n_882);
  nand g2553 (n_2320, A[46], n_883);
  nand g2554 (n_120, n_2318, n_2319, n_2320);
  xor g2558 (n_53, n_2321, n_886);
  nand g2561 (n_2324, A[46], n_886);
  nand g2562 (n_119, n_2322, n_2323, n_2324);
  xor g2564 (n_52, n_2185, A[44]);
  nand g2566 (n_2327, A[44], A[45]);
  nand g2568 (n_118, n_2136, n_2327, n_2328);
  nor g11 (n_2344, A[2], A[0]);
  nor g13 (n_2340, A[3], A[1]);
  nor g15 (n_2350, A[0], n_178);
  nand g16 (n_2345, A[0], n_178);
  nor g17 (n_2346, n_110, n_177);
  nand g18 (n_2347, n_110, n_177);
  nor g19 (n_2356, n_109, n_176);
  nand g20 (n_2351, n_109, n_176);
  nor g21 (n_2352, n_108, n_175);
  nand g22 (n_2353, n_108, n_175);
  nor g23 (n_2362, n_107, n_174);
  nand g24 (n_2357, n_107, n_174);
  nor g25 (n_2358, n_106, n_173);
  nand g26 (n_2359, n_106, n_173);
  nor g27 (n_2368, n_105, n_172);
  nand g28 (n_2363, n_105, n_172);
  nor g29 (n_2364, n_104, n_171);
  nand g30 (n_2365, n_104, n_171);
  nor g31 (n_2374, n_103, n_170);
  nand g32 (n_2369, n_103, n_170);
  nor g33 (n_2370, n_102, n_169);
  nand g34 (n_2371, n_102, n_169);
  nor g35 (n_2380, n_101, n_168);
  nand g36 (n_2375, n_101, n_168);
  nor g37 (n_2376, n_100, n_167);
  nand g38 (n_2377, n_100, n_167);
  nor g39 (n_2386, n_99, n_166);
  nand g40 (n_2381, n_99, n_166);
  nor g41 (n_2382, n_98, n_165);
  nand g42 (n_2383, n_98, n_165);
  nor g43 (n_2392, n_97, n_164);
  nand g44 (n_2387, n_97, n_164);
  nor g45 (n_2388, n_96, n_163);
  nand g46 (n_2389, n_96, n_163);
  nor g47 (n_2398, n_95, n_162);
  nand g48 (n_2393, n_95, n_162);
  nor g49 (n_2394, n_94, n_161);
  nand g50 (n_2395, n_94, n_161);
  nor g51 (n_2404, n_93, n_160);
  nand g52 (n_2399, n_93, n_160);
  nor g53 (n_2400, n_92, n_159);
  nand g54 (n_2401, n_92, n_159);
  nor g55 (n_2410, n_91, n_158);
  nand g56 (n_2405, n_91, n_158);
  nor g57 (n_2406, n_90, n_157);
  nand g58 (n_2407, n_90, n_157);
  nor g59 (n_2416, n_89, n_156);
  nand g60 (n_2411, n_89, n_156);
  nor g61 (n_2412, n_88, n_155);
  nand g62 (n_2413, n_88, n_155);
  nor g63 (n_2422, n_87, n_154);
  nand g64 (n_2417, n_87, n_154);
  nor g65 (n_2418, n_86, n_153);
  nand g66 (n_2419, n_86, n_153);
  nor g67 (n_2428, n_85, n_152);
  nand g68 (n_2423, n_85, n_152);
  nor g69 (n_2424, n_84, n_151);
  nand g70 (n_2425, n_84, n_151);
  nor g71 (n_2434, n_83, n_150);
  nand g72 (n_2429, n_83, n_150);
  nor g73 (n_2430, n_82, n_149);
  nand g74 (n_2431, n_82, n_149);
  nor g75 (n_2440, n_81, n_148);
  nand g76 (n_2435, n_81, n_148);
  nor g77 (n_2436, n_80, n_147);
  nand g78 (n_2437, n_80, n_147);
  nor g79 (n_2446, n_79, n_146);
  nand g80 (n_2441, n_79, n_146);
  nor g81 (n_2442, n_78, n_145);
  nand g82 (n_2443, n_78, n_145);
  nor g83 (n_2452, n_77, n_144);
  nand g84 (n_2447, n_77, n_144);
  nor g85 (n_2448, n_76, n_143);
  nand g86 (n_2449, n_76, n_143);
  nor g87 (n_2458, n_75, n_142);
  nand g88 (n_2453, n_75, n_142);
  nor g89 (n_2454, n_74, n_141);
  nand g90 (n_2455, n_74, n_141);
  nor g91 (n_2464, n_73, n_140);
  nand g92 (n_2459, n_73, n_140);
  nor g93 (n_2460, n_72, n_139);
  nand g94 (n_2461, n_72, n_139);
  nor g95 (n_2470, n_71, n_138);
  nand g96 (n_2465, n_71, n_138);
  nor g97 (n_2466, n_70, n_137);
  nand g98 (n_2467, n_70, n_137);
  nor g99 (n_2476, n_69, n_136);
  nand g100 (n_2471, n_69, n_136);
  nor g101 (n_2472, n_68, n_135);
  nand g102 (n_2473, n_68, n_135);
  nor g103 (n_2482, n_67, n_134);
  nand g104 (n_2477, n_67, n_134);
  nor g105 (n_2478, n_66, n_133);
  nand g106 (n_2479, n_66, n_133);
  nor g107 (n_2488, n_65, n_132);
  nand g108 (n_2483, n_65, n_132);
  nor g109 (n_2484, n_64, n_131);
  nand g110 (n_2485, n_64, n_131);
  nor g111 (n_2494, n_63, n_130);
  nand g112 (n_2489, n_63, n_130);
  nor g113 (n_2490, n_62, n_129);
  nand g114 (n_2491, n_62, n_129);
  nor g115 (n_2500, n_61, n_128);
  nand g116 (n_2495, n_61, n_128);
  nor g117 (n_2496, n_60, n_127);
  nand g118 (n_2497, n_60, n_127);
  nor g119 (n_2506, n_59, n_126);
  nand g120 (n_2501, n_59, n_126);
  nor g121 (n_2502, n_58, n_125);
  nand g122 (n_2503, n_58, n_125);
  nor g123 (n_2512, n_57, n_124);
  nand g124 (n_2507, n_57, n_124);
  nor g125 (n_2508, n_56, n_123);
  nand g126 (n_2509, n_56, n_123);
  nor g127 (n_2518, n_55, n_122);
  nand g128 (n_2513, n_55, n_122);
  nor g129 (n_2514, n_54, n_121);
  nand g130 (n_2515, n_54, n_121);
  nor g131 (n_2524, n_53, n_120);
  nand g132 (n_2519, n_53, n_120);
  nor g133 (n_2520, n_52, n_119);
  nand g134 (n_2521, n_52, n_119);
  nor g144 (n_2342, n_894, n_2340);
  nor g148 (n_2348, n_2345, n_2346);
  nor g151 (n_2541, n_2350, n_2346);
  nor g152 (n_2354, n_2351, n_2352);
  nor g155 (n_2535, n_2356, n_2352);
  nor g156 (n_2360, n_2357, n_2358);
  nor g159 (n_2548, n_2362, n_2358);
  nor g160 (n_2366, n_2363, n_2364);
  nor g163 (n_2542, n_2368, n_2364);
  nor g164 (n_2372, n_2369, n_2370);
  nor g167 (n_2555, n_2374, n_2370);
  nor g168 (n_2378, n_2375, n_2376);
  nor g171 (n_2549, n_2380, n_2376);
  nor g172 (n_2384, n_2381, n_2382);
  nor g175 (n_2562, n_2386, n_2382);
  nor g176 (n_2390, n_2387, n_2388);
  nor g179 (n_2556, n_2392, n_2388);
  nor g180 (n_2396, n_2393, n_2394);
  nor g183 (n_2569, n_2398, n_2394);
  nor g184 (n_2402, n_2399, n_2400);
  nor g187 (n_2563, n_2404, n_2400);
  nor g188 (n_2408, n_2405, n_2406);
  nor g191 (n_2576, n_2410, n_2406);
  nor g192 (n_2414, n_2411, n_2412);
  nor g195 (n_2570, n_2416, n_2412);
  nor g196 (n_2420, n_2417, n_2418);
  nor g199 (n_2583, n_2422, n_2418);
  nor g200 (n_2426, n_2423, n_2424);
  nor g203 (n_2577, n_2428, n_2424);
  nor g204 (n_2432, n_2429, n_2430);
  nor g207 (n_2590, n_2434, n_2430);
  nor g208 (n_2438, n_2435, n_2436);
  nor g211 (n_2584, n_2440, n_2436);
  nor g212 (n_2444, n_2441, n_2442);
  nor g215 (n_2597, n_2446, n_2442);
  nor g216 (n_2450, n_2447, n_2448);
  nor g219 (n_2591, n_2452, n_2448);
  nor g220 (n_2456, n_2453, n_2454);
  nor g223 (n_2604, n_2458, n_2454);
  nor g224 (n_2462, n_2459, n_2460);
  nor g227 (n_2598, n_2464, n_2460);
  nor g228 (n_2468, n_2465, n_2466);
  nor g231 (n_2611, n_2470, n_2466);
  nor g232 (n_2474, n_2471, n_2472);
  nor g235 (n_2605, n_2476, n_2472);
  nor g236 (n_2480, n_2477, n_2478);
  nor g239 (n_2618, n_2482, n_2478);
  nor g240 (n_2486, n_2483, n_2484);
  nor g243 (n_2612, n_2488, n_2484);
  nor g244 (n_2492, n_2489, n_2490);
  nor g247 (n_2625, n_2494, n_2490);
  nor g248 (n_2498, n_2495, n_2496);
  nor g251 (n_2619, n_2500, n_2496);
  nor g252 (n_2504, n_2501, n_2502);
  nor g255 (n_2632, n_2506, n_2502);
  nor g256 (n_2510, n_2507, n_2508);
  nor g259 (n_2626, n_2512, n_2508);
  nor g260 (n_2516, n_2513, n_2514);
  nor g263 (n_2639, n_2518, n_2514);
  nor g264 (n_2522, n_2519, n_2520);
  nor g267 (n_2633, n_2524, n_2520);
  nor g268 (n_2528, n_2525, n_2526);
  nor g271 (n_2772, n_2530, n_2526);
  nand g278 (n_2640, n_2541, n_2535);
  nand g283 (n_2650, n_2548, n_2542);
  nand g288 (n_2645, n_2555, n_2549);
  nand g293 (n_2656, n_2562, n_2556);
  nand g298 (n_2651, n_2569, n_2563);
  nand g303 (n_2662, n_2576, n_2570);
  nand g308 (n_2657, n_2583, n_2577);
  nand g313 (n_2668, n_2590, n_2584);
  nand g318 (n_2663, n_2597, n_2591);
  nand g323 (n_2674, n_2604, n_2598);
  nand g328 (n_2669, n_2611, n_2605);
  nand g333 (n_2680, n_2618, n_2612);
  nand g338 (n_2675, n_2625, n_2619);
  nand g343 (n_2686, n_2632, n_2626);
  nand g348 (n_2681, n_2639, n_2633);
  nand g351 (n_2688, n_2643, n_2644);
  nor g352 (n_2648, n_2645, n_2646);
  nor g355 (n_2687, n_2650, n_2645);
  nor g356 (n_2654, n_2651, n_2652);
  nor g359 (n_2697, n_2656, n_2651);
  nor g360 (n_2660, n_2657, n_2658);
  nor g363 (n_2691, n_2662, n_2657);
  nor g364 (n_2666, n_2663, n_2664);
  nor g367 (n_2704, n_2668, n_2663);
  nor g368 (n_2672, n_2669, n_2670);
  nor g371 (n_2698, n_2674, n_2669);
  nor g372 (n_2678, n_2675, n_2676);
  nor g375 (n_2711, n_2680, n_2675);
  nor g376 (n_2684, n_2681, n_2682);
  nor g379 (n_2705, n_2686, n_2681);
  nand g2576 (n_2690, n_2687, n_2688);
  nand g2577 (n_2713, n_2689, n_2690);
  nand g2582 (n_2712, n_2697, n_2691);
  nand g2587 (n_2722, n_2704, n_2698);
  nand g2592 (n_2717, n_2711, n_2705);
  nand g2595 (n_2724, n_2715, n_2716);
  nor g2596 (n_2720, n_2717, n_2718);
  nor g2599 (n_2723, n_2722, n_2717);
  nand g2600 (n_2726, n_2723, n_2724);
  nand g2601 (n_2773, n_2725, n_2726);
  nand g2604 (n_2731, n_2718, n_2728);
  nand g2605 (n_2729, n_2697, n_2713);
  nand g2606 (n_2737, n_2692, n_2729);
  nand g2607 (n_2730, n_2704, n_2724);
  nand g2608 (n_2742, n_2699, n_2730);
  nand g2609 (n_2732, n_2711, n_2731);
  nand g2610 (n_2747, n_2706, n_2732);
  nand g2613 (n_2752, n_2646, n_2734);
  nand g2616 (n_2755, n_2652, n_2736);
  nand g2619 (n_2758, n_2658, n_2739);
  nand g2622 (n_2761, n_2664, n_2741);
  nand g2625 (n_2764, n_2670, n_2744);
  nand g2628 (n_2767, n_2676, n_2746);
  nand g2631 (n_2770, n_2682, n_2749);
  nand g2633 (n_2780, n_2536, n_2750);
  nand g2634 (n_2751, n_2548, n_2688);
  nand g2635 (n_2785, n_2543, n_2751);
  nand g2636 (n_2753, n_2555, n_2752);
  nand g2637 (n_2790, n_2550, n_2753);
  nand g2638 (n_2754, n_2562, n_2713);
  nand g2639 (n_2795, n_2557, n_2754);
  nand g2640 (n_2756, n_2569, n_2755);
  nand g2641 (n_2800, n_2564, n_2756);
  nand g2642 (n_2757, n_2576, n_2737);
  nand g2643 (n_2805, n_2571, n_2757);
  nand g2644 (n_2759, n_2583, n_2758);
  nand g2645 (n_2810, n_2578, n_2759);
  nand g2646 (n_2760, n_2590, n_2724);
  nand g2647 (n_2815, n_2585, n_2760);
  nand g2648 (n_2762, n_2597, n_2761);
  nand g2649 (n_2820, n_2592, n_2762);
  nand g2650 (n_2763, n_2604, n_2742);
  nand g2651 (n_2825, n_2599, n_2763);
  nand g2652 (n_2765, n_2611, n_2764);
  nand g2653 (n_2830, n_2606, n_2765);
  nand g2654 (n_2766, n_2618, n_2731);
  nand g2655 (n_2835, n_2613, n_2766);
  nand g2656 (n_2768, n_2625, n_2767);
  nand g2657 (n_2840, n_2620, n_2768);
  nand g2658 (n_2769, n_2632, n_2747);
  nand g2659 (n_2845, n_2627, n_2769);
  nand g2660 (n_2771, n_2639, n_2770);
  nand g2661 (n_2850, n_2634, n_2771);
  nand g2662 (n_2775, n_2772, n_2773);
  nand g2663 (n_2856, n_2774, n_2775);
  nand g2669 (n_2866, n_2345, n_2779);
  nand g2672 (n_2870, n_2351, n_2782);
  nand g2675 (n_2874, n_2357, n_2784);
  nand g2678 (n_2878, n_2363, n_2787);
  nand g2681 (n_2882, n_2369, n_2789);
  nand g2684 (n_2886, n_2375, n_2792);
  nand g2687 (n_2890, n_2381, n_2794);
  nand g2690 (n_2894, n_2387, n_2797);
  nand g2693 (n_2898, n_2393, n_2799);
  nand g2696 (n_2902, n_2399, n_2802);
  nand g2699 (n_2906, n_2405, n_2804);
  nand g2702 (n_2910, n_2411, n_2807);
  nand g2705 (n_2914, n_2417, n_2809);
  nand g2708 (n_2918, n_2423, n_2812);
  nand g2711 (n_2922, n_2429, n_2814);
  nand g2714 (n_2926, n_2435, n_2817);
  nand g2717 (n_2930, n_2441, n_2819);
  nand g2720 (n_2934, n_2447, n_2822);
  nand g2723 (n_2938, n_2453, n_2824);
  nand g2726 (n_2942, n_2459, n_2827);
  nand g2729 (n_2946, n_2465, n_2829);
  nand g2732 (n_2950, n_2471, n_2832);
  nand g2735 (n_2954, n_2477, n_2834);
  nand g2738 (n_2958, n_2483, n_2837);
  nand g2741 (n_2962, n_2489, n_2839);
  nand g2744 (n_2966, n_2495, n_2842);
  nand g2747 (n_2970, n_2501, n_2844);
  nand g2750 (n_2974, n_2507, n_2847);
  nand g2753 (n_2978, n_2513, n_2849);
  nand g2756 (n_2982, n_2519, n_2852);
  nand g2759 (n_2986, n_2525, n_2854);
  xnor g2772 (Z[5], n_2866, n_2867);
  xnor g2774 (Z[6], n_2780, n_2868);
  xnor g2777 (Z[7], n_2870, n_2871);
  xnor g2779 (Z[8], n_2688, n_2872);
  xnor g2782 (Z[9], n_2874, n_2875);
  xnor g2784 (Z[10], n_2785, n_2876);
  xnor g2787 (Z[11], n_2878, n_2879);
  xnor g2789 (Z[12], n_2752, n_2880);
  xnor g2792 (Z[13], n_2882, n_2883);
  xnor g2794 (Z[14], n_2790, n_2884);
  xnor g2797 (Z[15], n_2886, n_2887);
  xnor g2799 (Z[16], n_2713, n_2888);
  xnor g2802 (Z[17], n_2890, n_2891);
  xnor g2804 (Z[18], n_2795, n_2892);
  xnor g2807 (Z[19], n_2894, n_2895);
  xnor g2809 (Z[20], n_2755, n_2896);
  xnor g2812 (Z[21], n_2898, n_2899);
  xnor g2814 (Z[22], n_2800, n_2900);
  xnor g2817 (Z[23], n_2902, n_2903);
  xnor g2819 (Z[24], n_2737, n_2904);
  xnor g2822 (Z[25], n_2906, n_2907);
  xnor g2824 (Z[26], n_2805, n_2908);
  xnor g2827 (Z[27], n_2910, n_2911);
  xnor g2829 (Z[28], n_2758, n_2912);
  xnor g2832 (Z[29], n_2914, n_2915);
  xnor g2834 (Z[30], n_2810, n_2916);
  xnor g2837 (Z[31], n_2918, n_2919);
  xnor g2839 (Z[32], n_2724, n_2920);
  xnor g2842 (Z[33], n_2922, n_2923);
  xnor g2844 (Z[34], n_2815, n_2924);
  xnor g2847 (Z[35], n_2926, n_2927);
  xnor g2849 (Z[36], n_2761, n_2928);
  xnor g2852 (Z[37], n_2930, n_2931);
  xnor g2854 (Z[38], n_2820, n_2932);
  xnor g2857 (Z[39], n_2934, n_2935);
  xnor g2859 (Z[40], n_2742, n_2936);
  xnor g2862 (Z[41], n_2938, n_2939);
  xnor g2864 (Z[42], n_2825, n_2940);
  xnor g2867 (Z[43], n_2942, n_2943);
  xnor g2869 (Z[44], n_2764, n_2944);
  xnor g2872 (Z[45], n_2946, n_2947);
  xnor g2874 (Z[46], n_2830, n_2948);
  xnor g2877 (Z[47], n_2950, n_2951);
  xnor g2879 (Z[48], n_2731, n_2952);
  xnor g2882 (Z[49], n_2954, n_2955);
  xnor g2884 (Z[50], n_2835, n_2956);
  xnor g2887 (Z[51], n_2958, n_2959);
  xnor g2889 (Z[52], n_2767, n_2960);
  xnor g2892 (Z[53], n_2962, n_2963);
  xnor g2894 (Z[54], n_2840, n_2964);
  xnor g2897 (Z[55], n_2966, n_2967);
  xnor g2899 (Z[56], n_2747, n_2968);
  xnor g2902 (Z[57], n_2970, n_2971);
  xnor g2904 (Z[58], n_2845, n_2972);
  xnor g2907 (Z[59], n_2974, n_2975);
  xnor g2909 (Z[60], n_2770, n_2976);
  xnor g2912 (Z[61], n_2978, n_2979);
  xnor g2914 (Z[62], n_2850, n_2980);
  xnor g2917 (Z[63], n_2982, n_2983);
  xnor g2919 (Z[64], n_2773, n_2984);
  xnor g2922 (Z[65], n_2986, n_2987);
  or g2938 (n_258, wc, wc0, n_110);
  not gc0 (wc0, n_894);
  not gc (wc, n_907);
  or g2939 (n_267, wc1, n_252, n_110);
  not gc1 (wc1, n_927);
  or g2940 (n_280, wc2, n_257, n_252);
  not gc2 (wc2, n_955);
  or g2941 (n_297, wc3, n_266, n_257);
  not gc3 (wc3, n_991);
  or g2942 (n_318, wc4, wc5, n_266);
  not gc5 (wc5, n_1034);
  not gc4 (wc4, n_1035);
  or g2943 (n_319, wc6, wc7, n_252);
  not gc7 (wc7, n_1038);
  not gc6 (wc6, n_1040);
  or g2944 (n_114, wc8, wc9, n_110);
  not gc9 (wc9, n_1040);
  not gc8 (wc8, n_1088);
  or g2945 (n_115, wc10, wc11, n_266);
  not gc11 (wc11, n_1090);
  not gc10 (wc10, n_1091);
  or g2946 (n_395, wc12, wc13, n_257);
  not gc13 (wc13, n_1091);
  not gc12 (wc12, n_1215);
  or g2947 (n_421, wc14, wc15, n_266);
  not gc15 (wc15, n_1155);
  not gc14 (wc14, n_1279);
  or g2948 (n_449, wc16, wc17, n_279);
  not gc17 (wc17, n_1219);
  not gc16 (wc16, n_1343);
  or g2949 (n_477, wc18, wc19, n_296);
  not gc19 (wc19, n_1148);
  not gc18 (wc18, n_1407);
  or g2950 (n_505, wc20, wc21, n_317);
  not gc21 (wc21, n_1212);
  not gc20 (wc20, n_1471);
  or g2951 (n_533, wc22, wc23, n_113);
  not gc23 (wc23, n_1276);
  not gc22 (wc22, n_1535);
  or g2952 (n_562, wc24, wc25, n_113);
  not gc25 (wc25, n_1598);
  not gc24 (wc24, n_1599);
  xnor g2953 (n_2073, A[47], A[33]);
  or g2954 (n_2074, wc26, A[47]);
  not gc26 (wc26, A[33]);
  or g2955 (n_2076, wc27, A[47]);
  not gc27 (wc27, A[31]);
  xnor g2956 (n_2113, A[34], A[32]);
  or g2957 (n_2114, A[32], wc28);
  not gc28 (wc28, A[34]);
  or g2958 (n_2136, wc29, A[47]);
  not gc29 (wc29, A[45]);
  xnor g2959 (n_2185, A[47], A[45]);
  or g2960 (n_2188, wc30, A[47]);
  not gc30 (wc30, A[41]);
  xnor g2961 (n_833, n_2165, A[44]);
  or g2962 (n_2215, wc31, A[44]);
  not gc31 (wc31, A[42]);
  or g2963 (n_2216, wc32, A[44]);
  not gc32 (wc32, A[36]);
  xnor g2965 (n_879, n_2305, A[46]);
  or g2966 (n_2307, wc33, A[46]);
  not gc33 (wc33, A[42]);
  or g2967 (n_2308, wc34, A[46]);
  not gc34 (wc34, A[44]);
  or g2968 (n_2082, wc35, A[47]);
  not gc35 (wc35, A[43]);
  xnor g2969 (n_2321, A[46], A[44]);
  or g2970 (n_2322, A[44], wc36);
  not gc36 (wc36, A[46]);
  or g2971 (n_2328, wc37, A[47]);
  not gc37 (wc37, A[44]);
  and g2972 (n_2526, wc38, A[47]);
  not gc38 (wc38, A[46]);
  or g2973 (n_2527, wc39, A[47]);
  not gc39 (wc39, A[46]);
  or g2974 (n_2172, A[46], wc40);
  not gc40 (wc40, n_807);
  xnor g2975 (n_853, n_748, n_2305);
  or g2976 (n_2255, A[44], wc41);
  not gc41 (wc41, n_748);
  or g2977 (n_2288, A[46], wc42);
  not gc42 (wc42, n_867);
  and g2978 (n_2533, wc43, n_891);
  not gc43 (wc43, n_2342);
  or g2980 (n_2860, n_2344, wc44);
  not gc44 (wc44, n_894);
  or g2981 (n_2863, n_2340, wc45);
  not gc45 (wc45, n_891);
  xnor g2982 (n_2081, A[47], A[43]);
  or g2983 (n_2084, wc46, A[47]);
  not gc46 (wc46, A[37]);
  or g2984 (n_2115, A[32], wc47);
  not gc47 (wc47, n_778);
  xnor g2985 (n_2169, n_806, A[46]);
  or g2986 (n_2170, A[46], wc48);
  not gc48 (wc48, n_806);
  xnor g2987 (n_2285, n_831, A[46]);
  or g2988 (n_2286, A[46], wc49);
  not gc49 (wc49, n_831);
  or g2989 (n_2323, A[44], wc50);
  not gc50 (wc50, n_886);
  and g2990 (n_2530, A[46], wc51);
  not gc51 (wc51, n_118);
  or g2991 (n_2525, A[46], wc52);
  not gc52 (wc52, n_118);
  or g2992 (n_2864, wc53, n_2350);
  not gc53 (wc53, n_2345);
  or g2993 (n_2987, wc54, n_2526);
  not gc54 (wc54, n_2527);
  and g2994 (n_2536, wc55, n_2347);
  not gc55 (wc55, n_2348);
  not g2995 (Z[2], n_2860);
  or g2996 (n_2867, wc56, n_2346);
  not gc56 (wc56, n_2347);
  or g2997 (n_2868, wc57, n_2356);
  not gc57 (wc57, n_2351);
  and g2998 (n_2538, wc58, n_2353);
  not gc58 (wc58, n_2354);
  and g2999 (n_2774, n_2527, wc59);
  not gc59 (wc59, n_2528);
  or g3002 (n_2871, wc60, n_2352);
  not gc60 (wc60, n_2353);
  or g3003 (n_2984, wc61, n_2530);
  not gc61 (wc61, n_2525);
  and g3004 (n_2543, wc62, n_2359);
  not gc62 (wc62, n_2360);
  and g3005 (n_2539, wc63, n_2535);
  not gc63 (wc63, n_2536);
  or g3006 (n_2750, n_2533, wc64);
  not gc64 (wc64, n_2541);
  or g3007 (n_2779, n_2350, n_2533);
  xor g3008 (Z[3], n_894, n_2863);
  xor g3009 (Z[4], n_2533, n_2864);
  or g3010 (n_2872, wc65, n_2362);
  not gc65 (wc65, n_2357);
  or g3011 (n_2875, wc66, n_2358);
  not gc66 (wc66, n_2359);
  and g3012 (n_2636, wc67, n_2521);
  not gc67 (wc67, n_2522);
  and g3013 (n_2643, wc68, n_2538);
  not gc68 (wc68, n_2539);
  or g3014 (n_2644, n_2640, n_2533);
  or g3015 (n_2876, wc69, n_2368);
  not gc69 (wc69, n_2363);
  or g3016 (n_2980, wc70, n_2524);
  not gc70 (wc70, n_2519);
  or g3017 (n_2983, wc71, n_2520);
  not gc71 (wc71, n_2521);
  and g3018 (n_2545, wc72, n_2365);
  not gc72 (wc72, n_2366);
  and g3019 (n_2550, wc73, n_2371);
  not gc73 (wc73, n_2372);
  or g3020 (n_2782, wc74, n_2356);
  not gc74 (wc74, n_2780);
  or g3021 (n_2879, wc75, n_2364);
  not gc75 (wc75, n_2365);
  or g3022 (n_2880, wc76, n_2374);
  not gc76 (wc76, n_2369);
  or g3023 (n_2883, wc77, n_2370);
  not gc77 (wc77, n_2371);
  or g3024 (n_2979, wc78, n_2514);
  not gc78 (wc78, n_2515);
  and g3025 (n_2552, wc79, n_2377);
  not gc79 (wc79, n_2378);
  and g3026 (n_2629, wc80, n_2509);
  not gc80 (wc80, n_2510);
  and g3027 (n_2634, wc81, n_2515);
  not gc81 (wc81, n_2516);
  and g3028 (n_2546, wc82, n_2542);
  not gc82 (wc82, n_2543);
  or g3029 (n_2784, wc83, n_2362);
  not gc83 (wc83, n_2688);
  or g3030 (n_2884, wc84, n_2380);
  not gc84 (wc84, n_2375);
  or g3031 (n_2887, wc85, n_2376);
  not gc85 (wc85, n_2377);
  or g3032 (n_2972, wc86, n_2512);
  not gc86 (wc86, n_2507);
  or g3033 (n_2975, wc87, n_2508);
  not gc87 (wc87, n_2509);
  or g3034 (n_2976, wc88, n_2518);
  not gc88 (wc88, n_2513);
  and g3035 (n_2557, wc89, n_2383);
  not gc89 (wc89, n_2384);
  and g3036 (n_2559, wc90, n_2389);
  not gc90 (wc90, n_2390);
  and g3037 (n_2646, wc91, n_2545);
  not gc91 (wc91, n_2546);
  and g3038 (n_2553, wc92, n_2549);
  not gc92 (wc92, n_2550);
  and g3039 (n_2637, wc93, n_2633);
  not gc93 (wc93, n_2634);
  or g3040 (n_2734, wc94, n_2650);
  not gc94 (wc94, n_2688);
  or g3041 (n_2888, wc95, n_2386);
  not gc95 (wc95, n_2381);
  or g3042 (n_2891, wc96, n_2382);
  not gc96 (wc96, n_2383);
  or g3043 (n_2892, wc97, n_2392);
  not gc97 (wc97, n_2387);
  or g3044 (n_2895, wc98, n_2388);
  not gc98 (wc98, n_2389);
  or g3045 (n_2896, wc99, n_2398);
  not gc99 (wc99, n_2393);
  or g3046 (n_2971, wc100, n_2502);
  not gc100 (wc100, n_2503);
  and g3047 (n_2564, wc101, n_2395);
  not gc101 (wc101, n_2396);
  and g3048 (n_2627, wc102, n_2503);
  not gc102 (wc102, n_2504);
  and g3049 (n_2647, wc103, n_2552);
  not gc103 (wc103, n_2553);
  and g3050 (n_2560, wc104, n_2556);
  not gc104 (wc104, n_2557);
  and g3051 (n_2683, wc105, n_2636);
  not gc105 (wc105, n_2637);
  or g3052 (n_2787, wc106, n_2368);
  not gc106 (wc106, n_2785);
  or g3053 (n_2899, wc107, n_2394);
  not gc107 (wc107, n_2395);
  or g3054 (n_2900, wc108, n_2404);
  not gc108 (wc108, n_2399);
  or g3055 (n_2967, wc109, n_2496);
  not gc109 (wc109, n_2497);
  or g3056 (n_2968, wc110, n_2506);
  not gc110 (wc110, n_2501);
  and g3057 (n_2566, wc111, n_2401);
  not gc111 (wc111, n_2402);
  and g3058 (n_2571, wc112, n_2407);
  not gc112 (wc112, n_2408);
  and g3059 (n_2573, wc113, n_2413);
  not gc113 (wc113, n_2414);
  and g3060 (n_2578, wc114, n_2419);
  not gc114 (wc114, n_2420);
  and g3061 (n_2580, wc115, n_2425);
  not gc115 (wc115, n_2426);
  and g3062 (n_2585, wc116, n_2431);
  not gc116 (wc116, n_2432);
  and g3063 (n_2587, wc117, n_2437);
  not gc117 (wc117, n_2438);
  and g3064 (n_2592, wc118, n_2443);
  not gc118 (wc118, n_2444);
  and g3065 (n_2594, wc119, n_2449);
  not gc119 (wc119, n_2450);
  and g3066 (n_2599, wc120, n_2455);
  not gc120 (wc120, n_2456);
  and g3067 (n_2601, wc121, n_2461);
  not gc121 (wc121, n_2462);
  and g3068 (n_2606, wc122, n_2467);
  not gc122 (wc122, n_2468);
  and g3069 (n_2608, wc123, n_2473);
  not gc123 (wc123, n_2474);
  and g3070 (n_2652, wc124, n_2559);
  not gc124 (wc124, n_2560);
  and g3071 (n_2630, wc125, n_2626);
  not gc125 (wc125, n_2627);
  or g3072 (n_2789, wc126, n_2374);
  not gc126 (wc126, n_2752);
  or g3073 (n_2903, wc127, n_2400);
  not gc127 (wc127, n_2401);
  or g3074 (n_2904, wc128, n_2410);
  not gc128 (wc128, n_2405);
  or g3075 (n_2907, wc129, n_2406);
  not gc129 (wc129, n_2407);
  or g3076 (n_2908, wc130, n_2416);
  not gc130 (wc130, n_2411);
  or g3077 (n_2911, wc131, n_2412);
  not gc131 (wc131, n_2413);
  or g3078 (n_2912, wc132, n_2422);
  not gc132 (wc132, n_2417);
  or g3079 (n_2915, wc133, n_2418);
  not gc133 (wc133, n_2419);
  or g3080 (n_2916, wc134, n_2428);
  not gc134 (wc134, n_2423);
  or g3081 (n_2919, wc135, n_2424);
  not gc135 (wc135, n_2425);
  or g3082 (n_2920, wc136, n_2434);
  not gc136 (wc136, n_2429);
  or g3083 (n_2923, wc137, n_2430);
  not gc137 (wc137, n_2431);
  or g3084 (n_2924, wc138, n_2440);
  not gc138 (wc138, n_2435);
  or g3085 (n_2927, wc139, n_2436);
  not gc139 (wc139, n_2437);
  or g3086 (n_2928, wc140, n_2446);
  not gc140 (wc140, n_2441);
  or g3087 (n_2931, wc141, n_2442);
  not gc141 (wc141, n_2443);
  or g3088 (n_2932, wc142, n_2452);
  not gc142 (wc142, n_2447);
  or g3089 (n_2935, wc143, n_2448);
  not gc143 (wc143, n_2449);
  or g3090 (n_2936, wc144, n_2458);
  not gc144 (wc144, n_2453);
  or g3091 (n_2939, wc145, n_2454);
  not gc145 (wc145, n_2455);
  or g3092 (n_2940, wc146, n_2464);
  not gc146 (wc146, n_2459);
  or g3093 (n_2943, wc147, n_2460);
  not gc147 (wc147, n_2461);
  or g3094 (n_2944, wc148, n_2470);
  not gc148 (wc148, n_2465);
  or g3095 (n_2947, wc149, n_2466);
  not gc149 (wc149, n_2467);
  or g3096 (n_2948, wc150, n_2476);
  not gc150 (wc150, n_2471);
  or g3097 (n_2951, wc151, n_2472);
  not gc151 (wc151, n_2473);
  or g3098 (n_2952, wc152, n_2482);
  not gc152 (wc152, n_2477);
  and g3099 (n_2613, wc153, n_2479);
  not gc153 (wc153, n_2480);
  and g3100 (n_2622, wc154, n_2497);
  not gc154 (wc154, n_2498);
  and g3101 (n_2567, wc155, n_2563);
  not gc155 (wc155, n_2564);
  and g3102 (n_2574, wc156, n_2570);
  not gc156 (wc156, n_2571);
  and g3103 (n_2581, wc157, n_2577);
  not gc157 (wc157, n_2578);
  and g3104 (n_2588, wc158, n_2584);
  not gc158 (wc158, n_2585);
  and g3105 (n_2595, wc159, n_2591);
  not gc159 (wc159, n_2592);
  and g3106 (n_2602, wc160, n_2598);
  not gc160 (wc160, n_2599);
  and g3107 (n_2609, wc161, n_2605);
  not gc161 (wc161, n_2606);
  and g3108 (n_2682, wc162, n_2629);
  not gc162 (wc162, n_2630);
  and g3109 (n_2689, n_2647, wc163);
  not gc163 (wc163, n_2648);
  or g3110 (n_2955, wc164, n_2478);
  not gc164 (wc164, n_2479);
  or g3111 (n_2956, wc165, n_2488);
  not gc165 (wc165, n_2483);
  or g3112 (n_2963, wc166, n_2490);
  not gc166 (wc166, n_2491);
  or g3113 (n_2964, wc167, n_2500);
  not gc167 (wc167, n_2495);
  and g3114 (n_2615, wc168, n_2485);
  not gc168 (wc168, n_2486);
  and g3115 (n_2620, wc169, n_2491);
  not gc169 (wc169, n_2492);
  and g3116 (n_2653, wc170, n_2566);
  not gc170 (wc170, n_2567);
  and g3117 (n_2658, wc171, n_2573);
  not gc171 (wc171, n_2574);
  and g3118 (n_2659, wc172, n_2580);
  not gc172 (wc172, n_2581);
  and g3119 (n_2664, wc173, n_2587);
  not gc173 (wc173, n_2588);
  and g3120 (n_2665, wc174, n_2594);
  not gc174 (wc174, n_2595);
  and g3121 (n_2670, wc175, n_2601);
  not gc175 (wc175, n_2602);
  and g3122 (n_2671, wc176, n_2608);
  not gc176 (wc176, n_2609);
  or g3123 (n_2792, wc177, n_2380);
  not gc177 (wc177, n_2790);
  or g3124 (n_2959, wc178, n_2484);
  not gc178 (wc178, n_2485);
  or g3125 (n_2960, wc179, n_2494);
  not gc179 (wc179, n_2489);
  and g3126 (n_2616, wc180, n_2612);
  not gc180 (wc180, n_2613);
  and g3127 (n_2623, wc181, n_2619);
  not gc181 (wc181, n_2620);
  and g3128 (n_2708, n_2683, wc182);
  not gc182 (wc182, n_2684);
  or g3129 (n_2736, wc183, n_2656);
  not gc183 (wc183, n_2713);
  or g3130 (n_2794, wc184, n_2386);
  not gc184 (wc184, n_2713);
  and g3131 (n_2676, wc185, n_2615);
  not gc185 (wc185, n_2616);
  and g3132 (n_2677, wc186, n_2622);
  not gc186 (wc186, n_2623);
  and g3133 (n_2692, n_2653, wc187);
  not gc187 (wc187, n_2654);
  and g3134 (n_2694, n_2659, wc188);
  not gc188 (wc188, n_2660);
  and g3135 (n_2699, n_2665, wc189);
  not gc189 (wc189, n_2666);
  and g3136 (n_2701, n_2671, wc190);
  not gc190 (wc190, n_2672);
  or g3137 (n_2716, n_2712, wc191);
  not gc191 (wc191, n_2713);
  and g3138 (n_2695, wc192, n_2691);
  not gc192 (wc192, n_2692);
  and g3139 (n_2702, wc193, n_2698);
  not gc193 (wc193, n_2699);
  or g3140 (n_2797, wc194, n_2392);
  not gc194 (wc194, n_2795);
  or g3141 (n_2799, wc195, n_2398);
  not gc195 (wc195, n_2755);
  and g3142 (n_2706, n_2677, wc196);
  not gc196 (wc196, n_2678);
  and g3143 (n_2715, wc197, n_2694);
  not gc197 (wc197, n_2695);
  and g3144 (n_2718, wc198, n_2701);
  not gc198 (wc198, n_2702);
  or g3145 (n_2739, wc199, n_2662);
  not gc199 (wc199, n_2737);
  or g3146 (n_2804, wc200, n_2410);
  not gc200 (wc200, n_2737);
  and g3147 (n_2709, wc201, n_2705);
  not gc201 (wc201, n_2706);
  or g3148 (n_2802, wc202, n_2404);
  not gc202 (wc202, n_2800);
  and g3149 (n_2719, wc203, n_2708);
  not gc203 (wc203, n_2709);
  or g3150 (n_2728, wc204, n_2722);
  not gc204 (wc204, n_2724);
  or g3151 (n_2741, wc205, n_2668);
  not gc205 (wc205, n_2724);
  or g3152 (n_2807, wc206, n_2416);
  not gc206 (wc206, n_2805);
  or g3153 (n_2809, wc207, n_2422);
  not gc207 (wc207, n_2758);
  or g3154 (n_2814, wc208, n_2434);
  not gc208 (wc208, n_2724);
  and g3155 (n_2725, n_2719, wc209);
  not gc209 (wc209, n_2720);
  or g3156 (n_2744, wc210, n_2674);
  not gc210 (wc210, n_2742);
  or g3157 (n_2746, wc211, n_2680);
  not gc211 (wc211, n_2731);
  or g3158 (n_2812, wc212, n_2428);
  not gc212 (wc212, n_2810);
  or g3159 (n_2817, wc213, n_2440);
  not gc213 (wc213, n_2815);
  or g3160 (n_2819, wc214, n_2446);
  not gc214 (wc214, n_2761);
  or g3161 (n_2824, wc215, n_2458);
  not gc215 (wc215, n_2742);
  or g3162 (n_2834, wc216, n_2482);
  not gc216 (wc216, n_2731);
  or g3163 (n_2749, wc217, n_2686);
  not gc217 (wc217, n_2747);
  or g3164 (n_2822, wc218, n_2452);
  not gc218 (wc218, n_2820);
  or g3165 (n_2827, wc219, n_2464);
  not gc219 (wc219, n_2825);
  or g3166 (n_2829, wc220, n_2470);
  not gc220 (wc220, n_2764);
  or g3167 (n_2837, wc221, n_2488);
  not gc221 (wc221, n_2835);
  or g3168 (n_2839, wc222, n_2494);
  not gc222 (wc222, n_2767);
  or g3169 (n_2844, wc223, n_2506);
  not gc223 (wc223, n_2747);
  or g3170 (n_2854, n_2530, wc224);
  not gc224 (wc224, n_2773);
  or g3171 (n_2832, wc225, n_2476);
  not gc225 (wc225, n_2830);
  or g3172 (n_2842, wc226, n_2500);
  not gc226 (wc226, n_2840);
  or g3173 (n_2847, wc227, n_2512);
  not gc227 (wc227, n_2845);
  or g3174 (n_2849, wc228, n_2518);
  not gc228 (wc228, n_2770);
  not g3175 (Z[66], n_2856);
  or g3176 (n_2852, wc229, n_2524);
  not gc229 (wc229, n_2850);
endmodule

module mult_signed_const_10729_GENERIC(A, Z);
  input [47:0] A;
  output [66:0] Z;
  wire [47:0] A;
  wire [66:0] Z;
  mult_signed_const_10729_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_11124_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [49:0] A;
  output [68:0] Z;
  wire [49:0] A;
  wire [68:0] Z;
  wire n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61;
  wire n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69;
  wire n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85;
  wire n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93;
  wire n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101;
  wire n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109;
  wire n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117;
  wire n_118, n_119, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_265, n_266, n_267, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_279;
  wire n_280, n_281, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_311;
  wire n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367;
  wire n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560;
  wire n_561, n_562, n_563, n_564, n_565, n_566, n_567, n_568;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_577, n_578, n_579, n_580, n_581, n_582, n_583, n_584;
  wire n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592;
  wire n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600;
  wire n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608;
  wire n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616;
  wire n_617, n_618, n_619, n_620, n_621, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_643, n_644, n_645, n_646, n_647, n_648;
  wire n_649, n_650, n_651, n_652, n_653, n_654, n_655, n_656;
  wire n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664;
  wire n_665, n_666, n_667, n_668, n_669, n_670, n_671, n_672;
  wire n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680;
  wire n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_691, n_692, n_693, n_694, n_695, n_696;
  wire n_697, n_698, n_699, n_700, n_701, n_702, n_703, n_704;
  wire n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736;
  wire n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_755, n_756, n_757, n_758, n_759, n_760;
  wire n_761, n_762, n_765, n_766, n_767, n_768, n_769, n_770;
  wire n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778;
  wire n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789;
  wire n_790, n_791, n_792, n_793, n_794, n_795, n_797, n_798;
  wire n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806;
  wire n_807, n_808, n_809, n_810, n_813, n_814, n_815, n_816;
  wire n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824;
  wire n_825, n_827, n_828, n_830, n_831, n_832, n_833, n_834;
  wire n_835, n_836, n_837, n_838, n_842, n_843, n_844, n_845;
  wire n_846, n_847, n_848, n_849, n_850, n_851, n_853, n_854;
  wire n_857, n_858, n_859, n_860, n_861, n_862, n_867, n_868;
  wire n_869, n_870, n_871, n_872, n_873, n_875, n_878, n_879;
  wire n_880, n_881, n_882, n_888, n_889, n_890, n_891, n_895;
  wire n_896, n_897, n_898, n_902, n_903, n_904, n_905, n_907;
  wire n_909, n_910, n_914, n_915, n_917, n_918, n_921, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932;
  wire n_933, n_934, n_936, n_937, n_938, n_939, n_943, n_944;
  wire n_945, n_946, n_947, n_948, n_949, n_950, n_952, n_954;
  wire n_955, n_956, n_957, n_958, n_959, n_960, n_962, n_964;
  wire n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_974;
  wire n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983;
  wire n_984, n_985, n_986, n_987, n_990, n_994, n_995, n_996;
  wire n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004;
  wire n_1005, n_1008, n_1009, n_1010, n_1012, n_1013, n_1014, n_1015;
  wire n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023;
  wire n_1024, n_1025, n_1026, n_1028, n_1029, n_1031, n_1032, n_1033;
  wire n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041;
  wire n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049;
  wire n_1051, n_1052, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059;
  wire n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067;
  wire n_1068, n_1071, n_1072, n_1073, n_1074, n_1076, n_1077, n_1078;
  wire n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086;
  wire n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094;
  wire n_1100, n_1101, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109;
  wire n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117;
  wire n_1118, n_1119, n_1120, n_1121, n_1123, n_1124, n_1126, n_1127;
  wire n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137;
  wire n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145;
  wire n_1146, n_1147, n_1148, n_1149, n_1150, n_1154, n_1155, n_1156;
  wire n_1157, n_1158, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165;
  wire n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173;
  wire n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181;
  wire n_1182, n_1183, n_1188, n_1189, n_1190, n_1192, n_1193, n_1194;
  wire n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202;
  wire n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210;
  wire n_1211, n_1212, n_1213, n_1214, n_1215, n_1220, n_1222, n_1224;
  wire n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240;
  wire n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1250;
  wire n_1251, n_1252, n_1253, n_1254, n_1256, n_1257, n_1258, n_1259;
  wire n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267;
  wire n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275;
  wire n_1276, n_1277, n_1278, n_1279, n_1282, n_1284, n_1285, n_1288;
  wire n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304;
  wire n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1314;
  wire n_1316, n_1317, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325;
  wire n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333;
  wire n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341;
  wire n_1342, n_1343, n_1344, n_1346, n_1348, n_1349, n_1352, n_1353;
  wire n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361;
  wire n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369;
  wire n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1378, n_1380;
  wire n_1381, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390;
  wire n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398;
  wire n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406;
  wire n_1407, n_1408, n_1409, n_1410, n_1412, n_1413, n_1416, n_1417;
  wire n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425;
  wire n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433;
  wire n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1442, n_1444;
  wire n_1445, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454;
  wire n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462;
  wire n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470;
  wire n_1471, n_1472, n_1474, n_1476, n_1477, n_1480, n_1481, n_1482;
  wire n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490;
  wire n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498;
  wire n_1499, n_1500, n_1501, n_1502, n_1503, n_1506, n_1508, n_1509;
  wire n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519;
  wire n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527;
  wire n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535;
  wire n_1536, n_1538, n_1540, n_1541, n_1544, n_1545, n_1546, n_1547;
  wire n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555;
  wire n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563;
  wire n_1564, n_1565, n_1566, n_1567, n_1570, n_1572, n_1573, n_1576;
  wire n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584;
  wire n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592;
  wire n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600;
  wire n_1601, n_1602, n_1604, n_1605, n_1608, n_1609, n_1610, n_1611;
  wire n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619;
  wire n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627;
  wire n_1628, n_1629, n_1630, n_1631, n_1634, n_1636, n_1637, n_1640;
  wire n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648;
  wire n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656;
  wire n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1666;
  wire n_1668, n_1669, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677;
  wire n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685;
  wire n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693;
  wire n_1694, n_1695, n_1698, n_1700, n_1701, n_1704, n_1705, n_1706;
  wire n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714;
  wire n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722;
  wire n_1723, n_1724, n_1725, n_1726, n_1727, n_1730, n_1732, n_1733;
  wire n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743;
  wire n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751;
  wire n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759;
  wire n_1762, n_1764, n_1765, n_1768, n_1769, n_1770, n_1771, n_1772;
  wire n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780;
  wire n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788;
  wire n_1789, n_1790, n_1791, n_1794, n_1796, n_1797, n_1800, n_1801;
  wire n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809;
  wire n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817;
  wire n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1826, n_1828;
  wire n_1829, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838;
  wire n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846;
  wire n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854;
  wire n_1855, n_1858, n_1860, n_1861, n_1864, n_1865, n_1866, n_1867;
  wire n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875;
  wire n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883;
  wire n_1884, n_1885, n_1886, n_1887, n_1890, n_1892, n_1893, n_1896;
  wire n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904;
  wire n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912;
  wire n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1922;
  wire n_1924, n_1925, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933;
  wire n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941;
  wire n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949;
  wire n_1950, n_1951, n_1954, n_1956, n_1957, n_1960, n_1961, n_1962;
  wire n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970;
  wire n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978;
  wire n_1979, n_1980, n_1981, n_1982, n_1983, n_1986, n_1988, n_1989;
  wire n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999;
  wire n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007;
  wire n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015;
  wire n_2018, n_2020, n_2021, n_2024, n_2025, n_2026, n_2027, n_2028;
  wire n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036;
  wire n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044;
  wire n_2045, n_2046, n_2047, n_2050, n_2052, n_2053, n_2056, n_2057;
  wire n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065;
  wire n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073;
  wire n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2082, n_2084;
  wire n_2085, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094;
  wire n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102;
  wire n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110;
  wire n_2111, n_2112, n_2113, n_2114, n_2116, n_2120, n_2121, n_2122;
  wire n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130;
  wire n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138;
  wire n_2139, n_2140, n_2141, n_2143, n_2144, n_2145, n_2146, n_2147;
  wire n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158;
  wire n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166;
  wire n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174;
  wire n_2175, n_2178, n_2180, n_2181, n_2183, n_2184, n_2185, n_2186;
  wire n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194;
  wire n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202;
  wire n_2203, n_2204, n_2205, n_2208, n_2212, n_2213, n_2214, n_2215;
  wire n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223;
  wire n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231;
  wire n_2236, n_2239, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247;
  wire n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255;
  wire n_2256, n_2257, n_2258, n_2259, n_2260, n_2264, n_2267, n_2268;
  wire n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277;
  wire n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2292, n_2294;
  wire n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302;
  wire n_2303, n_2304, n_2305, n_2306, n_2307, n_2314, n_2315, n_2316;
  wire n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324;
  wire n_2325, n_2326, n_2327, n_2336, n_2337, n_2338, n_2339, n_2340;
  wire n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2354;
  wire n_2355, n_2356, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363;
  wire n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377;
  wire n_2378, n_2379, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391;
  wire n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403;
  wire n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2416, n_2417;
  wire n_2418, n_2419, n_2421, n_2422, n_2423, n_2426, n_2427, n_2439;
  wire n_2441, n_2443, n_2444, n_2445, n_2446, n_2447, n_2449, n_2450;
  wire n_2451, n_2452, n_2453, n_2455, n_2456, n_2457, n_2458, n_2459;
  wire n_2461, n_2462, n_2463, n_2464, n_2465, n_2467, n_2468, n_2469;
  wire n_2470, n_2471, n_2473, n_2474, n_2475, n_2476, n_2477, n_2479;
  wire n_2480, n_2481, n_2482, n_2483, n_2485, n_2486, n_2487, n_2488;
  wire n_2489, n_2491, n_2492, n_2493, n_2494, n_2495, n_2497, n_2498;
  wire n_2499, n_2500, n_2501, n_2503, n_2504, n_2505, n_2506, n_2507;
  wire n_2509, n_2510, n_2511, n_2512, n_2513, n_2515, n_2516, n_2517;
  wire n_2518, n_2519, n_2521, n_2522, n_2523, n_2524, n_2525, n_2527;
  wire n_2528, n_2529, n_2530, n_2531, n_2533, n_2534, n_2535, n_2536;
  wire n_2537, n_2539, n_2540, n_2541, n_2542, n_2543, n_2545, n_2546;
  wire n_2547, n_2548, n_2549, n_2551, n_2552, n_2553, n_2554, n_2555;
  wire n_2557, n_2558, n_2559, n_2560, n_2561, n_2563, n_2564, n_2565;
  wire n_2566, n_2567, n_2569, n_2570, n_2571, n_2572, n_2573, n_2575;
  wire n_2576, n_2577, n_2578, n_2579, n_2581, n_2582, n_2583, n_2584;
  wire n_2585, n_2587, n_2588, n_2589, n_2590, n_2591, n_2593, n_2594;
  wire n_2595, n_2596, n_2597, n_2599, n_2600, n_2601, n_2602, n_2603;
  wire n_2605, n_2606, n_2607, n_2608, n_2609, n_2611, n_2612, n_2613;
  wire n_2614, n_2615, n_2617, n_2618, n_2619, n_2620, n_2621, n_2623;
  wire n_2624, n_2625, n_2626, n_2627, n_2629, n_2630, n_2631, n_2632;
  wire n_2633, n_2635, n_2638, n_2640, n_2641, n_2643, n_2644, n_2646;
  wire n_2647, n_2648, n_2650, n_2651, n_2653, n_2654, n_2655, n_2657;
  wire n_2658, n_2660, n_2661, n_2662, n_2664, n_2665, n_2667, n_2668;
  wire n_2669, n_2671, n_2672, n_2674, n_2675, n_2676, n_2678, n_2679;
  wire n_2681, n_2682, n_2683, n_2685, n_2686, n_2688, n_2689, n_2690;
  wire n_2692, n_2693, n_2695, n_2696, n_2697, n_2699, n_2700, n_2702;
  wire n_2703, n_2704, n_2706, n_2707, n_2709, n_2710, n_2711, n_2713;
  wire n_2714, n_2716, n_2717, n_2718, n_2720, n_2721, n_2723, n_2724;
  wire n_2725, n_2727, n_2728, n_2730, n_2731, n_2732, n_2734, n_2735;
  wire n_2737, n_2738, n_2739, n_2741, n_2742, n_2744, n_2745, n_2746;
  wire n_2748, n_2749, n_2751, n_2752, n_2755, n_2756, n_2757, n_2758;
  wire n_2759, n_2760, n_2762, n_2763, n_2764, n_2765, n_2766, n_2768;
  wire n_2769, n_2770, n_2771, n_2772, n_2774, n_2775, n_2776, n_2777;
  wire n_2778, n_2780, n_2781, n_2782, n_2783, n_2784, n_2786, n_2787;
  wire n_2788, n_2789, n_2790, n_2792, n_2793, n_2794, n_2795, n_2796;
  wire n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2806;
  wire n_2807, n_2809, n_2810, n_2811, n_2813, n_2814, n_2816, n_2817;
  wire n_2818, n_2820, n_2821, n_2823, n_2824, n_2825, n_2827, n_2828;
  wire n_2829, n_2830, n_2831, n_2832, n_2834, n_2835, n_2836, n_2837;
  wire n_2838, n_2840, n_2841, n_2842, n_2843, n_2844, n_2846, n_2848;
  wire n_2849, n_2851, n_2853, n_2854, n_2856, n_2858, n_2859, n_2861;
  wire n_2862, n_2863, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870;
  wire n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878;
  wire n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886;
  wire n_2887, n_2888, n_2889, n_2893, n_2894, n_2896, n_2898, n_2899;
  wire n_2901, n_2903, n_2904, n_2906, n_2908, n_2909, n_2911, n_2913;
  wire n_2914, n_2916, n_2918, n_2919, n_2921, n_2923, n_2924, n_2926;
  wire n_2928, n_2929, n_2931, n_2933, n_2934, n_2936, n_2938, n_2939;
  wire n_2941, n_2943, n_2944, n_2946, n_2948, n_2949, n_2951, n_2953;
  wire n_2954, n_2956, n_2958, n_2959, n_2961, n_2963, n_2964, n_2966;
  wire n_2968, n_2969, n_2971, n_2973, n_2977, n_2980, n_2981, n_2983;
  wire n_2984, n_2985, n_2987, n_2988, n_2989, n_2991, n_2992, n_2993;
  wire n_2995, n_2996, n_2997, n_2999, n_3000, n_3001, n_3003, n_3004;
  wire n_3005, n_3007, n_3008, n_3009, n_3011, n_3012, n_3013, n_3015;
  wire n_3016, n_3017, n_3019, n_3020, n_3021, n_3023, n_3024, n_3025;
  wire n_3027, n_3028, n_3029, n_3031, n_3032, n_3033, n_3035, n_3036;
  wire n_3037, n_3039, n_3040, n_3041, n_3043, n_3044, n_3045, n_3047;
  wire n_3048, n_3049, n_3051, n_3052, n_3053, n_3055, n_3056, n_3057;
  wire n_3059, n_3060, n_3061, n_3063, n_3064, n_3065, n_3067, n_3068;
  wire n_3069, n_3071, n_3072, n_3073, n_3075, n_3076, n_3077, n_3079;
  wire n_3080, n_3081, n_3083, n_3084, n_3085, n_3087, n_3088, n_3089;
  wire n_3091, n_3092, n_3093, n_3095, n_3096, n_3097, n_3099, n_3100;
  wire n_3101, n_3103, n_3104, n_3105, n_3107, n_3108;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g396 (n_184, A[4], A[0]);
  and g2 (n_114, A[4], A[0]);
  xor g397 (n_924, A[1], A[3]);
  xor g398 (n_183, n_924, A[5]);
  nand g3 (n_925, A[1], A[3]);
  nand g399 (n_926, A[5], A[3]);
  nand g400 (n_927, A[1], A[5]);
  nand g401 (n_113, n_925, n_926, n_927);
  xor g402 (n_259, A[6], A[4]);
  and g403 (n_260, A[6], A[4]);
  xor g404 (n_928, A[0], A[2]);
  xor g405 (n_182, n_928, n_259);
  nand g406 (n_929, A[0], A[2]);
  nand g4 (n_930, n_259, A[2]);
  nand g5 (n_931, A[0], n_259);
  nand g407 (n_112, n_929, n_930, n_931);
  xor g408 (n_932, A[1], A[7]);
  xor g409 (n_261, n_932, A[5]);
  nand g410 (n_933, A[1], A[7]);
  nand g411 (n_934, A[5], A[7]);
  nand g6 (n_263, n_933, n_934, n_927);
  xor g413 (n_936, A[3], n_260);
  xor g414 (n_181, n_936, n_261);
  nand g415 (n_937, A[3], n_260);
  nand g416 (n_938, n_261, n_260);
  nand g417 (n_939, A[3], n_261);
  nand g418 (n_111, n_937, n_938, n_939);
  xor g419 (n_262, A[8], A[6]);
  and g420 (n_265, A[8], A[6]);
  xor g422 (n_264, n_928, A[4]);
  nand g425 (n_943, A[2], A[4]);
  xor g427 (n_944, n_262, n_263);
  xor g428 (n_180, n_944, n_264);
  nand g429 (n_945, n_262, n_263);
  nand g430 (n_946, n_264, n_263);
  nand g431 (n_947, n_262, n_264);
  nand g432 (n_110, n_945, n_946, n_947);
  xor g433 (n_948, A[1], A[9]);
  xor g434 (n_267, n_948, A[3]);
  nand g435 (n_949, A[1], A[9]);
  nand g436 (n_950, A[3], A[9]);
  nand g438 (n_270, n_949, n_950, n_925);
  xor g439 (n_952, A[7], A[5]);
  xor g440 (n_268, n_952, n_265);
  nand g442 (n_954, n_265, A[5]);
  nand g443 (n_955, A[7], n_265);
  nand g444 (n_272, n_934, n_954, n_955);
  xor g445 (n_956, n_266, n_267);
  xor g446 (n_179, n_956, n_268);
  nand g447 (n_957, n_266, n_267);
  nand g448 (n_958, n_268, n_267);
  nand g449 (n_959, n_266, n_268);
  nand g450 (n_109, n_957, n_958, n_959);
  xor g451 (n_269, A[10], A[8]);
  and g452 (n_274, A[10], A[8]);
  xor g453 (n_960, A[4], A[2]);
  xor g454 (n_271, n_960, A[6]);
  nand g456 (n_962, A[6], A[2]);
  xor g459 (n_964, A[0], n_269);
  xor g460 (n_273, n_964, n_270);
  nand g461 (n_965, A[0], n_269);
  nand g462 (n_966, n_270, n_269);
  nand g463 (n_967, A[0], n_270);
  nand g464 (n_278, n_965, n_966, n_967);
  xor g465 (n_968, n_271, n_272);
  xor g466 (n_178, n_968, n_273);
  nand g467 (n_969, n_271, n_272);
  nand g468 (n_970, n_273, n_272);
  nand g469 (n_971, n_271, n_273);
  nand g470 (n_108, n_969, n_970, n_971);
  xor g472 (n_276, n_948, A[5]);
  nand g474 (n_974, A[5], A[9]);
  nand g476 (n_281, n_949, n_974, n_927);
  xor g477 (n_976, A[3], A[11]);
  xor g478 (n_277, n_976, A[7]);
  nand g479 (n_977, A[3], A[11]);
  nand g480 (n_978, A[7], A[11]);
  nand g481 (n_979, A[3], A[7]);
  nand g482 (n_282, n_977, n_978, n_979);
  xor g483 (n_980, n_274, n_275);
  xor g484 (n_279, n_980, n_276);
  nand g485 (n_981, n_274, n_275);
  nand g486 (n_982, n_276, n_275);
  nand g487 (n_983, n_274, n_276);
  nand g488 (n_286, n_981, n_982, n_983);
  xor g489 (n_984, n_277, n_278);
  xor g490 (n_177, n_984, n_279);
  nand g491 (n_985, n_277, n_278);
  nand g492 (n_986, n_279, n_278);
  nand g493 (n_987, n_277, n_279);
  nand g494 (n_107, n_985, n_986, n_987);
  xor g495 (n_280, A[12], A[10]);
  and g496 (n_287, A[12], A[10]);
  xor g498 (n_283, n_259, A[8]);
  nand g500 (n_990, A[8], A[4]);
  xor g504 (n_284, n_928, n_280);
  nand g506 (n_994, n_280, A[0]);
  nand g507 (n_995, A[2], n_280);
  nand g508 (n_291, n_929, n_994, n_995);
  xor g509 (n_996, n_281, n_282);
  xor g510 (n_285, n_996, n_283);
  nand g511 (n_997, n_281, n_282);
  nand g512 (n_998, n_283, n_282);
  nand g513 (n_999, n_281, n_283);
  nand g514 (n_293, n_997, n_998, n_999);
  xor g515 (n_1000, n_284, n_285);
  xor g516 (n_176, n_1000, n_286);
  nand g517 (n_1001, n_284, n_285);
  nand g518 (n_1002, n_286, n_285);
  nand g519 (n_1003, n_284, n_286);
  nand g520 (n_106, n_1001, n_1002, n_1003);
  xor g521 (n_1004, A[1], A[11]);
  xor g522 (n_290, n_1004, A[7]);
  nand g523 (n_1005, A[1], A[11]);
  nand g526 (n_296, n_1005, n_978, n_933);
  xor g527 (n_1008, A[5], A[13]);
  xor g528 (n_289, n_1008, A[3]);
  nand g529 (n_1009, A[5], A[13]);
  nand g530 (n_1010, A[3], A[13]);
  nand g532 (n_297, n_1009, n_1010, n_926);
  xor g533 (n_1012, A[9], n_287);
  xor g534 (n_292, n_1012, n_288);
  nand g535 (n_1013, A[9], n_287);
  nand g536 (n_1014, n_288, n_287);
  nand g537 (n_1015, A[9], n_288);
  nand g538 (n_300, n_1013, n_1014, n_1015);
  xor g539 (n_1016, n_289, n_290);
  xor g540 (n_294, n_1016, n_291);
  nand g541 (n_1017, n_289, n_290);
  nand g542 (n_1018, n_291, n_290);
  nand g543 (n_1019, n_289, n_291);
  nand g544 (n_302, n_1017, n_1018, n_1019);
  xor g545 (n_1020, n_292, n_293);
  xor g546 (n_175, n_1020, n_294);
  nand g547 (n_1021, n_292, n_293);
  nand g548 (n_1022, n_294, n_293);
  nand g549 (n_1023, n_292, n_294);
  nand g550 (n_105, n_1021, n_1022, n_1023);
  xor g551 (n_295, A[14], A[12]);
  and g552 (n_304, A[14], A[12]);
  xor g553 (n_1024, A[8], A[0]);
  xor g554 (n_299, n_1024, A[6]);
  nand g555 (n_1025, A[8], A[0]);
  nand g556 (n_1026, A[6], A[0]);
  xor g559 (n_1028, A[10], A[4]);
  xor g560 (n_298, n_1028, A[2]);
  nand g561 (n_1029, A[10], A[4]);
  nand g563 (n_1031, A[10], A[2]);
  nand g564 (n_306, n_1029, n_943, n_1031);
  xor g565 (n_1032, n_295, n_296);
  xor g566 (n_301, n_1032, n_297);
  nand g567 (n_1033, n_295, n_296);
  nand g568 (n_1034, n_297, n_296);
  nand g569 (n_1035, n_295, n_297);
  nand g570 (n_310, n_1033, n_1034, n_1035);
  xor g571 (n_1036, n_298, n_299);
  xor g572 (n_303, n_1036, n_300);
  nand g573 (n_1037, n_298, n_299);
  nand g574 (n_1038, n_300, n_299);
  nand g575 (n_1039, n_298, n_300);
  nand g576 (n_313, n_1037, n_1038, n_1039);
  xor g577 (n_1040, n_301, n_302);
  xor g578 (n_174, n_1040, n_303);
  nand g579 (n_1041, n_301, n_302);
  nand g580 (n_1042, n_303, n_302);
  nand g581 (n_1043, n_301, n_303);
  nand g582 (n_104, n_1041, n_1042, n_1043);
  xor g583 (n_1044, A[1], A[15]);
  xor g584 (n_307, n_1044, A[13]);
  nand g585 (n_1045, A[1], A[15]);
  nand g586 (n_1046, A[13], A[15]);
  nand g587 (n_1047, A[1], A[13]);
  nand g588 (n_315, n_1045, n_1046, n_1047);
  xor g589 (n_1048, A[9], A[7]);
  xor g590 (n_308, n_1048, A[11]);
  nand g591 (n_1049, A[9], A[7]);
  nand g593 (n_1051, A[9], A[11]);
  nand g594 (n_316, n_1049, n_978, n_1051);
  xor g595 (n_1052, A[5], A[3]);
  xor g596 (n_309, n_1052, n_304);
  nand g598 (n_1054, n_304, A[3]);
  nand g599 (n_1055, A[5], n_304);
  nand g600 (n_319, n_926, n_1054, n_1055);
  xor g601 (n_1056, n_305, n_306);
  xor g602 (n_311, n_1056, n_307);
  nand g603 (n_1057, n_305, n_306);
  nand g604 (n_1058, n_307, n_306);
  nand g605 (n_1059, n_305, n_307);
  nand g606 (n_321, n_1057, n_1058, n_1059);
  xor g607 (n_1060, n_308, n_309);
  xor g608 (n_312, n_1060, n_310);
  nand g609 (n_1061, n_308, n_309);
  nand g610 (n_1062, n_310, n_309);
  nand g611 (n_1063, n_308, n_310);
  nand g612 (n_323, n_1061, n_1062, n_1063);
  xor g613 (n_1064, n_311, n_312);
  xor g614 (n_173, n_1064, n_313);
  nand g615 (n_1065, n_311, n_312);
  nand g616 (n_1066, n_313, n_312);
  nand g617 (n_1067, n_311, n_313);
  nand g618 (n_103, n_1065, n_1066, n_1067);
  xor g619 (n_314, A[16], A[14]);
  and g620 (n_325, A[16], A[14]);
  xor g621 (n_1068, A[10], A[2]);
  xor g622 (n_318, n_1068, A[0]);
  nand g625 (n_1071, A[10], A[0]);
  nand g626 (n_326, n_1031, n_929, n_1071);
  xor g627 (n_1072, A[8], A[12]);
  xor g628 (n_317, n_1072, A[6]);
  nand g629 (n_1073, A[8], A[12]);
  nand g630 (n_1074, A[6], A[12]);
  xor g633 (n_1076, A[4], n_314);
  xor g634 (n_320, n_1076, n_315);
  nand g635 (n_1077, A[4], n_314);
  nand g636 (n_1078, n_315, n_314);
  nand g637 (n_1079, A[4], n_315);
  nand g638 (n_331, n_1077, n_1078, n_1079);
  xor g639 (n_1080, n_316, n_317);
  xor g640 (n_322, n_1080, n_318);
  nand g641 (n_1081, n_316, n_317);
  nand g642 (n_1082, n_318, n_317);
  nand g643 (n_1083, n_316, n_318);
  nand g644 (n_333, n_1081, n_1082, n_1083);
  xor g645 (n_1084, n_319, n_320);
  xor g646 (n_324, n_1084, n_321);
  nand g647 (n_1085, n_319, n_320);
  nand g648 (n_1086, n_321, n_320);
  nand g649 (n_1087, n_319, n_321);
  nand g650 (n_335, n_1085, n_1086, n_1087);
  xor g651 (n_1088, n_322, n_323);
  xor g652 (n_172, n_1088, n_324);
  nand g653 (n_1089, n_322, n_323);
  nand g654 (n_1090, n_324, n_323);
  nand g655 (n_1091, n_322, n_324);
  nand g656 (n_102, n_1089, n_1090, n_1091);
  xor g657 (n_1092, A[1], A[17]);
  xor g658 (n_329, n_1092, A[15]);
  nand g659 (n_1093, A[1], A[17]);
  nand g660 (n_1094, A[15], A[17]);
  nand g662 (n_338, n_1093, n_1094, n_1045);
  xor g664 (n_330, n_976, A[9]);
  nand g668 (n_340, n_977, n_1051, n_950);
  xor g669 (n_1100, A[13], A[7]);
  xor g670 (n_328, n_1100, A[5]);
  nand g671 (n_1101, A[13], A[7]);
  nand g674 (n_339, n_1101, n_934, n_1009);
  xor g675 (n_1104, n_325, n_326);
  xor g676 (n_332, n_1104, n_327);
  nand g677 (n_1105, n_325, n_326);
  nand g678 (n_1106, n_327, n_326);
  nand g679 (n_1107, n_325, n_327);
  nand g680 (n_344, n_1105, n_1106, n_1107);
  xor g681 (n_1108, n_328, n_329);
  xor g682 (n_334, n_1108, n_330);
  nand g683 (n_1109, n_328, n_329);
  nand g684 (n_1110, n_330, n_329);
  nand g685 (n_1111, n_328, n_330);
  nand g686 (n_346, n_1109, n_1110, n_1111);
  xor g687 (n_1112, n_331, n_332);
  xor g688 (n_336, n_1112, n_333);
  nand g689 (n_1113, n_331, n_332);
  nand g690 (n_1114, n_333, n_332);
  nand g691 (n_1115, n_331, n_333);
  nand g692 (n_348, n_1113, n_1114, n_1115);
  xor g693 (n_1116, n_334, n_335);
  xor g694 (n_171, n_1116, n_336);
  nand g695 (n_1117, n_334, n_335);
  nand g696 (n_1118, n_336, n_335);
  nand g697 (n_1119, n_334, n_336);
  nand g698 (n_101, n_1117, n_1118, n_1119);
  xor g699 (n_337, A[18], A[16]);
  and g700 (n_350, A[18], A[16]);
  xor g701 (n_1120, A[12], A[4]);
  xor g702 (n_341, n_1120, A[2]);
  nand g703 (n_1121, A[12], A[4]);
  nand g705 (n_1123, A[12], A[2]);
  nand g706 (n_351, n_1121, n_943, n_1123);
  xor g707 (n_1124, A[10], A[0]);
  xor g708 (n_342, n_1124, A[14]);
  nand g710 (n_1126, A[14], A[0]);
  nand g711 (n_1127, A[10], A[14]);
  nand g712 (n_115, n_1071, n_1126, n_1127);
  xor g714 (n_343, n_262, n_337);
  nand g716 (n_1130, n_337, A[6]);
  nand g717 (n_1131, A[8], n_337);
  xor g719 (n_1132, n_338, n_339);
  xor g720 (n_345, n_1132, n_340);
  nand g721 (n_1133, n_338, n_339);
  nand g722 (n_1134, n_340, n_339);
  nand g723 (n_1135, n_338, n_340);
  nand g724 (n_353, n_1133, n_1134, n_1135);
  xor g725 (n_1136, n_341, n_342);
  xor g726 (n_347, n_1136, n_343);
  nand g727 (n_1137, n_341, n_342);
  nand g728 (n_1138, n_343, n_342);
  nand g729 (n_1139, n_341, n_343);
  nand g730 (n_354, n_1137, n_1138, n_1139);
  xor g731 (n_1140, n_344, n_345);
  xor g732 (n_349, n_1140, n_346);
  nand g733 (n_1141, n_344, n_345);
  nand g734 (n_1142, n_346, n_345);
  nand g735 (n_1143, n_344, n_346);
  nand g736 (n_357, n_1141, n_1142, n_1143);
  xor g737 (n_1144, n_347, n_348);
  xor g738 (n_170, n_1144, n_349);
  nand g739 (n_1145, n_347, n_348);
  nand g740 (n_1146, n_349, n_348);
  nand g741 (n_1147, n_347, n_349);
  nand g742 (n_100, n_1145, n_1146, n_1147);
  xor g743 (n_1148, A[1], A[19]);
  xor g744 (n_117, n_1148, A[13]);
  nand g745 (n_1149, A[1], A[19]);
  nand g746 (n_1150, A[13], A[19]);
  nand g748 (n_359, n_1149, n_1150, n_1047);
  xor g750 (n_118, n_1052, A[17]);
  nand g752 (n_1154, A[17], A[3]);
  nand g753 (n_1155, A[5], A[17]);
  nand g754 (n_360, n_926, n_1154, n_1155);
  xor g755 (n_1156, A[11], A[15]);
  xor g756 (n_116, n_1156, A[9]);
  nand g757 (n_1157, A[11], A[15]);
  nand g758 (n_1158, A[9], A[15]);
  nand g760 (n_361, n_1157, n_1158, n_1051);
  xor g761 (n_1160, A[7], n_350);
  xor g762 (n_352, n_1160, n_351);
  nand g763 (n_1161, A[7], n_350);
  nand g764 (n_1162, n_351, n_350);
  nand g765 (n_1163, A[7], n_351);
  nand g766 (n_365, n_1161, n_1162, n_1163);
  xor g767 (n_1164, n_115, n_116);
  xor g768 (n_355, n_1164, n_117);
  nand g769 (n_1165, n_115, n_116);
  nand g770 (n_1166, n_117, n_116);
  nand g771 (n_1167, n_115, n_117);
  nand g772 (n_367, n_1165, n_1166, n_1167);
  xor g773 (n_1168, n_118, n_119);
  xor g774 (n_356, n_1168, n_352);
  nand g775 (n_1169, n_118, n_119);
  nand g776 (n_1170, n_352, n_119);
  nand g777 (n_1171, n_118, n_352);
  nand g778 (n_369, n_1169, n_1170, n_1171);
  xor g779 (n_1172, n_353, n_354);
  xor g780 (n_358, n_1172, n_355);
  nand g781 (n_1173, n_353, n_354);
  nand g782 (n_1174, n_355, n_354);
  nand g783 (n_1175, n_353, n_355);
  nand g784 (n_371, n_1173, n_1174, n_1175);
  xor g785 (n_1176, n_356, n_357);
  xor g786 (n_169, n_1176, n_358);
  nand g787 (n_1177, n_356, n_357);
  nand g788 (n_1178, n_358, n_357);
  nand g789 (n_1179, n_356, n_358);
  nand g790 (n_99, n_1177, n_1178, n_1179);
  xor g791 (n_1180, A[20], A[18]);
  xor g792 (n_363, n_1180, A[14]);
  nand g793 (n_1181, A[20], A[18]);
  nand g794 (n_1182, A[14], A[18]);
  nand g795 (n_1183, A[20], A[14]);
  nand g796 (n_373, n_1181, n_1182, n_1183);
  xor g798 (n_364, n_259, A[12]);
  xor g803 (n_1188, A[2], A[16]);
  xor g804 (n_362, n_1188, A[10]);
  nand g805 (n_1189, A[2], A[16]);
  nand g806 (n_1190, A[10], A[16]);
  nand g808 (n_375, n_1189, n_1190, n_1031);
  xor g809 (n_1192, A[8], n_359);
  xor g810 (n_366, n_1192, n_360);
  nand g811 (n_1193, A[8], n_359);
  nand g812 (n_1194, n_360, n_359);
  nand g813 (n_1195, A[8], n_360);
  nand g814 (n_379, n_1193, n_1194, n_1195);
  xor g815 (n_1196, n_361, n_362);
  xor g816 (n_368, n_1196, n_363);
  nand g817 (n_1197, n_361, n_362);
  nand g818 (n_1198, n_363, n_362);
  nand g819 (n_1199, n_361, n_363);
  nand g820 (n_381, n_1197, n_1198, n_1199);
  xor g821 (n_1200, n_364, n_365);
  xor g822 (n_370, n_1200, n_366);
  nand g823 (n_1201, n_364, n_365);
  nand g824 (n_1202, n_366, n_365);
  nand g825 (n_1203, n_364, n_366);
  nand g826 (n_383, n_1201, n_1202, n_1203);
  xor g827 (n_1204, n_367, n_368);
  xor g828 (n_372, n_1204, n_369);
  nand g829 (n_1205, n_367, n_368);
  nand g830 (n_1206, n_369, n_368);
  nand g831 (n_1207, n_367, n_369);
  nand g832 (n_385, n_1205, n_1206, n_1207);
  xor g833 (n_1208, n_370, n_371);
  xor g834 (n_168, n_1208, n_372);
  nand g835 (n_1209, n_370, n_371);
  nand g836 (n_1210, n_372, n_371);
  nand g837 (n_1211, n_370, n_372);
  nand g838 (n_98, n_1209, n_1210, n_1211);
  xor g839 (n_1212, A[21], A[19]);
  xor g840 (n_377, n_1212, A[15]);
  nand g841 (n_1213, A[21], A[19]);
  nand g842 (n_1214, A[15], A[19]);
  nand g843 (n_1215, A[21], A[15]);
  nand g844 (n_387, n_1213, n_1214, n_1215);
  xor g846 (n_378, n_952, A[13]);
  xor g851 (n_1220, A[3], A[17]);
  xor g852 (n_376, n_1220, A[11]);
  nand g854 (n_1222, A[11], A[17]);
  nand g856 (n_389, n_1154, n_1222, n_977);
  xor g857 (n_1224, A[9], n_373);
  xor g858 (n_380, n_1224, n_374);
  nand g859 (n_1225, A[9], n_373);
  nand g860 (n_1226, n_374, n_373);
  nand g861 (n_1227, A[9], n_374);
  nand g862 (n_393, n_1225, n_1226, n_1227);
  xor g863 (n_1228, n_375, n_376);
  xor g864 (n_382, n_1228, n_377);
  nand g865 (n_1229, n_375, n_376);
  nand g866 (n_1230, n_377, n_376);
  nand g867 (n_1231, n_375, n_377);
  nand g868 (n_395, n_1229, n_1230, n_1231);
  xor g869 (n_1232, n_378, n_379);
  xor g870 (n_384, n_1232, n_380);
  nand g871 (n_1233, n_378, n_379);
  nand g872 (n_1234, n_380, n_379);
  nand g873 (n_1235, n_378, n_380);
  nand g874 (n_397, n_1233, n_1234, n_1235);
  xor g875 (n_1236, n_381, n_382);
  xor g876 (n_386, n_1236, n_383);
  nand g877 (n_1237, n_381, n_382);
  nand g878 (n_1238, n_383, n_382);
  nand g879 (n_1239, n_381, n_383);
  nand g880 (n_400, n_1237, n_1238, n_1239);
  xor g881 (n_1240, n_384, n_385);
  xor g882 (n_167, n_1240, n_386);
  nand g883 (n_1241, n_384, n_385);
  nand g884 (n_1242, n_386, n_385);
  nand g885 (n_1243, n_384, n_386);
  nand g886 (n_97, n_1241, n_1242, n_1243);
  xor g887 (n_1244, A[22], A[20]);
  xor g888 (n_391, n_1244, A[16]);
  nand g889 (n_1245, A[22], A[20]);
  nand g890 (n_1246, A[16], A[20]);
  nand g891 (n_1247, A[22], A[16]);
  nand g892 (n_401, n_1245, n_1246, n_1247);
  xor g894 (n_392, n_262, A[14]);
  nand g896 (n_1250, A[14], A[6]);
  nand g897 (n_1251, A[8], A[14]);
  xor g899 (n_1252, A[4], A[18]);
  xor g900 (n_390, n_1252, A[12]);
  nand g901 (n_1253, A[4], A[18]);
  nand g902 (n_1254, A[12], A[18]);
  nand g904 (n_403, n_1253, n_1254, n_1121);
  xor g905 (n_1256, A[10], n_387);
  xor g906 (n_394, n_1256, n_339);
  nand g907 (n_1257, A[10], n_387);
  nand g908 (n_1258, n_339, n_387);
  nand g909 (n_1259, A[10], n_339);
  nand g910 (n_407, n_1257, n_1258, n_1259);
  xor g911 (n_1260, n_389, n_390);
  xor g912 (n_396, n_1260, n_391);
  nand g913 (n_1261, n_389, n_390);
  nand g914 (n_1262, n_391, n_390);
  nand g915 (n_1263, n_389, n_391);
  nand g916 (n_409, n_1261, n_1262, n_1263);
  xor g917 (n_1264, n_392, n_393);
  xor g918 (n_398, n_1264, n_394);
  nand g919 (n_1265, n_392, n_393);
  nand g920 (n_1266, n_394, n_393);
  nand g921 (n_1267, n_392, n_394);
  nand g922 (n_411, n_1265, n_1266, n_1267);
  xor g923 (n_1268, n_395, n_396);
  xor g924 (n_399, n_1268, n_397);
  nand g925 (n_1269, n_395, n_396);
  nand g926 (n_1270, n_397, n_396);
  nand g927 (n_1271, n_395, n_397);
  nand g928 (n_186, n_1269, n_1270, n_1271);
  xor g929 (n_1272, n_398, n_399);
  xor g930 (n_166, n_1272, n_400);
  nand g931 (n_1273, n_398, n_399);
  nand g932 (n_1274, n_400, n_399);
  nand g933 (n_1275, n_398, n_400);
  nand g934 (n_96, n_1273, n_1274, n_1275);
  xor g935 (n_1276, A[23], A[21]);
  xor g936 (n_405, n_1276, A[17]);
  nand g937 (n_1277, A[23], A[21]);
  nand g938 (n_1278, A[17], A[21]);
  nand g939 (n_1279, A[23], A[17]);
  nand g940 (n_413, n_1277, n_1278, n_1279);
  xor g942 (n_406, n_1048, A[15]);
  nand g944 (n_1282, A[15], A[7]);
  nand g946 (n_414, n_1049, n_1282, n_1158);
  xor g947 (n_1284, A[5], A[19]);
  xor g948 (n_404, n_1284, A[13]);
  nand g949 (n_1285, A[5], A[19]);
  nand g952 (n_415, n_1285, n_1150, n_1009);
  xor g953 (n_1288, A[11], n_401);
  xor g954 (n_408, n_1288, n_402);
  nand g955 (n_1289, A[11], n_401);
  nand g956 (n_1290, n_402, n_401);
  nand g957 (n_1291, A[11], n_402);
  nand g958 (n_419, n_1289, n_1290, n_1291);
  xor g959 (n_1292, n_403, n_404);
  xor g960 (n_410, n_1292, n_405);
  nand g961 (n_1293, n_403, n_404);
  nand g962 (n_1294, n_405, n_404);
  nand g963 (n_1295, n_403, n_405);
  nand g964 (n_421, n_1293, n_1294, n_1295);
  xor g965 (n_1296, n_406, n_407);
  xor g966 (n_412, n_1296, n_408);
  nand g967 (n_1297, n_406, n_407);
  nand g968 (n_1298, n_408, n_407);
  nand g969 (n_1299, n_406, n_408);
  nand g970 (n_423, n_1297, n_1298, n_1299);
  xor g971 (n_1300, n_409, n_410);
  xor g972 (n_185, n_1300, n_411);
  nand g973 (n_1301, n_409, n_410);
  nand g974 (n_1302, n_411, n_410);
  nand g975 (n_1303, n_409, n_411);
  nand g976 (n_426, n_1301, n_1302, n_1303);
  xor g977 (n_1304, n_412, n_185);
  xor g978 (n_165, n_1304, n_186);
  nand g979 (n_1305, n_412, n_185);
  nand g980 (n_1306, n_186, n_185);
  nand g981 (n_1307, n_412, n_186);
  nand g982 (n_95, n_1305, n_1306, n_1307);
  xor g983 (n_1308, A[24], A[22]);
  xor g984 (n_417, n_1308, A[18]);
  nand g985 (n_1309, A[24], A[22]);
  nand g986 (n_1310, A[18], A[22]);
  nand g987 (n_1311, A[24], A[18]);
  nand g988 (n_427, n_1309, n_1310, n_1311);
  xor g990 (n_418, n_269, A[16]);
  nand g992 (n_1314, A[16], A[8]);
  xor g995 (n_1316, A[6], A[20]);
  xor g996 (n_416, n_1316, A[14]);
  nand g997 (n_1317, A[6], A[20]);
  nand g1000 (n_429, n_1317, n_1183, n_1250);
  xor g1001 (n_1320, A[12], n_413);
  xor g1002 (n_420, n_1320, n_414);
  nand g1003 (n_1321, A[12], n_413);
  nand g1004 (n_1322, n_414, n_413);
  nand g1005 (n_1323, A[12], n_414);
  nand g1006 (n_433, n_1321, n_1322, n_1323);
  xor g1007 (n_1324, n_415, n_416);
  xor g1008 (n_422, n_1324, n_417);
  nand g1009 (n_1325, n_415, n_416);
  nand g1010 (n_1326, n_417, n_416);
  nand g1011 (n_1327, n_415, n_417);
  nand g1012 (n_435, n_1325, n_1326, n_1327);
  xor g1013 (n_1328, n_418, n_419);
  xor g1014 (n_424, n_1328, n_420);
  nand g1015 (n_1329, n_418, n_419);
  nand g1016 (n_1330, n_420, n_419);
  nand g1017 (n_1331, n_418, n_420);
  nand g1018 (n_437, n_1329, n_1330, n_1331);
  xor g1019 (n_1332, n_421, n_422);
  xor g1020 (n_425, n_1332, n_423);
  nand g1021 (n_1333, n_421, n_422);
  nand g1022 (n_1334, n_423, n_422);
  nand g1023 (n_1335, n_421, n_423);
  nand g1024 (n_440, n_1333, n_1334, n_1335);
  xor g1025 (n_1336, n_424, n_425);
  xor g1026 (n_164, n_1336, n_426);
  nand g1027 (n_1337, n_424, n_425);
  nand g1028 (n_1338, n_426, n_425);
  nand g1029 (n_1339, n_424, n_426);
  nand g1030 (n_94, n_1337, n_1338, n_1339);
  xor g1031 (n_1340, A[25], A[23]);
  xor g1032 (n_431, n_1340, A[19]);
  nand g1033 (n_1341, A[25], A[23]);
  nand g1034 (n_1342, A[19], A[23]);
  nand g1035 (n_1343, A[25], A[19]);
  nand g1036 (n_441, n_1341, n_1342, n_1343);
  xor g1037 (n_1344, A[11], A[9]);
  xor g1038 (n_432, n_1344, A[17]);
  nand g1040 (n_1346, A[17], A[9]);
  nand g1042 (n_442, n_1051, n_1346, n_1222);
  xor g1043 (n_1348, A[7], A[21]);
  xor g1044 (n_430, n_1348, A[15]);
  nand g1045 (n_1349, A[7], A[21]);
  nand g1048 (n_443, n_1349, n_1215, n_1282);
  xor g1049 (n_1352, A[13], n_427);
  xor g1050 (n_434, n_1352, n_428);
  nand g1051 (n_1353, A[13], n_427);
  nand g1052 (n_1354, n_428, n_427);
  nand g1053 (n_1355, A[13], n_428);
  nand g1054 (n_447, n_1353, n_1354, n_1355);
  xor g1055 (n_1356, n_429, n_430);
  xor g1056 (n_436, n_1356, n_431);
  nand g1057 (n_1357, n_429, n_430);
  nand g1058 (n_1358, n_431, n_430);
  nand g1059 (n_1359, n_429, n_431);
  nand g1060 (n_449, n_1357, n_1358, n_1359);
  xor g1061 (n_1360, n_432, n_433);
  xor g1062 (n_438, n_1360, n_434);
  nand g1063 (n_1361, n_432, n_433);
  nand g1064 (n_1362, n_434, n_433);
  nand g1065 (n_1363, n_432, n_434);
  nand g1066 (n_451, n_1361, n_1362, n_1363);
  xor g1067 (n_1364, n_435, n_436);
  xor g1068 (n_439, n_1364, n_437);
  nand g1069 (n_1365, n_435, n_436);
  nand g1070 (n_1366, n_437, n_436);
  nand g1071 (n_1367, n_435, n_437);
  nand g1072 (n_454, n_1365, n_1366, n_1367);
  xor g1073 (n_1368, n_438, n_439);
  xor g1074 (n_163, n_1368, n_440);
  nand g1075 (n_1369, n_438, n_439);
  nand g1076 (n_1370, n_440, n_439);
  nand g1077 (n_1371, n_438, n_440);
  nand g1078 (n_93, n_1369, n_1370, n_1371);
  xor g1079 (n_1372, A[26], A[24]);
  xor g1080 (n_445, n_1372, A[20]);
  nand g1081 (n_1373, A[26], A[24]);
  nand g1082 (n_1374, A[20], A[24]);
  nand g1083 (n_1375, A[26], A[20]);
  nand g1084 (n_455, n_1373, n_1374, n_1375);
  xor g1086 (n_446, n_280, A[18]);
  nand g1088 (n_1378, A[18], A[10]);
  xor g1091 (n_1380, A[8], A[22]);
  xor g1092 (n_444, n_1380, A[16]);
  nand g1093 (n_1381, A[8], A[22]);
  nand g1096 (n_457, n_1381, n_1247, n_1314);
  xor g1097 (n_1384, A[14], n_441);
  xor g1098 (n_448, n_1384, n_442);
  nand g1099 (n_1385, A[14], n_441);
  nand g1100 (n_1386, n_442, n_441);
  nand g1101 (n_1387, A[14], n_442);
  nand g1102 (n_461, n_1385, n_1386, n_1387);
  xor g1103 (n_1388, n_443, n_444);
  xor g1104 (n_450, n_1388, n_445);
  nand g1105 (n_1389, n_443, n_444);
  nand g1106 (n_1390, n_445, n_444);
  nand g1107 (n_1391, n_443, n_445);
  nand g1108 (n_463, n_1389, n_1390, n_1391);
  xor g1109 (n_1392, n_446, n_447);
  xor g1110 (n_452, n_1392, n_448);
  nand g1111 (n_1393, n_446, n_447);
  nand g1112 (n_1394, n_448, n_447);
  nand g1113 (n_1395, n_446, n_448);
  nand g1114 (n_465, n_1393, n_1394, n_1395);
  xor g1115 (n_1396, n_449, n_450);
  xor g1116 (n_453, n_1396, n_451);
  nand g1117 (n_1397, n_449, n_450);
  nand g1118 (n_1398, n_451, n_450);
  nand g1119 (n_1399, n_449, n_451);
  nand g1120 (n_468, n_1397, n_1398, n_1399);
  xor g1121 (n_1400, n_452, n_453);
  xor g1122 (n_162, n_1400, n_454);
  nand g1123 (n_1401, n_452, n_453);
  nand g1124 (n_1402, n_454, n_453);
  nand g1125 (n_1403, n_452, n_454);
  nand g1126 (n_92, n_1401, n_1402, n_1403);
  xor g1127 (n_1404, A[27], A[25]);
  xor g1128 (n_459, n_1404, A[21]);
  nand g1129 (n_1405, A[27], A[25]);
  nand g1130 (n_1406, A[21], A[25]);
  nand g1131 (n_1407, A[27], A[21]);
  nand g1132 (n_469, n_1405, n_1406, n_1407);
  xor g1133 (n_1408, A[13], A[11]);
  xor g1134 (n_460, n_1408, A[19]);
  nand g1135 (n_1409, A[13], A[11]);
  nand g1136 (n_1410, A[19], A[11]);
  nand g1138 (n_470, n_1409, n_1410, n_1150);
  xor g1139 (n_1412, A[9], A[23]);
  xor g1140 (n_458, n_1412, A[17]);
  nand g1141 (n_1413, A[9], A[23]);
  nand g1144 (n_471, n_1413, n_1279, n_1346);
  xor g1145 (n_1416, A[15], n_455);
  xor g1146 (n_462, n_1416, n_456);
  nand g1147 (n_1417, A[15], n_455);
  nand g1148 (n_1418, n_456, n_455);
  nand g1149 (n_1419, A[15], n_456);
  nand g1150 (n_475, n_1417, n_1418, n_1419);
  xor g1151 (n_1420, n_457, n_458);
  xor g1152 (n_464, n_1420, n_459);
  nand g1153 (n_1421, n_457, n_458);
  nand g1154 (n_1422, n_459, n_458);
  nand g1155 (n_1423, n_457, n_459);
  nand g1156 (n_477, n_1421, n_1422, n_1423);
  xor g1157 (n_1424, n_460, n_461);
  xor g1158 (n_466, n_1424, n_462);
  nand g1159 (n_1425, n_460, n_461);
  nand g1160 (n_1426, n_462, n_461);
  nand g1161 (n_1427, n_460, n_462);
  nand g1162 (n_479, n_1425, n_1426, n_1427);
  xor g1163 (n_1428, n_463, n_464);
  xor g1164 (n_467, n_1428, n_465);
  nand g1165 (n_1429, n_463, n_464);
  nand g1166 (n_1430, n_465, n_464);
  nand g1167 (n_1431, n_463, n_465);
  nand g1168 (n_482, n_1429, n_1430, n_1431);
  xor g1169 (n_1432, n_466, n_467);
  xor g1170 (n_161, n_1432, n_468);
  nand g1171 (n_1433, n_466, n_467);
  nand g1172 (n_1434, n_468, n_467);
  nand g1173 (n_1435, n_466, n_468);
  nand g1174 (n_91, n_1433, n_1434, n_1435);
  xor g1175 (n_1436, A[28], A[26]);
  xor g1176 (n_473, n_1436, A[22]);
  nand g1177 (n_1437, A[28], A[26]);
  nand g1178 (n_1438, A[22], A[26]);
  nand g1179 (n_1439, A[28], A[22]);
  nand g1180 (n_483, n_1437, n_1438, n_1439);
  xor g1182 (n_474, n_295, A[20]);
  nand g1184 (n_1442, A[20], A[12]);
  xor g1187 (n_1444, A[10], A[24]);
  xor g1188 (n_472, n_1444, A[18]);
  nand g1189 (n_1445, A[10], A[24]);
  nand g1192 (n_485, n_1445, n_1311, n_1378);
  xor g1193 (n_1448, A[16], n_469);
  xor g1194 (n_476, n_1448, n_470);
  nand g1195 (n_1449, A[16], n_469);
  nand g1196 (n_1450, n_470, n_469);
  nand g1197 (n_1451, A[16], n_470);
  nand g1198 (n_489, n_1449, n_1450, n_1451);
  xor g1199 (n_1452, n_471, n_472);
  xor g1200 (n_478, n_1452, n_473);
  nand g1201 (n_1453, n_471, n_472);
  nand g1202 (n_1454, n_473, n_472);
  nand g1203 (n_1455, n_471, n_473);
  nand g1204 (n_491, n_1453, n_1454, n_1455);
  xor g1205 (n_1456, n_474, n_475);
  xor g1206 (n_480, n_1456, n_476);
  nand g1207 (n_1457, n_474, n_475);
  nand g1208 (n_1458, n_476, n_475);
  nand g1209 (n_1459, n_474, n_476);
  nand g1210 (n_493, n_1457, n_1458, n_1459);
  xor g1211 (n_1460, n_477, n_478);
  xor g1212 (n_481, n_1460, n_479);
  nand g1213 (n_1461, n_477, n_478);
  nand g1214 (n_1462, n_479, n_478);
  nand g1215 (n_1463, n_477, n_479);
  nand g1216 (n_496, n_1461, n_1462, n_1463);
  xor g1217 (n_1464, n_480, n_481);
  xor g1218 (n_160, n_1464, n_482);
  nand g1219 (n_1465, n_480, n_481);
  nand g1220 (n_1466, n_482, n_481);
  nand g1221 (n_1467, n_480, n_482);
  nand g1222 (n_90, n_1465, n_1466, n_1467);
  xor g1223 (n_1468, A[29], A[27]);
  xor g1224 (n_487, n_1468, A[23]);
  nand g1225 (n_1469, A[29], A[27]);
  nand g1226 (n_1470, A[23], A[27]);
  nand g1227 (n_1471, A[29], A[23]);
  nand g1228 (n_497, n_1469, n_1470, n_1471);
  xor g1229 (n_1472, A[15], A[13]);
  xor g1230 (n_488, n_1472, A[21]);
  nand g1232 (n_1474, A[21], A[13]);
  nand g1234 (n_498, n_1046, n_1474, n_1215);
  xor g1235 (n_1476, A[11], A[25]);
  xor g1236 (n_486, n_1476, A[19]);
  nand g1237 (n_1477, A[11], A[25]);
  nand g1240 (n_499, n_1477, n_1343, n_1410);
  xor g1241 (n_1480, A[17], n_483);
  xor g1242 (n_490, n_1480, n_484);
  nand g1243 (n_1481, A[17], n_483);
  nand g1244 (n_1482, n_484, n_483);
  nand g1245 (n_1483, A[17], n_484);
  nand g1246 (n_503, n_1481, n_1482, n_1483);
  xor g1247 (n_1484, n_485, n_486);
  xor g1248 (n_492, n_1484, n_487);
  nand g1249 (n_1485, n_485, n_486);
  nand g1250 (n_1486, n_487, n_486);
  nand g1251 (n_1487, n_485, n_487);
  nand g1252 (n_505, n_1485, n_1486, n_1487);
  xor g1253 (n_1488, n_488, n_489);
  xor g1254 (n_494, n_1488, n_490);
  nand g1255 (n_1489, n_488, n_489);
  nand g1256 (n_1490, n_490, n_489);
  nand g1257 (n_1491, n_488, n_490);
  nand g1258 (n_507, n_1489, n_1490, n_1491);
  xor g1259 (n_1492, n_491, n_492);
  xor g1260 (n_495, n_1492, n_493);
  nand g1261 (n_1493, n_491, n_492);
  nand g1262 (n_1494, n_493, n_492);
  nand g1263 (n_1495, n_491, n_493);
  nand g1264 (n_510, n_1493, n_1494, n_1495);
  xor g1265 (n_1496, n_494, n_495);
  xor g1266 (n_159, n_1496, n_496);
  nand g1267 (n_1497, n_494, n_495);
  nand g1268 (n_1498, n_496, n_495);
  nand g1269 (n_1499, n_494, n_496);
  nand g1270 (n_89, n_1497, n_1498, n_1499);
  xor g1271 (n_1500, A[30], A[28]);
  xor g1272 (n_501, n_1500, A[24]);
  nand g1273 (n_1501, A[30], A[28]);
  nand g1274 (n_1502, A[24], A[28]);
  nand g1275 (n_1503, A[30], A[24]);
  nand g1276 (n_511, n_1501, n_1502, n_1503);
  xor g1278 (n_502, n_314, A[22]);
  nand g1280 (n_1506, A[22], A[14]);
  xor g1283 (n_1508, A[12], A[26]);
  xor g1284 (n_500, n_1508, A[20]);
  nand g1285 (n_1509, A[12], A[26]);
  nand g1288 (n_513, n_1509, n_1375, n_1442);
  xor g1289 (n_1512, A[18], n_497);
  xor g1290 (n_504, n_1512, n_498);
  nand g1291 (n_1513, A[18], n_497);
  nand g1292 (n_1514, n_498, n_497);
  nand g1293 (n_1515, A[18], n_498);
  nand g1294 (n_517, n_1513, n_1514, n_1515);
  xor g1295 (n_1516, n_499, n_500);
  xor g1296 (n_506, n_1516, n_501);
  nand g1297 (n_1517, n_499, n_500);
  nand g1298 (n_1518, n_501, n_500);
  nand g1299 (n_1519, n_499, n_501);
  nand g1300 (n_519, n_1517, n_1518, n_1519);
  xor g1301 (n_1520, n_502, n_503);
  xor g1302 (n_508, n_1520, n_504);
  nand g1303 (n_1521, n_502, n_503);
  nand g1304 (n_1522, n_504, n_503);
  nand g1305 (n_1523, n_502, n_504);
  nand g1306 (n_521, n_1521, n_1522, n_1523);
  xor g1307 (n_1524, n_505, n_506);
  xor g1308 (n_509, n_1524, n_507);
  nand g1309 (n_1525, n_505, n_506);
  nand g1310 (n_1526, n_507, n_506);
  nand g1311 (n_1527, n_505, n_507);
  nand g1312 (n_524, n_1525, n_1526, n_1527);
  xor g1313 (n_1528, n_508, n_509);
  xor g1314 (n_158, n_1528, n_510);
  nand g1315 (n_1529, n_508, n_509);
  nand g1316 (n_1530, n_510, n_509);
  nand g1317 (n_1531, n_508, n_510);
  nand g1318 (n_88, n_1529, n_1530, n_1531);
  xor g1319 (n_1532, A[31], A[29]);
  xor g1320 (n_515, n_1532, A[25]);
  nand g1321 (n_1533, A[31], A[29]);
  nand g1322 (n_1534, A[25], A[29]);
  nand g1323 (n_1535, A[31], A[25]);
  nand g1324 (n_525, n_1533, n_1534, n_1535);
  xor g1325 (n_1536, A[17], A[15]);
  xor g1326 (n_516, n_1536, A[23]);
  nand g1328 (n_1538, A[23], A[15]);
  nand g1330 (n_526, n_1094, n_1538, n_1279);
  xor g1331 (n_1540, A[13], A[27]);
  xor g1332 (n_514, n_1540, A[21]);
  nand g1333 (n_1541, A[13], A[27]);
  nand g1336 (n_527, n_1541, n_1407, n_1474);
  xor g1337 (n_1544, A[19], n_511);
  xor g1338 (n_518, n_1544, n_512);
  nand g1339 (n_1545, A[19], n_511);
  nand g1340 (n_1546, n_512, n_511);
  nand g1341 (n_1547, A[19], n_512);
  nand g1342 (n_531, n_1545, n_1546, n_1547);
  xor g1343 (n_1548, n_513, n_514);
  xor g1344 (n_520, n_1548, n_515);
  nand g1345 (n_1549, n_513, n_514);
  nand g1346 (n_1550, n_515, n_514);
  nand g1347 (n_1551, n_513, n_515);
  nand g1348 (n_533, n_1549, n_1550, n_1551);
  xor g1349 (n_1552, n_516, n_517);
  xor g1350 (n_522, n_1552, n_518);
  nand g1351 (n_1553, n_516, n_517);
  nand g1352 (n_1554, n_518, n_517);
  nand g1353 (n_1555, n_516, n_518);
  nand g1354 (n_535, n_1553, n_1554, n_1555);
  xor g1355 (n_1556, n_519, n_520);
  xor g1356 (n_523, n_1556, n_521);
  nand g1357 (n_1557, n_519, n_520);
  nand g1358 (n_1558, n_521, n_520);
  nand g1359 (n_1559, n_519, n_521);
  nand g1360 (n_538, n_1557, n_1558, n_1559);
  xor g1361 (n_1560, n_522, n_523);
  xor g1362 (n_157, n_1560, n_524);
  nand g1363 (n_1561, n_522, n_523);
  nand g1364 (n_1562, n_524, n_523);
  nand g1365 (n_1563, n_522, n_524);
  nand g1366 (n_87, n_1561, n_1562, n_1563);
  xor g1367 (n_1564, A[32], A[30]);
  xor g1368 (n_529, n_1564, A[26]);
  nand g1369 (n_1565, A[32], A[30]);
  nand g1370 (n_1566, A[26], A[30]);
  nand g1371 (n_1567, A[32], A[26]);
  nand g1372 (n_539, n_1565, n_1566, n_1567);
  xor g1374 (n_530, n_337, A[24]);
  nand g1376 (n_1570, A[24], A[16]);
  xor g1379 (n_1572, A[14], A[28]);
  xor g1380 (n_528, n_1572, A[22]);
  nand g1381 (n_1573, A[14], A[28]);
  nand g1384 (n_541, n_1573, n_1439, n_1506);
  xor g1385 (n_1576, A[20], n_525);
  xor g1386 (n_532, n_1576, n_526);
  nand g1387 (n_1577, A[20], n_525);
  nand g1388 (n_1578, n_526, n_525);
  nand g1389 (n_1579, A[20], n_526);
  nand g1390 (n_545, n_1577, n_1578, n_1579);
  xor g1391 (n_1580, n_527, n_528);
  xor g1392 (n_534, n_1580, n_529);
  nand g1393 (n_1581, n_527, n_528);
  nand g1394 (n_1582, n_529, n_528);
  nand g1395 (n_1583, n_527, n_529);
  nand g1396 (n_547, n_1581, n_1582, n_1583);
  xor g1397 (n_1584, n_530, n_531);
  xor g1398 (n_536, n_1584, n_532);
  nand g1399 (n_1585, n_530, n_531);
  nand g1400 (n_1586, n_532, n_531);
  nand g1401 (n_1587, n_530, n_532);
  nand g1402 (n_549, n_1585, n_1586, n_1587);
  xor g1403 (n_1588, n_533, n_534);
  xor g1404 (n_537, n_1588, n_535);
  nand g1405 (n_1589, n_533, n_534);
  nand g1406 (n_1590, n_535, n_534);
  nand g1407 (n_1591, n_533, n_535);
  nand g1408 (n_552, n_1589, n_1590, n_1591);
  xor g1409 (n_1592, n_536, n_537);
  xor g1410 (n_156, n_1592, n_538);
  nand g1411 (n_1593, n_536, n_537);
  nand g1412 (n_1594, n_538, n_537);
  nand g1413 (n_1595, n_536, n_538);
  nand g1414 (n_86, n_1593, n_1594, n_1595);
  xor g1415 (n_1596, A[33], A[31]);
  xor g1416 (n_543, n_1596, A[27]);
  nand g1417 (n_1597, A[33], A[31]);
  nand g1418 (n_1598, A[27], A[31]);
  nand g1419 (n_1599, A[33], A[27]);
  nand g1420 (n_553, n_1597, n_1598, n_1599);
  xor g1421 (n_1600, A[19], A[17]);
  xor g1422 (n_544, n_1600, A[25]);
  nand g1423 (n_1601, A[19], A[17]);
  nand g1424 (n_1602, A[25], A[17]);
  nand g1426 (n_554, n_1601, n_1602, n_1343);
  xor g1427 (n_1604, A[15], A[29]);
  xor g1428 (n_542, n_1604, A[23]);
  nand g1429 (n_1605, A[15], A[29]);
  nand g1432 (n_555, n_1605, n_1471, n_1538);
  xor g1433 (n_1608, A[21], n_539);
  xor g1434 (n_546, n_1608, n_540);
  nand g1435 (n_1609, A[21], n_539);
  nand g1436 (n_1610, n_540, n_539);
  nand g1437 (n_1611, A[21], n_540);
  nand g1438 (n_559, n_1609, n_1610, n_1611);
  xor g1439 (n_1612, n_541, n_542);
  xor g1440 (n_548, n_1612, n_543);
  nand g1441 (n_1613, n_541, n_542);
  nand g1442 (n_1614, n_543, n_542);
  nand g1443 (n_1615, n_541, n_543);
  nand g1444 (n_561, n_1613, n_1614, n_1615);
  xor g1445 (n_1616, n_544, n_545);
  xor g1446 (n_550, n_1616, n_546);
  nand g1447 (n_1617, n_544, n_545);
  nand g1448 (n_1618, n_546, n_545);
  nand g1449 (n_1619, n_544, n_546);
  nand g1450 (n_563, n_1617, n_1618, n_1619);
  xor g1451 (n_1620, n_547, n_548);
  xor g1452 (n_551, n_1620, n_549);
  nand g1453 (n_1621, n_547, n_548);
  nand g1454 (n_1622, n_549, n_548);
  nand g1455 (n_1623, n_547, n_549);
  nand g1456 (n_566, n_1621, n_1622, n_1623);
  xor g1457 (n_1624, n_550, n_551);
  xor g1458 (n_155, n_1624, n_552);
  nand g1459 (n_1625, n_550, n_551);
  nand g1460 (n_1626, n_552, n_551);
  nand g1461 (n_1627, n_550, n_552);
  nand g1462 (n_85, n_1625, n_1626, n_1627);
  xor g1463 (n_1628, A[34], A[32]);
  xor g1464 (n_557, n_1628, A[28]);
  nand g1465 (n_1629, A[34], A[32]);
  nand g1466 (n_1630, A[28], A[32]);
  nand g1467 (n_1631, A[34], A[28]);
  nand g1468 (n_567, n_1629, n_1630, n_1631);
  xor g1470 (n_558, n_1180, A[26]);
  nand g1472 (n_1634, A[26], A[18]);
  nand g1474 (n_568, n_1181, n_1634, n_1375);
  xor g1475 (n_1636, A[16], A[30]);
  xor g1476 (n_556, n_1636, A[24]);
  nand g1477 (n_1637, A[16], A[30]);
  nand g1480 (n_569, n_1637, n_1503, n_1570);
  xor g1481 (n_1640, A[22], n_553);
  xor g1482 (n_560, n_1640, n_554);
  nand g1483 (n_1641, A[22], n_553);
  nand g1484 (n_1642, n_554, n_553);
  nand g1485 (n_1643, A[22], n_554);
  nand g1486 (n_573, n_1641, n_1642, n_1643);
  xor g1487 (n_1644, n_555, n_556);
  xor g1488 (n_562, n_1644, n_557);
  nand g1489 (n_1645, n_555, n_556);
  nand g1490 (n_1646, n_557, n_556);
  nand g1491 (n_1647, n_555, n_557);
  nand g1492 (n_575, n_1645, n_1646, n_1647);
  xor g1493 (n_1648, n_558, n_559);
  xor g1494 (n_564, n_1648, n_560);
  nand g1495 (n_1649, n_558, n_559);
  nand g1496 (n_1650, n_560, n_559);
  nand g1497 (n_1651, n_558, n_560);
  nand g1498 (n_577, n_1649, n_1650, n_1651);
  xor g1499 (n_1652, n_561, n_562);
  xor g1500 (n_565, n_1652, n_563);
  nand g1501 (n_1653, n_561, n_562);
  nand g1502 (n_1654, n_563, n_562);
  nand g1503 (n_1655, n_561, n_563);
  nand g1504 (n_580, n_1653, n_1654, n_1655);
  xor g1505 (n_1656, n_564, n_565);
  xor g1506 (n_154, n_1656, n_566);
  nand g1507 (n_1657, n_564, n_565);
  nand g1508 (n_1658, n_566, n_565);
  nand g1509 (n_1659, n_564, n_566);
  nand g1510 (n_84, n_1657, n_1658, n_1659);
  xor g1511 (n_1660, A[35], A[33]);
  xor g1512 (n_571, n_1660, A[29]);
  nand g1513 (n_1661, A[35], A[33]);
  nand g1514 (n_1662, A[29], A[33]);
  nand g1515 (n_1663, A[35], A[29]);
  nand g1516 (n_581, n_1661, n_1662, n_1663);
  xor g1518 (n_572, n_1212, A[27]);
  nand g1520 (n_1666, A[27], A[19]);
  nand g1522 (n_582, n_1213, n_1666, n_1407);
  xor g1523 (n_1668, A[17], A[31]);
  xor g1524 (n_570, n_1668, A[25]);
  nand g1525 (n_1669, A[17], A[31]);
  nand g1528 (n_583, n_1669, n_1535, n_1602);
  xor g1529 (n_1672, A[23], n_567);
  xor g1530 (n_574, n_1672, n_568);
  nand g1531 (n_1673, A[23], n_567);
  nand g1532 (n_1674, n_568, n_567);
  nand g1533 (n_1675, A[23], n_568);
  nand g1534 (n_587, n_1673, n_1674, n_1675);
  xor g1535 (n_1676, n_569, n_570);
  xor g1536 (n_576, n_1676, n_571);
  nand g1537 (n_1677, n_569, n_570);
  nand g1538 (n_1678, n_571, n_570);
  nand g1539 (n_1679, n_569, n_571);
  nand g1540 (n_589, n_1677, n_1678, n_1679);
  xor g1541 (n_1680, n_572, n_573);
  xor g1542 (n_578, n_1680, n_574);
  nand g1543 (n_1681, n_572, n_573);
  nand g1544 (n_1682, n_574, n_573);
  nand g1545 (n_1683, n_572, n_574);
  nand g1546 (n_591, n_1681, n_1682, n_1683);
  xor g1547 (n_1684, n_575, n_576);
  xor g1548 (n_579, n_1684, n_577);
  nand g1549 (n_1685, n_575, n_576);
  nand g1550 (n_1686, n_577, n_576);
  nand g1551 (n_1687, n_575, n_577);
  nand g1552 (n_594, n_1685, n_1686, n_1687);
  xor g1553 (n_1688, n_578, n_579);
  xor g1554 (n_153, n_1688, n_580);
  nand g1555 (n_1689, n_578, n_579);
  nand g1556 (n_1690, n_580, n_579);
  nand g1557 (n_1691, n_578, n_580);
  nand g1558 (n_83, n_1689, n_1690, n_1691);
  xor g1559 (n_1692, A[36], A[34]);
  xor g1560 (n_585, n_1692, A[30]);
  nand g1561 (n_1693, A[36], A[34]);
  nand g1562 (n_1694, A[30], A[34]);
  nand g1563 (n_1695, A[36], A[30]);
  nand g1564 (n_595, n_1693, n_1694, n_1695);
  xor g1566 (n_586, n_1244, A[28]);
  nand g1568 (n_1698, A[28], A[20]);
  nand g1570 (n_596, n_1245, n_1698, n_1439);
  xor g1571 (n_1700, A[18], A[32]);
  xor g1572 (n_584, n_1700, A[26]);
  nand g1573 (n_1701, A[18], A[32]);
  nand g1576 (n_597, n_1701, n_1567, n_1634);
  xor g1577 (n_1704, A[24], n_581);
  xor g1578 (n_588, n_1704, n_582);
  nand g1579 (n_1705, A[24], n_581);
  nand g1580 (n_1706, n_582, n_581);
  nand g1581 (n_1707, A[24], n_582);
  nand g1582 (n_601, n_1705, n_1706, n_1707);
  xor g1583 (n_1708, n_583, n_584);
  xor g1584 (n_590, n_1708, n_585);
  nand g1585 (n_1709, n_583, n_584);
  nand g1586 (n_1710, n_585, n_584);
  nand g1587 (n_1711, n_583, n_585);
  nand g1588 (n_603, n_1709, n_1710, n_1711);
  xor g1589 (n_1712, n_586, n_587);
  xor g1590 (n_592, n_1712, n_588);
  nand g1591 (n_1713, n_586, n_587);
  nand g1592 (n_1714, n_588, n_587);
  nand g1593 (n_1715, n_586, n_588);
  nand g1594 (n_605, n_1713, n_1714, n_1715);
  xor g1595 (n_1716, n_589, n_590);
  xor g1596 (n_593, n_1716, n_591);
  nand g1597 (n_1717, n_589, n_590);
  nand g1598 (n_1718, n_591, n_590);
  nand g1599 (n_1719, n_589, n_591);
  nand g1600 (n_608, n_1717, n_1718, n_1719);
  xor g1601 (n_1720, n_592, n_593);
  xor g1602 (n_152, n_1720, n_594);
  nand g1603 (n_1721, n_592, n_593);
  nand g1604 (n_1722, n_594, n_593);
  nand g1605 (n_1723, n_592, n_594);
  nand g1606 (n_82, n_1721, n_1722, n_1723);
  xor g1607 (n_1724, A[37], A[35]);
  xor g1608 (n_599, n_1724, A[31]);
  nand g1609 (n_1725, A[37], A[35]);
  nand g1610 (n_1726, A[31], A[35]);
  nand g1611 (n_1727, A[37], A[31]);
  nand g1612 (n_609, n_1725, n_1726, n_1727);
  xor g1614 (n_600, n_1276, A[29]);
  nand g1616 (n_1730, A[29], A[21]);
  nand g1618 (n_610, n_1277, n_1730, n_1471);
  xor g1619 (n_1732, A[19], A[33]);
  xor g1620 (n_598, n_1732, A[27]);
  nand g1621 (n_1733, A[19], A[33]);
  nand g1624 (n_611, n_1733, n_1599, n_1666);
  xor g1625 (n_1736, A[25], n_595);
  xor g1626 (n_602, n_1736, n_596);
  nand g1627 (n_1737, A[25], n_595);
  nand g1628 (n_1738, n_596, n_595);
  nand g1629 (n_1739, A[25], n_596);
  nand g1630 (n_615, n_1737, n_1738, n_1739);
  xor g1631 (n_1740, n_597, n_598);
  xor g1632 (n_604, n_1740, n_599);
  nand g1633 (n_1741, n_597, n_598);
  nand g1634 (n_1742, n_599, n_598);
  nand g1635 (n_1743, n_597, n_599);
  nand g1636 (n_617, n_1741, n_1742, n_1743);
  xor g1637 (n_1744, n_600, n_601);
  xor g1638 (n_606, n_1744, n_602);
  nand g1639 (n_1745, n_600, n_601);
  nand g1640 (n_1746, n_602, n_601);
  nand g1641 (n_1747, n_600, n_602);
  nand g1642 (n_619, n_1745, n_1746, n_1747);
  xor g1643 (n_1748, n_603, n_604);
  xor g1644 (n_607, n_1748, n_605);
  nand g1645 (n_1749, n_603, n_604);
  nand g1646 (n_1750, n_605, n_604);
  nand g1647 (n_1751, n_603, n_605);
  nand g1648 (n_622, n_1749, n_1750, n_1751);
  xor g1649 (n_1752, n_606, n_607);
  xor g1650 (n_151, n_1752, n_608);
  nand g1651 (n_1753, n_606, n_607);
  nand g1652 (n_1754, n_608, n_607);
  nand g1653 (n_1755, n_606, n_608);
  nand g1654 (n_81, n_1753, n_1754, n_1755);
  xor g1655 (n_1756, A[38], A[36]);
  xor g1656 (n_613, n_1756, A[32]);
  nand g1657 (n_1757, A[38], A[36]);
  nand g1658 (n_1758, A[32], A[36]);
  nand g1659 (n_1759, A[38], A[32]);
  nand g1660 (n_623, n_1757, n_1758, n_1759);
  xor g1662 (n_614, n_1308, A[30]);
  nand g1664 (n_1762, A[30], A[22]);
  nand g1666 (n_624, n_1309, n_1762, n_1503);
  xor g1667 (n_1764, A[20], A[34]);
  xor g1668 (n_612, n_1764, A[28]);
  nand g1669 (n_1765, A[20], A[34]);
  nand g1672 (n_625, n_1765, n_1631, n_1698);
  xor g1673 (n_1768, A[26], n_609);
  xor g1674 (n_616, n_1768, n_610);
  nand g1675 (n_1769, A[26], n_609);
  nand g1676 (n_1770, n_610, n_609);
  nand g1677 (n_1771, A[26], n_610);
  nand g1678 (n_629, n_1769, n_1770, n_1771);
  xor g1679 (n_1772, n_611, n_612);
  xor g1680 (n_618, n_1772, n_613);
  nand g1681 (n_1773, n_611, n_612);
  nand g1682 (n_1774, n_613, n_612);
  nand g1683 (n_1775, n_611, n_613);
  nand g1684 (n_631, n_1773, n_1774, n_1775);
  xor g1685 (n_1776, n_614, n_615);
  xor g1686 (n_620, n_1776, n_616);
  nand g1687 (n_1777, n_614, n_615);
  nand g1688 (n_1778, n_616, n_615);
  nand g1689 (n_1779, n_614, n_616);
  nand g1690 (n_633, n_1777, n_1778, n_1779);
  xor g1691 (n_1780, n_617, n_618);
  xor g1692 (n_621, n_1780, n_619);
  nand g1693 (n_1781, n_617, n_618);
  nand g1694 (n_1782, n_619, n_618);
  nand g1695 (n_1783, n_617, n_619);
  nand g1696 (n_636, n_1781, n_1782, n_1783);
  xor g1697 (n_1784, n_620, n_621);
  xor g1698 (n_150, n_1784, n_622);
  nand g1699 (n_1785, n_620, n_621);
  nand g1700 (n_1786, n_622, n_621);
  nand g1701 (n_1787, n_620, n_622);
  nand g1702 (n_80, n_1785, n_1786, n_1787);
  xor g1703 (n_1788, A[39], A[37]);
  xor g1704 (n_627, n_1788, A[33]);
  nand g1705 (n_1789, A[39], A[37]);
  nand g1706 (n_1790, A[33], A[37]);
  nand g1707 (n_1791, A[39], A[33]);
  nand g1708 (n_637, n_1789, n_1790, n_1791);
  xor g1710 (n_628, n_1340, A[31]);
  nand g1712 (n_1794, A[31], A[23]);
  nand g1714 (n_638, n_1341, n_1794, n_1535);
  xor g1715 (n_1796, A[21], A[35]);
  xor g1716 (n_626, n_1796, A[29]);
  nand g1717 (n_1797, A[21], A[35]);
  nand g1720 (n_639, n_1797, n_1663, n_1730);
  xor g1721 (n_1800, A[27], n_623);
  xor g1722 (n_630, n_1800, n_624);
  nand g1723 (n_1801, A[27], n_623);
  nand g1724 (n_1802, n_624, n_623);
  nand g1725 (n_1803, A[27], n_624);
  nand g1726 (n_643, n_1801, n_1802, n_1803);
  xor g1727 (n_1804, n_625, n_626);
  xor g1728 (n_632, n_1804, n_627);
  nand g1729 (n_1805, n_625, n_626);
  nand g1730 (n_1806, n_627, n_626);
  nand g1731 (n_1807, n_625, n_627);
  nand g1732 (n_645, n_1805, n_1806, n_1807);
  xor g1733 (n_1808, n_628, n_629);
  xor g1734 (n_634, n_1808, n_630);
  nand g1735 (n_1809, n_628, n_629);
  nand g1736 (n_1810, n_630, n_629);
  nand g1737 (n_1811, n_628, n_630);
  nand g1738 (n_647, n_1809, n_1810, n_1811);
  xor g1739 (n_1812, n_631, n_632);
  xor g1740 (n_635, n_1812, n_633);
  nand g1741 (n_1813, n_631, n_632);
  nand g1742 (n_1814, n_633, n_632);
  nand g1743 (n_1815, n_631, n_633);
  nand g1744 (n_650, n_1813, n_1814, n_1815);
  xor g1745 (n_1816, n_634, n_635);
  xor g1746 (n_149, n_1816, n_636);
  nand g1747 (n_1817, n_634, n_635);
  nand g1748 (n_1818, n_636, n_635);
  nand g1749 (n_1819, n_634, n_636);
  nand g1750 (n_79, n_1817, n_1818, n_1819);
  xor g1751 (n_1820, A[40], A[38]);
  xor g1752 (n_641, n_1820, A[34]);
  nand g1753 (n_1821, A[40], A[38]);
  nand g1754 (n_1822, A[34], A[38]);
  nand g1755 (n_1823, A[40], A[34]);
  nand g1756 (n_651, n_1821, n_1822, n_1823);
  xor g1758 (n_642, n_1372, A[32]);
  nand g1760 (n_1826, A[32], A[24]);
  nand g1762 (n_652, n_1373, n_1826, n_1567);
  xor g1763 (n_1828, A[22], A[36]);
  xor g1764 (n_640, n_1828, A[30]);
  nand g1765 (n_1829, A[22], A[36]);
  nand g1768 (n_653, n_1829, n_1695, n_1762);
  xor g1769 (n_1832, A[28], n_637);
  xor g1770 (n_644, n_1832, n_638);
  nand g1771 (n_1833, A[28], n_637);
  nand g1772 (n_1834, n_638, n_637);
  nand g1773 (n_1835, A[28], n_638);
  nand g1774 (n_657, n_1833, n_1834, n_1835);
  xor g1775 (n_1836, n_639, n_640);
  xor g1776 (n_646, n_1836, n_641);
  nand g1777 (n_1837, n_639, n_640);
  nand g1778 (n_1838, n_641, n_640);
  nand g1779 (n_1839, n_639, n_641);
  nand g1780 (n_659, n_1837, n_1838, n_1839);
  xor g1781 (n_1840, n_642, n_643);
  xor g1782 (n_648, n_1840, n_644);
  nand g1783 (n_1841, n_642, n_643);
  nand g1784 (n_1842, n_644, n_643);
  nand g1785 (n_1843, n_642, n_644);
  nand g1786 (n_661, n_1841, n_1842, n_1843);
  xor g1787 (n_1844, n_645, n_646);
  xor g1788 (n_649, n_1844, n_647);
  nand g1789 (n_1845, n_645, n_646);
  nand g1790 (n_1846, n_647, n_646);
  nand g1791 (n_1847, n_645, n_647);
  nand g1792 (n_664, n_1845, n_1846, n_1847);
  xor g1793 (n_1848, n_648, n_649);
  xor g1794 (n_148, n_1848, n_650);
  nand g1795 (n_1849, n_648, n_649);
  nand g1796 (n_1850, n_650, n_649);
  nand g1797 (n_1851, n_648, n_650);
  nand g1798 (n_78, n_1849, n_1850, n_1851);
  xor g1799 (n_1852, A[41], A[39]);
  xor g1800 (n_655, n_1852, A[35]);
  nand g1801 (n_1853, A[41], A[39]);
  nand g1802 (n_1854, A[35], A[39]);
  nand g1803 (n_1855, A[41], A[35]);
  nand g1804 (n_665, n_1853, n_1854, n_1855);
  xor g1806 (n_656, n_1404, A[33]);
  nand g1808 (n_1858, A[33], A[25]);
  nand g1810 (n_666, n_1405, n_1858, n_1599);
  xor g1811 (n_1860, A[23], A[37]);
  xor g1812 (n_654, n_1860, A[31]);
  nand g1813 (n_1861, A[23], A[37]);
  nand g1816 (n_667, n_1861, n_1727, n_1794);
  xor g1817 (n_1864, A[29], n_651);
  xor g1818 (n_658, n_1864, n_652);
  nand g1819 (n_1865, A[29], n_651);
  nand g1820 (n_1866, n_652, n_651);
  nand g1821 (n_1867, A[29], n_652);
  nand g1822 (n_671, n_1865, n_1866, n_1867);
  xor g1823 (n_1868, n_653, n_654);
  xor g1824 (n_660, n_1868, n_655);
  nand g1825 (n_1869, n_653, n_654);
  nand g1826 (n_1870, n_655, n_654);
  nand g1827 (n_1871, n_653, n_655);
  nand g1828 (n_673, n_1869, n_1870, n_1871);
  xor g1829 (n_1872, n_656, n_657);
  xor g1830 (n_662, n_1872, n_658);
  nand g1831 (n_1873, n_656, n_657);
  nand g1832 (n_1874, n_658, n_657);
  nand g1833 (n_1875, n_656, n_658);
  nand g1834 (n_675, n_1873, n_1874, n_1875);
  xor g1835 (n_1876, n_659, n_660);
  xor g1836 (n_663, n_1876, n_661);
  nand g1837 (n_1877, n_659, n_660);
  nand g1838 (n_1878, n_661, n_660);
  nand g1839 (n_1879, n_659, n_661);
  nand g1840 (n_678, n_1877, n_1878, n_1879);
  xor g1841 (n_1880, n_662, n_663);
  xor g1842 (n_147, n_1880, n_664);
  nand g1843 (n_1881, n_662, n_663);
  nand g1844 (n_1882, n_664, n_663);
  nand g1845 (n_1883, n_662, n_664);
  nand g1846 (n_77, n_1881, n_1882, n_1883);
  xor g1847 (n_1884, A[42], A[40]);
  xor g1848 (n_669, n_1884, A[36]);
  nand g1849 (n_1885, A[42], A[40]);
  nand g1850 (n_1886, A[36], A[40]);
  nand g1851 (n_1887, A[42], A[36]);
  nand g1852 (n_679, n_1885, n_1886, n_1887);
  xor g1854 (n_670, n_1436, A[34]);
  nand g1856 (n_1890, A[34], A[26]);
  nand g1858 (n_680, n_1437, n_1890, n_1631);
  xor g1859 (n_1892, A[24], A[38]);
  xor g1860 (n_668, n_1892, A[32]);
  nand g1861 (n_1893, A[24], A[38]);
  nand g1864 (n_681, n_1893, n_1759, n_1826);
  xor g1865 (n_1896, A[30], n_665);
  xor g1866 (n_672, n_1896, n_666);
  nand g1867 (n_1897, A[30], n_665);
  nand g1868 (n_1898, n_666, n_665);
  nand g1869 (n_1899, A[30], n_666);
  nand g1870 (n_685, n_1897, n_1898, n_1899);
  xor g1871 (n_1900, n_667, n_668);
  xor g1872 (n_674, n_1900, n_669);
  nand g1873 (n_1901, n_667, n_668);
  nand g1874 (n_1902, n_669, n_668);
  nand g1875 (n_1903, n_667, n_669);
  nand g1876 (n_687, n_1901, n_1902, n_1903);
  xor g1877 (n_1904, n_670, n_671);
  xor g1878 (n_676, n_1904, n_672);
  nand g1879 (n_1905, n_670, n_671);
  nand g1880 (n_1906, n_672, n_671);
  nand g1881 (n_1907, n_670, n_672);
  nand g1882 (n_689, n_1905, n_1906, n_1907);
  xor g1883 (n_1908, n_673, n_674);
  xor g1884 (n_677, n_1908, n_675);
  nand g1885 (n_1909, n_673, n_674);
  nand g1886 (n_1910, n_675, n_674);
  nand g1887 (n_1911, n_673, n_675);
  nand g1888 (n_692, n_1909, n_1910, n_1911);
  xor g1889 (n_1912, n_676, n_677);
  xor g1890 (n_146, n_1912, n_678);
  nand g1891 (n_1913, n_676, n_677);
  nand g1892 (n_1914, n_678, n_677);
  nand g1893 (n_1915, n_676, n_678);
  nand g1894 (n_76, n_1913, n_1914, n_1915);
  xor g1895 (n_1916, A[43], A[41]);
  xor g1896 (n_683, n_1916, A[37]);
  nand g1897 (n_1917, A[43], A[41]);
  nand g1898 (n_1918, A[37], A[41]);
  nand g1899 (n_1919, A[43], A[37]);
  nand g1900 (n_693, n_1917, n_1918, n_1919);
  xor g1902 (n_684, n_1468, A[35]);
  nand g1904 (n_1922, A[35], A[27]);
  nand g1906 (n_694, n_1469, n_1922, n_1663);
  xor g1907 (n_1924, A[25], A[39]);
  xor g1908 (n_682, n_1924, A[33]);
  nand g1909 (n_1925, A[25], A[39]);
  nand g1912 (n_695, n_1925, n_1791, n_1858);
  xor g1913 (n_1928, A[31], n_679);
  xor g1914 (n_686, n_1928, n_680);
  nand g1915 (n_1929, A[31], n_679);
  nand g1916 (n_1930, n_680, n_679);
  nand g1917 (n_1931, A[31], n_680);
  nand g1918 (n_699, n_1929, n_1930, n_1931);
  xor g1919 (n_1932, n_681, n_682);
  xor g1920 (n_688, n_1932, n_683);
  nand g1921 (n_1933, n_681, n_682);
  nand g1922 (n_1934, n_683, n_682);
  nand g1923 (n_1935, n_681, n_683);
  nand g1924 (n_701, n_1933, n_1934, n_1935);
  xor g1925 (n_1936, n_684, n_685);
  xor g1926 (n_690, n_1936, n_686);
  nand g1927 (n_1937, n_684, n_685);
  nand g1928 (n_1938, n_686, n_685);
  nand g1929 (n_1939, n_684, n_686);
  nand g1930 (n_703, n_1937, n_1938, n_1939);
  xor g1931 (n_1940, n_687, n_688);
  xor g1932 (n_691, n_1940, n_689);
  nand g1933 (n_1941, n_687, n_688);
  nand g1934 (n_1942, n_689, n_688);
  nand g1935 (n_1943, n_687, n_689);
  nand g1936 (n_706, n_1941, n_1942, n_1943);
  xor g1937 (n_1944, n_690, n_691);
  xor g1938 (n_145, n_1944, n_692);
  nand g1939 (n_1945, n_690, n_691);
  nand g1940 (n_1946, n_692, n_691);
  nand g1941 (n_1947, n_690, n_692);
  nand g1942 (n_75, n_1945, n_1946, n_1947);
  xor g1943 (n_1948, A[44], A[42]);
  xor g1944 (n_697, n_1948, A[38]);
  nand g1945 (n_1949, A[44], A[42]);
  nand g1946 (n_1950, A[38], A[42]);
  nand g1947 (n_1951, A[44], A[38]);
  nand g1948 (n_707, n_1949, n_1950, n_1951);
  xor g1950 (n_698, n_1500, A[36]);
  nand g1952 (n_1954, A[36], A[28]);
  nand g1954 (n_708, n_1501, n_1954, n_1695);
  xor g1955 (n_1956, A[26], A[40]);
  xor g1956 (n_696, n_1956, A[34]);
  nand g1957 (n_1957, A[26], A[40]);
  nand g1960 (n_709, n_1957, n_1823, n_1890);
  xor g1961 (n_1960, A[32], n_693);
  xor g1962 (n_700, n_1960, n_694);
  nand g1963 (n_1961, A[32], n_693);
  nand g1964 (n_1962, n_694, n_693);
  nand g1965 (n_1963, A[32], n_694);
  nand g1966 (n_713, n_1961, n_1962, n_1963);
  xor g1967 (n_1964, n_695, n_696);
  xor g1968 (n_702, n_1964, n_697);
  nand g1969 (n_1965, n_695, n_696);
  nand g1970 (n_1966, n_697, n_696);
  nand g1971 (n_1967, n_695, n_697);
  nand g1972 (n_715, n_1965, n_1966, n_1967);
  xor g1973 (n_1968, n_698, n_699);
  xor g1974 (n_704, n_1968, n_700);
  nand g1975 (n_1969, n_698, n_699);
  nand g1976 (n_1970, n_700, n_699);
  nand g1977 (n_1971, n_698, n_700);
  nand g1978 (n_717, n_1969, n_1970, n_1971);
  xor g1979 (n_1972, n_701, n_702);
  xor g1980 (n_705, n_1972, n_703);
  nand g1981 (n_1973, n_701, n_702);
  nand g1982 (n_1974, n_703, n_702);
  nand g1983 (n_1975, n_701, n_703);
  nand g1984 (n_720, n_1973, n_1974, n_1975);
  xor g1985 (n_1976, n_704, n_705);
  xor g1986 (n_144, n_1976, n_706);
  nand g1987 (n_1977, n_704, n_705);
  nand g1988 (n_1978, n_706, n_705);
  nand g1989 (n_1979, n_704, n_706);
  nand g1990 (n_74, n_1977, n_1978, n_1979);
  xor g1991 (n_1980, A[45], A[43]);
  xor g1992 (n_711, n_1980, A[39]);
  nand g1993 (n_1981, A[45], A[43]);
  nand g1994 (n_1982, A[39], A[43]);
  nand g1995 (n_1983, A[45], A[39]);
  nand g1996 (n_721, n_1981, n_1982, n_1983);
  xor g1998 (n_712, n_1532, A[37]);
  nand g2000 (n_1986, A[37], A[29]);
  nand g2002 (n_722, n_1533, n_1986, n_1727);
  xor g2003 (n_1988, A[27], A[41]);
  xor g2004 (n_710, n_1988, A[35]);
  nand g2005 (n_1989, A[27], A[41]);
  nand g2008 (n_723, n_1989, n_1855, n_1922);
  xor g2009 (n_1992, A[33], n_707);
  xor g2010 (n_714, n_1992, n_708);
  nand g2011 (n_1993, A[33], n_707);
  nand g2012 (n_1994, n_708, n_707);
  nand g2013 (n_1995, A[33], n_708);
  nand g2014 (n_727, n_1993, n_1994, n_1995);
  xor g2015 (n_1996, n_709, n_710);
  xor g2016 (n_716, n_1996, n_711);
  nand g2017 (n_1997, n_709, n_710);
  nand g2018 (n_1998, n_711, n_710);
  nand g2019 (n_1999, n_709, n_711);
  nand g2020 (n_729, n_1997, n_1998, n_1999);
  xor g2021 (n_2000, n_712, n_713);
  xor g2022 (n_718, n_2000, n_714);
  nand g2023 (n_2001, n_712, n_713);
  nand g2024 (n_2002, n_714, n_713);
  nand g2025 (n_2003, n_712, n_714);
  nand g2026 (n_731, n_2001, n_2002, n_2003);
  xor g2027 (n_2004, n_715, n_716);
  xor g2028 (n_719, n_2004, n_717);
  nand g2029 (n_2005, n_715, n_716);
  nand g2030 (n_2006, n_717, n_716);
  nand g2031 (n_2007, n_715, n_717);
  nand g2032 (n_734, n_2005, n_2006, n_2007);
  xor g2033 (n_2008, n_718, n_719);
  xor g2034 (n_143, n_2008, n_720);
  nand g2035 (n_2009, n_718, n_719);
  nand g2036 (n_2010, n_720, n_719);
  nand g2037 (n_2011, n_718, n_720);
  nand g2038 (n_73, n_2009, n_2010, n_2011);
  xor g2039 (n_2012, A[46], A[44]);
  xor g2040 (n_725, n_2012, A[40]);
  nand g2041 (n_2013, A[46], A[44]);
  nand g2042 (n_2014, A[40], A[44]);
  nand g2043 (n_2015, A[46], A[40]);
  nand g2044 (n_735, n_2013, n_2014, n_2015);
  xor g2046 (n_726, n_1564, A[38]);
  nand g2048 (n_2018, A[38], A[30]);
  nand g2050 (n_736, n_1565, n_2018, n_1759);
  xor g2051 (n_2020, A[28], A[42]);
  xor g2052 (n_724, n_2020, A[36]);
  nand g2053 (n_2021, A[28], A[42]);
  nand g2056 (n_737, n_2021, n_1887, n_1954);
  xor g2057 (n_2024, A[34], n_721);
  xor g2058 (n_728, n_2024, n_722);
  nand g2059 (n_2025, A[34], n_721);
  nand g2060 (n_2026, n_722, n_721);
  nand g2061 (n_2027, A[34], n_722);
  nand g2062 (n_741, n_2025, n_2026, n_2027);
  xor g2063 (n_2028, n_723, n_724);
  xor g2064 (n_730, n_2028, n_725);
  nand g2065 (n_2029, n_723, n_724);
  nand g2066 (n_2030, n_725, n_724);
  nand g2067 (n_2031, n_723, n_725);
  nand g2068 (n_743, n_2029, n_2030, n_2031);
  xor g2069 (n_2032, n_726, n_727);
  xor g2070 (n_732, n_2032, n_728);
  nand g2071 (n_2033, n_726, n_727);
  nand g2072 (n_2034, n_728, n_727);
  nand g2073 (n_2035, n_726, n_728);
  nand g2074 (n_745, n_2033, n_2034, n_2035);
  xor g2075 (n_2036, n_729, n_730);
  xor g2076 (n_733, n_2036, n_731);
  nand g2077 (n_2037, n_729, n_730);
  nand g2078 (n_2038, n_731, n_730);
  nand g2079 (n_2039, n_729, n_731);
  nand g2080 (n_748, n_2037, n_2038, n_2039);
  xor g2081 (n_2040, n_732, n_733);
  xor g2082 (n_142, n_2040, n_734);
  nand g2083 (n_2041, n_732, n_733);
  nand g2084 (n_2042, n_734, n_733);
  nand g2085 (n_2043, n_732, n_734);
  nand g2086 (n_72, n_2041, n_2042, n_2043);
  xor g2087 (n_2044, A[47], A[45]);
  xor g2088 (n_739, n_2044, A[41]);
  nand g2089 (n_2045, A[47], A[45]);
  nand g2090 (n_2046, A[41], A[45]);
  nand g2091 (n_2047, A[47], A[41]);
  nand g2092 (n_749, n_2045, n_2046, n_2047);
  xor g2094 (n_740, n_1596, A[39]);
  nand g2096 (n_2050, A[39], A[31]);
  nand g2098 (n_750, n_1597, n_2050, n_1791);
  xor g2099 (n_2052, A[29], A[43]);
  xor g2100 (n_738, n_2052, A[37]);
  nand g2101 (n_2053, A[29], A[43]);
  nand g2104 (n_751, n_2053, n_1919, n_1986);
  xor g2105 (n_2056, A[35], n_735);
  xor g2106 (n_742, n_2056, n_736);
  nand g2107 (n_2057, A[35], n_735);
  nand g2108 (n_2058, n_736, n_735);
  nand g2109 (n_2059, A[35], n_736);
  nand g2110 (n_755, n_2057, n_2058, n_2059);
  xor g2111 (n_2060, n_737, n_738);
  xor g2112 (n_744, n_2060, n_739);
  nand g2113 (n_2061, n_737, n_738);
  nand g2114 (n_2062, n_739, n_738);
  nand g2115 (n_2063, n_737, n_739);
  nand g2116 (n_757, n_2061, n_2062, n_2063);
  xor g2117 (n_2064, n_740, n_741);
  xor g2118 (n_746, n_2064, n_742);
  nand g2119 (n_2065, n_740, n_741);
  nand g2120 (n_2066, n_742, n_741);
  nand g2121 (n_2067, n_740, n_742);
  nand g2122 (n_759, n_2065, n_2066, n_2067);
  xor g2123 (n_2068, n_743, n_744);
  xor g2124 (n_747, n_2068, n_745);
  nand g2125 (n_2069, n_743, n_744);
  nand g2126 (n_2070, n_745, n_744);
  nand g2127 (n_2071, n_743, n_745);
  nand g2128 (n_762, n_2069, n_2070, n_2071);
  xor g2129 (n_2072, n_746, n_747);
  xor g2130 (n_141, n_2072, n_748);
  nand g2131 (n_2073, n_746, n_747);
  nand g2132 (n_2074, n_748, n_747);
  nand g2133 (n_2075, n_746, n_748);
  nand g2134 (n_71, n_2073, n_2074, n_2075);
  xor g2135 (n_2076, A[48], A[46]);
  xor g2136 (n_753, n_2076, A[42]);
  nand g2137 (n_2077, A[48], A[46]);
  nand g2138 (n_2078, A[42], A[46]);
  nand g2139 (n_2079, A[48], A[42]);
  nand g2140 (n_766, n_2077, n_2078, n_2079);
  xor g2142 (n_754, n_1628, A[40]);
  nand g2144 (n_2082, A[40], A[32]);
  nand g2146 (n_767, n_1629, n_2082, n_1823);
  xor g2147 (n_2084, A[30], A[44]);
  xor g2148 (n_752, n_2084, A[38]);
  nand g2149 (n_2085, A[30], A[44]);
  nand g2152 (n_765, n_2085, n_1951, n_2018);
  xor g2153 (n_2088, A[36], n_749);
  xor g2154 (n_756, n_2088, n_750);
  nand g2155 (n_2089, A[36], n_749);
  nand g2156 (n_2090, n_750, n_749);
  nand g2157 (n_2091, A[36], n_750);
  nand g2158 (n_771, n_2089, n_2090, n_2091);
  xor g2159 (n_2092, n_751, n_752);
  xor g2160 (n_758, n_2092, n_753);
  nand g2161 (n_2093, n_751, n_752);
  nand g2162 (n_2094, n_753, n_752);
  nand g2163 (n_2095, n_751, n_753);
  nand g2164 (n_773, n_2093, n_2094, n_2095);
  xor g2165 (n_2096, n_754, n_755);
  xor g2166 (n_760, n_2096, n_756);
  nand g2167 (n_2097, n_754, n_755);
  nand g2168 (n_2098, n_756, n_755);
  nand g2169 (n_2099, n_754, n_756);
  nand g2170 (n_775, n_2097, n_2098, n_2099);
  xor g2171 (n_2100, n_757, n_758);
  xor g2172 (n_761, n_2100, n_759);
  nand g2173 (n_2101, n_757, n_758);
  nand g2174 (n_2102, n_759, n_758);
  nand g2175 (n_2103, n_757, n_759);
  nand g2176 (n_778, n_2101, n_2102, n_2103);
  xor g2177 (n_2104, n_760, n_761);
  xor g2178 (n_140, n_2104, n_762);
  nand g2179 (n_2105, n_760, n_761);
  nand g2180 (n_2106, n_762, n_761);
  nand g2181 (n_2107, n_760, n_762);
  nand g2182 (n_70, n_2105, n_2106, n_2107);
  xor g2185 (n_2108, A[49], A[43]);
  xor g2186 (n_769, n_2108, A[35]);
  nand g2187 (n_2109, A[49], A[43]);
  nand g2188 (n_2110, A[35], A[43]);
  nand g2189 (n_2111, A[49], A[35]);
  nand g2190 (n_783, n_2109, n_2110, n_2111);
  xor g2191 (n_2112, A[33], A[47]);
  xor g2192 (n_770, n_2112, A[31]);
  nand g2193 (n_2113, A[33], A[47]);
  nand g2194 (n_2114, A[31], A[47]);
  nand g2196 (n_784, n_2113, n_2114, n_1597);
  xor g2197 (n_2116, A[41], A[45]);
  xor g2198 (n_768, n_2116, A[39]);
  nand g2202 (n_782, n_2046, n_1983, n_1853);
  xor g2203 (n_2120, A[37], n_765);
  xor g2204 (n_772, n_2120, n_766);
  nand g2205 (n_2121, A[37], n_765);
  nand g2206 (n_2122, n_766, n_765);
  nand g2207 (n_2123, A[37], n_766);
  nand g2208 (n_788, n_2121, n_2122, n_2123);
  xor g2209 (n_2124, n_767, n_768);
  xor g2210 (n_774, n_2124, n_769);
  nand g2211 (n_2125, n_767, n_768);
  nand g2212 (n_2126, n_769, n_768);
  nand g2213 (n_2127, n_767, n_769);
  nand g2214 (n_790, n_2125, n_2126, n_2127);
  xor g2215 (n_2128, n_770, n_771);
  xor g2216 (n_776, n_2128, n_772);
  nand g2217 (n_2129, n_770, n_771);
  nand g2218 (n_2130, n_772, n_771);
  nand g2219 (n_2131, n_770, n_772);
  nand g2220 (n_792, n_2129, n_2130, n_2131);
  xor g2221 (n_2132, n_773, n_774);
  xor g2222 (n_777, n_2132, n_775);
  nand g2223 (n_2133, n_773, n_774);
  nand g2224 (n_2134, n_775, n_774);
  nand g2225 (n_2135, n_773, n_775);
  nand g2226 (n_795, n_2133, n_2134, n_2135);
  xor g2227 (n_2136, n_776, n_777);
  xor g2228 (n_139, n_2136, n_778);
  nand g2229 (n_2137, n_776, n_777);
  nand g2230 (n_2138, n_778, n_777);
  nand g2231 (n_2139, n_776, n_778);
  nand g2232 (n_69, n_2137, n_2138, n_2139);
  xor g2235 (n_2140, A[42], A[34]);
  xor g2236 (n_786, n_2140, A[32]);
  nand g2237 (n_2141, A[42], A[34]);
  nand g2239 (n_2143, A[42], A[32]);
  nand g2240 (n_797, n_2141, n_1629, n_2143);
  xor g2241 (n_2144, A[49], A[48]);
  xor g2242 (n_787, n_2144, A[40]);
  nand g2243 (n_2145, A[49], A[48]);
  nand g2244 (n_2146, A[40], A[48]);
  nand g2245 (n_2147, A[49], A[40]);
  nand g2246 (n_798, n_2145, n_2146, n_2147);
  xor g2248 (n_785, n_2012, A[38]);
  nand g2251 (n_2151, A[46], A[38]);
  nand g2252 (n_799, n_2013, n_1951, n_2151);
  xor g2253 (n_2152, A[36], n_782);
  xor g2254 (n_789, n_2152, n_783);
  nand g2255 (n_2153, A[36], n_782);
  nand g2256 (n_2154, n_783, n_782);
  nand g2257 (n_2155, A[36], n_783);
  nand g2258 (n_803, n_2153, n_2154, n_2155);
  xor g2259 (n_2156, n_784, n_785);
  xor g2260 (n_791, n_2156, n_786);
  nand g2261 (n_2157, n_784, n_785);
  nand g2262 (n_2158, n_786, n_785);
  nand g2263 (n_2159, n_784, n_786);
  nand g2264 (n_805, n_2157, n_2158, n_2159);
  xor g2265 (n_2160, n_787, n_788);
  xor g2266 (n_793, n_2160, n_789);
  nand g2267 (n_2161, n_787, n_788);
  nand g2268 (n_2162, n_789, n_788);
  nand g2269 (n_2163, n_787, n_789);
  nand g2270 (n_807, n_2161, n_2162, n_2163);
  xor g2271 (n_2164, n_790, n_791);
  xor g2272 (n_794, n_2164, n_792);
  nand g2273 (n_2165, n_790, n_791);
  nand g2274 (n_2166, n_792, n_791);
  nand g2275 (n_2167, n_790, n_792);
  nand g2276 (n_810, n_2165, n_2166, n_2167);
  xor g2277 (n_2168, n_793, n_794);
  xor g2278 (n_138, n_2168, n_795);
  nand g2279 (n_2169, n_793, n_794);
  nand g2280 (n_2170, n_795, n_794);
  nand g2281 (n_2171, n_793, n_795);
  nand g2282 (n_68, n_2169, n_2170, n_2171);
  xor g2284 (n_801, n_2172, A[43]);
  nand g2286 (n_2174, A[43], A[47]);
  nand g2288 (n_813, n_2173, n_2174, n_2175);
  xor g2290 (n_802, n_1660, A[41]);
  nand g2292 (n_2178, A[41], A[33]);
  nand g2294 (n_814, n_1661, n_2178, n_1855);
  xor g2296 (n_800, n_2180, A[39]);
  nand g2300 (n_815, n_2181, n_1983, n_2183);
  xor g2301 (n_2184, A[37], n_797);
  xor g2302 (n_804, n_2184, n_798);
  nand g2303 (n_2185, A[37], n_797);
  nand g2304 (n_2186, n_798, n_797);
  nand g2305 (n_2187, A[37], n_798);
  nand g2306 (n_819, n_2185, n_2186, n_2187);
  xor g2307 (n_2188, n_799, n_800);
  xor g2308 (n_806, n_2188, n_801);
  nand g2309 (n_2189, n_799, n_800);
  nand g2310 (n_2190, n_801, n_800);
  nand g2311 (n_2191, n_799, n_801);
  nand g2312 (n_821, n_2189, n_2190, n_2191);
  xor g2313 (n_2192, n_802, n_803);
  xor g2314 (n_808, n_2192, n_804);
  nand g2315 (n_2193, n_802, n_803);
  nand g2316 (n_2194, n_804, n_803);
  nand g2317 (n_2195, n_802, n_804);
  nand g2318 (n_823, n_2193, n_2194, n_2195);
  xor g2319 (n_2196, n_805, n_806);
  xor g2320 (n_809, n_2196, n_807);
  nand g2321 (n_2197, n_805, n_806);
  nand g2322 (n_2198, n_807, n_806);
  nand g2323 (n_2199, n_805, n_807);
  nand g2324 (n_825, n_2197, n_2198, n_2199);
  xor g2325 (n_2200, n_808, n_809);
  xor g2326 (n_137, n_2200, n_810);
  nand g2327 (n_2201, n_808, n_809);
  nand g2328 (n_2202, n_810, n_809);
  nand g2329 (n_2203, n_808, n_810);
  nand g2330 (n_67, n_2201, n_2202, n_2203);
  xor g2333 (n_2204, A[46], A[34]);
  xor g2334 (n_817, n_2204, A[42]);
  nand g2335 (n_2205, A[46], A[34]);
  nand g2338 (n_828, n_2205, n_2141, n_2078);
  xor g2339 (n_2208, A[40], A[44]);
  xor g2340 (n_816, n_2208, A[38]);
  nand g2344 (n_827, n_2014, n_1951, n_1821);
  xor g2346 (n_818, n_2212, n_813);
  nand g2349 (n_2215, A[36], n_813);
  nand g2350 (n_832, n_2213, n_2214, n_2215);
  xor g2351 (n_2216, n_814, n_815);
  xor g2352 (n_820, n_2216, n_816);
  nand g2353 (n_2217, n_814, n_815);
  nand g2354 (n_2218, n_816, n_815);
  nand g2355 (n_2219, n_814, n_816);
  nand g2356 (n_834, n_2217, n_2218, n_2219);
  xor g2357 (n_2220, n_817, n_818);
  xor g2358 (n_822, n_2220, n_819);
  nand g2359 (n_2221, n_817, n_818);
  nand g2360 (n_2222, n_819, n_818);
  nand g2361 (n_2223, n_817, n_819);
  nand g2362 (n_835, n_2221, n_2222, n_2223);
  xor g2363 (n_2224, n_820, n_821);
  xor g2364 (n_824, n_2224, n_822);
  nand g2365 (n_2225, n_820, n_821);
  nand g2366 (n_2226, n_822, n_821);
  nand g2367 (n_2227, n_820, n_822);
  nand g2368 (n_838, n_2225, n_2226, n_2227);
  xor g2369 (n_2228, n_823, n_824);
  xor g2370 (n_136, n_2228, n_825);
  nand g2371 (n_2229, n_823, n_824);
  nand g2372 (n_2230, n_825, n_824);
  nand g2373 (n_2231, n_823, n_825);
  nand g2374 (n_66, n_2229, n_2230, n_2231);
  xor g2381 (n_2236, A[35], A[41]);
  xor g2382 (n_830, n_2236, A[45]);
  nand g2385 (n_2239, A[35], A[45]);
  nand g2386 (n_842, n_1855, n_2046, n_2239);
  xor g2388 (n_831, n_1788, A[48]);
  nand g2390 (n_2242, A[48], A[37]);
  nand g2391 (n_2243, A[39], A[48]);
  nand g2392 (n_845, n_1789, n_2242, n_2243);
  xor g2393 (n_2244, n_827, n_828);
  xor g2394 (n_833, n_2244, n_801);
  nand g2395 (n_2245, n_827, n_828);
  nand g2396 (n_2246, n_801, n_828);
  nand g2397 (n_2247, n_827, n_801);
  nand g2398 (n_847, n_2245, n_2246, n_2247);
  xor g2399 (n_2248, n_830, n_831);
  xor g2400 (n_836, n_2248, n_832);
  nand g2401 (n_2249, n_830, n_831);
  nand g2402 (n_2250, n_832, n_831);
  nand g2403 (n_2251, n_830, n_832);
  nand g2404 (n_849, n_2249, n_2250, n_2251);
  xor g2405 (n_2252, n_833, n_834);
  xor g2406 (n_837, n_2252, n_835);
  nand g2407 (n_2253, n_833, n_834);
  nand g2408 (n_2254, n_835, n_834);
  nand g2409 (n_2255, n_833, n_835);
  nand g2410 (n_851, n_2253, n_2254, n_2255);
  xor g2411 (n_2256, n_836, n_837);
  xor g2412 (n_135, n_2256, n_838);
  nand g2413 (n_2257, n_836, n_837);
  nand g2414 (n_2258, n_838, n_837);
  nand g2415 (n_2259, n_836, n_838);
  nand g2416 (n_134, n_2257, n_2258, n_2259);
  xor g2419 (n_2260, A[46], A[42]);
  xor g2420 (n_844, n_2260, A[40]);
  nand g2424 (n_853, n_2078, n_1885, n_2015);
  xor g2425 (n_2264, A[44], A[38]);
  xor g2426 (n_843, n_2264, A[36]);
  nand g2429 (n_2267, A[44], A[36]);
  nand g2430 (n_854, n_1951, n_1757, n_2267);
  xor g2432 (n_846, n_2268, n_842);
  nand g2434 (n_2270, n_842, n_813);
  nand g2436 (n_858, n_2214, n_2270, n_2271);
  xor g2437 (n_2272, n_843, n_844);
  xor g2438 (n_848, n_2272, n_845);
  nand g2439 (n_2273, n_843, n_844);
  nand g2440 (n_2274, n_845, n_844);
  nand g2441 (n_2275, n_843, n_845);
  nand g2442 (n_859, n_2273, n_2274, n_2275);
  xor g2443 (n_2276, n_846, n_847);
  xor g2444 (n_850, n_2276, n_848);
  nand g2445 (n_2277, n_846, n_847);
  nand g2446 (n_2278, n_848, n_847);
  nand g2447 (n_2279, n_846, n_848);
  nand g2448 (n_862, n_2277, n_2278, n_2279);
  xor g2449 (n_2280, n_849, n_850);
  xor g2450 (n_65, n_2280, n_851);
  nand g2451 (n_2281, n_849, n_850);
  nand g2452 (n_2282, n_851, n_850);
  nand g2453 (n_2283, n_849, n_851);
  nand g2454 (n_64, n_2281, n_2282, n_2283);
  xor g2467 (n_2292, A[37], A[48]);
  xor g2468 (n_857, n_2292, n_853);
  nand g2470 (n_2294, n_853, A[48]);
  nand g2471 (n_2295, A[37], n_853);
  nand g2472 (n_869, n_2242, n_2294, n_2295);
  xor g2473 (n_2296, n_854, n_768);
  xor g2474 (n_860, n_2296, n_801);
  nand g2475 (n_2297, n_854, n_768);
  nand g2476 (n_2298, n_801, n_768);
  nand g2477 (n_2299, n_854, n_801);
  nand g2478 (n_870, n_2297, n_2298, n_2299);
  xor g2479 (n_2300, n_857, n_858);
  xor g2480 (n_861, n_2300, n_859);
  nand g2481 (n_2301, n_857, n_858);
  nand g2482 (n_2302, n_859, n_858);
  nand g2483 (n_2303, n_857, n_859);
  nand g2484 (n_873, n_2301, n_2302, n_2303);
  xor g2485 (n_2304, n_860, n_861);
  xor g2486 (n_133, n_2304, n_862);
  nand g2487 (n_2305, n_860, n_861);
  nand g2488 (n_2306, n_862, n_861);
  nand g2489 (n_2307, n_860, n_862);
  nand g2490 (n_63, n_2305, n_2306, n_2307);
  xor g2494 (n_867, n_1884, A[48]);
  nand g2498 (n_875, n_1885, n_2146, n_2079);
  nand g2504 (n_878, n_1951, n_2314, n_2315);
  xor g2505 (n_2316, n_782, n_813);
  xor g2506 (n_871, n_2316, n_867);
  nand g2507 (n_2317, n_782, n_813);
  nand g2508 (n_2318, n_867, n_813);
  nand g2509 (n_2319, n_782, n_867);
  nand g2510 (n_880, n_2317, n_2318, n_2319);
  xor g2511 (n_2320, n_868, n_869);
  xor g2512 (n_872, n_2320, n_870);
  nand g2513 (n_2321, n_868, n_869);
  nand g2514 (n_2322, n_870, n_869);
  nand g2515 (n_2323, n_868, n_870);
  nand g2516 (n_882, n_2321, n_2322, n_2323);
  xor g2517 (n_2324, n_871, n_872);
  xor g2518 (n_132, n_2324, n_873);
  nand g2519 (n_2325, n_871, n_872);
  nand g2520 (n_2326, n_873, n_872);
  nand g2521 (n_2327, n_871, n_873);
  nand g2522 (n_62, n_2325, n_2326, n_2327);
  xor g2535 (n_2336, A[46], n_875);
  xor g2536 (n_879, n_2336, n_768);
  nand g2537 (n_2337, A[46], n_875);
  nand g2538 (n_2338, n_768, n_875);
  nand g2539 (n_2339, A[46], n_768);
  nand g2540 (n_889, n_2337, n_2338, n_2339);
  xor g2541 (n_2340, n_801, n_878);
  xor g2542 (n_881, n_2340, n_879);
  nand g2543 (n_2341, n_801, n_878);
  nand g2544 (n_2342, n_879, n_878);
  nand g2545 (n_2343, n_801, n_879);
  nand g2546 (n_891, n_2341, n_2342, n_2343);
  xor g2547 (n_2344, n_880, n_881);
  xor g2548 (n_131, n_2344, n_882);
  nand g2549 (n_2345, n_880, n_881);
  nand g2550 (n_2346, n_882, n_881);
  nand g2551 (n_2347, n_880, n_882);
  nand g2552 (n_61, n_2345, n_2346, n_2347);
  nand g2565 (n_2355, A[44], n_782);
  nand g2566 (n_896, n_2314, n_2354, n_2355);
  xor g2567 (n_2356, n_813, n_867);
  xor g2568 (n_890, n_2356, n_888);
  nand g2570 (n_2358, n_888, n_867);
  nand g2571 (n_2359, n_813, n_888);
  nand g2572 (n_898, n_2318, n_2358, n_2359);
  xor g2573 (n_2360, n_889, n_890);
  xor g2574 (n_130, n_2360, n_891);
  nand g2575 (n_2361, n_889, n_890);
  nand g2576 (n_2362, n_891, n_890);
  nand g2577 (n_2363, n_889, n_891);
  nand g2578 (n_129, n_2361, n_2362, n_2363);
  xor g2586 (n_895, n_2116, A[46]);
  nand g2588 (n_2370, A[46], A[45]);
  nand g2589 (n_2371, A[41], A[46]);
  nand g2590 (n_903, n_2046, n_2370, n_2371);
  xor g2591 (n_2372, n_875, n_801);
  xor g2592 (n_897, n_2372, n_895);
  nand g2593 (n_2373, n_875, n_801);
  nand g2594 (n_2374, n_895, n_801);
  nand g2595 (n_2375, n_875, n_895);
  nand g2596 (n_905, n_2373, n_2374, n_2375);
  xor g2597 (n_2376, n_896, n_897);
  xor g2598 (n_60, n_2376, n_898);
  nand g2599 (n_2377, n_896, n_897);
  nand g2600 (n_2378, n_898, n_897);
  nand g2601 (n_2379, n_896, n_898);
  nand g2602 (n_128, n_2377, n_2378, n_2379);
  xor g2606 (n_902, n_2260, A[44]);
  nand g2610 (n_907, n_2078, n_2013, n_1949);
  xor g2612 (n_904, n_2268, n_902);
  nand g2614 (n_2386, n_902, n_813);
  nand g2616 (n_910, n_2214, n_2386, n_2387);
  xor g2617 (n_2388, n_903, n_904);
  xor g2618 (n_59, n_2388, n_905);
  nand g2619 (n_2389, n_903, n_904);
  nand g2620 (n_2390, n_905, n_904);
  nand g2621 (n_2391, n_903, n_905);
  nand g2622 (n_127, n_2389, n_2390, n_2391);
  xor g2629 (n_2396, A[45], A[48]);
  xor g2630 (n_909, n_2396, n_907);
  nand g2631 (n_2397, A[45], A[48]);
  nand g2632 (n_2398, n_907, A[48]);
  nand g2633 (n_2399, A[45], n_907);
  nand g2634 (n_915, n_2397, n_2398, n_2399);
  xor g2635 (n_2400, n_801, n_909);
  xor g2636 (n_58, n_2400, n_910);
  nand g2637 (n_2401, n_801, n_909);
  nand g2638 (n_2402, n_910, n_909);
  nand g2639 (n_2403, n_801, n_910);
  nand g2640 (n_126, n_2401, n_2402, n_2403);
  nand g2648 (n_918, n_2013, n_2406, n_2407);
  xor g2649 (n_2408, n_813, n_914);
  xor g2650 (n_57, n_2408, n_915);
  nand g2651 (n_2409, n_813, n_914);
  nand g2652 (n_2410, n_915, n_914);
  nand g2653 (n_2411, n_813, n_915);
  nand g2654 (n_125, n_2409, n_2410, n_2411);
  xor g2656 (n_917, n_2172, A[45]);
  nand g2660 (n_921, n_2173, n_2045, n_2181);
  xor g2661 (n_2416, A[48], n_917);
  xor g2662 (n_56, n_2416, n_918);
  nand g2663 (n_2417, A[48], n_917);
  nand g2664 (n_2418, n_918, n_917);
  nand g2665 (n_2419, A[48], n_918);
  nand g2666 (n_124, n_2417, n_2418, n_2419);
  nand g2673 (n_2423, A[48], n_921);
  nand g2674 (n_123, n_2421, n_2422, n_2423);
  xor g2676 (n_54, n_2172, A[46]);
  nand g2678 (n_2426, A[46], A[47]);
  nand g2680 (n_122, n_2173, n_2426, n_2427);
  nor g11 (n_2443, A[2], A[0]);
  nor g13 (n_2439, A[1], A[3]);
  nor g15 (n_2449, A[2], n_184);
  nand g16 (n_2444, A[2], n_184);
  nor g17 (n_2445, n_114, n_183);
  nand g18 (n_2446, n_114, n_183);
  nor g19 (n_2455, n_113, n_182);
  nand g20 (n_2450, n_113, n_182);
  nor g21 (n_2451, n_112, n_181);
  nand g22 (n_2452, n_112, n_181);
  nor g23 (n_2461, n_111, n_180);
  nand g24 (n_2456, n_111, n_180);
  nor g25 (n_2457, n_110, n_179);
  nand g26 (n_2458, n_110, n_179);
  nor g27 (n_2467, n_109, n_178);
  nand g28 (n_2462, n_109, n_178);
  nor g29 (n_2463, n_108, n_177);
  nand g30 (n_2464, n_108, n_177);
  nor g31 (n_2473, n_107, n_176);
  nand g32 (n_2468, n_107, n_176);
  nor g33 (n_2469, n_106, n_175);
  nand g34 (n_2470, n_106, n_175);
  nor g35 (n_2479, n_105, n_174);
  nand g36 (n_2474, n_105, n_174);
  nor g37 (n_2475, n_104, n_173);
  nand g38 (n_2476, n_104, n_173);
  nor g39 (n_2485, n_103, n_172);
  nand g40 (n_2480, n_103, n_172);
  nor g41 (n_2481, n_102, n_171);
  nand g42 (n_2482, n_102, n_171);
  nor g43 (n_2491, n_101, n_170);
  nand g44 (n_2486, n_101, n_170);
  nor g45 (n_2487, n_100, n_169);
  nand g46 (n_2488, n_100, n_169);
  nor g47 (n_2497, n_99, n_168);
  nand g48 (n_2492, n_99, n_168);
  nor g49 (n_2493, n_98, n_167);
  nand g50 (n_2494, n_98, n_167);
  nor g51 (n_2503, n_97, n_166);
  nand g52 (n_2498, n_97, n_166);
  nor g53 (n_2499, n_96, n_165);
  nand g54 (n_2500, n_96, n_165);
  nor g55 (n_2509, n_95, n_164);
  nand g56 (n_2504, n_95, n_164);
  nor g57 (n_2505, n_94, n_163);
  nand g58 (n_2506, n_94, n_163);
  nor g59 (n_2515, n_93, n_162);
  nand g60 (n_2510, n_93, n_162);
  nor g61 (n_2511, n_92, n_161);
  nand g62 (n_2512, n_92, n_161);
  nor g63 (n_2521, n_91, n_160);
  nand g64 (n_2516, n_91, n_160);
  nor g65 (n_2517, n_90, n_159);
  nand g66 (n_2518, n_90, n_159);
  nor g67 (n_2527, n_89, n_158);
  nand g68 (n_2522, n_89, n_158);
  nor g69 (n_2523, n_88, n_157);
  nand g70 (n_2524, n_88, n_157);
  nor g71 (n_2533, n_87, n_156);
  nand g72 (n_2528, n_87, n_156);
  nor g73 (n_2529, n_86, n_155);
  nand g74 (n_2530, n_86, n_155);
  nor g75 (n_2539, n_85, n_154);
  nand g76 (n_2534, n_85, n_154);
  nor g77 (n_2535, n_84, n_153);
  nand g78 (n_2536, n_84, n_153);
  nor g79 (n_2545, n_83, n_152);
  nand g80 (n_2540, n_83, n_152);
  nor g81 (n_2541, n_82, n_151);
  nand g82 (n_2542, n_82, n_151);
  nor g83 (n_2551, n_81, n_150);
  nand g84 (n_2546, n_81, n_150);
  nor g85 (n_2547, n_80, n_149);
  nand g86 (n_2548, n_80, n_149);
  nor g87 (n_2557, n_79, n_148);
  nand g88 (n_2552, n_79, n_148);
  nor g89 (n_2553, n_78, n_147);
  nand g90 (n_2554, n_78, n_147);
  nor g91 (n_2563, n_77, n_146);
  nand g92 (n_2558, n_77, n_146);
  nor g93 (n_2559, n_76, n_145);
  nand g94 (n_2560, n_76, n_145);
  nor g95 (n_2569, n_75, n_144);
  nand g96 (n_2564, n_75, n_144);
  nor g97 (n_2565, n_74, n_143);
  nand g98 (n_2566, n_74, n_143);
  nor g99 (n_2575, n_73, n_142);
  nand g100 (n_2570, n_73, n_142);
  nor g101 (n_2571, n_72, n_141);
  nand g102 (n_2572, n_72, n_141);
  nor g103 (n_2581, n_71, n_140);
  nand g104 (n_2576, n_71, n_140);
  nor g105 (n_2577, n_70, n_139);
  nand g106 (n_2578, n_70, n_139);
  nor g107 (n_2587, n_69, n_138);
  nand g108 (n_2582, n_69, n_138);
  nor g109 (n_2583, n_68, n_137);
  nand g110 (n_2584, n_68, n_137);
  nor g111 (n_2593, n_67, n_136);
  nand g112 (n_2588, n_67, n_136);
  nor g113 (n_2589, n_66, n_135);
  nand g114 (n_2590, n_66, n_135);
  nor g115 (n_2599, n_65, n_134);
  nand g116 (n_2594, n_65, n_134);
  nor g117 (n_2595, n_64, n_133);
  nand g118 (n_2596, n_64, n_133);
  nor g119 (n_2605, n_63, n_132);
  nand g120 (n_2600, n_63, n_132);
  nor g121 (n_2601, n_62, n_131);
  nand g122 (n_2602, n_62, n_131);
  nor g123 (n_2611, n_61, n_130);
  nand g124 (n_2606, n_61, n_130);
  nor g125 (n_2607, n_60, n_129);
  nand g126 (n_2608, n_60, n_129);
  nor g127 (n_2617, n_59, n_128);
  nand g128 (n_2612, n_59, n_128);
  nor g129 (n_2613, n_58, n_127);
  nand g130 (n_2614, n_58, n_127);
  nor g131 (n_2623, n_57, n_126);
  nand g132 (n_2618, n_57, n_126);
  nor g133 (n_2619, n_56, n_125);
  nand g134 (n_2620, n_56, n_125);
  nor g135 (n_2629, n_55, n_124);
  nand g136 (n_2624, n_55, n_124);
  nor g137 (n_2625, n_54, n_123);
  nand g138 (n_2626, n_54, n_123);
  nor g148 (n_2441, n_929, n_2439);
  nor g152 (n_2447, n_2444, n_2445);
  nor g155 (n_2646, n_2449, n_2445);
  nor g156 (n_2453, n_2450, n_2451);
  nor g159 (n_2640, n_2455, n_2451);
  nor g160 (n_2459, n_2456, n_2457);
  nor g163 (n_2653, n_2461, n_2457);
  nor g164 (n_2465, n_2462, n_2463);
  nor g167 (n_2647, n_2467, n_2463);
  nor g168 (n_2471, n_2468, n_2469);
  nor g171 (n_2660, n_2473, n_2469);
  nor g172 (n_2477, n_2474, n_2475);
  nor g175 (n_2654, n_2479, n_2475);
  nor g176 (n_2483, n_2480, n_2481);
  nor g179 (n_2667, n_2485, n_2481);
  nor g180 (n_2489, n_2486, n_2487);
  nor g183 (n_2661, n_2491, n_2487);
  nor g184 (n_2495, n_2492, n_2493);
  nor g187 (n_2674, n_2497, n_2493);
  nor g188 (n_2501, n_2498, n_2499);
  nor g191 (n_2668, n_2503, n_2499);
  nor g192 (n_2507, n_2504, n_2505);
  nor g195 (n_2681, n_2509, n_2505);
  nor g196 (n_2513, n_2510, n_2511);
  nor g199 (n_2675, n_2515, n_2511);
  nor g200 (n_2519, n_2516, n_2517);
  nor g203 (n_2688, n_2521, n_2517);
  nor g204 (n_2525, n_2522, n_2523);
  nor g207 (n_2682, n_2527, n_2523);
  nor g208 (n_2531, n_2528, n_2529);
  nor g211 (n_2695, n_2533, n_2529);
  nor g212 (n_2537, n_2534, n_2535);
  nor g215 (n_2689, n_2539, n_2535);
  nor g216 (n_2543, n_2540, n_2541);
  nor g219 (n_2702, n_2545, n_2541);
  nor g220 (n_2549, n_2546, n_2547);
  nor g223 (n_2696, n_2551, n_2547);
  nor g224 (n_2555, n_2552, n_2553);
  nor g227 (n_2709, n_2557, n_2553);
  nor g228 (n_2561, n_2558, n_2559);
  nor g231 (n_2703, n_2563, n_2559);
  nor g232 (n_2567, n_2564, n_2565);
  nor g235 (n_2716, n_2569, n_2565);
  nor g236 (n_2573, n_2570, n_2571);
  nor g239 (n_2710, n_2575, n_2571);
  nor g240 (n_2579, n_2576, n_2577);
  nor g243 (n_2723, n_2581, n_2577);
  nor g244 (n_2585, n_2582, n_2583);
  nor g247 (n_2717, n_2587, n_2583);
  nor g248 (n_2591, n_2588, n_2589);
  nor g251 (n_2730, n_2593, n_2589);
  nor g252 (n_2597, n_2594, n_2595);
  nor g255 (n_2724, n_2599, n_2595);
  nor g256 (n_2603, n_2600, n_2601);
  nor g259 (n_2737, n_2605, n_2601);
  nor g260 (n_2609, n_2606, n_2607);
  nor g263 (n_2731, n_2611, n_2607);
  nor g264 (n_2615, n_2612, n_2613);
  nor g267 (n_2744, n_2617, n_2613);
  nor g268 (n_2621, n_2618, n_2619);
  nor g271 (n_2738, n_2623, n_2619);
  nor g272 (n_2627, n_2624, n_2625);
  nor g275 (n_2751, n_2629, n_2625);
  nor g276 (n_2633, n_2630, n_2631);
  nor g279 (n_2745, n_2635, n_2631);
  nand g286 (n_2752, n_2646, n_2640);
  nand g291 (n_2762, n_2653, n_2647);
  nand g296 (n_2757, n_2660, n_2654);
  nand g301 (n_2768, n_2667, n_2661);
  nand g306 (n_2763, n_2674, n_2668);
  nand g311 (n_2774, n_2681, n_2675);
  nand g316 (n_2769, n_2688, n_2682);
  nand g321 (n_2780, n_2695, n_2689);
  nand g326 (n_2775, n_2702, n_2696);
  nand g331 (n_2786, n_2709, n_2703);
  nand g336 (n_2781, n_2716, n_2710);
  nand g341 (n_2792, n_2723, n_2717);
  nand g346 (n_2787, n_2730, n_2724);
  nand g351 (n_2798, n_2737, n_2731);
  nand g356 (n_2793, n_2744, n_2738);
  nand g361 (n_2862, n_2751, n_2745);
  nand g364 (n_2800, n_2755, n_2756);
  nor g365 (n_2760, n_2757, n_2758);
  nor g368 (n_2799, n_2762, n_2757);
  nor g369 (n_2766, n_2763, n_2764);
  nor g372 (n_2809, n_2768, n_2763);
  nor g373 (n_2772, n_2769, n_2770);
  nor g376 (n_2803, n_2774, n_2769);
  nor g377 (n_2778, n_2775, n_2776);
  nor g380 (n_2816, n_2780, n_2775);
  nor g381 (n_2784, n_2781, n_2782);
  nor g384 (n_2810, n_2786, n_2781);
  nor g385 (n_2790, n_2787, n_2788);
  nor g388 (n_2823, n_2792, n_2787);
  nor g389 (n_2796, n_2793, n_2794);
  nor g392 (n_2817, n_2798, n_2793);
  nand g393 (n_2802, n_2799, n_2800);
  nand g394 (n_2825, n_2801, n_2802);
  nand g2691 (n_2824, n_2809, n_2803);
  nand g2696 (n_2834, n_2816, n_2810);
  nand g2701 (n_2829, n_2823, n_2817);
  nand g2704 (n_2836, n_2827, n_2828);
  nor g2705 (n_2832, n_2829, n_2830);
  nor g2708 (n_2835, n_2834, n_2829);
  nand g2709 (n_2838, n_2835, n_2836);
  nand g2710 (n_2863, n_2837, n_2838);
  nand g2713 (n_2843, n_2830, n_2840);
  nand g2714 (n_2841, n_2809, n_2825);
  nand g2715 (n_2849, n_2804, n_2841);
  nand g2716 (n_2842, n_2816, n_2836);
  nand g2717 (n_2854, n_2811, n_2842);
  nand g2718 (n_2844, n_2823, n_2843);
  nand g2719 (n_2859, n_2818, n_2844);
  nand g2722 (n_2869, n_2758, n_2846);
  nand g2725 (n_2872, n_2764, n_2848);
  nand g2728 (n_2875, n_2770, n_2851);
  nand g2731 (n_2878, n_2776, n_2853);
  nand g2734 (n_2881, n_2782, n_2856);
  nand g2737 (n_2884, n_2788, n_2858);
  nand g2740 (n_2887, n_2794, n_2861);
  nand g2743 (n_2973, n_2865, n_2866);
  nand g2745 (n_2894, n_2641, n_2867);
  nand g2746 (n_2868, n_2653, n_2800);
  nand g2747 (n_2899, n_2648, n_2868);
  nand g2748 (n_2870, n_2660, n_2869);
  nand g2749 (n_2904, n_2655, n_2870);
  nand g2750 (n_2871, n_2667, n_2825);
  nand g2751 (n_2909, n_2662, n_2871);
  nand g2752 (n_2873, n_2674, n_2872);
  nand g2753 (n_2914, n_2669, n_2873);
  nand g2754 (n_2874, n_2681, n_2849);
  nand g2755 (n_2919, n_2676, n_2874);
  nand g2756 (n_2876, n_2688, n_2875);
  nand g2757 (n_2924, n_2683, n_2876);
  nand g2758 (n_2877, n_2695, n_2836);
  nand g2759 (n_2929, n_2690, n_2877);
  nand g2760 (n_2879, n_2702, n_2878);
  nand g2761 (n_2934, n_2697, n_2879);
  nand g2762 (n_2880, n_2709, n_2854);
  nand g2763 (n_2939, n_2704, n_2880);
  nand g2764 (n_2882, n_2716, n_2881);
  nand g2765 (n_2944, n_2711, n_2882);
  nand g2766 (n_2883, n_2723, n_2843);
  nand g2767 (n_2949, n_2718, n_2883);
  nand g2768 (n_2885, n_2730, n_2884);
  nand g2769 (n_2954, n_2725, n_2885);
  nand g2770 (n_2886, n_2737, n_2859);
  nand g2771 (n_2959, n_2732, n_2886);
  nand g2772 (n_2888, n_2744, n_2887);
  nand g2773 (n_2964, n_2739, n_2888);
  nand g2774 (n_2889, n_2751, n_2863);
  nand g2775 (n_2969, n_2746, n_2889);
  nand g2781 (n_2983, n_2444, n_2893);
  nand g2784 (n_2987, n_2450, n_2896);
  nand g2787 (n_2991, n_2456, n_2898);
  nand g2790 (n_2995, n_2462, n_2901);
  nand g2793 (n_2999, n_2468, n_2903);
  nand g2796 (n_3003, n_2474, n_2906);
  nand g2799 (n_3007, n_2480, n_2908);
  nand g2802 (n_3011, n_2486, n_2911);
  nand g2805 (n_3015, n_2492, n_2913);
  nand g2808 (n_3019, n_2498, n_2916);
  nand g2811 (n_3023, n_2504, n_2918);
  nand g2814 (n_3027, n_2510, n_2921);
  nand g2817 (n_3031, n_2516, n_2923);
  nand g2820 (n_3035, n_2522, n_2926);
  nand g2823 (n_3039, n_2528, n_2928);
  nand g2826 (n_3043, n_2534, n_2931);
  nand g2829 (n_3047, n_2540, n_2933);
  nand g2832 (n_3051, n_2546, n_2936);
  nand g2835 (n_3055, n_2552, n_2938);
  nand g2838 (n_3059, n_2558, n_2941);
  nand g2841 (n_3063, n_2564, n_2943);
  nand g2844 (n_3067, n_2570, n_2946);
  nand g2847 (n_3071, n_2576, n_2948);
  nand g2850 (n_3075, n_2582, n_2951);
  nand g2853 (n_3079, n_2588, n_2953);
  nand g2856 (n_3083, n_2594, n_2956);
  nand g2859 (n_3087, n_2600, n_2958);
  nand g2862 (n_3091, n_2606, n_2961);
  nand g2865 (n_3095, n_2612, n_2963);
  nand g2868 (n_3099, n_2618, n_2966);
  nand g2871 (n_3103, n_2624, n_2968);
  nand g2874 (n_3107, n_2630, n_2971);
  xnor g2887 (Z[5], n_2983, n_2984);
  xnor g2889 (Z[6], n_2894, n_2985);
  xnor g2892 (Z[7], n_2987, n_2988);
  xnor g2894 (Z[8], n_2800, n_2989);
  xnor g2897 (Z[9], n_2991, n_2992);
  xnor g2899 (Z[10], n_2899, n_2993);
  xnor g2902 (Z[11], n_2995, n_2996);
  xnor g2904 (Z[12], n_2869, n_2997);
  xnor g2907 (Z[13], n_2999, n_3000);
  xnor g2909 (Z[14], n_2904, n_3001);
  xnor g2912 (Z[15], n_3003, n_3004);
  xnor g2914 (Z[16], n_2825, n_3005);
  xnor g2917 (Z[17], n_3007, n_3008);
  xnor g2919 (Z[18], n_2909, n_3009);
  xnor g2922 (Z[19], n_3011, n_3012);
  xnor g2924 (Z[20], n_2872, n_3013);
  xnor g2927 (Z[21], n_3015, n_3016);
  xnor g2929 (Z[22], n_2914, n_3017);
  xnor g2932 (Z[23], n_3019, n_3020);
  xnor g2934 (Z[24], n_2849, n_3021);
  xnor g2937 (Z[25], n_3023, n_3024);
  xnor g2939 (Z[26], n_2919, n_3025);
  xnor g2942 (Z[27], n_3027, n_3028);
  xnor g2944 (Z[28], n_2875, n_3029);
  xnor g2947 (Z[29], n_3031, n_3032);
  xnor g2949 (Z[30], n_2924, n_3033);
  xnor g2952 (Z[31], n_3035, n_3036);
  xnor g2954 (Z[32], n_2836, n_3037);
  xnor g2957 (Z[33], n_3039, n_3040);
  xnor g2959 (Z[34], n_2929, n_3041);
  xnor g2962 (Z[35], n_3043, n_3044);
  xnor g2964 (Z[36], n_2878, n_3045);
  xnor g2967 (Z[37], n_3047, n_3048);
  xnor g2969 (Z[38], n_2934, n_3049);
  xnor g2972 (Z[39], n_3051, n_3052);
  xnor g2974 (Z[40], n_2854, n_3053);
  xnor g2977 (Z[41], n_3055, n_3056);
  xnor g2979 (Z[42], n_2939, n_3057);
  xnor g2982 (Z[43], n_3059, n_3060);
  xnor g2984 (Z[44], n_2881, n_3061);
  xnor g2987 (Z[45], n_3063, n_3064);
  xnor g2989 (Z[46], n_2944, n_3065);
  xnor g2992 (Z[47], n_3067, n_3068);
  xnor g2994 (Z[48], n_2843, n_3069);
  xnor g2997 (Z[49], n_3071, n_3072);
  xnor g2999 (Z[50], n_2949, n_3073);
  xnor g3002 (Z[51], n_3075, n_3076);
  xnor g3004 (Z[52], n_2884, n_3077);
  xnor g3007 (Z[53], n_3079, n_3080);
  xnor g3009 (Z[54], n_2954, n_3081);
  xnor g3012 (Z[55], n_3083, n_3084);
  xnor g3014 (Z[56], n_2859, n_3085);
  xnor g3017 (Z[57], n_3087, n_3088);
  xnor g3019 (Z[58], n_2959, n_3089);
  xnor g3022 (Z[59], n_3091, n_3092);
  xnor g3024 (Z[60], n_2887, n_3093);
  xnor g3027 (Z[61], n_3095, n_3096);
  xnor g3029 (Z[62], n_2964, n_3097);
  xnor g3032 (Z[63], n_3099, n_3100);
  xnor g3034 (Z[64], n_2863, n_3101);
  xnor g3037 (Z[65], n_3103, n_3104);
  xnor g3039 (Z[66], n_2969, n_3105);
  xnor g3042 (Z[67], n_3107, n_3108);
  or g3057 (n_266, wc, wc0, n_114);
  not gc0 (wc0, n_929);
  not gc (wc, n_943);
  or g3058 (n_275, wc1, wc2, n_260);
  not gc2 (wc2, n_943);
  not gc1 (wc1, n_962);
  or g3059 (n_288, wc3, n_265, n_260);
  not gc3 (wc3, n_990);
  or g3060 (n_305, wc4, wc5, n_265);
  not gc5 (wc5, n_1025);
  not gc4 (wc4, n_1026);
  or g3061 (n_327, wc6, wc7, n_265);
  not gc7 (wc7, n_1073);
  not gc6 (wc6, n_1074);
  or g3062 (n_374, wc8, wc9, n_260);
  not gc9 (wc9, n_1074);
  not gc8 (wc8, n_1121);
  or g3063 (n_402, wc10, wc11, n_265);
  not gc11 (wc11, n_1250);
  not gc10 (wc10, n_1251);
  or g3064 (n_428, wc12, wc13, n_274);
  not gc13 (wc13, n_1190);
  not gc12 (wc12, n_1314);
  or g3065 (n_456, wc14, wc15, n_287);
  not gc15 (wc15, n_1254);
  not gc14 (wc14, n_1378);
  or g3066 (n_484, wc16, wc17, n_304);
  not gc17 (wc17, n_1183);
  not gc16 (wc16, n_1442);
  or g3067 (n_512, wc18, wc19, n_325);
  not gc19 (wc19, n_1247);
  not gc18 (wc18, n_1506);
  or g3068 (n_540, wc20, wc21, n_350);
  not gc21 (wc21, n_1311);
  not gc20 (wc20, n_1570);
  xnor g3069 (n_2172, A[49], A[47]);
  or g3070 (n_2173, wc22, A[49]);
  not gc22 (wc22, A[47]);
  or g3071 (n_2175, wc23, A[49]);
  not gc23 (wc23, A[43]);
  xnor g3072 (n_2212, A[48], A[36]);
  or g3073 (n_2213, wc24, A[48]);
  not gc24 (wc24, A[36]);
  xnor g3074 (n_868, n_2264, A[46]);
  or g3075 (n_2314, wc25, A[46]);
  not gc25 (wc25, A[44]);
  or g3076 (n_2315, wc26, A[46]);
  not gc26 (wc26, A[38]);
  xnor g3078 (n_914, n_2012, A[48]);
  or g3079 (n_2406, wc27, A[48]);
  not gc27 (wc27, A[44]);
  or g3080 (n_2407, wc28, A[48]);
  not gc28 (wc28, A[46]);
  or g3081 (n_2181, wc29, A[49]);
  not gc29 (wc29, A[45]);
  or g3083 (n_2421, A[46], wc30);
  not gc30 (wc30, A[48]);
  or g3084 (n_2427, wc31, A[49]);
  not gc31 (wc31, A[46]);
  and g3085 (n_2631, wc32, A[49]);
  not gc32 (wc32, A[48]);
  or g3086 (n_2632, wc33, A[49]);
  not gc33 (wc33, A[48]);
  or g3087 (n_119, wc34, wc35, n_265);
  not gc35 (wc35, n_1130);
  not gc34 (wc34, n_1131);
  or g3088 (n_2271, A[48], wc36);
  not gc36 (wc36, n_842);
  xnor g3089 (n_888, n_2012, n_782);
  or g3090 (n_2354, A[46], wc37);
  not gc37 (wc37, n_782);
  or g3091 (n_2387, A[48], wc38);
  not gc38 (wc38, n_902);
  and g3092 (n_2638, wc39, n_925);
  not gc39 (wc39, n_2441);
  or g3094 (n_2977, n_2443, wc40);
  not gc40 (wc40, n_929);
  or g3095 (n_2980, n_2439, wc41);
  not gc41 (wc41, n_925);
  xnor g3096 (n_2180, A[49], A[45]);
  or g3097 (n_2183, wc42, A[49]);
  not gc42 (wc42, A[39]);
  or g3098 (n_2214, A[48], wc43);
  not gc43 (wc43, n_813);
  xnor g3099 (n_2268, n_813, A[48]);
  xnor g3100 (n_55, n_2076, n_921);
  or g3101 (n_2422, A[46], wc44);
  not gc44 (wc44, n_921);
  and g3102 (n_2635, A[48], wc45);
  not gc45 (wc45, n_122);
  or g3103 (n_2630, A[48], wc46);
  not gc46 (wc46, n_122);
  or g3104 (n_2981, wc47, n_2449);
  not gc47 (wc47, n_2444);
  or g3105 (n_3108, wc48, n_2631);
  not gc48 (wc48, n_2632);
  and g3106 (n_2641, wc49, n_2446);
  not gc49 (wc49, n_2447);
  not g3107 (Z[2], n_2977);
  or g3108 (n_2984, wc50, n_2445);
  not gc50 (wc50, n_2446);
  or g3109 (n_2985, wc51, n_2455);
  not gc51 (wc51, n_2450);
  and g3110 (n_2643, wc52, n_2452);
  not gc52 (wc52, n_2453);
  and g3111 (n_2748, n_2632, wc53);
  not gc53 (wc53, n_2633);
  or g3114 (n_2988, wc54, n_2451);
  not gc54 (wc54, n_2452);
  or g3115 (n_3105, wc55, n_2635);
  not gc55 (wc55, n_2630);
  and g3116 (n_2648, wc56, n_2458);
  not gc56 (wc56, n_2459);
  and g3117 (n_2644, wc57, n_2640);
  not gc57 (wc57, n_2641);
  or g3118 (n_2867, n_2638, wc58);
  not gc58 (wc58, n_2646);
  or g3119 (n_2893, n_2449, n_2638);
  xor g3120 (Z[3], n_929, n_2980);
  xor g3121 (Z[4], n_2638, n_2981);
  or g3122 (n_2989, wc59, n_2461);
  not gc59 (wc59, n_2456);
  or g3123 (n_2992, wc60, n_2457);
  not gc60 (wc60, n_2458);
  and g3124 (n_2746, wc61, n_2626);
  not gc61 (wc61, n_2627);
  and g3125 (n_2755, wc62, n_2643);
  not gc62 (wc62, n_2644);
  or g3126 (n_2756, n_2752, n_2638);
  or g3127 (n_2993, wc63, n_2467);
  not gc63 (wc63, n_2462);
  or g3128 (n_3101, wc64, n_2629);
  not gc64 (wc64, n_2624);
  or g3129 (n_3104, wc65, n_2625);
  not gc65 (wc65, n_2626);
  and g3130 (n_2650, wc66, n_2464);
  not gc66 (wc66, n_2465);
  and g3131 (n_2655, wc67, n_2470);
  not gc67 (wc67, n_2471);
  and g3132 (n_2749, wc68, n_2745);
  not gc68 (wc68, n_2746);
  or g3133 (n_2896, wc69, n_2455);
  not gc69 (wc69, n_2894);
  or g3134 (n_2996, wc70, n_2463);
  not gc70 (wc70, n_2464);
  or g3135 (n_2997, wc71, n_2473);
  not gc71 (wc71, n_2468);
  or g3136 (n_3000, wc72, n_2469);
  not gc72 (wc72, n_2470);
  or g3137 (n_3100, wc73, n_2619);
  not gc73 (wc73, n_2620);
  and g3138 (n_2657, wc74, n_2476);
  not gc74 (wc74, n_2477);
  and g3139 (n_2739, wc75, n_2614);
  not gc75 (wc75, n_2615);
  and g3140 (n_2741, wc76, n_2620);
  not gc76 (wc76, n_2621);
  and g3141 (n_2651, wc77, n_2647);
  not gc77 (wc77, n_2648);
  and g3142 (n_2865, wc78, n_2748);
  not gc78 (wc78, n_2749);
  or g3143 (n_2898, wc79, n_2461);
  not gc79 (wc79, n_2800);
  or g3144 (n_3001, wc80, n_2479);
  not gc80 (wc80, n_2474);
  or g3145 (n_3004, wc81, n_2475);
  not gc81 (wc81, n_2476);
  or g3146 (n_3093, wc82, n_2617);
  not gc82 (wc82, n_2612);
  or g3147 (n_3096, wc83, n_2613);
  not gc83 (wc83, n_2614);
  or g3148 (n_3097, wc84, n_2623);
  not gc84 (wc84, n_2618);
  and g3149 (n_2662, wc85, n_2482);
  not gc85 (wc85, n_2483);
  and g3150 (n_2664, wc86, n_2488);
  not gc86 (wc86, n_2489);
  and g3151 (n_2758, wc87, n_2650);
  not gc87 (wc87, n_2651);
  and g3152 (n_2658, wc88, n_2654);
  not gc88 (wc88, n_2655);
  and g3153 (n_2742, wc89, n_2738);
  not gc89 (wc89, n_2739);
  or g3154 (n_2846, wc90, n_2762);
  not gc90 (wc90, n_2800);
  or g3155 (n_3005, wc91, n_2485);
  not gc91 (wc91, n_2480);
  or g3156 (n_3008, wc92, n_2481);
  not gc92 (wc92, n_2482);
  or g3157 (n_3009, wc93, n_2491);
  not gc93 (wc93, n_2486);
  or g3158 (n_3012, wc94, n_2487);
  not gc94 (wc94, n_2488);
  or g3159 (n_3013, wc95, n_2497);
  not gc95 (wc95, n_2492);
  or g3160 (n_3092, wc96, n_2607);
  not gc96 (wc96, n_2608);
  and g3161 (n_2669, wc97, n_2494);
  not gc97 (wc97, n_2495);
  and g3162 (n_2732, wc98, n_2602);
  not gc98 (wc98, n_2603);
  and g3163 (n_2734, wc99, n_2608);
  not gc99 (wc99, n_2609);
  and g3164 (n_2759, wc100, n_2657);
  not gc100 (wc100, n_2658);
  and g3165 (n_2665, wc101, n_2661);
  not gc101 (wc101, n_2662);
  and g3166 (n_2795, wc102, n_2741);
  not gc102 (wc102, n_2742);
  or g3167 (n_2901, wc103, n_2467);
  not gc103 (wc103, n_2899);
  or g3168 (n_3016, wc104, n_2493);
  not gc104 (wc104, n_2494);
  or g3169 (n_3017, wc105, n_2503);
  not gc105 (wc105, n_2498);
  or g3170 (n_3085, wc106, n_2605);
  not gc106 (wc106, n_2600);
  or g3171 (n_3088, wc107, n_2601);
  not gc107 (wc107, n_2602);
  or g3172 (n_3089, wc108, n_2611);
  not gc108 (wc108, n_2606);
  and g3173 (n_2671, wc109, n_2500);
  not gc109 (wc109, n_2501);
  and g3174 (n_2676, wc110, n_2506);
  not gc110 (wc110, n_2507);
  and g3175 (n_2678, wc111, n_2512);
  not gc111 (wc111, n_2513);
  and g3176 (n_2683, wc112, n_2518);
  not gc112 (wc112, n_2519);
  and g3177 (n_2685, wc113, n_2524);
  not gc113 (wc113, n_2525);
  and g3178 (n_2690, wc114, n_2530);
  not gc114 (wc114, n_2531);
  and g3179 (n_2692, wc115, n_2536);
  not gc115 (wc115, n_2537);
  and g3180 (n_2697, wc116, n_2542);
  not gc116 (wc116, n_2543);
  and g3181 (n_2699, wc117, n_2548);
  not gc117 (wc117, n_2549);
  and g3182 (n_2704, wc118, n_2554);
  not gc118 (wc118, n_2555);
  and g3183 (n_2706, wc119, n_2560);
  not gc119 (wc119, n_2561);
  and g3184 (n_2711, wc120, n_2566);
  not gc120 (wc120, n_2567);
  and g3185 (n_2713, wc121, n_2572);
  not gc121 (wc121, n_2573);
  and g3186 (n_2718, wc122, n_2578);
  not gc122 (wc122, n_2579);
  and g3187 (n_2764, wc123, n_2664);
  not gc123 (wc123, n_2665);
  and g3188 (n_2735, wc124, n_2731);
  not gc124 (wc124, n_2732);
  or g3189 (n_2903, wc125, n_2473);
  not gc125 (wc125, n_2869);
  or g3190 (n_3020, wc126, n_2499);
  not gc126 (wc126, n_2500);
  or g3191 (n_3021, wc127, n_2509);
  not gc127 (wc127, n_2504);
  or g3192 (n_3024, wc128, n_2505);
  not gc128 (wc128, n_2506);
  or g3193 (n_3025, wc129, n_2515);
  not gc129 (wc129, n_2510);
  or g3194 (n_3028, wc130, n_2511);
  not gc130 (wc130, n_2512);
  or g3195 (n_3029, wc131, n_2521);
  not gc131 (wc131, n_2516);
  or g3196 (n_3032, wc132, n_2517);
  not gc132 (wc132, n_2518);
  or g3197 (n_3033, wc133, n_2527);
  not gc133 (wc133, n_2522);
  or g3198 (n_3036, wc134, n_2523);
  not gc134 (wc134, n_2524);
  or g3199 (n_3037, wc135, n_2533);
  not gc135 (wc135, n_2528);
  or g3200 (n_3040, wc136, n_2529);
  not gc136 (wc136, n_2530);
  or g3201 (n_3041, wc137, n_2539);
  not gc137 (wc137, n_2534);
  or g3202 (n_3044, wc138, n_2535);
  not gc138 (wc138, n_2536);
  or g3203 (n_3045, wc139, n_2545);
  not gc139 (wc139, n_2540);
  or g3204 (n_3048, wc140, n_2541);
  not gc140 (wc140, n_2542);
  or g3205 (n_3049, wc141, n_2551);
  not gc141 (wc141, n_2546);
  or g3206 (n_3052, wc142, n_2547);
  not gc142 (wc142, n_2548);
  or g3207 (n_3053, wc143, n_2557);
  not gc143 (wc143, n_2552);
  or g3208 (n_3056, wc144, n_2553);
  not gc144 (wc144, n_2554);
  or g3209 (n_3057, wc145, n_2563);
  not gc145 (wc145, n_2558);
  or g3210 (n_3060, wc146, n_2559);
  not gc146 (wc146, n_2560);
  or g3211 (n_3061, wc147, n_2569);
  not gc147 (wc147, n_2564);
  or g3212 (n_3064, wc148, n_2565);
  not gc148 (wc148, n_2566);
  or g3213 (n_3065, wc149, n_2575);
  not gc149 (wc149, n_2570);
  or g3214 (n_3068, wc150, n_2571);
  not gc150 (wc150, n_2572);
  or g3215 (n_3069, wc151, n_2581);
  not gc151 (wc151, n_2576);
  or g3216 (n_3072, wc152, n_2577);
  not gc152 (wc152, n_2578);
  or g3217 (n_3073, wc153, n_2587);
  not gc153 (wc153, n_2582);
  and g3218 (n_2720, wc154, n_2584);
  not gc154 (wc154, n_2585);
  and g3219 (n_2672, wc155, n_2668);
  not gc155 (wc155, n_2669);
  and g3220 (n_2679, wc156, n_2675);
  not gc156 (wc156, n_2676);
  and g3221 (n_2686, wc157, n_2682);
  not gc157 (wc157, n_2683);
  and g3222 (n_2693, wc158, n_2689);
  not gc158 (wc158, n_2690);
  and g3223 (n_2700, wc159, n_2696);
  not gc159 (wc159, n_2697);
  and g3224 (n_2707, wc160, n_2703);
  not gc160 (wc160, n_2704);
  and g3225 (n_2714, wc161, n_2710);
  not gc161 (wc161, n_2711);
  and g3226 (n_2794, wc162, n_2734);
  not gc162 (wc162, n_2735);
  and g3227 (n_2801, n_2759, wc163);
  not gc163 (wc163, n_2760);
  or g3228 (n_3076, wc164, n_2583);
  not gc164 (wc164, n_2584);
  or g3229 (n_3077, wc165, n_2593);
  not gc165 (wc165, n_2588);
  and g3230 (n_2725, wc166, n_2590);
  not gc166 (wc166, n_2591);
  and g3231 (n_2765, wc167, n_2671);
  not gc167 (wc167, n_2672);
  and g3232 (n_2770, wc168, n_2678);
  not gc168 (wc168, n_2679);
  and g3233 (n_2771, wc169, n_2685);
  not gc169 (wc169, n_2686);
  and g3234 (n_2776, wc170, n_2692);
  not gc170 (wc170, n_2693);
  and g3235 (n_2777, wc171, n_2699);
  not gc171 (wc171, n_2700);
  and g3236 (n_2782, wc172, n_2706);
  not gc172 (wc172, n_2707);
  and g3237 (n_2783, wc173, n_2713);
  not gc173 (wc173, n_2714);
  and g3238 (n_2721, wc174, n_2717);
  not gc174 (wc174, n_2718);
  or g3239 (n_2906, wc175, n_2479);
  not gc175 (wc175, n_2904);
  or g3240 (n_3080, wc176, n_2589);
  not gc176 (wc176, n_2590);
  or g3241 (n_3081, wc177, n_2599);
  not gc177 (wc177, n_2594);
  and g3242 (n_2727, wc178, n_2596);
  not gc178 (wc178, n_2597);
  and g3243 (n_2788, wc179, n_2720);
  not gc179 (wc179, n_2721);
  and g3244 (n_2820, n_2795, wc180);
  not gc180 (wc180, n_2796);
  or g3245 (n_2848, wc181, n_2768);
  not gc181 (wc181, n_2825);
  or g3246 (n_2908, wc182, n_2485);
  not gc182 (wc182, n_2825);
  or g3247 (n_3084, wc183, n_2595);
  not gc183 (wc183, n_2596);
  and g3248 (n_2728, wc184, n_2724);
  not gc184 (wc184, n_2725);
  and g3249 (n_2804, n_2765, wc185);
  not gc185 (wc185, n_2766);
  and g3250 (n_2806, n_2771, wc186);
  not gc186 (wc186, n_2772);
  and g3251 (n_2811, n_2777, wc187);
  not gc187 (wc187, n_2778);
  and g3252 (n_2813, n_2783, wc188);
  not gc188 (wc188, n_2784);
  or g3253 (n_2828, n_2824, wc189);
  not gc189 (wc189, n_2825);
  and g3254 (n_2789, wc190, n_2727);
  not gc190 (wc190, n_2728);
  and g3255 (n_2807, wc191, n_2803);
  not gc191 (wc191, n_2804);
  and g3256 (n_2814, wc192, n_2810);
  not gc192 (wc192, n_2811);
  or g3257 (n_2911, wc193, n_2491);
  not gc193 (wc193, n_2909);
  or g3258 (n_2913, wc194, n_2497);
  not gc194 (wc194, n_2872);
  and g3259 (n_2827, wc195, n_2806);
  not gc195 (wc195, n_2807);
  and g3260 (n_2830, wc196, n_2813);
  not gc196 (wc196, n_2814);
  or g3261 (n_2851, wc197, n_2774);
  not gc197 (wc197, n_2849);
  or g3262 (n_2918, wc198, n_2509);
  not gc198 (wc198, n_2849);
  and g3263 (n_2818, n_2789, wc199);
  not gc199 (wc199, n_2790);
  or g3264 (n_2916, wc200, n_2503);
  not gc200 (wc200, n_2914);
  and g3265 (n_2821, wc201, n_2817);
  not gc201 (wc201, n_2818);
  or g3266 (n_2840, wc202, n_2834);
  not gc202 (wc202, n_2836);
  or g3267 (n_2853, wc203, n_2780);
  not gc203 (wc203, n_2836);
  or g3268 (n_2921, wc204, n_2515);
  not gc204 (wc204, n_2919);
  or g3269 (n_2923, wc205, n_2521);
  not gc205 (wc205, n_2875);
  or g3270 (n_2928, wc206, n_2533);
  not gc206 (wc206, n_2836);
  and g3271 (n_2831, wc207, n_2820);
  not gc207 (wc207, n_2821);
  or g3272 (n_2856, wc208, n_2786);
  not gc208 (wc208, n_2854);
  or g3273 (n_2858, wc209, n_2792);
  not gc209 (wc209, n_2843);
  or g3274 (n_2926, wc210, n_2527);
  not gc210 (wc210, n_2924);
  or g3275 (n_2931, wc211, n_2539);
  not gc211 (wc211, n_2929);
  or g3276 (n_2933, wc212, n_2545);
  not gc212 (wc212, n_2878);
  or g3277 (n_2938, wc213, n_2557);
  not gc213 (wc213, n_2854);
  or g3278 (n_2948, wc214, n_2581);
  not gc214 (wc214, n_2843);
  and g3279 (n_2837, n_2831, wc215);
  not gc215 (wc215, n_2832);
  or g3280 (n_2861, wc216, n_2798);
  not gc216 (wc216, n_2859);
  or g3281 (n_2936, wc217, n_2551);
  not gc217 (wc217, n_2934);
  or g3282 (n_2941, wc218, n_2563);
  not gc218 (wc218, n_2939);
  or g3283 (n_2943, wc219, n_2569);
  not gc219 (wc219, n_2881);
  or g3284 (n_2951, wc220, n_2587);
  not gc220 (wc220, n_2949);
  or g3285 (n_2953, wc221, n_2593);
  not gc221 (wc221, n_2884);
  or g3286 (n_2958, wc222, n_2605);
  not gc222 (wc222, n_2859);
  or g3287 (n_2866, wc223, n_2862);
  not gc223 (wc223, n_2863);
  or g3288 (n_2968, wc224, n_2629);
  not gc224 (wc224, n_2863);
  or g3289 (n_2946, wc225, n_2575);
  not gc225 (wc225, n_2944);
  or g3290 (n_2956, wc226, n_2599);
  not gc226 (wc226, n_2954);
  or g3291 (n_2961, wc227, n_2611);
  not gc227 (wc227, n_2959);
  or g3292 (n_2963, wc228, n_2617);
  not gc228 (wc228, n_2887);
  or g3293 (n_2971, n_2635, wc229);
  not gc229 (wc229, n_2969);
  not g3294 (Z[68], n_2973);
  or g3295 (n_2966, wc230, n_2623);
  not gc230 (wc230, n_2964);
endmodule

module mult_signed_const_11124_GENERIC(A, Z);
  input [49:0] A;
  output [68:0] Z;
  wire [49:0] A;
  wire [68:0] Z;
  mult_signed_const_11124_GENERIC_REAL g1(.A ({A[49:2], A[0], A[0]}),
       .Z (Z));
endmodule

module mult_signed_const_11527_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [50:0] A;
  output [69:0] Z;
  wire [50:0] A;
  wire [69:0] Z;
  wire n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62;
  wire n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78;
  wire n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_263, n_264, n_265;
  wire n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_279, n_280, n_281;
  wire n_282, n_283, n_286, n_287, n_288, n_289, n_290, n_292;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_330, n_331, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_368, n_369, n_370, n_371;
  wire n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379;
  wire n_380, n_381, n_383, n_384, n_385, n_386, n_387, n_388;
  wire n_389, n_390, n_391, n_393, n_394, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_530;
  wire n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538;
  wire n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_563;
  wire n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571;
  wire n_572, n_573, n_575, n_577, n_578, n_579, n_580, n_581;
  wire n_582, n_583, n_584, n_585, n_586, n_587, n_589, n_590;
  wire n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598;
  wire n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606;
  wire n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_615;
  wire n_616, n_617, n_618, n_619, n_620, n_621, n_622, n_623;
  wire n_624, n_625, n_626, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_642;
  wire n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650;
  wire n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658;
  wire n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666;
  wire n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674;
  wire n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682;
  wire n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690;
  wire n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698;
  wire n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706;
  wire n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714;
  wire n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722;
  wire n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730;
  wire n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738;
  wire n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746;
  wire n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754;
  wire n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762;
  wire n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770;
  wire n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778;
  wire n_779, n_780, n_783, n_784, n_785, n_786, n_787, n_788;
  wire n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796;
  wire n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807;
  wire n_808, n_809, n_810, n_811, n_812, n_813, n_815, n_816;
  wire n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824;
  wire n_825, n_826, n_827, n_828, n_831, n_832, n_833, n_834;
  wire n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842;
  wire n_843, n_845, n_846, n_848, n_849, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_860, n_861, n_862, n_863;
  wire n_864, n_865, n_866, n_867, n_868, n_869, n_871, n_872;
  wire n_875, n_876, n_877, n_878, n_879, n_880, n_885, n_886;
  wire n_887, n_888, n_889, n_890, n_891, n_893, n_896, n_897;
  wire n_898, n_899, n_900, n_906, n_907, n_908, n_909, n_913;
  wire n_914, n_915, n_916, n_920, n_921, n_922, n_923, n_925;
  wire n_927, n_928, n_932, n_933, n_935, n_936, n_939, n_942;
  wire n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950;
  wire n_951, n_953, n_954, n_955, n_956, n_957, n_958, n_959;
  wire n_962, n_963, n_964, n_965, n_966, n_967, n_969, n_970;
  wire n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979;
  wire n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_994, n_995, n_997, n_998, n_999;
  wire n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007;
  wire n_1008, n_1009, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017;
  wire n_1018, n_1019, n_1020, n_1021, n_1026, n_1027, n_1028, n_1030;
  wire n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039;
  wire n_1040, n_1041, n_1045, n_1046, n_1047, n_1050, n_1051, n_1052;
  wire n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060;
  wire n_1061, n_1062, n_1063, n_1065, n_1066, n_1067, n_1068, n_1072;
  wire n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080;
  wire n_1081, n_1082, n_1083, n_1084, n_1085, n_1092, n_1093, n_1094;
  wire n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102;
  wire n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1114;
  wire n_1115, n_1118, n_1119, n_1120, n_1122, n_1123, n_1124, n_1125;
  wire n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133;
  wire n_1134, n_1135, n_1136, n_1137, n_1141, n_1142, n_1143, n_1144;
  wire n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155;
  wire n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163;
  wire n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1172, n_1173;
  wire n_1174, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184;
  wire n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192;
  wire n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200;
  wire n_1201, n_1206, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215;
  wire n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223;
  wire n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231;
  wire n_1233, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248;
  wire n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264;
  wire n_1265, n_1266, n_1268, n_1270, n_1271, n_1273, n_1274, n_1275;
  wire n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283;
  wire n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291;
  wire n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1302;
  wire n_1303, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311;
  wire n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319;
  wire n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327;
  wire n_1328, n_1330, n_1331, n_1334, n_1335, n_1336, n_1337, n_1338;
  wire n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346;
  wire n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354;
  wire n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1362, n_1363;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381;
  wire n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
  wire n_1396, n_1397, n_1398, n_1402, n_1403, n_1404, n_1405, n_1406;
  wire n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414;
  wire n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1428;
  wire n_1429, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440;
  wire n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448;
  wire n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456;
  wire n_1457, n_1460, n_1461, n_1465, n_1466, n_1467, n_1468, n_1469;
  wire n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477;
  wire n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485;
  wire n_1486, n_1487, n_1488, n_1489, n_1492, n_1493, n_1497, n_1498;
  wire n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506;
  wire n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514;
  wire n_1515, n_1516, n_1517, n_1525, n_1526, n_1527, n_1528, n_1530;
  wire n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538;
  wire n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546;
  wire n_1547, n_1548, n_1549, n_1557, n_1558, n_1559, n_1560, n_1562;
  wire n_1563, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571;
  wire n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579;
  wire n_1580, n_1581, n_1582, n_1583, n_1588, n_1589, n_1590, n_1591;
  wire n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600;
  wire n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608;
  wire n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1620;
  wire n_1621, n_1622, n_1623, n_1625, n_1626, n_1627, n_1628, n_1629;
  wire n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637;
  wire n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645;
  wire n_1646, n_1647, n_1650, n_1651, n_1652, n_1653, n_1658, n_1659;
  wire n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667;
  wire n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675;
  wire n_1676, n_1677, n_1678, n_1679, n_1682, n_1683, n_1684, n_1685;
  wire n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697;
  wire n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705;
  wire n_1706, n_1707, n_1708, n_1709, n_1714, n_1715, n_1716, n_1717;
  wire n_1718, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726;
  wire n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734;
  wire n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1746;
  wire n_1747, n_1748, n_1749, n_1750, n_1752, n_1753, n_1754, n_1755;
  wire n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763;
  wire n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771;
  wire n_1772, n_1773, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
  wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1810, n_1811;
  wire n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819;
  wire n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
  wire n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836;
  wire n_1837, n_1841, n_1842, n_1844, n_1845, n_1846, n_1847, n_1848;
  wire n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856;
  wire n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864;
  wire n_1865, n_1866, n_1867, n_1868, n_1869, n_1873, n_1874, n_1876;
  wire n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884;
  wire n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892;
  wire n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900;
  wire n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1909;
  wire n_1910, n_1912, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919;
  wire n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927;
  wire n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935;
  wire n_1936, n_1937, n_1938, n_1939, n_1941, n_1942, n_1944, n_1946;
  wire n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954;
  wire n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962;
  wire n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1972, n_1974;
  wire n_1975, n_1976, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983;
  wire n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991;
  wire n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999;
  wire n_2000, n_2004, n_2006, n_2007, n_2008, n_2010, n_2011, n_2012;
  wire n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020;
  wire n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028;
  wire n_2029, n_2030, n_2031, n_2032, n_2034, n_2036, n_2037, n_2038;
  wire n_2039, n_2040, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047;
  wire n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055;
  wire n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063;
  wire n_2064, n_2066, n_2068, n_2069, n_2070, n_2071, n_2072, n_2074;
  wire n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082;
  wire n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090;
  wire n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2102;
  wire n_2104, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112;
  wire n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120;
  wire n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128;
  wire n_2129, n_2134, n_2136, n_2138, n_2139, n_2140, n_2141, n_2142;
  wire n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150;
  wire n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158;
  wire n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2166, n_2170;
  wire n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178;
  wire n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186;
  wire n_2187, n_2188, n_2189, n_2190, n_2191, n_2193, n_2194, n_2195;
  wire n_2196, n_2197, n_2198, n_2199, n_2201, n_2202, n_2203, n_2204;
  wire n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212;
  wire n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220;
  wire n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2228, n_2230;
  wire n_2231, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239;
  wire n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247;
  wire n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255;
  wire n_2258, n_2259, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266;
  wire n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274;
  wire n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2286;
  wire n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296;
  wire n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304;
  wire n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2314, n_2317;
  wire n_2318, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326;
  wire n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2342;
  wire n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351;
  wire n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2364;
  wire n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372;
  wire n_2373, n_2374, n_2375, n_2376, n_2377, n_2386, n_2387, n_2388;
  wire n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396;
  wire n_2397, n_2404, n_2405, n_2406, n_2408, n_2409, n_2410, n_2411;
  wire n_2412, n_2413, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425;
  wire n_2426, n_2427, n_2428, n_2429, n_2436, n_2437, n_2438, n_2439;
  wire n_2440, n_2441, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451;
  wire n_2452, n_2453, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461;
  wire n_2466, n_2467, n_2468, n_2469, n_2471, n_2472, n_2473, n_2476;
  wire n_2477, n_2489, n_2491, n_2493, n_2494, n_2495, n_2496, n_2497;
  wire n_2499, n_2500, n_2501, n_2502, n_2503, n_2505, n_2506, n_2507;
  wire n_2508, n_2509, n_2511, n_2512, n_2513, n_2514, n_2515, n_2517;
  wire n_2518, n_2519, n_2520, n_2521, n_2523, n_2524, n_2525, n_2526;
  wire n_2527, n_2529, n_2530, n_2531, n_2532, n_2533, n_2535, n_2536;
  wire n_2537, n_2538, n_2539, n_2541, n_2542, n_2543, n_2544, n_2545;
  wire n_2547, n_2548, n_2549, n_2550, n_2551, n_2553, n_2554, n_2555;
  wire n_2556, n_2557, n_2559, n_2560, n_2561, n_2562, n_2563, n_2565;
  wire n_2566, n_2567, n_2568, n_2569, n_2571, n_2572, n_2573, n_2574;
  wire n_2575, n_2577, n_2578, n_2579, n_2580, n_2581, n_2583, n_2584;
  wire n_2585, n_2586, n_2587, n_2589, n_2590, n_2591, n_2592, n_2593;
  wire n_2595, n_2596, n_2597, n_2598, n_2599, n_2601, n_2602, n_2603;
  wire n_2604, n_2605, n_2607, n_2608, n_2609, n_2610, n_2611, n_2613;
  wire n_2614, n_2615, n_2616, n_2617, n_2619, n_2620, n_2621, n_2622;
  wire n_2623, n_2625, n_2626, n_2627, n_2628, n_2629, n_2631, n_2632;
  wire n_2633, n_2634, n_2635, n_2637, n_2638, n_2639, n_2640, n_2641;
  wire n_2643, n_2644, n_2645, n_2646, n_2647, n_2649, n_2650, n_2651;
  wire n_2652, n_2653, n_2655, n_2656, n_2657, n_2658, n_2659, n_2661;
  wire n_2662, n_2663, n_2664, n_2665, n_2667, n_2668, n_2669, n_2670;
  wire n_2671, n_2673, n_2674, n_2675, n_2676, n_2677, n_2679, n_2680;
  wire n_2681, n_2682, n_2683, n_2685, n_2686, n_2689, n_2692, n_2694;
  wire n_2695, n_2697, n_2698, n_2700, n_2701, n_2702, n_2704, n_2705;
  wire n_2707, n_2708, n_2709, n_2711, n_2712, n_2714, n_2715, n_2716;
  wire n_2718, n_2719, n_2721, n_2722, n_2723, n_2725, n_2726, n_2728;
  wire n_2729, n_2730, n_2732, n_2733, n_2735, n_2736, n_2737, n_2739;
  wire n_2740, n_2742, n_2743, n_2744, n_2746, n_2747, n_2749, n_2750;
  wire n_2751, n_2753, n_2754, n_2756, n_2757, n_2758, n_2760, n_2761;
  wire n_2763, n_2764, n_2765, n_2767, n_2768, n_2770, n_2771, n_2772;
  wire n_2774, n_2775, n_2777, n_2778, n_2779, n_2781, n_2782, n_2784;
  wire n_2785, n_2786, n_2788, n_2789, n_2791, n_2792, n_2793, n_2795;
  wire n_2796, n_2798, n_2799, n_2800, n_2802, n_2803, n_2805, n_2806;
  wire n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2816, n_2817;
  wire n_2818, n_2819, n_2820, n_2822, n_2823, n_2824, n_2825, n_2826;
  wire n_2828, n_2829, n_2830, n_2831, n_2832, n_2834, n_2835, n_2836;
  wire n_2837, n_2838, n_2840, n_2841, n_2842, n_2843, n_2844, n_2846;
  wire n_2847, n_2848, n_2849, n_2850, n_2852, n_2853, n_2854, n_2855;
  wire n_2856, n_2857, n_2858, n_2860, n_2861, n_2863, n_2864, n_2865;
  wire n_2867, n_2868, n_2870, n_2871, n_2872, n_2874, n_2875, n_2877;
  wire n_2878, n_2879, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886;
  wire n_2888, n_2889, n_2890, n_2891, n_2892, n_2894, n_2895, n_2896;
  wire n_2897, n_2898, n_2900, n_2902, n_2903, n_2905, n_2907, n_2908;
  wire n_2910, n_2912, n_2913, n_2915, n_2916, n_2917, n_2919, n_2920;
  wire n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928;
  wire n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936;
  wire n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944;
  wire n_2948, n_2949, n_2951, n_2953, n_2954, n_2956, n_2958, n_2959;
  wire n_2961, n_2963, n_2964, n_2966, n_2968, n_2969, n_2971, n_2973;
  wire n_2974, n_2976, n_2978, n_2979, n_2981, n_2983, n_2984, n_2986;
  wire n_2988, n_2989, n_2991, n_2993, n_2994, n_2996, n_2998, n_2999;
  wire n_3001, n_3003, n_3004, n_3006, n_3008, n_3009, n_3011, n_3013;
  wire n_3014, n_3016, n_3018, n_3019, n_3021, n_3023, n_3024, n_3026;
  wire n_3028, n_3030, n_3033, n_3034, n_3036, n_3037, n_3038, n_3040;
  wire n_3041, n_3042, n_3044, n_3045, n_3046, n_3048, n_3049, n_3050;
  wire n_3052, n_3053, n_3054, n_3056, n_3057, n_3058, n_3060, n_3061;
  wire n_3062, n_3064, n_3065, n_3066, n_3068, n_3069, n_3070, n_3072;
  wire n_3073, n_3074, n_3076, n_3077, n_3078, n_3080, n_3081, n_3082;
  wire n_3084, n_3085, n_3086, n_3088, n_3089, n_3090, n_3092, n_3093;
  wire n_3094, n_3096, n_3097, n_3098, n_3100, n_3101, n_3102, n_3104;
  wire n_3105, n_3106, n_3108, n_3109, n_3110, n_3112, n_3113, n_3114;
  wire n_3116, n_3117, n_3118, n_3120, n_3121, n_3122, n_3124, n_3125;
  wire n_3126, n_3128, n_3129, n_3130, n_3132, n_3133, n_3134, n_3136;
  wire n_3137, n_3138, n_3140, n_3141, n_3142, n_3144, n_3145, n_3146;
  wire n_3148, n_3149, n_3150, n_3152, n_3153, n_3154, n_3156, n_3157;
  wire n_3158, n_3160, n_3161, n_3162, n_3164;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g404 (n_187, A[4], A[0]);
  and g2 (n_116, A[4], A[0]);
  xor g405 (n_942, A[5], A[3]);
  xor g406 (n_186, n_942, A[1]);
  nand g3 (n_943, A[5], A[3]);
  nand g407 (n_944, A[1], A[3]);
  nand g408 (n_945, A[5], A[1]);
  nand g409 (n_115, n_943, n_944, n_945);
  xor g410 (n_263, A[6], A[4]);
  and g411 (n_264, A[6], A[4]);
  xor g412 (n_946, A[0], A[2]);
  xor g413 (n_185, n_946, n_263);
  nand g414 (n_947, A[0], A[2]);
  nand g4 (n_948, n_263, A[2]);
  nand g5 (n_949, A[0], n_263);
  nand g415 (n_114, n_947, n_948, n_949);
  xor g416 (n_950, A[7], A[5]);
  xor g417 (n_265, n_950, A[1]);
  nand g418 (n_951, A[7], A[5]);
  nand g420 (n_953, A[7], A[1]);
  nand g6 (n_267, n_951, n_945, n_953);
  xor g421 (n_954, A[3], n_264);
  xor g422 (n_184, n_954, n_265);
  nand g423 (n_955, A[3], n_264);
  nand g424 (n_956, n_265, n_264);
  nand g425 (n_957, A[3], n_265);
  nand g426 (n_113, n_955, n_956, n_957);
  xor g427 (n_266, A[8], A[6]);
  and g428 (n_269, A[8], A[6]);
  xor g429 (n_958, A[4], A[2]);
  xor g430 (n_268, n_958, A[0]);
  nand g431 (n_959, A[4], A[2]);
  xor g435 (n_962, n_266, n_267);
  xor g436 (n_183, n_962, n_268);
  nand g437 (n_963, n_266, n_267);
  nand g438 (n_964, n_268, n_267);
  nand g439 (n_965, n_266, n_268);
  nand g440 (n_112, n_963, n_964, n_965);
  xor g441 (n_966, A[9], A[7]);
  xor g442 (n_270, n_966, A[5]);
  nand g443 (n_967, A[9], A[7]);
  nand g445 (n_969, A[9], A[5]);
  nand g446 (n_274, n_967, n_951, n_969);
  xor g447 (n_970, A[3], A[1]);
  xor g448 (n_272, n_970, n_269);
  nand g450 (n_972, n_269, A[1]);
  nand g451 (n_973, A[3], n_269);
  nand g452 (n_275, n_944, n_972, n_973);
  xor g453 (n_974, n_270, n_271);
  xor g454 (n_182, n_974, n_272);
  nand g455 (n_975, n_270, n_271);
  nand g456 (n_976, n_272, n_271);
  nand g457 (n_977, n_270, n_272);
  nand g458 (n_111, n_975, n_976, n_977);
  xor g459 (n_273, A[8], A[4]);
  and g460 (n_278, A[8], A[4]);
  xor g461 (n_978, A[6], A[10]);
  xor g462 (n_276, n_978, A[2]);
  nand g463 (n_979, A[6], A[10]);
  nand g464 (n_980, A[2], A[10]);
  nand g465 (n_981, A[6], A[2]);
  nand g466 (n_280, n_979, n_980, n_981);
  xor g467 (n_982, A[0], n_273);
  xor g468 (n_277, n_982, n_274);
  nand g469 (n_983, A[0], n_273);
  nand g470 (n_984, n_274, n_273);
  nand g471 (n_985, A[0], n_274);
  nand g472 (n_282, n_983, n_984, n_985);
  xor g473 (n_986, n_275, n_276);
  xor g474 (n_181, n_986, n_277);
  nand g475 (n_987, n_275, n_276);
  nand g476 (n_988, n_277, n_276);
  nand g477 (n_989, n_275, n_277);
  nand g478 (n_110, n_987, n_988, n_989);
  xor g479 (n_990, A[9], A[5]);
  xor g480 (n_279, n_990, A[7]);
  xor g485 (n_994, A[11], A[3]);
  xor g486 (n_281, n_994, A[1]);
  nand g487 (n_995, A[11], A[3]);
  nand g489 (n_997, A[11], A[1]);
  nand g490 (n_286, n_995, n_944, n_997);
  xor g491 (n_998, n_278, n_279);
  xor g492 (n_283, n_998, n_280);
  nand g493 (n_999, n_278, n_279);
  nand g494 (n_1000, n_280, n_279);
  nand g495 (n_1001, n_278, n_280);
  nand g496 (n_289, n_999, n_1000, n_1001);
  xor g497 (n_1002, n_281, n_282);
  xor g498 (n_180, n_1002, n_283);
  nand g499 (n_1003, n_281, n_282);
  nand g500 (n_1004, n_283, n_282);
  nand g501 (n_1005, n_281, n_283);
  nand g502 (n_109, n_1003, n_1004, n_1005);
  xor g505 (n_1006, A[4], A[10]);
  xor g506 (n_287, n_1006, A[12]);
  nand g507 (n_1007, A[4], A[10]);
  nand g508 (n_1008, A[12], A[10]);
  nand g509 (n_1009, A[4], A[12]);
  nand g510 (n_292, n_1007, n_1008, n_1009);
  xor g512 (n_288, n_946, n_266);
  nand g514 (n_1012, n_266, A[0]);
  nand g515 (n_1013, A[2], n_266);
  nand g516 (n_295, n_947, n_1012, n_1013);
  xor g517 (n_1014, n_274, n_286);
  xor g518 (n_290, n_1014, n_287);
  nand g519 (n_1015, n_274, n_286);
  nand g520 (n_1016, n_287, n_286);
  nand g521 (n_1017, n_274, n_287);
  nand g522 (n_297, n_1015, n_1016, n_1017);
  xor g523 (n_1018, n_288, n_289);
  xor g524 (n_179, n_1018, n_290);
  nand g525 (n_1019, n_288, n_289);
  nand g526 (n_1020, n_290, n_289);
  nand g527 (n_1021, n_288, n_290);
  nand g528 (n_108, n_1019, n_1020, n_1021);
  xor g535 (n_1026, A[11], A[13]);
  xor g536 (n_294, n_1026, A[3]);
  nand g537 (n_1027, A[11], A[13]);
  nand g538 (n_1028, A[3], A[13]);
  nand g540 (n_301, n_1027, n_1028, n_995);
  xor g541 (n_1030, A[1], n_269);
  xor g542 (n_296, n_1030, n_292);
  nand g544 (n_1032, n_292, n_269);
  nand g545 (n_1033, A[1], n_292);
  nand g546 (n_304, n_972, n_1032, n_1033);
  xor g547 (n_1034, n_270, n_294);
  xor g548 (n_298, n_1034, n_295);
  nand g549 (n_1035, n_270, n_294);
  nand g550 (n_1036, n_295, n_294);
  nand g551 (n_1037, n_270, n_295);
  nand g552 (n_306, n_1035, n_1036, n_1037);
  xor g553 (n_1038, n_296, n_297);
  xor g554 (n_178, n_1038, n_298);
  nand g555 (n_1039, n_296, n_297);
  nand g556 (n_1040, n_298, n_297);
  nand g557 (n_1041, n_296, n_298);
  nand g558 (n_107, n_1039, n_1040, n_1041);
  xor g559 (n_299, A[14], A[8]);
  and g560 (n_308, A[14], A[8]);
  xor g562 (n_302, n_263, A[12]);
  nand g565 (n_1045, A[6], A[12]);
  xor g567 (n_1046, A[0], A[10]);
  xor g568 (n_303, n_1046, A[2]);
  nand g569 (n_1047, A[0], A[10]);
  nand g572 (n_309, n_1047, n_980, n_947);
  xor g573 (n_1050, n_299, n_274);
  xor g574 (n_305, n_1050, n_301);
  nand g575 (n_1051, n_299, n_274);
  nand g576 (n_1052, n_301, n_274);
  nand g577 (n_1053, n_299, n_301);
  nand g578 (n_314, n_1051, n_1052, n_1053);
  xor g579 (n_1054, n_302, n_303);
  xor g580 (n_307, n_1054, n_304);
  nand g581 (n_1055, n_302, n_303);
  nand g582 (n_1056, n_304, n_303);
  nand g583 (n_1057, n_302, n_304);
  nand g584 (n_317, n_1055, n_1056, n_1057);
  xor g585 (n_1058, n_305, n_306);
  xor g586 (n_177, n_1058, n_307);
  nand g587 (n_1059, n_305, n_306);
  nand g588 (n_1060, n_307, n_306);
  nand g589 (n_1061, n_305, n_307);
  nand g590 (n_106, n_1059, n_1060, n_1061);
  xor g591 (n_1062, A[15], A[9]);
  xor g592 (n_311, n_1062, A[7]);
  nand g593 (n_1063, A[15], A[9]);
  nand g595 (n_1065, A[15], A[7]);
  nand g596 (n_319, n_1063, n_967, n_1065);
  xor g597 (n_1066, A[5], A[13]);
  xor g598 (n_313, n_1066, A[1]);
  nand g599 (n_1067, A[5], A[13]);
  nand g600 (n_1068, A[1], A[13]);
  nand g602 (n_320, n_1067, n_1068, n_945);
  xor g604 (n_312, n_994, n_308);
  nand g606 (n_1072, n_308, A[3]);
  nand g607 (n_1073, A[11], n_308);
  nand g608 (n_322, n_995, n_1072, n_1073);
  xor g609 (n_1074, n_309, n_310);
  xor g610 (n_315, n_1074, n_311);
  nand g611 (n_1075, n_309, n_310);
  nand g612 (n_1076, n_311, n_310);
  nand g613 (n_1077, n_309, n_311);
  nand g614 (n_325, n_1075, n_1076, n_1077);
  xor g615 (n_1078, n_312, n_313);
  xor g616 (n_316, n_1078, n_314);
  nand g617 (n_1079, n_312, n_313);
  nand g618 (n_1080, n_314, n_313);
  nand g619 (n_1081, n_312, n_314);
  nand g620 (n_328, n_1079, n_1080, n_1081);
  xor g621 (n_1082, n_315, n_316);
  xor g622 (n_176, n_1082, n_317);
  nand g623 (n_1083, n_315, n_316);
  nand g624 (n_1084, n_317, n_316);
  nand g625 (n_1085, n_315, n_317);
  nand g626 (n_105, n_1083, n_1084, n_1085);
  xor g630 (n_321, n_263, A[10]);
  xor g636 (n_323, n_946, A[16]);
  nand g638 (n_1092, A[16], A[0]);
  nand g639 (n_1093, A[2], A[16]);
  nand g640 (n_331, n_947, n_1092, n_1093);
  xor g641 (n_1094, A[12], n_299);
  xor g642 (n_324, n_1094, n_319);
  nand g643 (n_1095, A[12], n_299);
  nand g644 (n_1096, n_319, n_299);
  nand g645 (n_1097, A[12], n_319);
  nand g646 (n_335, n_1095, n_1096, n_1097);
  xor g647 (n_1098, n_320, n_321);
  xor g648 (n_326, n_1098, n_322);
  nand g649 (n_1099, n_320, n_321);
  nand g650 (n_1100, n_322, n_321);
  nand g651 (n_1101, n_320, n_322);
  nand g652 (n_337, n_1099, n_1100, n_1101);
  xor g653 (n_1102, n_323, n_324);
  xor g654 (n_327, n_1102, n_325);
  nand g655 (n_1103, n_323, n_324);
  nand g656 (n_1104, n_325, n_324);
  nand g657 (n_1105, n_323, n_325);
  nand g658 (n_339, n_1103, n_1104, n_1105);
  xor g659 (n_1106, n_326, n_327);
  xor g660 (n_175, n_1106, n_328);
  nand g661 (n_1107, n_326, n_327);
  nand g662 (n_1108, n_328, n_327);
  nand g663 (n_1109, n_326, n_328);
  nand g664 (n_104, n_1107, n_1108, n_1109);
  xor g671 (n_1114, A[5], A[11]);
  xor g672 (n_334, n_1114, A[3]);
  nand g673 (n_1115, A[5], A[11]);
  nand g676 (n_343, n_1115, n_995, n_943);
  xor g677 (n_1118, A[1], A[17]);
  xor g678 (n_333, n_1118, A[13]);
  nand g679 (n_1119, A[1], A[17]);
  nand g680 (n_1120, A[13], A[17]);
  nand g682 (n_344, n_1119, n_1120, n_1068);
  xor g683 (n_1122, n_308, n_330);
  xor g684 (n_336, n_1122, n_331);
  nand g685 (n_1123, n_308, n_330);
  nand g686 (n_1124, n_331, n_330);
  nand g687 (n_1125, n_308, n_331);
  nand g688 (n_348, n_1123, n_1124, n_1125);
  xor g689 (n_1126, n_311, n_333);
  xor g690 (n_338, n_1126, n_334);
  nand g691 (n_1127, n_311, n_333);
  nand g692 (n_1128, n_334, n_333);
  nand g693 (n_1129, n_311, n_334);
  nand g694 (n_350, n_1127, n_1128, n_1129);
  xor g695 (n_1130, n_335, n_336);
  xor g696 (n_340, n_1130, n_337);
  nand g697 (n_1131, n_335, n_336);
  nand g698 (n_1132, n_337, n_336);
  nand g699 (n_1133, n_335, n_337);
  nand g700 (n_352, n_1131, n_1132, n_1133);
  xor g701 (n_1134, n_338, n_339);
  xor g702 (n_174, n_1134, n_340);
  nand g703 (n_1135, n_338, n_339);
  nand g704 (n_1136, n_340, n_339);
  nand g705 (n_1137, n_338, n_340);
  nand g706 (n_103, n_1135, n_1136, n_1137);
  xor g707 (n_341, A[18], A[4]);
  and g708 (n_354, A[18], A[4]);
  xor g710 (n_345, n_299, A[6]);
  nand g713 (n_1141, A[14], A[6]);
  xor g715 (n_1142, A[16], A[12]);
  xor g716 (n_346, n_1142, A[2]);
  nand g717 (n_1143, A[16], A[12]);
  nand g718 (n_1144, A[2], A[12]);
  nand g720 (n_357, n_1143, n_1144, n_1093);
  xor g722 (n_347, n_1046, n_341);
  nand g724 (n_1148, n_341, A[0]);
  nand g725 (n_1149, A[10], n_341);
  nand g726 (n_119, n_1047, n_1148, n_1149);
  xor g727 (n_1150, n_319, n_343);
  xor g728 (n_349, n_1150, n_344);
  nand g729 (n_1151, n_319, n_343);
  nand g730 (n_1152, n_344, n_343);
  nand g731 (n_1153, n_319, n_344);
  nand g732 (n_121, n_1151, n_1152, n_1153);
  xor g733 (n_1154, n_345, n_346);
  xor g734 (n_351, n_1154, n_347);
  nand g735 (n_1155, n_345, n_346);
  nand g736 (n_1156, n_347, n_346);
  nand g737 (n_1157, n_345, n_347);
  nand g738 (n_359, n_1155, n_1156, n_1157);
  xor g739 (n_1158, n_348, n_349);
  xor g740 (n_353, n_1158, n_350);
  nand g741 (n_1159, n_348, n_349);
  nand g742 (n_1160, n_350, n_349);
  nand g743 (n_1161, n_348, n_350);
  nand g744 (n_361, n_1159, n_1160, n_1161);
  xor g745 (n_1162, n_351, n_352);
  xor g746 (n_173, n_1162, n_353);
  nand g747 (n_1163, n_351, n_352);
  nand g748 (n_1164, n_353, n_352);
  nand g749 (n_1165, n_351, n_353);
  nand g750 (n_102, n_1163, n_1164, n_1165);
  xor g751 (n_1166, A[19], A[5]);
  xor g752 (n_356, n_1166, A[15]);
  nand g753 (n_1167, A[19], A[5]);
  nand g754 (n_1168, A[15], A[5]);
  nand g755 (n_1169, A[19], A[15]);
  nand g756 (n_363, n_1167, n_1168, n_1169);
  xor g758 (n_117, n_966, A[17]);
  nand g760 (n_1172, A[17], A[7]);
  nand g761 (n_1173, A[9], A[17]);
  nand g762 (n_366, n_967, n_1172, n_1173);
  xor g763 (n_1174, A[13], A[3]);
  xor g764 (n_118, n_1174, A[11]);
  xor g769 (n_1178, A[1], n_354);
  xor g770 (n_120, n_1178, n_355);
  nand g771 (n_1179, A[1], n_354);
  nand g772 (n_1180, n_355, n_354);
  nand g773 (n_1181, A[1], n_355);
  nand g774 (n_369, n_1179, n_1180, n_1181);
  xor g775 (n_1182, n_356, n_357);
  xor g776 (n_358, n_1182, n_117);
  nand g777 (n_1183, n_356, n_357);
  nand g778 (n_1184, n_117, n_357);
  nand g779 (n_1185, n_356, n_117);
  nand g780 (n_370, n_1183, n_1184, n_1185);
  xor g781 (n_1186, n_118, n_119);
  xor g782 (n_360, n_1186, n_120);
  nand g783 (n_1187, n_118, n_119);
  nand g784 (n_1188, n_120, n_119);
  nand g785 (n_1189, n_118, n_120);
  nand g786 (n_373, n_1187, n_1188, n_1189);
  xor g787 (n_1190, n_121, n_358);
  xor g788 (n_362, n_1190, n_359);
  nand g789 (n_1191, n_121, n_358);
  nand g790 (n_1192, n_359, n_358);
  nand g791 (n_1193, n_121, n_359);
  nand g792 (n_375, n_1191, n_1192, n_1193);
  xor g793 (n_1194, n_360, n_361);
  xor g794 (n_172, n_1194, n_362);
  nand g795 (n_1195, n_360, n_361);
  nand g796 (n_1196, n_362, n_361);
  nand g797 (n_1197, n_360, n_362);
  nand g798 (n_101, n_1195, n_1196, n_1197);
  xor g799 (n_1198, A[20], A[18]);
  xor g800 (n_364, n_1198, A[14]);
  nand g801 (n_1199, A[20], A[18]);
  nand g802 (n_1200, A[14], A[18]);
  nand g803 (n_1201, A[20], A[14]);
  nand g804 (n_377, n_1199, n_1200, n_1201);
  xor g806 (n_365, n_263, A[8]);
  xor g811 (n_1206, A[12], A[2]);
  xor g812 (n_368, n_1206, A[10]);
  nand g816 (n_381, n_1144, n_980, n_1008);
  xor g817 (n_1210, A[16], n_363);
  xor g818 (n_371, n_1210, n_364);
  nand g819 (n_1211, A[16], n_363);
  nand g820 (n_1212, n_364, n_363);
  nand g821 (n_1213, A[16], n_364);
  nand g822 (n_385, n_1211, n_1212, n_1213);
  xor g823 (n_1214, n_365, n_366);
  xor g824 (n_372, n_1214, n_301);
  nand g825 (n_1215, n_365, n_366);
  nand g826 (n_1216, n_301, n_366);
  nand g827 (n_1217, n_365, n_301);
  nand g828 (n_383, n_1215, n_1216, n_1217);
  xor g829 (n_1218, n_368, n_369);
  xor g830 (n_374, n_1218, n_370);
  nand g831 (n_1219, n_368, n_369);
  nand g832 (n_1220, n_370, n_369);
  nand g833 (n_1221, n_368, n_370);
  nand g834 (n_387, n_1219, n_1220, n_1221);
  xor g835 (n_1222, n_371, n_372);
  xor g836 (n_376, n_1222, n_373);
  nand g837 (n_1223, n_371, n_372);
  nand g838 (n_1224, n_373, n_372);
  nand g839 (n_1225, n_371, n_373);
  nand g840 (n_389, n_1223, n_1224, n_1225);
  xor g841 (n_1226, n_374, n_375);
  xor g842 (n_171, n_1226, n_376);
  nand g843 (n_1227, n_374, n_375);
  nand g844 (n_1228, n_376, n_375);
  nand g845 (n_1229, n_374, n_376);
  nand g846 (n_100, n_1227, n_1228, n_1229);
  xor g847 (n_1230, A[21], A[19]);
  xor g848 (n_379, n_1230, A[15]);
  nand g849 (n_1231, A[21], A[19]);
  nand g851 (n_1233, A[21], A[15]);
  nand g852 (n_391, n_1231, n_1169, n_1233);
  xor g854 (n_380, n_950, A[9]);
  xor g865 (n_1242, A[17], n_377);
  xor g866 (n_384, n_1242, n_378);
  nand g867 (n_1243, A[17], n_377);
  nand g868 (n_1244, n_378, n_377);
  nand g869 (n_1245, A[17], n_378);
  nand g870 (n_397, n_1243, n_1244, n_1245);
  xor g871 (n_1246, n_379, n_380);
  xor g872 (n_386, n_1246, n_381);
  nand g873 (n_1247, n_379, n_380);
  nand g874 (n_1248, n_381, n_380);
  nand g875 (n_1249, n_379, n_381);
  nand g876 (n_398, n_1247, n_1248, n_1249);
  xor g877 (n_1250, n_118, n_383);
  xor g878 (n_388, n_1250, n_384);
  nand g879 (n_1251, n_118, n_383);
  nand g880 (n_1252, n_384, n_383);
  nand g881 (n_1253, n_118, n_384);
  nand g882 (n_402, n_1251, n_1252, n_1253);
  xor g883 (n_1254, n_385, n_386);
  xor g884 (n_390, n_1254, n_387);
  nand g885 (n_1255, n_385, n_386);
  nand g886 (n_1256, n_387, n_386);
  nand g887 (n_1257, n_385, n_387);
  nand g888 (n_404, n_1255, n_1256, n_1257);
  xor g889 (n_1258, n_388, n_389);
  xor g890 (n_170, n_1258, n_390);
  nand g891 (n_1259, n_388, n_389);
  nand g892 (n_1260, n_390, n_389);
  nand g893 (n_1261, n_388, n_390);
  nand g894 (n_99, n_1259, n_1260, n_1261);
  xor g895 (n_1262, A[22], A[20]);
  xor g896 (n_393, n_1262, A[8]);
  nand g897 (n_1263, A[22], A[20]);
  nand g898 (n_1264, A[8], A[20]);
  nand g899 (n_1265, A[22], A[8]);
  nand g900 (n_405, n_1263, n_1264, n_1265);
  xor g901 (n_1266, A[6], A[14]);
  xor g902 (n_394, n_1266, A[4]);
  nand g904 (n_1268, A[4], A[14]);
  xor g907 (n_1270, A[18], A[16]);
  xor g908 (n_396, n_1270, A[12]);
  nand g909 (n_1271, A[18], A[16]);
  nand g911 (n_1273, A[18], A[12]);
  nand g912 (n_409, n_1271, n_1143, n_1273);
  xor g913 (n_1274, A[10], n_391);
  xor g914 (n_399, n_1274, n_274);
  nand g915 (n_1275, A[10], n_391);
  nand g916 (n_1276, n_274, n_391);
  nand g917 (n_1277, A[10], n_274);
  nand g918 (n_411, n_1275, n_1276, n_1277);
  xor g919 (n_1278, n_393, n_394);
  xor g920 (n_400, n_1278, n_301);
  nand g921 (n_1279, n_393, n_394);
  nand g922 (n_1280, n_301, n_394);
  nand g923 (n_1281, n_393, n_301);
  nand g924 (n_412, n_1279, n_1280, n_1281);
  xor g925 (n_1282, n_396, n_397);
  xor g926 (n_401, n_1282, n_398);
  nand g927 (n_1283, n_396, n_397);
  nand g928 (n_1284, n_398, n_397);
  nand g929 (n_1285, n_396, n_398);
  nand g930 (n_416, n_1283, n_1284, n_1285);
  xor g931 (n_1286, n_399, n_400);
  xor g932 (n_403, n_1286, n_401);
  nand g933 (n_1287, n_399, n_400);
  nand g934 (n_1288, n_401, n_400);
  nand g935 (n_1289, n_399, n_401);
  nand g936 (n_418, n_1287, n_1288, n_1289);
  xor g937 (n_1290, n_402, n_403);
  xor g938 (n_169, n_1290, n_404);
  nand g939 (n_1291, n_402, n_403);
  nand g940 (n_1292, n_404, n_403);
  nand g941 (n_1293, n_402, n_404);
  nand g942 (n_98, n_1291, n_1292, n_1293);
  xor g943 (n_1294, A[23], A[21]);
  xor g944 (n_407, n_1294, A[9]);
  nand g945 (n_1295, A[23], A[21]);
  nand g946 (n_1296, A[9], A[21]);
  nand g947 (n_1297, A[23], A[9]);
  nand g948 (n_188, n_1295, n_1296, n_1297);
  xor g949 (n_1298, A[7], A[15]);
  xor g950 (n_408, n_1298, A[5]);
  nand g954 (n_189, n_1065, n_1168, n_951);
  xor g955 (n_1302, A[19], A[17]);
  xor g956 (n_410, n_1302, A[13]);
  nand g957 (n_1303, A[19], A[17]);
  nand g959 (n_1305, A[19], A[13]);
  nand g960 (n_420, n_1303, n_1120, n_1305);
  xor g961 (n_1306, A[11], n_405);
  xor g962 (n_413, n_1306, n_406);
  nand g963 (n_1307, A[11], n_405);
  nand g964 (n_1308, n_406, n_405);
  nand g965 (n_1309, A[11], n_406);
  nand g966 (n_423, n_1307, n_1308, n_1309);
  xor g967 (n_1310, n_407, n_408);
  xor g968 (n_414, n_1310, n_409);
  nand g969 (n_1311, n_407, n_408);
  nand g970 (n_1312, n_409, n_408);
  nand g971 (n_1313, n_407, n_409);
  nand g972 (n_424, n_1311, n_1312, n_1313);
  xor g973 (n_1314, n_410, n_411);
  xor g974 (n_415, n_1314, n_412);
  nand g975 (n_1315, n_410, n_411);
  nand g976 (n_1316, n_412, n_411);
  nand g977 (n_1317, n_410, n_412);
  nand g978 (n_428, n_1315, n_1316, n_1317);
  xor g979 (n_1318, n_413, n_414);
  xor g980 (n_417, n_1318, n_415);
  nand g981 (n_1319, n_413, n_414);
  nand g982 (n_1320, n_415, n_414);
  nand g983 (n_1321, n_413, n_415);
  nand g984 (n_430, n_1319, n_1320, n_1321);
  xor g985 (n_1322, n_416, n_417);
  xor g986 (n_168, n_1322, n_418);
  nand g987 (n_1323, n_416, n_417);
  nand g988 (n_1324, n_418, n_417);
  nand g989 (n_1325, n_416, n_418);
  nand g990 (n_97, n_1323, n_1324, n_1325);
  xor g991 (n_1326, A[22], A[18]);
  xor g992 (n_419, n_1326, A[8]);
  nand g993 (n_1327, A[22], A[18]);
  nand g994 (n_1328, A[8], A[18]);
  nand g996 (n_431, n_1327, n_1328, n_1265);
  xor g997 (n_1330, A[6], A[20]);
  xor g998 (n_421, n_1330, A[14]);
  nand g999 (n_1331, A[6], A[20]);
  nand g1002 (n_432, n_1331, n_1201, n_1141);
  xor g1003 (n_1334, A[10], A[24]);
  xor g1004 (n_422, n_1334, A[16]);
  nand g1005 (n_1335, A[10], A[24]);
  nand g1006 (n_1336, A[16], A[24]);
  nand g1007 (n_1337, A[10], A[16]);
  nand g1008 (n_434, n_1335, n_1336, n_1337);
  xor g1009 (n_1338, A[12], n_188);
  xor g1010 (n_425, n_1338, n_189);
  nand g1011 (n_1339, A[12], n_188);
  nand g1012 (n_1340, n_189, n_188);
  nand g1013 (n_1341, A[12], n_189);
  nand g1014 (n_437, n_1339, n_1340, n_1341);
  xor g1015 (n_1342, n_419, n_420);
  xor g1016 (n_426, n_1342, n_421);
  nand g1017 (n_1343, n_419, n_420);
  nand g1018 (n_1344, n_421, n_420);
  nand g1019 (n_1345, n_419, n_421);
  nand g1020 (n_438, n_1343, n_1344, n_1345);
  xor g1021 (n_1346, n_422, n_423);
  xor g1022 (n_427, n_1346, n_424);
  nand g1023 (n_1347, n_422, n_423);
  nand g1024 (n_1348, n_424, n_423);
  nand g1025 (n_1349, n_422, n_424);
  nand g1026 (n_442, n_1347, n_1348, n_1349);
  xor g1027 (n_1350, n_425, n_426);
  xor g1028 (n_429, n_1350, n_427);
  nand g1029 (n_1351, n_425, n_426);
  nand g1030 (n_1352, n_427, n_426);
  nand g1031 (n_1353, n_425, n_427);
  nand g1032 (n_444, n_1351, n_1352, n_1353);
  xor g1033 (n_1354, n_428, n_429);
  xor g1034 (n_167, n_1354, n_430);
  nand g1035 (n_1355, n_428, n_429);
  nand g1036 (n_1356, n_430, n_429);
  nand g1037 (n_1357, n_428, n_430);
  nand g1038 (n_96, n_1355, n_1356, n_1357);
  xor g1039 (n_1358, A[23], A[19]);
  xor g1040 (n_433, n_1358, A[9]);
  nand g1041 (n_1359, A[23], A[19]);
  nand g1042 (n_1360, A[9], A[19]);
  nand g1044 (n_445, n_1359, n_1360, n_1297);
  xor g1045 (n_1362, A[7], A[21]);
  xor g1046 (n_435, n_1362, A[15]);
  nand g1047 (n_1363, A[7], A[21]);
  nand g1050 (n_446, n_1363, n_1233, n_1065);
  xor g1051 (n_1366, A[11], A[25]);
  xor g1052 (n_436, n_1366, A[17]);
  nand g1053 (n_1367, A[11], A[25]);
  nand g1054 (n_1368, A[17], A[25]);
  nand g1055 (n_1369, A[11], A[17]);
  nand g1056 (n_449, n_1367, n_1368, n_1369);
  xor g1057 (n_1370, A[13], n_431);
  xor g1058 (n_439, n_1370, n_432);
  nand g1059 (n_1371, A[13], n_431);
  nand g1060 (n_1372, n_432, n_431);
  nand g1061 (n_1373, A[13], n_432);
  nand g1062 (n_451, n_1371, n_1372, n_1373);
  xor g1063 (n_1374, n_433, n_434);
  xor g1064 (n_440, n_1374, n_435);
  nand g1065 (n_1375, n_433, n_434);
  nand g1066 (n_1376, n_435, n_434);
  nand g1067 (n_1377, n_433, n_435);
  nand g1068 (n_452, n_1375, n_1376, n_1377);
  xor g1069 (n_1378, n_436, n_437);
  xor g1070 (n_441, n_1378, n_438);
  nand g1071 (n_1379, n_436, n_437);
  nand g1072 (n_1380, n_438, n_437);
  nand g1073 (n_1381, n_436, n_438);
  nand g1074 (n_456, n_1379, n_1380, n_1381);
  xor g1075 (n_1382, n_439, n_440);
  xor g1076 (n_443, n_1382, n_441);
  nand g1077 (n_1383, n_439, n_440);
  nand g1078 (n_1384, n_441, n_440);
  nand g1079 (n_1385, n_439, n_441);
  nand g1080 (n_458, n_1383, n_1384, n_1385);
  xor g1081 (n_1386, n_442, n_443);
  xor g1082 (n_166, n_1386, n_444);
  nand g1083 (n_1387, n_442, n_443);
  nand g1084 (n_1388, n_444, n_443);
  nand g1085 (n_1389, n_442, n_444);
  nand g1086 (n_95, n_1387, n_1388, n_1389);
  xor g1088 (n_447, n_1262, A[18]);
  nand g1092 (n_459, n_1263, n_1199, n_1327);
  xor g1094 (n_448, n_299, A[24]);
  nand g1096 (n_1396, A[24], A[14]);
  nand g1097 (n_1397, A[8], A[24]);
  xor g1099 (n_1398, A[12], A[10]);
  xor g1100 (n_450, n_1398, A[16]);
  nand g1104 (n_463, n_1008, n_1337, n_1143);
  xor g1105 (n_1402, A[26], n_445);
  xor g1106 (n_453, n_1402, n_446);
  nand g1107 (n_1403, A[26], n_445);
  nand g1108 (n_1404, n_446, n_445);
  nand g1109 (n_1405, A[26], n_446);
  nand g1110 (n_465, n_1403, n_1404, n_1405);
  xor g1111 (n_1406, n_447, n_448);
  xor g1112 (n_454, n_1406, n_449);
  nand g1113 (n_1407, n_447, n_448);
  nand g1114 (n_1408, n_449, n_448);
  nand g1115 (n_1409, n_447, n_449);
  nand g1116 (n_466, n_1407, n_1408, n_1409);
  xor g1117 (n_1410, n_450, n_451);
  xor g1118 (n_455, n_1410, n_452);
  nand g1119 (n_1411, n_450, n_451);
  nand g1120 (n_1412, n_452, n_451);
  nand g1121 (n_1413, n_450, n_452);
  nand g1122 (n_470, n_1411, n_1412, n_1413);
  xor g1123 (n_1414, n_453, n_454);
  xor g1124 (n_457, n_1414, n_455);
  nand g1125 (n_1415, n_453, n_454);
  nand g1126 (n_1416, n_455, n_454);
  nand g1127 (n_1417, n_453, n_455);
  nand g1128 (n_472, n_1415, n_1416, n_1417);
  xor g1129 (n_1418, n_456, n_457);
  xor g1130 (n_165, n_1418, n_458);
  nand g1131 (n_1419, n_456, n_457);
  nand g1132 (n_1420, n_458, n_457);
  nand g1133 (n_1421, n_456, n_458);
  nand g1134 (n_94, n_1419, n_1420, n_1421);
  xor g1136 (n_460, n_1294, A[19]);
  nand g1140 (n_473, n_1295, n_1231, n_1359);
  xor g1142 (n_461, n_1062, A[25]);
  nand g1144 (n_1428, A[25], A[15]);
  nand g1145 (n_1429, A[9], A[25]);
  nand g1146 (n_476, n_1063, n_1428, n_1429);
  xor g1148 (n_464, n_1026, A[17]);
  nand g1152 (n_477, n_1027, n_1369, n_1120);
  xor g1153 (n_1434, A[27], n_459);
  xor g1154 (n_467, n_1434, n_460);
  nand g1155 (n_1435, A[27], n_459);
  nand g1156 (n_1436, n_460, n_459);
  nand g1157 (n_1437, A[27], n_460);
  nand g1158 (n_480, n_1435, n_1436, n_1437);
  xor g1159 (n_1438, n_461, n_462);
  xor g1160 (n_468, n_1438, n_463);
  nand g1161 (n_1439, n_461, n_462);
  nand g1162 (n_1440, n_463, n_462);
  nand g1163 (n_1441, n_461, n_463);
  nand g1164 (n_479, n_1439, n_1440, n_1441);
  xor g1165 (n_1442, n_464, n_465);
  xor g1166 (n_469, n_1442, n_466);
  nand g1167 (n_1443, n_464, n_465);
  nand g1168 (n_1444, n_466, n_465);
  nand g1169 (n_1445, n_464, n_466);
  nand g1170 (n_483, n_1443, n_1444, n_1445);
  xor g1171 (n_1446, n_467, n_468);
  xor g1172 (n_471, n_1446, n_469);
  nand g1173 (n_1447, n_467, n_468);
  nand g1174 (n_1448, n_469, n_468);
  nand g1175 (n_1449, n_467, n_469);
  nand g1176 (n_486, n_1447, n_1448, n_1449);
  xor g1177 (n_1450, n_470, n_471);
  xor g1178 (n_164, n_1450, n_472);
  nand g1179 (n_1451, n_470, n_471);
  nand g1180 (n_1452, n_472, n_471);
  nand g1181 (n_1453, n_470, n_472);
  nand g1182 (n_93, n_1451, n_1452, n_1453);
  xor g1183 (n_1454, A[28], A[22]);
  xor g1184 (n_474, n_1454, A[14]);
  nand g1185 (n_1455, A[28], A[22]);
  nand g1186 (n_1456, A[14], A[22]);
  nand g1187 (n_1457, A[28], A[14]);
  nand g1188 (n_487, n_1455, n_1456, n_1457);
  xor g1190 (n_475, n_1198, A[26]);
  nand g1192 (n_1460, A[26], A[18]);
  nand g1193 (n_1461, A[20], A[26]);
  nand g1194 (n_490, n_1199, n_1460, n_1461);
  xor g1196 (n_478, n_1398, A[24]);
  nand g1199 (n_1465, A[12], A[24]);
  nand g1200 (n_491, n_1008, n_1335, n_1465);
  xor g1201 (n_1466, A[16], n_473);
  xor g1202 (n_481, n_1466, n_474);
  nand g1203 (n_1467, A[16], n_473);
  nand g1204 (n_1468, n_474, n_473);
  nand g1205 (n_1469, A[16], n_474);
  nand g1206 (n_494, n_1467, n_1468, n_1469);
  xor g1207 (n_1470, n_475, n_476);
  xor g1208 (n_482, n_1470, n_477);
  nand g1209 (n_1471, n_475, n_476);
  nand g1210 (n_1472, n_477, n_476);
  nand g1211 (n_1473, n_475, n_477);
  nand g1212 (n_493, n_1471, n_1472, n_1473);
  xor g1213 (n_1474, n_478, n_479);
  xor g1214 (n_484, n_1474, n_480);
  nand g1215 (n_1475, n_478, n_479);
  nand g1216 (n_1476, n_480, n_479);
  nand g1217 (n_1477, n_478, n_480);
  nand g1218 (n_497, n_1475, n_1476, n_1477);
  xor g1219 (n_1478, n_481, n_482);
  xor g1220 (n_485, n_1478, n_483);
  nand g1221 (n_1479, n_481, n_482);
  nand g1222 (n_1480, n_483, n_482);
  nand g1223 (n_1481, n_481, n_483);
  nand g1224 (n_500, n_1479, n_1480, n_1481);
  xor g1225 (n_1482, n_484, n_485);
  xor g1226 (n_163, n_1482, n_486);
  nand g1227 (n_1483, n_484, n_485);
  nand g1228 (n_1484, n_486, n_485);
  nand g1229 (n_1485, n_484, n_486);
  nand g1230 (n_92, n_1483, n_1484, n_1485);
  xor g1231 (n_1486, A[29], A[23]);
  xor g1232 (n_488, n_1486, A[15]);
  nand g1233 (n_1487, A[29], A[23]);
  nand g1234 (n_1488, A[15], A[23]);
  nand g1235 (n_1489, A[29], A[15]);
  nand g1236 (n_501, n_1487, n_1488, n_1489);
  xor g1238 (n_489, n_1230, A[27]);
  nand g1240 (n_1492, A[27], A[19]);
  nand g1241 (n_1493, A[21], A[27]);
  nand g1242 (n_504, n_1231, n_1492, n_1493);
  xor g1244 (n_492, n_1026, A[25]);
  nand g1247 (n_1497, A[13], A[25]);
  nand g1248 (n_503, n_1027, n_1367, n_1497);
  xor g1249 (n_1498, A[17], n_487);
  xor g1250 (n_495, n_1498, n_488);
  nand g1251 (n_1499, A[17], n_487);
  nand g1252 (n_1500, n_488, n_487);
  nand g1253 (n_1501, A[17], n_488);
  nand g1254 (n_508, n_1499, n_1500, n_1501);
  xor g1255 (n_1502, n_489, n_490);
  xor g1256 (n_496, n_1502, n_491);
  nand g1257 (n_1503, n_489, n_490);
  nand g1258 (n_1504, n_491, n_490);
  nand g1259 (n_1505, n_489, n_491);
  nand g1260 (n_507, n_1503, n_1504, n_1505);
  xor g1261 (n_1506, n_492, n_493);
  xor g1262 (n_498, n_1506, n_494);
  nand g1263 (n_1507, n_492, n_493);
  nand g1264 (n_1508, n_494, n_493);
  nand g1265 (n_1509, n_492, n_494);
  nand g1266 (n_511, n_1507, n_1508, n_1509);
  xor g1267 (n_1510, n_495, n_496);
  xor g1268 (n_499, n_1510, n_497);
  nand g1269 (n_1511, n_495, n_496);
  nand g1270 (n_1512, n_497, n_496);
  nand g1271 (n_1513, n_495, n_497);
  nand g1272 (n_514, n_1511, n_1512, n_1513);
  xor g1273 (n_1514, n_498, n_499);
  xor g1274 (n_162, n_1514, n_500);
  nand g1275 (n_1515, n_498, n_499);
  nand g1276 (n_1516, n_500, n_499);
  nand g1277 (n_1517, n_498, n_500);
  nand g1278 (n_91, n_1515, n_1516, n_1517);
  xor g1286 (n_505, n_1198, A[16]);
  nand g1289 (n_1525, A[20], A[16]);
  nand g1290 (n_518, n_1199, n_1271, n_1525);
  xor g1291 (n_1526, A[24], A[30]);
  xor g1292 (n_506, n_1526, A[12]);
  nand g1293 (n_1527, A[24], A[30]);
  nand g1294 (n_1528, A[12], A[30]);
  nand g1296 (n_517, n_1527, n_1528, n_1465);
  xor g1297 (n_1530, A[26], n_501);
  xor g1298 (n_509, n_1530, n_474);
  nand g1299 (n_1531, A[26], n_501);
  nand g1300 (n_1532, n_474, n_501);
  nand g1301 (n_1533, A[26], n_474);
  nand g1302 (n_522, n_1531, n_1532, n_1533);
  xor g1303 (n_1534, n_503, n_504);
  xor g1304 (n_510, n_1534, n_505);
  nand g1305 (n_1535, n_503, n_504);
  nand g1306 (n_1536, n_505, n_504);
  nand g1307 (n_1537, n_503, n_505);
  nand g1308 (n_521, n_1535, n_1536, n_1537);
  xor g1309 (n_1538, n_506, n_507);
  xor g1310 (n_512, n_1538, n_508);
  nand g1311 (n_1539, n_506, n_507);
  nand g1312 (n_1540, n_508, n_507);
  nand g1313 (n_1541, n_506, n_508);
  nand g1314 (n_525, n_1539, n_1540, n_1541);
  xor g1315 (n_1542, n_509, n_510);
  xor g1316 (n_513, n_1542, n_511);
  nand g1317 (n_1543, n_509, n_510);
  nand g1318 (n_1544, n_511, n_510);
  nand g1319 (n_1545, n_509, n_511);
  nand g1320 (n_528, n_1543, n_1544, n_1545);
  xor g1321 (n_1546, n_512, n_513);
  xor g1322 (n_161, n_1546, n_514);
  nand g1323 (n_1547, n_512, n_513);
  nand g1324 (n_1548, n_514, n_513);
  nand g1325 (n_1549, n_512, n_514);
  nand g1326 (n_90, n_1547, n_1548, n_1549);
  xor g1334 (n_519, n_1230, A[17]);
  nand g1337 (n_1557, A[21], A[17]);
  nand g1338 (n_532, n_1231, n_1303, n_1557);
  xor g1339 (n_1558, A[25], A[31]);
  xor g1340 (n_520, n_1558, A[13]);
  nand g1341 (n_1559, A[25], A[31]);
  nand g1342 (n_1560, A[13], A[31]);
  nand g1344 (n_531, n_1559, n_1560, n_1497);
  xor g1345 (n_1562, A[27], n_487);
  xor g1346 (n_523, n_1562, n_488);
  nand g1347 (n_1563, A[27], n_487);
  nand g1349 (n_1565, A[27], n_488);
  nand g1350 (n_536, n_1563, n_1500, n_1565);
  xor g1351 (n_1566, n_517, n_518);
  xor g1352 (n_524, n_1566, n_519);
  nand g1353 (n_1567, n_517, n_518);
  nand g1354 (n_1568, n_519, n_518);
  nand g1355 (n_1569, n_517, n_519);
  nand g1356 (n_535, n_1567, n_1568, n_1569);
  xor g1357 (n_1570, n_520, n_521);
  xor g1358 (n_526, n_1570, n_522);
  nand g1359 (n_1571, n_520, n_521);
  nand g1360 (n_1572, n_522, n_521);
  nand g1361 (n_1573, n_520, n_522);
  nand g1362 (n_539, n_1571, n_1572, n_1573);
  xor g1363 (n_1574, n_523, n_524);
  xor g1364 (n_527, n_1574, n_525);
  nand g1365 (n_1575, n_523, n_524);
  nand g1366 (n_1576, n_525, n_524);
  nand g1367 (n_1577, n_523, n_525);
  nand g1368 (n_542, n_1575, n_1576, n_1577);
  xor g1369 (n_1578, n_526, n_527);
  xor g1370 (n_160, n_1578, n_528);
  nand g1371 (n_1579, n_526, n_527);
  nand g1372 (n_1580, n_528, n_527);
  nand g1373 (n_1581, n_526, n_528);
  nand g1374 (n_89, n_1579, n_1580, n_1581);
  xor g1375 (n_1582, A[28], A[18]);
  xor g1376 (n_530, n_1582, A[14]);
  nand g1377 (n_1583, A[28], A[18]);
  nand g1380 (n_543, n_1583, n_1200, n_1457);
  xor g1382 (n_533, n_1262, A[30]);
  nand g1384 (n_1588, A[30], A[20]);
  nand g1385 (n_1589, A[22], A[30]);
  nand g1386 (n_546, n_1263, n_1588, n_1589);
  xor g1387 (n_1590, A[26], A[16]);
  xor g1388 (n_534, n_1590, A[24]);
  nand g1389 (n_1591, A[26], A[16]);
  nand g1391 (n_1593, A[26], A[24]);
  nand g1392 (n_545, n_1591, n_1336, n_1593);
  xor g1393 (n_1594, A[32], n_501);
  xor g1394 (n_537, n_1594, n_530);
  nand g1395 (n_1595, A[32], n_501);
  nand g1396 (n_1596, n_530, n_501);
  nand g1397 (n_1597, A[32], n_530);
  nand g1398 (n_550, n_1595, n_1596, n_1597);
  xor g1399 (n_1598, n_531, n_532);
  xor g1400 (n_538, n_1598, n_533);
  nand g1401 (n_1599, n_531, n_532);
  nand g1402 (n_1600, n_533, n_532);
  nand g1403 (n_1601, n_531, n_533);
  nand g1404 (n_549, n_1599, n_1600, n_1601);
  xor g1405 (n_1602, n_534, n_535);
  xor g1406 (n_540, n_1602, n_536);
  nand g1407 (n_1603, n_534, n_535);
  nand g1408 (n_1604, n_536, n_535);
  nand g1409 (n_1605, n_534, n_536);
  nand g1410 (n_553, n_1603, n_1604, n_1605);
  xor g1411 (n_1606, n_537, n_538);
  xor g1412 (n_541, n_1606, n_539);
  nand g1413 (n_1607, n_537, n_538);
  nand g1414 (n_1608, n_539, n_538);
  nand g1415 (n_1609, n_537, n_539);
  nand g1416 (n_556, n_1607, n_1608, n_1609);
  xor g1417 (n_1610, n_540, n_541);
  xor g1418 (n_159, n_1610, n_542);
  nand g1419 (n_1611, n_540, n_541);
  nand g1420 (n_1612, n_542, n_541);
  nand g1421 (n_1613, n_540, n_542);
  nand g1422 (n_88, n_1611, n_1612, n_1613);
  xor g1423 (n_1614, A[29], A[19]);
  xor g1424 (n_544, n_1614, A[15]);
  nand g1425 (n_1615, A[29], A[19]);
  nand g1428 (n_557, n_1615, n_1169, n_1489);
  xor g1430 (n_547, n_1294, A[31]);
  nand g1432 (n_1620, A[31], A[21]);
  nand g1433 (n_1621, A[23], A[31]);
  nand g1434 (n_559, n_1295, n_1620, n_1621);
  xor g1435 (n_1622, A[27], A[17]);
  xor g1436 (n_548, n_1622, A[25]);
  nand g1437 (n_1623, A[27], A[17]);
  nand g1439 (n_1625, A[27], A[25]);
  nand g1440 (n_560, n_1623, n_1368, n_1625);
  xor g1441 (n_1626, A[33], n_543);
  xor g1442 (n_551, n_1626, n_544);
  nand g1443 (n_1627, A[33], n_543);
  nand g1444 (n_1628, n_544, n_543);
  nand g1445 (n_1629, A[33], n_544);
  nand g1446 (n_563, n_1627, n_1628, n_1629);
  xor g1447 (n_1630, n_545, n_546);
  xor g1448 (n_552, n_1630, n_547);
  nand g1449 (n_1631, n_545, n_546);
  nand g1450 (n_1632, n_547, n_546);
  nand g1451 (n_1633, n_545, n_547);
  nand g1452 (n_564, n_1631, n_1632, n_1633);
  xor g1453 (n_1634, n_548, n_549);
  xor g1454 (n_554, n_1634, n_550);
  nand g1455 (n_1635, n_548, n_549);
  nand g1456 (n_1636, n_550, n_549);
  nand g1457 (n_1637, n_548, n_550);
  nand g1458 (n_567, n_1635, n_1636, n_1637);
  xor g1459 (n_1638, n_551, n_552);
  xor g1460 (n_555, n_1638, n_553);
  nand g1461 (n_1639, n_551, n_552);
  nand g1462 (n_1640, n_553, n_552);
  nand g1463 (n_1641, n_551, n_553);
  nand g1464 (n_570, n_1639, n_1640, n_1641);
  xor g1465 (n_1642, n_554, n_555);
  xor g1466 (n_158, n_1642, n_556);
  nand g1467 (n_1643, n_554, n_555);
  nand g1468 (n_1644, n_556, n_555);
  nand g1469 (n_1645, n_554, n_556);
  nand g1470 (n_87, n_1643, n_1644, n_1645);
  xor g1471 (n_1646, A[28], A[20]);
  xor g1472 (n_558, n_1646, A[18]);
  nand g1473 (n_1647, A[28], A[20]);
  nand g1476 (n_571, n_1647, n_1199, n_1583);
  xor g1477 (n_1650, A[22], A[32]);
  xor g1478 (n_561, n_1650, A[34]);
  nand g1479 (n_1651, A[22], A[32]);
  nand g1480 (n_1652, A[34], A[32]);
  nand g1481 (n_1653, A[22], A[34]);
  nand g1482 (n_573, n_1651, n_1652, n_1653);
  xor g1489 (n_1658, A[30], n_557);
  xor g1490 (n_565, n_1658, n_558);
  nand g1491 (n_1659, A[30], n_557);
  nand g1492 (n_1660, n_558, n_557);
  nand g1493 (n_1661, A[30], n_558);
  nand g1494 (n_577, n_1659, n_1660, n_1661);
  xor g1495 (n_1662, n_559, n_560);
  xor g1496 (n_566, n_1662, n_561);
  nand g1497 (n_1663, n_559, n_560);
  nand g1498 (n_1664, n_561, n_560);
  nand g1499 (n_1665, n_559, n_561);
  nand g1500 (n_580, n_1663, n_1664, n_1665);
  xor g1501 (n_1666, n_534, n_563);
  xor g1502 (n_568, n_1666, n_564);
  nand g1503 (n_1667, n_534, n_563);
  nand g1504 (n_1668, n_564, n_563);
  nand g1505 (n_1669, n_534, n_564);
  nand g1506 (n_581, n_1667, n_1668, n_1669);
  xor g1507 (n_1670, n_565, n_566);
  xor g1508 (n_569, n_1670, n_567);
  nand g1509 (n_1671, n_565, n_566);
  nand g1510 (n_1672, n_567, n_566);
  nand g1511 (n_1673, n_565, n_567);
  nand g1512 (n_584, n_1671, n_1672, n_1673);
  xor g1513 (n_1674, n_568, n_569);
  xor g1514 (n_157, n_1674, n_570);
  nand g1515 (n_1675, n_568, n_569);
  nand g1516 (n_1676, n_570, n_569);
  nand g1517 (n_1677, n_568, n_570);
  nand g1518 (n_86, n_1675, n_1676, n_1677);
  xor g1519 (n_1678, A[29], A[21]);
  xor g1520 (n_572, n_1678, A[19]);
  nand g1521 (n_1679, A[29], A[21]);
  nand g1524 (n_585, n_1679, n_1231, n_1615);
  xor g1525 (n_1682, A[23], A[33]);
  xor g1526 (n_575, n_1682, A[35]);
  nand g1527 (n_1683, A[23], A[33]);
  nand g1528 (n_1684, A[35], A[33]);
  nand g1529 (n_1685, A[23], A[35]);
  nand g1530 (n_587, n_1683, n_1684, n_1685);
  xor g1537 (n_1690, A[31], n_571);
  xor g1538 (n_578, n_1690, n_572);
  nand g1539 (n_1691, A[31], n_571);
  nand g1540 (n_1692, n_572, n_571);
  nand g1541 (n_1693, A[31], n_572);
  nand g1542 (n_591, n_1691, n_1692, n_1693);
  xor g1543 (n_1694, n_573, n_545);
  xor g1544 (n_579, n_1694, n_575);
  nand g1545 (n_1695, n_573, n_545);
  nand g1546 (n_1696, n_575, n_545);
  nand g1547 (n_1697, n_573, n_575);
  nand g1548 (n_594, n_1695, n_1696, n_1697);
  xor g1549 (n_1698, n_548, n_577);
  xor g1550 (n_582, n_1698, n_578);
  nand g1551 (n_1699, n_548, n_577);
  nand g1552 (n_1700, n_578, n_577);
  nand g1553 (n_1701, n_548, n_578);
  nand g1554 (n_595, n_1699, n_1700, n_1701);
  xor g1555 (n_1702, n_579, n_580);
  xor g1556 (n_583, n_1702, n_581);
  nand g1557 (n_1703, n_579, n_580);
  nand g1558 (n_1704, n_581, n_580);
  nand g1559 (n_1705, n_579, n_581);
  nand g1560 (n_598, n_1703, n_1704, n_1705);
  xor g1561 (n_1706, n_582, n_583);
  xor g1562 (n_156, n_1706, n_584);
  nand g1563 (n_1707, n_582, n_583);
  nand g1564 (n_1708, n_584, n_583);
  nand g1565 (n_1709, n_582, n_584);
  nand g1566 (n_85, n_1707, n_1708, n_1709);
  xor g1568 (n_586, n_1454, A[20]);
  nand g1572 (n_599, n_1455, n_1263, n_1647);
  xor g1573 (n_1714, A[18], A[30]);
  xor g1574 (n_590, n_1714, A[36]);
  nand g1575 (n_1715, A[18], A[30]);
  nand g1576 (n_1716, A[36], A[30]);
  nand g1577 (n_1717, A[18], A[36]);
  nand g1578 (n_601, n_1715, n_1716, n_1717);
  xor g1579 (n_1718, A[34], A[32]);
  xor g1580 (n_589, n_1718, A[26]);
  nand g1582 (n_1720, A[26], A[32]);
  nand g1583 (n_1721, A[34], A[26]);
  nand g1584 (n_602, n_1652, n_1720, n_1721);
  xor g1585 (n_1722, A[24], n_585);
  xor g1586 (n_592, n_1722, n_586);
  nand g1587 (n_1723, A[24], n_585);
  nand g1588 (n_1724, n_586, n_585);
  nand g1589 (n_1725, A[24], n_586);
  nand g1590 (n_605, n_1723, n_1724, n_1725);
  xor g1591 (n_1726, n_587, n_560);
  xor g1592 (n_593, n_1726, n_589);
  nand g1593 (n_1727, n_587, n_560);
  nand g1594 (n_1728, n_589, n_560);
  nand g1595 (n_1729, n_587, n_589);
  nand g1596 (n_608, n_1727, n_1728, n_1729);
  xor g1597 (n_1730, n_590, n_591);
  xor g1598 (n_596, n_1730, n_592);
  nand g1599 (n_1731, n_590, n_591);
  nand g1600 (n_1732, n_592, n_591);
  nand g1601 (n_1733, n_590, n_592);
  nand g1602 (n_609, n_1731, n_1732, n_1733);
  xor g1603 (n_1734, n_593, n_594);
  xor g1604 (n_597, n_1734, n_595);
  nand g1605 (n_1735, n_593, n_594);
  nand g1606 (n_1736, n_595, n_594);
  nand g1607 (n_1737, n_593, n_595);
  nand g1608 (n_612, n_1735, n_1736, n_1737);
  xor g1609 (n_1738, n_596, n_597);
  xor g1610 (n_155, n_1738, n_598);
  nand g1611 (n_1739, n_596, n_597);
  nand g1612 (n_1740, n_598, n_597);
  nand g1613 (n_1741, n_596, n_598);
  nand g1614 (n_84, n_1739, n_1740, n_1741);
  xor g1616 (n_600, n_1486, A[21]);
  nand g1620 (n_613, n_1487, n_1295, n_1679);
  xor g1621 (n_1746, A[19], A[31]);
  xor g1622 (n_604, n_1746, A[37]);
  nand g1623 (n_1747, A[19], A[31]);
  nand g1624 (n_1748, A[37], A[31]);
  nand g1625 (n_1749, A[19], A[37]);
  nand g1626 (n_615, n_1747, n_1748, n_1749);
  xor g1627 (n_1750, A[35], A[33]);
  xor g1628 (n_603, n_1750, A[27]);
  nand g1630 (n_1752, A[27], A[33]);
  nand g1631 (n_1753, A[35], A[27]);
  nand g1632 (n_616, n_1684, n_1752, n_1753);
  xor g1633 (n_1754, A[25], n_599);
  xor g1634 (n_606, n_1754, n_600);
  nand g1635 (n_1755, A[25], n_599);
  nand g1636 (n_1756, n_600, n_599);
  nand g1637 (n_1757, A[25], n_600);
  nand g1638 (n_619, n_1755, n_1756, n_1757);
  xor g1639 (n_1758, n_601, n_602);
  xor g1640 (n_607, n_1758, n_603);
  nand g1641 (n_1759, n_601, n_602);
  nand g1642 (n_1760, n_603, n_602);
  nand g1643 (n_1761, n_601, n_603);
  nand g1644 (n_622, n_1759, n_1760, n_1761);
  xor g1645 (n_1762, n_604, n_605);
  xor g1646 (n_610, n_1762, n_606);
  nand g1647 (n_1763, n_604, n_605);
  nand g1648 (n_1764, n_606, n_605);
  nand g1649 (n_1765, n_604, n_606);
  nand g1650 (n_623, n_1763, n_1764, n_1765);
  xor g1651 (n_1766, n_607, n_608);
  xor g1652 (n_611, n_1766, n_609);
  nand g1653 (n_1767, n_607, n_608);
  nand g1654 (n_1768, n_609, n_608);
  nand g1655 (n_1769, n_607, n_609);
  nand g1656 (n_626, n_1767, n_1768, n_1769);
  xor g1657 (n_1770, n_610, n_611);
  xor g1658 (n_154, n_1770, n_612);
  nand g1659 (n_1771, n_610, n_611);
  nand g1660 (n_1772, n_612, n_611);
  nand g1661 (n_1773, n_610, n_612);
  nand g1662 (n_83, n_1771, n_1772, n_1773);
  xor g1669 (n_1778, A[36], A[24]);
  xor g1670 (n_618, n_1778, A[32]);
  nand g1671 (n_1779, A[36], A[24]);
  nand g1672 (n_1780, A[32], A[24]);
  nand g1673 (n_1781, A[36], A[32]);
  nand g1674 (n_629, n_1779, n_1780, n_1781);
  xor g1675 (n_1782, A[30], A[38]);
  xor g1676 (n_617, n_1782, A[34]);
  nand g1677 (n_1783, A[30], A[38]);
  nand g1678 (n_1784, A[34], A[38]);
  nand g1679 (n_1785, A[30], A[34]);
  nand g1680 (n_630, n_1783, n_1784, n_1785);
  xor g1681 (n_1786, A[26], n_613);
  xor g1682 (n_620, n_1786, n_586);
  nand g1683 (n_1787, A[26], n_613);
  nand g1684 (n_1788, n_586, n_613);
  nand g1685 (n_1789, A[26], n_586);
  nand g1686 (n_633, n_1787, n_1788, n_1789);
  xor g1687 (n_1790, n_615, n_616);
  xor g1688 (n_621, n_1790, n_617);
  nand g1689 (n_1791, n_615, n_616);
  nand g1690 (n_1792, n_617, n_616);
  nand g1691 (n_1793, n_615, n_617);
  nand g1692 (n_636, n_1791, n_1792, n_1793);
  xor g1693 (n_1794, n_618, n_619);
  xor g1694 (n_624, n_1794, n_620);
  nand g1695 (n_1795, n_618, n_619);
  nand g1696 (n_1796, n_620, n_619);
  nand g1697 (n_1797, n_618, n_620);
  nand g1698 (n_637, n_1795, n_1796, n_1797);
  xor g1699 (n_1798, n_621, n_622);
  xor g1700 (n_625, n_1798, n_623);
  nand g1701 (n_1799, n_621, n_622);
  nand g1702 (n_1800, n_623, n_622);
  nand g1703 (n_1801, n_621, n_623);
  nand g1704 (n_640, n_1799, n_1800, n_1801);
  xor g1705 (n_1802, n_624, n_625);
  xor g1706 (n_153, n_1802, n_626);
  nand g1707 (n_1803, n_624, n_625);
  nand g1708 (n_1804, n_626, n_625);
  nand g1709 (n_1805, n_624, n_626);
  nand g1710 (n_82, n_1803, n_1804, n_1805);
  xor g1717 (n_1810, A[37], A[25]);
  xor g1718 (n_632, n_1810, A[33]);
  nand g1719 (n_1811, A[37], A[25]);
  nand g1720 (n_1812, A[33], A[25]);
  nand g1721 (n_1813, A[37], A[33]);
  nand g1722 (n_643, n_1811, n_1812, n_1813);
  xor g1723 (n_1814, A[31], A[39]);
  xor g1724 (n_631, n_1814, A[35]);
  nand g1725 (n_1815, A[31], A[39]);
  nand g1726 (n_1816, A[35], A[39]);
  nand g1727 (n_1817, A[31], A[35]);
  nand g1728 (n_644, n_1815, n_1816, n_1817);
  xor g1729 (n_1818, A[27], n_599);
  xor g1730 (n_634, n_1818, n_600);
  nand g1731 (n_1819, A[27], n_599);
  nand g1733 (n_1821, A[27], n_600);
  nand g1734 (n_647, n_1819, n_1756, n_1821);
  xor g1735 (n_1822, n_629, n_630);
  xor g1736 (n_635, n_1822, n_631);
  nand g1737 (n_1823, n_629, n_630);
  nand g1738 (n_1824, n_631, n_630);
  nand g1739 (n_1825, n_629, n_631);
  nand g1740 (n_650, n_1823, n_1824, n_1825);
  xor g1741 (n_1826, n_632, n_633);
  xor g1742 (n_638, n_1826, n_634);
  nand g1743 (n_1827, n_632, n_633);
  nand g1744 (n_1828, n_634, n_633);
  nand g1745 (n_1829, n_632, n_634);
  nand g1746 (n_651, n_1827, n_1828, n_1829);
  xor g1747 (n_1830, n_635, n_636);
  xor g1748 (n_639, n_1830, n_637);
  nand g1749 (n_1831, n_635, n_636);
  nand g1750 (n_1832, n_637, n_636);
  nand g1751 (n_1833, n_635, n_637);
  nand g1752 (n_654, n_1831, n_1832, n_1833);
  xor g1753 (n_1834, n_638, n_639);
  xor g1754 (n_152, n_1834, n_640);
  nand g1755 (n_1835, n_638, n_639);
  nand g1756 (n_1836, n_640, n_639);
  nand g1757 (n_1837, n_638, n_640);
  nand g1758 (n_81, n_1835, n_1836, n_1837);
  xor g1760 (n_642, n_1454, A[34]);
  nand g1763 (n_1841, A[28], A[34]);
  nand g1764 (n_656, n_1455, n_1653, n_1841);
  xor g1765 (n_1842, A[26], A[24]);
  xor g1766 (n_646, n_1842, A[38]);
  nand g1768 (n_1844, A[38], A[24]);
  nand g1769 (n_1845, A[26], A[38]);
  nand g1770 (n_657, n_1593, n_1844, n_1845);
  xor g1771 (n_1846, A[32], A[40]);
  xor g1772 (n_645, n_1846, A[30]);
  nand g1773 (n_1847, A[32], A[40]);
  nand g1774 (n_1848, A[30], A[40]);
  nand g1775 (n_1849, A[32], A[30]);
  nand g1776 (n_658, n_1847, n_1848, n_1849);
  xor g1777 (n_1850, A[36], n_613);
  xor g1778 (n_648, n_1850, n_642);
  nand g1779 (n_1851, A[36], n_613);
  nand g1780 (n_1852, n_642, n_613);
  nand g1781 (n_1853, A[36], n_642);
  nand g1782 (n_661, n_1851, n_1852, n_1853);
  xor g1783 (n_1854, n_643, n_644);
  xor g1784 (n_649, n_1854, n_645);
  nand g1785 (n_1855, n_643, n_644);
  nand g1786 (n_1856, n_645, n_644);
  nand g1787 (n_1857, n_643, n_645);
  nand g1788 (n_663, n_1855, n_1856, n_1857);
  xor g1789 (n_1858, n_646, n_647);
  xor g1790 (n_652, n_1858, n_648);
  nand g1791 (n_1859, n_646, n_647);
  nand g1792 (n_1860, n_648, n_647);
  nand g1793 (n_1861, n_646, n_648);
  nand g1794 (n_665, n_1859, n_1860, n_1861);
  xor g1795 (n_1862, n_649, n_650);
  xor g1796 (n_653, n_1862, n_651);
  nand g1797 (n_1863, n_649, n_650);
  nand g1798 (n_1864, n_651, n_650);
  nand g1799 (n_1865, n_649, n_651);
  nand g1800 (n_668, n_1863, n_1864, n_1865);
  xor g1801 (n_1866, n_652, n_653);
  xor g1802 (n_151, n_1866, n_654);
  nand g1803 (n_1867, n_652, n_653);
  nand g1804 (n_1868, n_654, n_653);
  nand g1805 (n_1869, n_652, n_654);
  nand g1806 (n_80, n_1867, n_1868, n_1869);
  xor g1808 (n_655, n_1486, A[35]);
  nand g1811 (n_1873, A[29], A[35]);
  nand g1812 (n_669, n_1487, n_1685, n_1873);
  xor g1813 (n_1874, A[27], A[25]);
  xor g1814 (n_660, n_1874, A[39]);
  nand g1816 (n_1876, A[39], A[25]);
  nand g1817 (n_1877, A[27], A[39]);
  nand g1818 (n_670, n_1625, n_1876, n_1877);
  xor g1819 (n_1878, A[33], A[41]);
  xor g1820 (n_659, n_1878, A[31]);
  nand g1821 (n_1879, A[33], A[41]);
  nand g1822 (n_1880, A[31], A[41]);
  nand g1823 (n_1881, A[33], A[31]);
  nand g1824 (n_671, n_1879, n_1880, n_1881);
  xor g1825 (n_1882, A[37], n_655);
  xor g1826 (n_664, n_1882, n_656);
  nand g1827 (n_1883, A[37], n_655);
  nand g1828 (n_1884, n_656, n_655);
  nand g1829 (n_1885, A[37], n_656);
  nand g1830 (n_675, n_1883, n_1884, n_1885);
  xor g1831 (n_1886, n_657, n_658);
  xor g1832 (n_662, n_1886, n_659);
  nand g1833 (n_1887, n_657, n_658);
  nand g1834 (n_1888, n_659, n_658);
  nand g1835 (n_1889, n_657, n_659);
  nand g1836 (n_677, n_1887, n_1888, n_1889);
  xor g1837 (n_1890, n_660, n_661);
  xor g1838 (n_666, n_1890, n_662);
  nand g1839 (n_1891, n_660, n_661);
  nand g1840 (n_1892, n_662, n_661);
  nand g1841 (n_1893, n_660, n_662);
  nand g1842 (n_679, n_1891, n_1892, n_1893);
  xor g1843 (n_1894, n_663, n_664);
  xor g1844 (n_667, n_1894, n_665);
  nand g1845 (n_1895, n_663, n_664);
  nand g1846 (n_1896, n_665, n_664);
  nand g1847 (n_1897, n_663, n_665);
  nand g1848 (n_681, n_1895, n_1896, n_1897);
  xor g1849 (n_1898, n_666, n_667);
  xor g1850 (n_150, n_1898, n_668);
  nand g1851 (n_1899, n_666, n_667);
  nand g1852 (n_1900, n_668, n_667);
  nand g1853 (n_1901, n_666, n_668);
  nand g1854 (n_79, n_1899, n_1900, n_1901);
  xor g1855 (n_1902, A[28], A[42]);
  xor g1856 (n_673, n_1902, A[40]);
  nand g1857 (n_1903, A[28], A[42]);
  nand g1858 (n_1904, A[40], A[42]);
  nand g1859 (n_1905, A[28], A[40]);
  nand g1860 (n_683, n_1903, n_1904, n_1905);
  xor g1861 (n_1906, A[36], A[26]);
  xor g1862 (n_674, n_1906, A[34]);
  nand g1863 (n_1907, A[36], A[26]);
  nand g1865 (n_1909, A[36], A[34]);
  nand g1866 (n_684, n_1907, n_1721, n_1909);
  xor g1867 (n_1910, A[24], A[38]);
  xor g1868 (n_672, n_1910, A[32]);
  nand g1870 (n_1912, A[32], A[38]);
  nand g1872 (n_685, n_1844, n_1912, n_1780);
  xor g1873 (n_1914, A[30], n_669);
  xor g1874 (n_676, n_1914, n_670);
  nand g1875 (n_1915, A[30], n_669);
  nand g1876 (n_1916, n_670, n_669);
  nand g1877 (n_1917, A[30], n_670);
  nand g1878 (n_689, n_1915, n_1916, n_1917);
  xor g1879 (n_1918, n_671, n_672);
  xor g1880 (n_678, n_1918, n_673);
  nand g1881 (n_1919, n_671, n_672);
  nand g1882 (n_1920, n_673, n_672);
  nand g1883 (n_1921, n_671, n_673);
  nand g1884 (n_691, n_1919, n_1920, n_1921);
  xor g1885 (n_1922, n_674, n_675);
  xor g1886 (n_680, n_1922, n_676);
  nand g1887 (n_1923, n_674, n_675);
  nand g1888 (n_1924, n_676, n_675);
  nand g1889 (n_1925, n_674, n_676);
  nand g1890 (n_693, n_1923, n_1924, n_1925);
  xor g1891 (n_1926, n_677, n_678);
  xor g1892 (n_682, n_1926, n_679);
  nand g1893 (n_1927, n_677, n_678);
  nand g1894 (n_1928, n_679, n_678);
  nand g1895 (n_1929, n_677, n_679);
  nand g1896 (n_696, n_1927, n_1928, n_1929);
  xor g1897 (n_1930, n_680, n_681);
  xor g1898 (n_149, n_1930, n_682);
  nand g1899 (n_1931, n_680, n_681);
  nand g1900 (n_1932, n_682, n_681);
  nand g1901 (n_1933, n_680, n_682);
  nand g1902 (n_78, n_1931, n_1932, n_1933);
  xor g1903 (n_1934, A[29], A[43]);
  xor g1904 (n_687, n_1934, A[41]);
  nand g1905 (n_1935, A[29], A[43]);
  nand g1906 (n_1936, A[41], A[43]);
  nand g1907 (n_1937, A[29], A[41]);
  nand g1908 (n_697, n_1935, n_1936, n_1937);
  xor g1909 (n_1938, A[37], A[27]);
  xor g1910 (n_688, n_1938, A[35]);
  nand g1911 (n_1939, A[37], A[27]);
  nand g1913 (n_1941, A[37], A[35]);
  nand g1914 (n_698, n_1939, n_1753, n_1941);
  xor g1915 (n_1942, A[25], A[39]);
  xor g1916 (n_686, n_1942, A[33]);
  nand g1918 (n_1944, A[33], A[39]);
  nand g1920 (n_699, n_1876, n_1944, n_1812);
  xor g1921 (n_1946, A[31], n_683);
  xor g1922 (n_690, n_1946, n_684);
  nand g1923 (n_1947, A[31], n_683);
  nand g1924 (n_1948, n_684, n_683);
  nand g1925 (n_1949, A[31], n_684);
  nand g1926 (n_703, n_1947, n_1948, n_1949);
  xor g1927 (n_1950, n_685, n_686);
  xor g1928 (n_692, n_1950, n_687);
  nand g1929 (n_1951, n_685, n_686);
  nand g1930 (n_1952, n_687, n_686);
  nand g1931 (n_1953, n_685, n_687);
  nand g1932 (n_705, n_1951, n_1952, n_1953);
  xor g1933 (n_1954, n_688, n_689);
  xor g1934 (n_694, n_1954, n_690);
  nand g1935 (n_1955, n_688, n_689);
  nand g1936 (n_1956, n_690, n_689);
  nand g1937 (n_1957, n_688, n_690);
  nand g1938 (n_707, n_1955, n_1956, n_1957);
  xor g1939 (n_1958, n_691, n_692);
  xor g1940 (n_695, n_1958, n_693);
  nand g1941 (n_1959, n_691, n_692);
  nand g1942 (n_1960, n_693, n_692);
  nand g1943 (n_1961, n_691, n_693);
  nand g1944 (n_710, n_1959, n_1960, n_1961);
  xor g1945 (n_1962, n_694, n_695);
  xor g1946 (n_148, n_1962, n_696);
  nand g1947 (n_1963, n_694, n_695);
  nand g1948 (n_1964, n_696, n_695);
  nand g1949 (n_1965, n_694, n_696);
  nand g1950 (n_77, n_1963, n_1964, n_1965);
  xor g1951 (n_1966, A[28], A[44]);
  xor g1952 (n_701, n_1966, A[42]);
  nand g1953 (n_1967, A[28], A[44]);
  nand g1954 (n_1968, A[42], A[44]);
  nand g1956 (n_711, n_1967, n_1968, n_1903);
  xor g1958 (n_702, n_1782, A[36]);
  nand g1960 (n_1972, A[36], A[38]);
  nand g1962 (n_712, n_1783, n_1972, n_1716);
  xor g1963 (n_1974, A[26], A[40]);
  xor g1964 (n_700, n_1974, A[34]);
  nand g1965 (n_1975, A[26], A[40]);
  nand g1966 (n_1976, A[34], A[40]);
  nand g1968 (n_713, n_1975, n_1976, n_1721);
  xor g1969 (n_1978, A[32], n_697);
  xor g1970 (n_704, n_1978, n_698);
  nand g1971 (n_1979, A[32], n_697);
  nand g1972 (n_1980, n_698, n_697);
  nand g1973 (n_1981, A[32], n_698);
  nand g1974 (n_717, n_1979, n_1980, n_1981);
  xor g1975 (n_1982, n_699, n_700);
  xor g1976 (n_706, n_1982, n_701);
  nand g1977 (n_1983, n_699, n_700);
  nand g1978 (n_1984, n_701, n_700);
  nand g1979 (n_1985, n_699, n_701);
  nand g1980 (n_719, n_1983, n_1984, n_1985);
  xor g1981 (n_1986, n_702, n_703);
  xor g1982 (n_708, n_1986, n_704);
  nand g1983 (n_1987, n_702, n_703);
  nand g1984 (n_1988, n_704, n_703);
  nand g1985 (n_1989, n_702, n_704);
  nand g1986 (n_721, n_1987, n_1988, n_1989);
  xor g1987 (n_1990, n_705, n_706);
  xor g1988 (n_709, n_1990, n_707);
  nand g1989 (n_1991, n_705, n_706);
  nand g1990 (n_1992, n_707, n_706);
  nand g1991 (n_1993, n_705, n_707);
  nand g1992 (n_724, n_1991, n_1992, n_1993);
  xor g1993 (n_1994, n_708, n_709);
  xor g1994 (n_147, n_1994, n_710);
  nand g1995 (n_1995, n_708, n_709);
  nand g1996 (n_1996, n_710, n_709);
  nand g1997 (n_1997, n_708, n_710);
  nand g1998 (n_76, n_1995, n_1996, n_1997);
  xor g1999 (n_1998, A[29], A[45]);
  xor g2000 (n_715, n_1998, A[43]);
  nand g2001 (n_1999, A[29], A[45]);
  nand g2002 (n_2000, A[43], A[45]);
  nand g2004 (n_725, n_1999, n_2000, n_1935);
  xor g2006 (n_716, n_1814, A[37]);
  nand g2008 (n_2004, A[37], A[39]);
  nand g2010 (n_726, n_1815, n_2004, n_1748);
  xor g2011 (n_2006, A[27], A[41]);
  xor g2012 (n_714, n_2006, A[35]);
  nand g2013 (n_2007, A[27], A[41]);
  nand g2014 (n_2008, A[35], A[41]);
  nand g2016 (n_727, n_2007, n_2008, n_1753);
  xor g2017 (n_2010, A[33], n_711);
  xor g2018 (n_718, n_2010, n_712);
  nand g2019 (n_2011, A[33], n_711);
  nand g2020 (n_2012, n_712, n_711);
  nand g2021 (n_2013, A[33], n_712);
  nand g2022 (n_731, n_2011, n_2012, n_2013);
  xor g2023 (n_2014, n_713, n_714);
  xor g2024 (n_720, n_2014, n_715);
  nand g2025 (n_2015, n_713, n_714);
  nand g2026 (n_2016, n_715, n_714);
  nand g2027 (n_2017, n_713, n_715);
  nand g2028 (n_733, n_2015, n_2016, n_2017);
  xor g2029 (n_2018, n_716, n_717);
  xor g2030 (n_722, n_2018, n_718);
  nand g2031 (n_2019, n_716, n_717);
  nand g2032 (n_2020, n_718, n_717);
  nand g2033 (n_2021, n_716, n_718);
  nand g2034 (n_735, n_2019, n_2020, n_2021);
  xor g2035 (n_2022, n_719, n_720);
  xor g2036 (n_723, n_2022, n_721);
  nand g2037 (n_2023, n_719, n_720);
  nand g2038 (n_2024, n_721, n_720);
  nand g2039 (n_2025, n_719, n_721);
  nand g2040 (n_738, n_2023, n_2024, n_2025);
  xor g2041 (n_2026, n_722, n_723);
  xor g2042 (n_146, n_2026, n_724);
  nand g2043 (n_2027, n_722, n_723);
  nand g2044 (n_2028, n_724, n_723);
  nand g2045 (n_2029, n_722, n_724);
  nand g2046 (n_75, n_2027, n_2028, n_2029);
  xor g2047 (n_2030, A[28], A[46]);
  xor g2048 (n_729, n_2030, A[40]);
  nand g2049 (n_2031, A[28], A[46]);
  nand g2050 (n_2032, A[40], A[46]);
  nand g2052 (n_739, n_2031, n_2032, n_1905);
  xor g2053 (n_2034, A[32], A[30]);
  xor g2054 (n_730, n_2034, A[44]);
  nand g2056 (n_2036, A[44], A[30]);
  nand g2057 (n_2037, A[32], A[44]);
  nand g2058 (n_740, n_1849, n_2036, n_2037);
  xor g2059 (n_2038, A[38], A[42]);
  xor g2060 (n_728, n_2038, A[36]);
  nand g2061 (n_2039, A[38], A[42]);
  nand g2062 (n_2040, A[36], A[42]);
  nand g2064 (n_741, n_2039, n_2040, n_1972);
  xor g2065 (n_2042, A[34], n_725);
  xor g2066 (n_732, n_2042, n_726);
  nand g2067 (n_2043, A[34], n_725);
  nand g2068 (n_2044, n_726, n_725);
  nand g2069 (n_2045, A[34], n_726);
  nand g2070 (n_745, n_2043, n_2044, n_2045);
  xor g2071 (n_2046, n_727, n_728);
  xor g2072 (n_734, n_2046, n_729);
  nand g2073 (n_2047, n_727, n_728);
  nand g2074 (n_2048, n_729, n_728);
  nand g2075 (n_2049, n_727, n_729);
  nand g2076 (n_747, n_2047, n_2048, n_2049);
  xor g2077 (n_2050, n_730, n_731);
  xor g2078 (n_736, n_2050, n_732);
  nand g2079 (n_2051, n_730, n_731);
  nand g2080 (n_2052, n_732, n_731);
  nand g2081 (n_2053, n_730, n_732);
  nand g2082 (n_749, n_2051, n_2052, n_2053);
  xor g2083 (n_2054, n_733, n_734);
  xor g2084 (n_737, n_2054, n_735);
  nand g2085 (n_2055, n_733, n_734);
  nand g2086 (n_2056, n_735, n_734);
  nand g2087 (n_2057, n_733, n_735);
  nand g2088 (n_752, n_2055, n_2056, n_2057);
  xor g2089 (n_2058, n_736, n_737);
  xor g2090 (n_145, n_2058, n_738);
  nand g2091 (n_2059, n_736, n_737);
  nand g2092 (n_2060, n_738, n_737);
  nand g2093 (n_2061, n_736, n_738);
  nand g2094 (n_74, n_2059, n_2060, n_2061);
  xor g2095 (n_2062, A[29], A[47]);
  xor g2096 (n_743, n_2062, A[41]);
  nand g2097 (n_2063, A[29], A[47]);
  nand g2098 (n_2064, A[41], A[47]);
  nand g2100 (n_753, n_2063, n_2064, n_1937);
  xor g2101 (n_2066, A[33], A[31]);
  xor g2102 (n_744, n_2066, A[45]);
  nand g2104 (n_2068, A[45], A[31]);
  nand g2105 (n_2069, A[33], A[45]);
  nand g2106 (n_754, n_1881, n_2068, n_2069);
  xor g2107 (n_2070, A[39], A[43]);
  xor g2108 (n_742, n_2070, A[37]);
  nand g2109 (n_2071, A[39], A[43]);
  nand g2110 (n_2072, A[37], A[43]);
  nand g2112 (n_755, n_2071, n_2072, n_2004);
  xor g2113 (n_2074, A[35], n_739);
  xor g2114 (n_746, n_2074, n_740);
  nand g2115 (n_2075, A[35], n_739);
  nand g2116 (n_2076, n_740, n_739);
  nand g2117 (n_2077, A[35], n_740);
  nand g2118 (n_759, n_2075, n_2076, n_2077);
  xor g2119 (n_2078, n_741, n_742);
  xor g2120 (n_748, n_2078, n_743);
  nand g2121 (n_2079, n_741, n_742);
  nand g2122 (n_2080, n_743, n_742);
  nand g2123 (n_2081, n_741, n_743);
  nand g2124 (n_761, n_2079, n_2080, n_2081);
  xor g2125 (n_2082, n_744, n_745);
  xor g2126 (n_750, n_2082, n_746);
  nand g2127 (n_2083, n_744, n_745);
  nand g2128 (n_2084, n_746, n_745);
  nand g2129 (n_2085, n_744, n_746);
  nand g2130 (n_763, n_2083, n_2084, n_2085);
  xor g2131 (n_2086, n_747, n_748);
  xor g2132 (n_751, n_2086, n_749);
  nand g2133 (n_2087, n_747, n_748);
  nand g2134 (n_2088, n_749, n_748);
  nand g2135 (n_2089, n_747, n_749);
  nand g2136 (n_766, n_2087, n_2088, n_2089);
  xor g2137 (n_2090, n_750, n_751);
  xor g2138 (n_144, n_2090, n_752);
  nand g2139 (n_2091, n_750, n_751);
  nand g2140 (n_2092, n_752, n_751);
  nand g2141 (n_2093, n_750, n_752);
  nand g2142 (n_73, n_2091, n_2092, n_2093);
  xor g2143 (n_2094, A[48], A[46]);
  xor g2144 (n_757, n_2094, A[42]);
  nand g2145 (n_2095, A[48], A[46]);
  nand g2146 (n_2096, A[42], A[46]);
  nand g2147 (n_2097, A[48], A[42]);
  nand g2148 (n_767, n_2095, n_2096, n_2097);
  xor g2150 (n_758, n_1718, A[40]);
  nand g2154 (n_768, n_1652, n_1847, n_1976);
  xor g2155 (n_2102, A[30], A[44]);
  xor g2156 (n_756, n_2102, A[38]);
  nand g2158 (n_2104, A[38], A[44]);
  nand g2160 (n_769, n_2036, n_2104, n_1783);
  xor g2161 (n_2106, A[36], n_753);
  xor g2162 (n_760, n_2106, n_754);
  nand g2163 (n_2107, A[36], n_753);
  nand g2164 (n_2108, n_754, n_753);
  nand g2165 (n_2109, A[36], n_754);
  nand g2166 (n_773, n_2107, n_2108, n_2109);
  xor g2167 (n_2110, n_755, n_756);
  xor g2168 (n_762, n_2110, n_757);
  nand g2169 (n_2111, n_755, n_756);
  nand g2170 (n_2112, n_757, n_756);
  nand g2171 (n_2113, n_755, n_757);
  nand g2172 (n_775, n_2111, n_2112, n_2113);
  xor g2173 (n_2114, n_758, n_759);
  xor g2174 (n_764, n_2114, n_760);
  nand g2175 (n_2115, n_758, n_759);
  nand g2176 (n_2116, n_760, n_759);
  nand g2177 (n_2117, n_758, n_760);
  nand g2178 (n_777, n_2115, n_2116, n_2117);
  xor g2179 (n_2118, n_761, n_762);
  xor g2180 (n_765, n_2118, n_763);
  nand g2181 (n_2119, n_761, n_762);
  nand g2182 (n_2120, n_763, n_762);
  nand g2183 (n_2121, n_761, n_763);
  nand g2184 (n_780, n_2119, n_2120, n_2121);
  xor g2185 (n_2122, n_764, n_765);
  xor g2186 (n_143, n_2122, n_766);
  nand g2187 (n_2123, n_764, n_765);
  nand g2188 (n_2124, n_766, n_765);
  nand g2189 (n_2125, n_764, n_766);
  nand g2190 (n_72, n_2123, n_2124, n_2125);
  xor g2191 (n_2126, A[49], A[47]);
  xor g2192 (n_771, n_2126, A[43]);
  nand g2193 (n_2127, A[49], A[47]);
  nand g2194 (n_2128, A[43], A[47]);
  nand g2195 (n_2129, A[49], A[43]);
  nand g2196 (n_784, n_2127, n_2128, n_2129);
  xor g2198 (n_772, n_1750, A[41]);
  nand g2202 (n_785, n_1684, n_1879, n_2008);
  xor g2203 (n_2134, A[31], A[45]);
  xor g2204 (n_770, n_2134, A[39]);
  nand g2206 (n_2136, A[39], A[45]);
  nand g2208 (n_783, n_2068, n_2136, n_1815);
  xor g2209 (n_2138, A[37], n_767);
  xor g2210 (n_774, n_2138, n_768);
  nand g2211 (n_2139, A[37], n_767);
  nand g2212 (n_2140, n_768, n_767);
  nand g2213 (n_2141, A[37], n_768);
  nand g2214 (n_789, n_2139, n_2140, n_2141);
  xor g2215 (n_2142, n_769, n_770);
  xor g2216 (n_776, n_2142, n_771);
  nand g2217 (n_2143, n_769, n_770);
  nand g2218 (n_2144, n_771, n_770);
  nand g2219 (n_2145, n_769, n_771);
  nand g2220 (n_791, n_2143, n_2144, n_2145);
  xor g2221 (n_2146, n_772, n_773);
  xor g2222 (n_778, n_2146, n_774);
  nand g2223 (n_2147, n_772, n_773);
  nand g2224 (n_2148, n_774, n_773);
  nand g2225 (n_2149, n_772, n_774);
  nand g2226 (n_793, n_2147, n_2148, n_2149);
  xor g2227 (n_2150, n_775, n_776);
  xor g2228 (n_779, n_2150, n_777);
  nand g2229 (n_2151, n_775, n_776);
  nand g2230 (n_2152, n_777, n_776);
  nand g2231 (n_2153, n_775, n_777);
  nand g2232 (n_796, n_2151, n_2152, n_2153);
  xor g2233 (n_2154, n_778, n_779);
  xor g2234 (n_142, n_2154, n_780);
  nand g2235 (n_2155, n_778, n_779);
  nand g2236 (n_2156, n_780, n_779);
  nand g2237 (n_2157, n_778, n_780);
  nand g2238 (n_71, n_2155, n_2156, n_2157);
  xor g2241 (n_2158, A[50], A[44]);
  xor g2242 (n_787, n_2158, A[36]);
  nand g2243 (n_2159, A[50], A[44]);
  nand g2244 (n_2160, A[36], A[44]);
  nand g2245 (n_2161, A[50], A[36]);
  nand g2246 (n_801, n_2159, n_2160, n_2161);
  xor g2247 (n_2162, A[34], A[48]);
  xor g2248 (n_788, n_2162, A[32]);
  nand g2249 (n_2163, A[34], A[48]);
  nand g2250 (n_2164, A[32], A[48]);
  nand g2252 (n_802, n_2163, n_2164, n_1652);
  xor g2253 (n_2166, A[42], A[46]);
  xor g2254 (n_786, n_2166, A[40]);
  nand g2258 (n_800, n_2096, n_2032, n_1904);
  xor g2259 (n_2170, A[38], n_783);
  xor g2260 (n_790, n_2170, n_784);
  nand g2261 (n_2171, A[38], n_783);
  nand g2262 (n_2172, n_784, n_783);
  nand g2263 (n_2173, A[38], n_784);
  nand g2264 (n_806, n_2171, n_2172, n_2173);
  xor g2265 (n_2174, n_785, n_786);
  xor g2266 (n_792, n_2174, n_787);
  nand g2267 (n_2175, n_785, n_786);
  nand g2268 (n_2176, n_787, n_786);
  nand g2269 (n_2177, n_785, n_787);
  nand g2270 (n_808, n_2175, n_2176, n_2177);
  xor g2271 (n_2178, n_788, n_789);
  xor g2272 (n_794, n_2178, n_790);
  nand g2273 (n_2179, n_788, n_789);
  nand g2274 (n_2180, n_790, n_789);
  nand g2275 (n_2181, n_788, n_790);
  nand g2276 (n_810, n_2179, n_2180, n_2181);
  xor g2277 (n_2182, n_791, n_792);
  xor g2278 (n_795, n_2182, n_793);
  nand g2279 (n_2183, n_791, n_792);
  nand g2280 (n_2184, n_793, n_792);
  nand g2281 (n_2185, n_791, n_793);
  nand g2282 (n_813, n_2183, n_2184, n_2185);
  xor g2283 (n_2186, n_794, n_795);
  xor g2284 (n_141, n_2186, n_796);
  nand g2285 (n_2187, n_794, n_795);
  nand g2286 (n_2188, n_796, n_795);
  nand g2287 (n_2189, n_794, n_796);
  nand g2288 (n_70, n_2187, n_2188, n_2189);
  xor g2291 (n_2190, A[43], A[35]);
  xor g2292 (n_804, n_2190, A[33]);
  nand g2293 (n_2191, A[43], A[35]);
  nand g2295 (n_2193, A[43], A[33]);
  nand g2296 (n_815, n_2191, n_1684, n_2193);
  xor g2297 (n_2194, A[50], A[49]);
  xor g2298 (n_805, n_2194, A[41]);
  nand g2299 (n_2195, A[50], A[49]);
  nand g2300 (n_2196, A[41], A[49]);
  nand g2301 (n_2197, A[50], A[41]);
  nand g2302 (n_816, n_2195, n_2196, n_2197);
  xor g2303 (n_2198, A[47], A[45]);
  xor g2304 (n_803, n_2198, A[39]);
  nand g2305 (n_2199, A[47], A[45]);
  nand g2307 (n_2201, A[47], A[39]);
  nand g2308 (n_817, n_2199, n_2136, n_2201);
  xor g2309 (n_2202, A[37], n_800);
  xor g2310 (n_807, n_2202, n_801);
  nand g2311 (n_2203, A[37], n_800);
  nand g2312 (n_2204, n_801, n_800);
  nand g2313 (n_2205, A[37], n_801);
  nand g2314 (n_821, n_2203, n_2204, n_2205);
  xor g2315 (n_2206, n_802, n_803);
  xor g2316 (n_809, n_2206, n_804);
  nand g2317 (n_2207, n_802, n_803);
  nand g2318 (n_2208, n_804, n_803);
  nand g2319 (n_2209, n_802, n_804);
  nand g2320 (n_823, n_2207, n_2208, n_2209);
  xor g2321 (n_2210, n_805, n_806);
  xor g2322 (n_811, n_2210, n_807);
  nand g2323 (n_2211, n_805, n_806);
  nand g2324 (n_2212, n_807, n_806);
  nand g2325 (n_2213, n_805, n_807);
  nand g2326 (n_825, n_2211, n_2212, n_2213);
  xor g2327 (n_2214, n_808, n_809);
  xor g2328 (n_812, n_2214, n_810);
  nand g2329 (n_2215, n_808, n_809);
  nand g2330 (n_2216, n_810, n_809);
  nand g2331 (n_2217, n_808, n_810);
  nand g2332 (n_828, n_2215, n_2216, n_2217);
  xor g2333 (n_2218, n_811, n_812);
  xor g2334 (n_140, n_2218, n_813);
  nand g2335 (n_2219, n_811, n_812);
  nand g2336 (n_2220, n_813, n_812);
  nand g2337 (n_2221, n_811, n_813);
  nand g2338 (n_69, n_2219, n_2220, n_2221);
  xor g2340 (n_819, n_2222, A[44]);
  nand g2342 (n_2224, A[44], A[48]);
  nand g2344 (n_831, n_2223, n_2224, n_2225);
  xor g2345 (n_2226, A[36], A[34]);
  xor g2346 (n_820, n_2226, A[42]);
  nand g2348 (n_2228, A[42], A[34]);
  nand g2350 (n_832, n_1909, n_2228, n_2040);
  xor g2352 (n_818, n_2230, A[40]);
  nand g2356 (n_833, n_2231, n_2032, n_2233);
  xor g2357 (n_2234, A[38], n_815);
  xor g2358 (n_822, n_2234, n_816);
  nand g2359 (n_2235, A[38], n_815);
  nand g2360 (n_2236, n_816, n_815);
  nand g2361 (n_2237, A[38], n_816);
  nand g2362 (n_837, n_2235, n_2236, n_2237);
  xor g2363 (n_2238, n_817, n_818);
  xor g2364 (n_824, n_2238, n_819);
  nand g2365 (n_2239, n_817, n_818);
  nand g2366 (n_2240, n_819, n_818);
  nand g2367 (n_2241, n_817, n_819);
  nand g2368 (n_839, n_2239, n_2240, n_2241);
  xor g2369 (n_2242, n_820, n_821);
  xor g2370 (n_826, n_2242, n_822);
  nand g2371 (n_2243, n_820, n_821);
  nand g2372 (n_2244, n_822, n_821);
  nand g2373 (n_2245, n_820, n_822);
  nand g2374 (n_841, n_2243, n_2244, n_2245);
  xor g2375 (n_2246, n_823, n_824);
  xor g2376 (n_827, n_2246, n_825);
  nand g2377 (n_2247, n_823, n_824);
  nand g2378 (n_2248, n_825, n_824);
  nand g2379 (n_2249, n_823, n_825);
  nand g2380 (n_843, n_2247, n_2248, n_2249);
  xor g2381 (n_2250, n_826, n_827);
  xor g2382 (n_139, n_2250, n_828);
  nand g2383 (n_2251, n_826, n_827);
  nand g2384 (n_2252, n_828, n_827);
  nand g2385 (n_2253, n_826, n_828);
  nand g2386 (n_68, n_2251, n_2252, n_2253);
  xor g2389 (n_2254, A[47], A[35]);
  xor g2390 (n_835, n_2254, A[43]);
  nand g2391 (n_2255, A[47], A[35]);
  nand g2394 (n_846, n_2255, n_2191, n_2128);
  xor g2395 (n_2258, A[41], A[45]);
  xor g2396 (n_834, n_2258, A[39]);
  nand g2397 (n_2259, A[41], A[45]);
  nand g2399 (n_2261, A[41], A[39]);
  nand g2400 (n_845, n_2259, n_2136, n_2261);
  xor g2402 (n_836, n_2262, n_831);
  nand g2405 (n_2265, A[37], n_831);
  nand g2406 (n_850, n_2263, n_2264, n_2265);
  xor g2407 (n_2266, n_832, n_833);
  xor g2408 (n_838, n_2266, n_834);
  nand g2409 (n_2267, n_832, n_833);
  nand g2410 (n_2268, n_834, n_833);
  nand g2411 (n_2269, n_832, n_834);
  nand g2412 (n_852, n_2267, n_2268, n_2269);
  xor g2413 (n_2270, n_835, n_836);
  xor g2414 (n_840, n_2270, n_837);
  nand g2415 (n_2271, n_835, n_836);
  nand g2416 (n_2272, n_837, n_836);
  nand g2417 (n_2273, n_835, n_837);
  nand g2418 (n_853, n_2271, n_2272, n_2273);
  xor g2419 (n_2274, n_838, n_839);
  xor g2420 (n_842, n_2274, n_840);
  nand g2421 (n_2275, n_838, n_839);
  nand g2422 (n_2276, n_840, n_839);
  nand g2423 (n_2277, n_838, n_840);
  nand g2424 (n_856, n_2275, n_2276, n_2277);
  xor g2425 (n_2278, n_841, n_842);
  xor g2426 (n_138, n_2278, n_843);
  nand g2427 (n_2279, n_841, n_842);
  nand g2428 (n_2280, n_843, n_842);
  nand g2429 (n_2281, n_841, n_843);
  nand g2430 (n_67, n_2279, n_2280, n_2281);
  xor g2437 (n_2286, A[36], A[42]);
  xor g2438 (n_848, n_2286, A[46]);
  nand g2441 (n_2289, A[36], A[46]);
  nand g2442 (n_860, n_2040, n_2096, n_2289);
  xor g2443 (n_2290, A[40], A[38]);
  xor g2444 (n_849, n_2290, A[49]);
  nand g2445 (n_2291, A[40], A[38]);
  nand g2446 (n_2292, A[49], A[38]);
  nand g2447 (n_2293, A[40], A[49]);
  nand g2448 (n_863, n_2291, n_2292, n_2293);
  xor g2449 (n_2294, n_845, n_846);
  xor g2450 (n_851, n_2294, n_819);
  nand g2451 (n_2295, n_845, n_846);
  nand g2452 (n_2296, n_819, n_846);
  nand g2453 (n_2297, n_845, n_819);
  nand g2454 (n_865, n_2295, n_2296, n_2297);
  xor g2455 (n_2298, n_848, n_849);
  xor g2456 (n_854, n_2298, n_850);
  nand g2457 (n_2299, n_848, n_849);
  nand g2458 (n_2300, n_850, n_849);
  nand g2459 (n_2301, n_848, n_850);
  nand g2460 (n_867, n_2299, n_2300, n_2301);
  xor g2461 (n_2302, n_851, n_852);
  xor g2462 (n_855, n_2302, n_853);
  nand g2463 (n_2303, n_851, n_852);
  nand g2464 (n_2304, n_853, n_852);
  nand g2465 (n_2305, n_851, n_853);
  nand g2466 (n_869, n_2303, n_2304, n_2305);
  xor g2467 (n_2306, n_854, n_855);
  xor g2468 (n_137, n_2306, n_856);
  nand g2469 (n_2307, n_854, n_855);
  nand g2470 (n_2308, n_856, n_855);
  nand g2471 (n_2309, n_854, n_856);
  nand g2472 (n_136, n_2307, n_2308, n_2309);
  xor g2475 (n_2310, A[47], A[43]);
  xor g2476 (n_862, n_2310, A[41]);
  nand g2480 (n_871, n_2128, n_1936, n_2064);
  xor g2481 (n_2314, A[45], A[39]);
  xor g2482 (n_861, n_2314, A[37]);
  nand g2485 (n_2317, A[45], A[37]);
  nand g2486 (n_872, n_2136, n_2004, n_2317);
  xor g2488 (n_864, n_2318, n_860);
  nand g2490 (n_2320, n_860, n_831);
  nand g2492 (n_876, n_2264, n_2320, n_2321);
  xor g2493 (n_2322, n_861, n_862);
  xor g2494 (n_866, n_2322, n_863);
  nand g2495 (n_2323, n_861, n_862);
  nand g2496 (n_2324, n_863, n_862);
  nand g2497 (n_2325, n_861, n_863);
  nand g2498 (n_877, n_2323, n_2324, n_2325);
  xor g2499 (n_2326, n_864, n_865);
  xor g2500 (n_868, n_2326, n_866);
  nand g2501 (n_2327, n_864, n_865);
  nand g2502 (n_2328, n_866, n_865);
  nand g2503 (n_2329, n_864, n_866);
  nand g2504 (n_880, n_2327, n_2328, n_2329);
  xor g2505 (n_2330, n_867, n_868);
  xor g2506 (n_66, n_2330, n_869);
  nand g2507 (n_2331, n_867, n_868);
  nand g2508 (n_2332, n_869, n_868);
  nand g2509 (n_2333, n_867, n_869);
  nand g2510 (n_65, n_2331, n_2332, n_2333);
  xor g2523 (n_2342, A[38], A[49]);
  xor g2524 (n_875, n_2342, n_871);
  nand g2526 (n_2344, n_871, A[49]);
  nand g2527 (n_2345, A[38], n_871);
  nand g2528 (n_887, n_2292, n_2344, n_2345);
  xor g2529 (n_2346, n_872, n_786);
  xor g2530 (n_878, n_2346, n_819);
  nand g2531 (n_2347, n_872, n_786);
  nand g2532 (n_2348, n_819, n_786);
  nand g2533 (n_2349, n_872, n_819);
  nand g2534 (n_888, n_2347, n_2348, n_2349);
  xor g2535 (n_2350, n_875, n_876);
  xor g2536 (n_879, n_2350, n_877);
  nand g2537 (n_2351, n_875, n_876);
  nand g2538 (n_2352, n_877, n_876);
  nand g2539 (n_2353, n_875, n_877);
  nand g2540 (n_891, n_2351, n_2352, n_2353);
  xor g2541 (n_2354, n_878, n_879);
  xor g2542 (n_135, n_2354, n_880);
  nand g2543 (n_2355, n_878, n_879);
  nand g2544 (n_2356, n_880, n_879);
  nand g2545 (n_2357, n_878, n_880);
  nand g2546 (n_64, n_2355, n_2356, n_2357);
  xor g2549 (n_2358, A[43], A[41]);
  xor g2550 (n_885, n_2358, A[49]);
  nand g2554 (n_893, n_1936, n_2196, n_2129);
  nand g2560 (n_896, n_2136, n_2364, n_2365);
  xor g2561 (n_2366, n_800, n_831);
  xor g2562 (n_889, n_2366, n_885);
  nand g2563 (n_2367, n_800, n_831);
  nand g2564 (n_2368, n_885, n_831);
  nand g2565 (n_2369, n_800, n_885);
  nand g2566 (n_898, n_2367, n_2368, n_2369);
  xor g2567 (n_2370, n_886, n_887);
  xor g2568 (n_890, n_2370, n_888);
  nand g2569 (n_2371, n_886, n_887);
  nand g2570 (n_2372, n_888, n_887);
  nand g2571 (n_2373, n_886, n_888);
  nand g2572 (n_900, n_2371, n_2372, n_2373);
  xor g2573 (n_2374, n_889, n_890);
  xor g2574 (n_134, n_2374, n_891);
  nand g2575 (n_2375, n_889, n_890);
  nand g2576 (n_2376, n_891, n_890);
  nand g2577 (n_2377, n_889, n_891);
  nand g2578 (n_63, n_2375, n_2376, n_2377);
  xor g2591 (n_2386, A[47], n_893);
  xor g2592 (n_897, n_2386, n_786);
  nand g2593 (n_2387, A[47], n_893);
  nand g2594 (n_2388, n_786, n_893);
  nand g2595 (n_2389, A[47], n_786);
  nand g2596 (n_907, n_2387, n_2388, n_2389);
  xor g2597 (n_2390, n_819, n_896);
  xor g2598 (n_899, n_2390, n_897);
  nand g2599 (n_2391, n_819, n_896);
  nand g2600 (n_2392, n_897, n_896);
  nand g2601 (n_2393, n_819, n_897);
  nand g2602 (n_909, n_2391, n_2392, n_2393);
  xor g2603 (n_2394, n_898, n_899);
  xor g2604 (n_133, n_2394, n_900);
  nand g2605 (n_2395, n_898, n_899);
  nand g2606 (n_2396, n_900, n_899);
  nand g2607 (n_2397, n_898, n_900);
  nand g2608 (n_62, n_2395, n_2396, n_2397);
  nand g2621 (n_2405, A[45], n_800);
  nand g2622 (n_914, n_2364, n_2404, n_2405);
  xor g2623 (n_2406, n_831, n_885);
  xor g2624 (n_908, n_2406, n_906);
  nand g2626 (n_2408, n_906, n_885);
  nand g2627 (n_2409, n_831, n_906);
  nand g2628 (n_916, n_2368, n_2408, n_2409);
  xor g2629 (n_2410, n_907, n_908);
  xor g2630 (n_132, n_2410, n_909);
  nand g2631 (n_2411, n_907, n_908);
  nand g2632 (n_2412, n_909, n_908);
  nand g2633 (n_2413, n_907, n_909);
  nand g2634 (n_131, n_2411, n_2412, n_2413);
  xor g2642 (n_913, n_2166, A[47]);
  nand g2644 (n_2420, A[47], A[46]);
  nand g2645 (n_2421, A[42], A[47]);
  nand g2646 (n_921, n_2096, n_2420, n_2421);
  xor g2647 (n_2422, n_893, n_819);
  xor g2648 (n_915, n_2422, n_913);
  nand g2649 (n_2423, n_893, n_819);
  nand g2650 (n_2424, n_913, n_819);
  nand g2651 (n_2425, n_893, n_913);
  nand g2652 (n_923, n_2423, n_2424, n_2425);
  xor g2653 (n_2426, n_914, n_915);
  xor g2654 (n_61, n_2426, n_916);
  nand g2655 (n_2427, n_914, n_915);
  nand g2656 (n_2428, n_916, n_915);
  nand g2657 (n_2429, n_914, n_916);
  nand g2658 (n_130, n_2427, n_2428, n_2429);
  xor g2662 (n_920, n_2310, A[45]);
  nand g2666 (n_925, n_2128, n_2199, n_2000);
  xor g2668 (n_922, n_2318, n_920);
  nand g2670 (n_2436, n_920, n_831);
  nand g2672 (n_928, n_2264, n_2436, n_2437);
  xor g2673 (n_2438, n_921, n_922);
  xor g2674 (n_60, n_2438, n_923);
  nand g2675 (n_2439, n_921, n_922);
  nand g2676 (n_2440, n_923, n_922);
  nand g2677 (n_2441, n_921, n_923);
  nand g2678 (n_129, n_2439, n_2440, n_2441);
  xor g2685 (n_2446, A[46], A[49]);
  xor g2686 (n_927, n_2446, n_925);
  nand g2687 (n_2447, A[46], A[49]);
  nand g2688 (n_2448, n_925, A[49]);
  nand g2689 (n_2449, A[46], n_925);
  nand g2690 (n_933, n_2447, n_2448, n_2449);
  xor g2691 (n_2450, n_819, n_927);
  xor g2692 (n_59, n_2450, n_928);
  nand g2693 (n_2451, n_819, n_927);
  nand g2694 (n_2452, n_928, n_927);
  nand g2695 (n_2453, n_819, n_928);
  nand g2696 (n_128, n_2451, n_2452, n_2453);
  nand g2704 (n_936, n_2199, n_2456, n_2457);
  xor g2705 (n_2458, n_831, n_932);
  xor g2706 (n_58, n_2458, n_933);
  nand g2707 (n_2459, n_831, n_932);
  nand g2708 (n_2460, n_933, n_932);
  nand g2709 (n_2461, n_831, n_933);
  nand g2710 (n_127, n_2459, n_2460, n_2461);
  xor g2712 (n_935, n_2222, A[46]);
  nand g2716 (n_939, n_2223, n_2095, n_2231);
  xor g2717 (n_2466, A[49], n_935);
  xor g2718 (n_57, n_2466, n_936);
  nand g2719 (n_2467, A[49], n_935);
  nand g2720 (n_2468, n_936, n_935);
  nand g2721 (n_2469, A[49], n_936);
  nand g2722 (n_126, n_2467, n_2468, n_2469);
  nand g2729 (n_2473, A[49], n_939);
  nand g2730 (n_125, n_2471, n_2472, n_2473);
  xor g2732 (n_55, n_2222, A[47]);
  nand g2734 (n_2476, A[47], A[48]);
  nand g2736 (n_124, n_2223, n_2476, n_2477);
  nor g11 (n_2493, A[2], A[0]);
  nor g13 (n_2489, A[3], A[1]);
  nor g15 (n_2499, A[2], n_187);
  nand g16 (n_2494, A[2], n_187);
  nor g17 (n_2495, n_116, n_186);
  nand g18 (n_2496, n_116, n_186);
  nor g19 (n_2505, n_115, n_185);
  nand g20 (n_2500, n_115, n_185);
  nor g21 (n_2501, n_114, n_184);
  nand g22 (n_2502, n_114, n_184);
  nor g23 (n_2511, n_113, n_183);
  nand g24 (n_2506, n_113, n_183);
  nor g25 (n_2507, n_112, n_182);
  nand g26 (n_2508, n_112, n_182);
  nor g27 (n_2517, n_111, n_181);
  nand g28 (n_2512, n_111, n_181);
  nor g29 (n_2513, n_110, n_180);
  nand g30 (n_2514, n_110, n_180);
  nor g31 (n_2523, n_109, n_179);
  nand g32 (n_2518, n_109, n_179);
  nor g33 (n_2519, n_108, n_178);
  nand g34 (n_2520, n_108, n_178);
  nor g35 (n_2529, n_107, n_177);
  nand g36 (n_2524, n_107, n_177);
  nor g37 (n_2525, n_106, n_176);
  nand g38 (n_2526, n_106, n_176);
  nor g39 (n_2535, n_105, n_175);
  nand g40 (n_2530, n_105, n_175);
  nor g41 (n_2531, n_104, n_174);
  nand g42 (n_2532, n_104, n_174);
  nor g43 (n_2541, n_103, n_173);
  nand g44 (n_2536, n_103, n_173);
  nor g45 (n_2537, n_102, n_172);
  nand g46 (n_2538, n_102, n_172);
  nor g47 (n_2547, n_101, n_171);
  nand g48 (n_2542, n_101, n_171);
  nor g49 (n_2543, n_100, n_170);
  nand g50 (n_2544, n_100, n_170);
  nor g51 (n_2553, n_99, n_169);
  nand g52 (n_2548, n_99, n_169);
  nor g53 (n_2549, n_98, n_168);
  nand g54 (n_2550, n_98, n_168);
  nor g55 (n_2559, n_97, n_167);
  nand g56 (n_2554, n_97, n_167);
  nor g57 (n_2555, n_96, n_166);
  nand g58 (n_2556, n_96, n_166);
  nor g59 (n_2565, n_95, n_165);
  nand g60 (n_2560, n_95, n_165);
  nor g61 (n_2561, n_94, n_164);
  nand g62 (n_2562, n_94, n_164);
  nor g63 (n_2571, n_93, n_163);
  nand g64 (n_2566, n_93, n_163);
  nor g65 (n_2567, n_92, n_162);
  nand g66 (n_2568, n_92, n_162);
  nor g67 (n_2577, n_91, n_161);
  nand g68 (n_2572, n_91, n_161);
  nor g69 (n_2573, n_90, n_160);
  nand g70 (n_2574, n_90, n_160);
  nor g71 (n_2583, n_89, n_159);
  nand g72 (n_2578, n_89, n_159);
  nor g73 (n_2579, n_88, n_158);
  nand g74 (n_2580, n_88, n_158);
  nor g75 (n_2589, n_87, n_157);
  nand g76 (n_2584, n_87, n_157);
  nor g77 (n_2585, n_86, n_156);
  nand g78 (n_2586, n_86, n_156);
  nor g79 (n_2595, n_85, n_155);
  nand g80 (n_2590, n_85, n_155);
  nor g81 (n_2591, n_84, n_154);
  nand g82 (n_2592, n_84, n_154);
  nor g83 (n_2601, n_83, n_153);
  nand g84 (n_2596, n_83, n_153);
  nor g85 (n_2597, n_82, n_152);
  nand g86 (n_2598, n_82, n_152);
  nor g87 (n_2607, n_81, n_151);
  nand g88 (n_2602, n_81, n_151);
  nor g89 (n_2603, n_80, n_150);
  nand g90 (n_2604, n_80, n_150);
  nor g91 (n_2613, n_79, n_149);
  nand g92 (n_2608, n_79, n_149);
  nor g93 (n_2609, n_78, n_148);
  nand g94 (n_2610, n_78, n_148);
  nor g95 (n_2619, n_77, n_147);
  nand g96 (n_2614, n_77, n_147);
  nor g97 (n_2615, n_76, n_146);
  nand g98 (n_2616, n_76, n_146);
  nor g99 (n_2625, n_75, n_145);
  nand g100 (n_2620, n_75, n_145);
  nor g101 (n_2621, n_74, n_144);
  nand g102 (n_2622, n_74, n_144);
  nor g103 (n_2631, n_73, n_143);
  nand g104 (n_2626, n_73, n_143);
  nor g105 (n_2627, n_72, n_142);
  nand g106 (n_2628, n_72, n_142);
  nor g107 (n_2637, n_71, n_141);
  nand g108 (n_2632, n_71, n_141);
  nor g109 (n_2633, n_70, n_140);
  nand g110 (n_2634, n_70, n_140);
  nor g111 (n_2643, n_69, n_139);
  nand g112 (n_2638, n_69, n_139);
  nor g113 (n_2639, n_68, n_138);
  nand g114 (n_2640, n_68, n_138);
  nor g115 (n_2649, n_67, n_137);
  nand g116 (n_2644, n_67, n_137);
  nor g117 (n_2645, n_66, n_136);
  nand g118 (n_2646, n_66, n_136);
  nor g119 (n_2655, n_65, n_135);
  nand g120 (n_2650, n_65, n_135);
  nor g121 (n_2651, n_64, n_134);
  nand g122 (n_2652, n_64, n_134);
  nor g123 (n_2661, n_63, n_133);
  nand g124 (n_2656, n_63, n_133);
  nor g125 (n_2657, n_62, n_132);
  nand g126 (n_2658, n_62, n_132);
  nor g127 (n_2667, n_61, n_131);
  nand g128 (n_2662, n_61, n_131);
  nor g129 (n_2663, n_60, n_130);
  nand g130 (n_2664, n_60, n_130);
  nor g131 (n_2673, n_59, n_129);
  nand g132 (n_2668, n_59, n_129);
  nor g133 (n_2669, n_58, n_128);
  nand g134 (n_2670, n_58, n_128);
  nor g135 (n_2679, n_57, n_127);
  nand g136 (n_2674, n_57, n_127);
  nor g137 (n_2675, n_56, n_126);
  nand g138 (n_2676, n_56, n_126);
  nor g139 (n_2685, n_55, n_125);
  nand g140 (n_2680, n_55, n_125);
  nor g150 (n_2491, n_947, n_2489);
  nor g154 (n_2497, n_2494, n_2495);
  nor g157 (n_2700, n_2499, n_2495);
  nor g158 (n_2503, n_2500, n_2501);
  nor g161 (n_2694, n_2505, n_2501);
  nor g162 (n_2509, n_2506, n_2507);
  nor g165 (n_2707, n_2511, n_2507);
  nor g166 (n_2515, n_2512, n_2513);
  nor g169 (n_2701, n_2517, n_2513);
  nor g170 (n_2521, n_2518, n_2519);
  nor g173 (n_2714, n_2523, n_2519);
  nor g174 (n_2527, n_2524, n_2525);
  nor g177 (n_2708, n_2529, n_2525);
  nor g178 (n_2533, n_2530, n_2531);
  nor g181 (n_2721, n_2535, n_2531);
  nor g182 (n_2539, n_2536, n_2537);
  nor g185 (n_2715, n_2541, n_2537);
  nor g186 (n_2545, n_2542, n_2543);
  nor g189 (n_2728, n_2547, n_2543);
  nor g190 (n_2551, n_2548, n_2549);
  nor g193 (n_2722, n_2553, n_2549);
  nor g194 (n_2557, n_2554, n_2555);
  nor g197 (n_2735, n_2559, n_2555);
  nor g198 (n_2563, n_2560, n_2561);
  nor g201 (n_2729, n_2565, n_2561);
  nor g202 (n_2569, n_2566, n_2567);
  nor g205 (n_2742, n_2571, n_2567);
  nor g206 (n_2575, n_2572, n_2573);
  nor g209 (n_2736, n_2577, n_2573);
  nor g210 (n_2581, n_2578, n_2579);
  nor g213 (n_2749, n_2583, n_2579);
  nor g214 (n_2587, n_2584, n_2585);
  nor g217 (n_2743, n_2589, n_2585);
  nor g218 (n_2593, n_2590, n_2591);
  nor g221 (n_2756, n_2595, n_2591);
  nor g222 (n_2599, n_2596, n_2597);
  nor g225 (n_2750, n_2601, n_2597);
  nor g226 (n_2605, n_2602, n_2603);
  nor g229 (n_2763, n_2607, n_2603);
  nor g230 (n_2611, n_2608, n_2609);
  nor g233 (n_2757, n_2613, n_2609);
  nor g234 (n_2617, n_2614, n_2615);
  nor g237 (n_2770, n_2619, n_2615);
  nor g238 (n_2623, n_2620, n_2621);
  nor g241 (n_2764, n_2625, n_2621);
  nor g242 (n_2629, n_2626, n_2627);
  nor g245 (n_2777, n_2631, n_2627);
  nor g246 (n_2635, n_2632, n_2633);
  nor g249 (n_2771, n_2637, n_2633);
  nor g250 (n_2641, n_2638, n_2639);
  nor g253 (n_2784, n_2643, n_2639);
  nor g254 (n_2647, n_2644, n_2645);
  nor g257 (n_2778, n_2649, n_2645);
  nor g258 (n_2653, n_2650, n_2651);
  nor g261 (n_2791, n_2655, n_2651);
  nor g262 (n_2659, n_2656, n_2657);
  nor g265 (n_2785, n_2661, n_2657);
  nor g266 (n_2665, n_2662, n_2663);
  nor g269 (n_2798, n_2667, n_2663);
  nor g270 (n_2671, n_2668, n_2669);
  nor g273 (n_2792, n_2673, n_2669);
  nor g274 (n_2677, n_2674, n_2675);
  nor g277 (n_2805, n_2679, n_2675);
  nor g278 (n_2683, n_2680, n_2681);
  nor g281 (n_2799, n_2685, n_2681);
  nand g292 (n_2806, n_2700, n_2694);
  nand g297 (n_2816, n_2707, n_2701);
  nand g302 (n_2811, n_2714, n_2708);
  nand g307 (n_2822, n_2721, n_2715);
  nand g312 (n_2817, n_2728, n_2722);
  nand g317 (n_2828, n_2735, n_2729);
  nand g322 (n_2823, n_2742, n_2736);
  nand g327 (n_2834, n_2749, n_2743);
  nand g332 (n_2829, n_2756, n_2750);
  nand g337 (n_2840, n_2763, n_2757);
  nand g342 (n_2835, n_2770, n_2764);
  nand g347 (n_2846, n_2777, n_2771);
  nand g352 (n_2841, n_2784, n_2778);
  nand g357 (n_2852, n_2791, n_2785);
  nand g362 (n_2847, n_2798, n_2792);
  nand g367 (n_2916, n_2805, n_2799);
  nand g370 (n_2854, n_2809, n_2810);
  nor g371 (n_2814, n_2811, n_2812);
  nor g374 (n_2853, n_2816, n_2811);
  nor g375 (n_2820, n_2817, n_2818);
  nor g378 (n_2863, n_2822, n_2817);
  nor g379 (n_2826, n_2823, n_2824);
  nor g382 (n_2857, n_2828, n_2823);
  nor g383 (n_2832, n_2829, n_2830);
  nor g386 (n_2870, n_2834, n_2829);
  nor g387 (n_2838, n_2835, n_2836);
  nor g390 (n_2864, n_2840, n_2835);
  nor g391 (n_2844, n_2841, n_2842);
  nor g394 (n_2877, n_2846, n_2841);
  nor g395 (n_2850, n_2847, n_2848);
  nor g398 (n_2871, n_2852, n_2847);
  nand g399 (n_2856, n_2853, n_2854);
  nand g400 (n_2879, n_2855, n_2856);
  nand g2745 (n_2878, n_2863, n_2857);
  nand g2750 (n_2888, n_2870, n_2864);
  nand g2755 (n_2883, n_2877, n_2871);
  nand g2758 (n_2890, n_2881, n_2882);
  nor g2759 (n_2886, n_2883, n_2884);
  nor g2762 (n_2889, n_2888, n_2883);
  nand g2763 (n_2892, n_2889, n_2890);
  nand g2764 (n_2917, n_2891, n_2892);
  nand g2767 (n_2897, n_2884, n_2894);
  nand g2768 (n_2895, n_2863, n_2879);
  nand g2769 (n_2903, n_2858, n_2895);
  nand g2770 (n_2896, n_2870, n_2890);
  nand g2771 (n_2908, n_2865, n_2896);
  nand g2772 (n_2898, n_2877, n_2897);
  nand g2773 (n_2913, n_2872, n_2898);
  nand g2776 (n_2923, n_2812, n_2900);
  nand g2779 (n_2926, n_2818, n_2902);
  nand g2782 (n_2929, n_2824, n_2905);
  nand g2785 (n_2932, n_2830, n_2907);
  nand g2788 (n_2935, n_2836, n_2910);
  nand g2791 (n_2938, n_2842, n_2912);
  nand g2794 (n_2941, n_2848, n_2915);
  nand g2797 (n_2944, n_2919, n_2920);
  nand g2799 (n_2949, n_2695, n_2921);
  nand g2800 (n_2922, n_2707, n_2854);
  nand g2801 (n_2954, n_2702, n_2922);
  nand g2802 (n_2924, n_2714, n_2923);
  nand g2803 (n_2959, n_2709, n_2924);
  nand g2804 (n_2925, n_2721, n_2879);
  nand g2805 (n_2964, n_2716, n_2925);
  nand g2806 (n_2927, n_2728, n_2926);
  nand g2807 (n_2969, n_2723, n_2927);
  nand g2808 (n_2928, n_2735, n_2903);
  nand g2809 (n_2974, n_2730, n_2928);
  nand g2810 (n_2930, n_2742, n_2929);
  nand g2811 (n_2979, n_2737, n_2930);
  nand g2812 (n_2931, n_2749, n_2890);
  nand g2813 (n_2984, n_2744, n_2931);
  nand g2814 (n_2933, n_2756, n_2932);
  nand g2815 (n_2989, n_2751, n_2933);
  nand g2816 (n_2934, n_2763, n_2908);
  nand g2817 (n_2994, n_2758, n_2934);
  nand g2818 (n_2936, n_2770, n_2935);
  nand g2819 (n_2999, n_2765, n_2936);
  nand g2820 (n_2937, n_2777, n_2897);
  nand g2821 (n_3004, n_2772, n_2937);
  nand g2822 (n_2939, n_2784, n_2938);
  nand g2823 (n_3009, n_2779, n_2939);
  nand g2824 (n_2940, n_2791, n_2913);
  nand g2825 (n_3014, n_2786, n_2940);
  nand g2826 (n_2942, n_2798, n_2941);
  nand g2827 (n_3019, n_2793, n_2942);
  nand g2828 (n_2943, n_2805, n_2917);
  nand g2829 (n_3024, n_2800, n_2943);
  nand g2835 (n_3036, n_2494, n_2948);
  nand g2838 (n_3040, n_2500, n_2951);
  nand g2841 (n_3044, n_2506, n_2953);
  nand g2844 (n_3048, n_2512, n_2956);
  nand g2847 (n_3052, n_2518, n_2958);
  nand g2850 (n_3056, n_2524, n_2961);
  nand g2853 (n_3060, n_2530, n_2963);
  nand g2856 (n_3064, n_2536, n_2966);
  nand g2859 (n_3068, n_2542, n_2968);
  nand g2862 (n_3072, n_2548, n_2971);
  nand g2865 (n_3076, n_2554, n_2973);
  nand g2868 (n_3080, n_2560, n_2976);
  nand g2871 (n_3084, n_2566, n_2978);
  nand g2874 (n_3088, n_2572, n_2981);
  nand g2877 (n_3092, n_2578, n_2983);
  nand g2880 (n_3096, n_2584, n_2986);
  nand g2883 (n_3100, n_2590, n_2988);
  nand g2886 (n_3104, n_2596, n_2991);
  nand g2889 (n_3108, n_2602, n_2993);
  nand g2892 (n_3112, n_2608, n_2996);
  nand g2895 (n_3116, n_2614, n_2998);
  nand g2898 (n_3120, n_2620, n_3001);
  nand g2901 (n_3124, n_2626, n_3003);
  nand g2904 (n_3128, n_2632, n_3006);
  nand g2907 (n_3132, n_2638, n_3008);
  nand g2910 (n_3136, n_2644, n_3011);
  nand g2913 (n_3140, n_2650, n_3013);
  nand g2916 (n_3144, n_2656, n_3016);
  nand g2919 (n_3148, n_2662, n_3018);
  nand g2922 (n_3152, n_2668, n_3021);
  nand g2925 (n_3156, n_2674, n_3023);
  nand g2928 (n_3160, n_2680, n_3026);
  nand g2931 (n_3164, n_2686, n_3028);
  xnor g2943 (Z[5], n_3036, n_3037);
  xnor g2945 (Z[6], n_2949, n_3038);
  xnor g2948 (Z[7], n_3040, n_3041);
  xnor g2950 (Z[8], n_2854, n_3042);
  xnor g2953 (Z[9], n_3044, n_3045);
  xnor g2955 (Z[10], n_2954, n_3046);
  xnor g2958 (Z[11], n_3048, n_3049);
  xnor g2960 (Z[12], n_2923, n_3050);
  xnor g2963 (Z[13], n_3052, n_3053);
  xnor g2965 (Z[14], n_2959, n_3054);
  xnor g2968 (Z[15], n_3056, n_3057);
  xnor g2970 (Z[16], n_2879, n_3058);
  xnor g2973 (Z[17], n_3060, n_3061);
  xnor g2975 (Z[18], n_2964, n_3062);
  xnor g2978 (Z[19], n_3064, n_3065);
  xnor g2980 (Z[20], n_2926, n_3066);
  xnor g2983 (Z[21], n_3068, n_3069);
  xnor g2985 (Z[22], n_2969, n_3070);
  xnor g2988 (Z[23], n_3072, n_3073);
  xnor g2990 (Z[24], n_2903, n_3074);
  xnor g2993 (Z[25], n_3076, n_3077);
  xnor g2995 (Z[26], n_2974, n_3078);
  xnor g2998 (Z[27], n_3080, n_3081);
  xnor g3000 (Z[28], n_2929, n_3082);
  xnor g3003 (Z[29], n_3084, n_3085);
  xnor g3005 (Z[30], n_2979, n_3086);
  xnor g3008 (Z[31], n_3088, n_3089);
  xnor g3010 (Z[32], n_2890, n_3090);
  xnor g3013 (Z[33], n_3092, n_3093);
  xnor g3015 (Z[34], n_2984, n_3094);
  xnor g3018 (Z[35], n_3096, n_3097);
  xnor g3020 (Z[36], n_2932, n_3098);
  xnor g3023 (Z[37], n_3100, n_3101);
  xnor g3025 (Z[38], n_2989, n_3102);
  xnor g3028 (Z[39], n_3104, n_3105);
  xnor g3030 (Z[40], n_2908, n_3106);
  xnor g3033 (Z[41], n_3108, n_3109);
  xnor g3035 (Z[42], n_2994, n_3110);
  xnor g3038 (Z[43], n_3112, n_3113);
  xnor g3040 (Z[44], n_2935, n_3114);
  xnor g3043 (Z[45], n_3116, n_3117);
  xnor g3045 (Z[46], n_2999, n_3118);
  xnor g3048 (Z[47], n_3120, n_3121);
  xnor g3050 (Z[48], n_2897, n_3122);
  xnor g3053 (Z[49], n_3124, n_3125);
  xnor g3055 (Z[50], n_3004, n_3126);
  xnor g3058 (Z[51], n_3128, n_3129);
  xnor g3060 (Z[52], n_2938, n_3130);
  xnor g3063 (Z[53], n_3132, n_3133);
  xnor g3065 (Z[54], n_3009, n_3134);
  xnor g3068 (Z[55], n_3136, n_3137);
  xnor g3070 (Z[56], n_2913, n_3138);
  xnor g3073 (Z[57], n_3140, n_3141);
  xnor g3075 (Z[58], n_3014, n_3142);
  xnor g3078 (Z[59], n_3144, n_3145);
  xnor g3080 (Z[60], n_2941, n_3146);
  xnor g3083 (Z[61], n_3148, n_3149);
  xnor g3085 (Z[62], n_3019, n_3150);
  xnor g3088 (Z[63], n_3152, n_3153);
  xnor g3090 (Z[64], n_2917, n_3154);
  xnor g3093 (Z[65], n_3156, n_3157);
  xnor g3095 (Z[66], n_3024, n_3158);
  xnor g3098 (Z[67], n_3160, n_3161);
  xnor g3100 (Z[68], n_2944, n_3162);
  or g3113 (n_271, wc, wc0, n_116);
  not gc0 (wc0, n_947);
  not gc (wc, n_959);
  or g3114 (n_310, wc1, wc2, n_264);
  not gc2 (wc2, n_1009);
  not gc1 (wc1, n_1045);
  or g3115 (n_330, wc3, wc4, n_264);
  not gc4 (wc4, n_979);
  not gc3 (wc3, n_1007);
  or g3116 (n_355, wc5, n_308, n_269);
  not gc5 (wc5, n_1141);
  or g3117 (n_378, n_264, n_269, n_278);
  or g3118 (n_406, wc6, wc7, n_264);
  not gc7 (wc7, n_1141);
  not gc6 (wc6, n_1268);
  or g3119 (n_462, wc8, wc9, n_308);
  not gc9 (wc9, n_1396);
  not gc8 (wc8, n_1397);
  xnor g3120 (n_2222, A[50], A[48]);
  or g3121 (n_2223, wc10, A[50]);
  not gc10 (wc10, A[48]);
  or g3122 (n_2225, wc11, A[50]);
  not gc11 (wc11, A[44]);
  xnor g3123 (n_2262, A[49], A[37]);
  or g3124 (n_2263, wc12, A[49]);
  not gc12 (wc12, A[37]);
  xnor g3125 (n_886, n_2314, A[47]);
  or g3126 (n_2364, wc13, A[47]);
  not gc13 (wc13, A[45]);
  or g3127 (n_2365, wc14, A[47]);
  not gc14 (wc14, A[39]);
  xnor g3129 (n_932, n_2198, A[49]);
  or g3130 (n_2456, wc15, A[49]);
  not gc15 (wc15, A[45]);
  or g3131 (n_2457, wc16, A[49]);
  not gc16 (wc16, A[47]);
  or g3132 (n_2231, wc17, A[50]);
  not gc17 (wc17, A[46]);
  or g3134 (n_2471, A[47], wc18);
  not gc18 (wc18, A[49]);
  or g3135 (n_2477, wc19, A[50]);
  not gc19 (wc19, A[47]);
  and g3136 (n_2689, wc20, A[50]);
  not gc20 (wc20, A[49]);
  or g3137 (n_2686, wc21, A[50]);
  not gc21 (wc21, A[49]);
  or g3138 (n_2321, A[49], wc22);
  not gc22 (wc22, n_860);
  xnor g3139 (n_906, n_800, n_2198);
  or g3140 (n_2404, A[47], wc23);
  not gc23 (wc23, n_800);
  or g3141 (n_2437, A[49], wc24);
  not gc24 (wc24, n_920);
  and g3142 (n_2692, wc25, n_944);
  not gc25 (wc25, n_2491);
  or g3144 (n_3030, n_2493, wc26);
  not gc26 (wc26, n_947);
  or g3145 (n_3033, n_2489, wc27);
  not gc27 (wc27, n_944);
  xnor g3146 (n_2230, A[50], A[46]);
  or g3147 (n_2233, wc28, A[50]);
  not gc28 (wc28, A[40]);
  or g3148 (n_2264, A[49], wc29);
  not gc29 (wc29, n_831);
  xnor g3149 (n_2318, n_831, A[49]);
  xnor g3150 (n_56, n_2126, n_939);
  or g3151 (n_2472, A[47], wc30);
  not gc30 (wc30, n_939);
  and g3152 (n_2681, A[49], wc31);
  not gc31 (wc31, n_124);
  or g3153 (n_2682, A[49], wc32);
  not gc32 (wc32, n_124);
  or g3154 (n_3034, wc33, n_2499);
  not gc33 (wc33, n_2494);
  or g3155 (n_3162, wc34, n_2689);
  not gc34 (wc34, n_2686);
  and g3156 (n_2695, wc35, n_2496);
  not gc35 (wc35, n_2497);
  not g3157 (Z[2], n_3030);
  or g3158 (n_3037, wc36, n_2495);
  not gc36 (wc36, n_2496);
  or g3159 (n_3038, wc37, n_2505);
  not gc37 (wc37, n_2500);
  and g3160 (n_2697, wc38, n_2502);
  not gc38 (wc38, n_2503);
  or g3163 (n_3041, wc39, n_2501);
  not gc39 (wc39, n_2502);
  or g3164 (n_3161, wc40, n_2681);
  not gc40 (wc40, n_2682);
  and g3165 (n_2702, wc41, n_2508);
  not gc41 (wc41, n_2509);
  and g3166 (n_2698, wc42, n_2694);
  not gc42 (wc42, n_2695);
  or g3167 (n_2921, n_2692, wc43);
  not gc43 (wc43, n_2700);
  or g3168 (n_2948, n_2499, n_2692);
  xor g3169 (Z[3], n_947, n_3033);
  xor g3170 (Z[4], n_2692, n_3034);
  or g3171 (n_3042, wc44, n_2511);
  not gc44 (wc44, n_2506);
  or g3172 (n_3045, wc45, n_2507);
  not gc45 (wc45, n_2508);
  and g3173 (n_2802, n_2682, wc46);
  not gc46 (wc46, n_2683);
  and g3174 (n_2809, wc47, n_2697);
  not gc47 (wc47, n_2698);
  or g3175 (n_2810, n_2806, n_2692);
  or g3176 (n_3046, wc48, n_2517);
  not gc48 (wc48, n_2512);
  or g3177 (n_3157, wc49, n_2675);
  not gc49 (wc49, n_2676);
  or g3178 (n_3158, wc50, n_2685);
  not gc50 (wc50, n_2680);
  and g3179 (n_2704, wc51, n_2514);
  not gc51 (wc51, n_2515);
  and g3180 (n_2709, wc52, n_2520);
  not gc52 (wc52, n_2521);
  and g3181 (n_2800, wc53, n_2676);
  not gc53 (wc53, n_2677);
  or g3182 (n_2951, wc54, n_2505);
  not gc54 (wc54, n_2949);
  or g3183 (n_3049, wc55, n_2513);
  not gc55 (wc55, n_2514);
  or g3184 (n_3050, wc56, n_2523);
  not gc56 (wc56, n_2518);
  or g3185 (n_3053, wc57, n_2519);
  not gc57 (wc57, n_2520);
  or g3186 (n_3154, wc58, n_2679);
  not gc58 (wc58, n_2674);
  and g3187 (n_2711, wc59, n_2526);
  not gc59 (wc59, n_2527);
  and g3188 (n_2795, wc60, n_2670);
  not gc60 (wc60, n_2671);
  and g3189 (n_2705, wc61, n_2701);
  not gc61 (wc61, n_2702);
  and g3190 (n_2803, wc62, n_2799);
  not gc62 (wc62, n_2800);
  or g3191 (n_2953, wc63, n_2511);
  not gc63 (wc63, n_2854);
  or g3192 (n_3054, wc64, n_2529);
  not gc64 (wc64, n_2524);
  or g3193 (n_3057, wc65, n_2525);
  not gc65 (wc65, n_2526);
  or g3194 (n_3149, wc66, n_2663);
  not gc66 (wc66, n_2664);
  or g3195 (n_3150, wc67, n_2673);
  not gc67 (wc67, n_2668);
  or g3196 (n_3153, wc68, n_2669);
  not gc68 (wc68, n_2670);
  and g3197 (n_2716, wc69, n_2532);
  not gc69 (wc69, n_2533);
  and g3198 (n_2793, wc70, n_2664);
  not gc70 (wc70, n_2665);
  and g3199 (n_2812, wc71, n_2704);
  not gc71 (wc71, n_2705);
  and g3200 (n_2712, wc72, n_2708);
  not gc72 (wc72, n_2709);
  and g3201 (n_2919, wc73, n_2802);
  not gc73 (wc73, n_2803);
  or g3202 (n_2900, wc74, n_2816);
  not gc74 (wc74, n_2854);
  or g3203 (n_3058, wc75, n_2535);
  not gc75 (wc75, n_2530);
  or g3204 (n_3061, wc76, n_2531);
  not gc76 (wc76, n_2532);
  or g3205 (n_3066, wc77, n_2547);
  not gc77 (wc77, n_2542);
  or g3206 (n_3146, wc78, n_2667);
  not gc78 (wc78, n_2662);
  and g3207 (n_2718, wc79, n_2538);
  not gc79 (wc79, n_2539);
  and g3208 (n_2723, wc80, n_2544);
  not gc80 (wc80, n_2545);
  and g3209 (n_2788, wc81, n_2658);
  not gc81 (wc81, n_2659);
  and g3210 (n_2813, wc82, n_2711);
  not gc82 (wc82, n_2712);
  and g3211 (n_2796, wc83, n_2792);
  not gc83 (wc83, n_2793);
  or g3212 (n_2956, wc84, n_2517);
  not gc84 (wc84, n_2954);
  or g3213 (n_3062, wc85, n_2541);
  not gc85 (wc85, n_2536);
  or g3214 (n_3065, wc86, n_2537);
  not gc86 (wc86, n_2538);
  or g3215 (n_3069, wc87, n_2543);
  not gc87 (wc87, n_2544);
  or g3216 (n_3070, wc88, n_2553);
  not gc88 (wc88, n_2548);
  or g3217 (n_3141, wc89, n_2651);
  not gc89 (wc89, n_2652);
  or g3218 (n_3142, wc90, n_2661);
  not gc90 (wc90, n_2656);
  or g3219 (n_3145, wc91, n_2657);
  not gc91 (wc91, n_2658);
  and g3220 (n_2725, wc92, n_2550);
  not gc92 (wc92, n_2551);
  and g3221 (n_2730, wc93, n_2556);
  not gc93 (wc93, n_2557);
  and g3222 (n_2732, wc94, n_2562);
  not gc94 (wc94, n_2563);
  and g3223 (n_2737, wc95, n_2568);
  not gc95 (wc95, n_2569);
  and g3224 (n_2739, wc96, n_2574);
  not gc96 (wc96, n_2575);
  and g3225 (n_2744, wc97, n_2580);
  not gc97 (wc97, n_2581);
  and g3226 (n_2746, wc98, n_2586);
  not gc98 (wc98, n_2587);
  and g3227 (n_2751, wc99, n_2592);
  not gc99 (wc99, n_2593);
  and g3228 (n_2753, wc100, n_2598);
  not gc100 (wc100, n_2599);
  and g3229 (n_2758, wc101, n_2604);
  not gc101 (wc101, n_2605);
  and g3230 (n_2760, wc102, n_2610);
  not gc102 (wc102, n_2611);
  and g3231 (n_2765, wc103, n_2616);
  not gc103 (wc103, n_2617);
  and g3232 (n_2767, wc104, n_2622);
  not gc104 (wc104, n_2623);
  and g3233 (n_2772, wc105, n_2628);
  not gc105 (wc105, n_2629);
  and g3234 (n_2774, wc106, n_2634);
  not gc106 (wc106, n_2635);
  and g3235 (n_2719, wc107, n_2715);
  not gc107 (wc107, n_2716);
  and g3236 (n_2849, wc108, n_2795);
  not gc108 (wc108, n_2796);
  or g3237 (n_2958, wc109, n_2523);
  not gc109 (wc109, n_2923);
  or g3238 (n_3073, wc110, n_2549);
  not gc110 (wc110, n_2550);
  or g3239 (n_3074, wc111, n_2559);
  not gc111 (wc111, n_2554);
  or g3240 (n_3077, wc112, n_2555);
  not gc112 (wc112, n_2556);
  or g3241 (n_3078, wc113, n_2565);
  not gc113 (wc113, n_2560);
  or g3242 (n_3081, wc114, n_2561);
  not gc114 (wc114, n_2562);
  or g3243 (n_3082, wc115, n_2571);
  not gc115 (wc115, n_2566);
  or g3244 (n_3085, wc116, n_2567);
  not gc116 (wc116, n_2568);
  or g3245 (n_3086, wc117, n_2577);
  not gc117 (wc117, n_2572);
  or g3246 (n_3089, wc118, n_2573);
  not gc118 (wc118, n_2574);
  or g3247 (n_3090, wc119, n_2583);
  not gc119 (wc119, n_2578);
  or g3248 (n_3093, wc120, n_2579);
  not gc120 (wc120, n_2580);
  or g3249 (n_3094, wc121, n_2589);
  not gc121 (wc121, n_2584);
  or g3250 (n_3097, wc122, n_2585);
  not gc122 (wc122, n_2586);
  or g3251 (n_3098, wc123, n_2595);
  not gc123 (wc123, n_2590);
  or g3252 (n_3101, wc124, n_2591);
  not gc124 (wc124, n_2592);
  or g3253 (n_3102, wc125, n_2601);
  not gc125 (wc125, n_2596);
  or g3254 (n_3105, wc126, n_2597);
  not gc126 (wc126, n_2598);
  or g3255 (n_3106, wc127, n_2607);
  not gc127 (wc127, n_2602);
  or g3256 (n_3109, wc128, n_2603);
  not gc128 (wc128, n_2604);
  or g3257 (n_3110, wc129, n_2613);
  not gc129 (wc129, n_2608);
  or g3258 (n_3113, wc130, n_2609);
  not gc130 (wc130, n_2610);
  or g3259 (n_3114, wc131, n_2619);
  not gc131 (wc131, n_2614);
  or g3260 (n_3117, wc132, n_2615);
  not gc132 (wc132, n_2616);
  or g3261 (n_3118, wc133, n_2625);
  not gc133 (wc133, n_2620);
  or g3262 (n_3121, wc134, n_2621);
  not gc134 (wc134, n_2622);
  or g3263 (n_3122, wc135, n_2631);
  not gc135 (wc135, n_2626);
  or g3264 (n_3125, wc136, n_2627);
  not gc136 (wc136, n_2628);
  or g3265 (n_3126, wc137, n_2637);
  not gc137 (wc137, n_2632);
  or g3266 (n_3129, wc138, n_2633);
  not gc138 (wc138, n_2634);
  and g3267 (n_2779, wc139, n_2640);
  not gc139 (wc139, n_2641);
  and g3268 (n_2818, wc140, n_2718);
  not gc140 (wc140, n_2719);
  and g3269 (n_2726, wc141, n_2722);
  not gc141 (wc141, n_2723);
  and g3270 (n_2733, wc142, n_2729);
  not gc142 (wc142, n_2730);
  and g3271 (n_2740, wc143, n_2736);
  not gc143 (wc143, n_2737);
  and g3272 (n_2747, wc144, n_2743);
  not gc144 (wc144, n_2744);
  and g3273 (n_2754, wc145, n_2750);
  not gc145 (wc145, n_2751);
  and g3274 (n_2761, wc146, n_2757);
  not gc146 (wc146, n_2758);
  and g3275 (n_2768, wc147, n_2764);
  not gc147 (wc147, n_2765);
  and g3276 (n_2775, wc148, n_2771);
  not gc148 (wc148, n_2772);
  and g3277 (n_2855, n_2813, wc149);
  not gc149 (wc149, n_2814);
  or g3278 (n_3130, wc150, n_2643);
  not gc150 (wc150, n_2638);
  or g3279 (n_3133, wc151, n_2639);
  not gc151 (wc151, n_2640);
  and g3280 (n_2781, wc152, n_2646);
  not gc152 (wc152, n_2647);
  and g3281 (n_2819, wc153, n_2725);
  not gc153 (wc153, n_2726);
  and g3282 (n_2824, wc154, n_2732);
  not gc154 (wc154, n_2733);
  and g3283 (n_2825, wc155, n_2739);
  not gc155 (wc155, n_2740);
  and g3284 (n_2830, wc156, n_2746);
  not gc156 (wc156, n_2747);
  and g3285 (n_2831, wc157, n_2753);
  not gc157 (wc157, n_2754);
  and g3286 (n_2836, wc158, n_2760);
  not gc158 (wc158, n_2761);
  and g3287 (n_2837, wc159, n_2767);
  not gc159 (wc159, n_2768);
  and g3288 (n_2842, wc160, n_2774);
  not gc160 (wc160, n_2775);
  or g3289 (n_2961, wc161, n_2529);
  not gc161 (wc161, n_2959);
  or g3290 (n_3134, wc162, n_2649);
  not gc162 (wc162, n_2644);
  or g3291 (n_3137, wc163, n_2645);
  not gc163 (wc163, n_2646);
  and g3292 (n_2786, wc164, n_2652);
  not gc164 (wc164, n_2653);
  and g3293 (n_2782, wc165, n_2778);
  not gc165 (wc165, n_2779);
  or g3294 (n_2902, wc166, n_2822);
  not gc166 (wc166, n_2879);
  or g3295 (n_2963, wc167, n_2535);
  not gc167 (wc167, n_2879);
  or g3296 (n_3138, wc168, n_2655);
  not gc168 (wc168, n_2650);
  and g3297 (n_2843, wc169, n_2781);
  not gc169 (wc169, n_2782);
  and g3298 (n_2789, wc170, n_2785);
  not gc170 (wc170, n_2786);
  and g3299 (n_2858, n_2819, wc171);
  not gc171 (wc171, n_2820);
  and g3300 (n_2860, n_2825, wc172);
  not gc172 (wc172, n_2826);
  and g3301 (n_2865, n_2831, wc173);
  not gc173 (wc173, n_2832);
  and g3302 (n_2867, n_2837, wc174);
  not gc174 (wc174, n_2838);
  or g3303 (n_2882, n_2878, wc175);
  not gc175 (wc175, n_2879);
  and g3304 (n_2848, wc176, n_2788);
  not gc176 (wc176, n_2789);
  and g3305 (n_2861, wc177, n_2857);
  not gc177 (wc177, n_2858);
  and g3306 (n_2868, wc178, n_2864);
  not gc178 (wc178, n_2865);
  or g3307 (n_2966, wc179, n_2541);
  not gc179 (wc179, n_2964);
  or g3308 (n_2968, wc180, n_2547);
  not gc180 (wc180, n_2926);
  and g3309 (n_2872, n_2843, wc181);
  not gc181 (wc181, n_2844);
  and g3310 (n_2881, wc182, n_2860);
  not gc182 (wc182, n_2861);
  and g3311 (n_2884, wc183, n_2867);
  not gc183 (wc183, n_2868);
  or g3312 (n_2905, wc184, n_2828);
  not gc184 (wc184, n_2903);
  or g3313 (n_2973, wc185, n_2559);
  not gc185 (wc185, n_2903);
  and g3314 (n_2874, n_2849, wc186);
  not gc186 (wc186, n_2850);
  and g3315 (n_2875, wc187, n_2871);
  not gc187 (wc187, n_2872);
  or g3316 (n_2971, wc188, n_2553);
  not gc188 (wc188, n_2969);
  or g3317 (n_2894, wc189, n_2888);
  not gc189 (wc189, n_2890);
  or g3318 (n_2907, wc190, n_2834);
  not gc190 (wc190, n_2890);
  or g3319 (n_2976, wc191, n_2565);
  not gc191 (wc191, n_2974);
  or g3320 (n_2978, wc192, n_2571);
  not gc192 (wc192, n_2929);
  or g3321 (n_2983, wc193, n_2583);
  not gc193 (wc193, n_2890);
  and g3322 (n_2885, wc194, n_2874);
  not gc194 (wc194, n_2875);
  or g3323 (n_2910, wc195, n_2840);
  not gc195 (wc195, n_2908);
  or g3324 (n_2912, wc196, n_2846);
  not gc196 (wc196, n_2897);
  or g3325 (n_2981, wc197, n_2577);
  not gc197 (wc197, n_2979);
  or g3326 (n_2986, wc198, n_2589);
  not gc198 (wc198, n_2984);
  or g3327 (n_2988, wc199, n_2595);
  not gc199 (wc199, n_2932);
  or g3328 (n_2993, wc200, n_2607);
  not gc200 (wc200, n_2908);
  or g3329 (n_3003, wc201, n_2631);
  not gc201 (wc201, n_2897);
  and g3330 (n_2891, n_2885, wc202);
  not gc202 (wc202, n_2886);
  or g3331 (n_2915, wc203, n_2852);
  not gc203 (wc203, n_2913);
  or g3332 (n_2991, wc204, n_2601);
  not gc204 (wc204, n_2989);
  or g3333 (n_2996, wc205, n_2613);
  not gc205 (wc205, n_2994);
  or g3334 (n_2998, wc206, n_2619);
  not gc206 (wc206, n_2935);
  or g3335 (n_3006, wc207, n_2637);
  not gc207 (wc207, n_3004);
  or g3336 (n_3008, wc208, n_2643);
  not gc208 (wc208, n_2938);
  or g3337 (n_3013, wc209, n_2655);
  not gc209 (wc209, n_2913);
  or g3338 (n_2920, wc210, n_2916);
  not gc210 (wc210, n_2917);
  or g3339 (n_3023, wc211, n_2679);
  not gc211 (wc211, n_2917);
  or g3340 (n_3001, wc212, n_2625);
  not gc212 (wc212, n_2999);
  or g3341 (n_3011, wc213, n_2649);
  not gc213 (wc213, n_3009);
  or g3342 (n_3016, wc214, n_2661);
  not gc214 (wc214, n_3014);
  or g3343 (n_3018, wc215, n_2667);
  not gc215 (wc215, n_2941);
  or g3344 (n_3026, wc216, n_2685);
  not gc216 (wc216, n_3024);
  or g3345 (n_3028, n_2689, wc217);
  not gc217 (wc217, n_2944);
  or g3346 (n_3021, wc218, n_2673);
  not gc218 (wc218, n_3019);
  not g3347 (Z[69], n_3164);
endmodule

module mult_signed_const_11527_GENERIC(A, Z);
  input [50:0] A;
  output [69:0] Z;
  wire [50:0] A;
  wire [69:0] Z;
  mult_signed_const_11527_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_11946_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [52:0] A;
  output [71:0] Z;
  wire [52:0] A;
  wire [71:0] Z;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285;
  wire n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381;
  wire n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389;
  wire n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397;
  wire n_398, n_399, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502;
  wire n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510;
  wire n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518;
  wire n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526;
  wire n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550;
  wire n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558;
  wire n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566;
  wire n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574;
  wire n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582;
  wire n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590;
  wire n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598;
  wire n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606;
  wire n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614;
  wire n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622;
  wire n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630;
  wire n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638;
  wire n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646;
  wire n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654;
  wire n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662;
  wire n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670;
  wire n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678;
  wire n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686;
  wire n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694;
  wire n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702;
  wire n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710;
  wire n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718;
  wire n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726;
  wire n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734;
  wire n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758;
  wire n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766;
  wire n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774;
  wire n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782;
  wire n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790;
  wire n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798;
  wire n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806;
  wire n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814;
  wire n_815, n_816, n_819, n_820, n_821, n_822, n_823, n_824;
  wire n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832;
  wire n_837, n_838, n_839, n_840, n_842, n_843, n_844, n_845;
  wire n_846, n_847, n_848, n_849, n_851, n_852, n_853, n_855;
  wire n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864;
  wire n_867, n_868, n_872, n_873, n_874, n_875, n_876, n_877;
  wire n_878, n_879, n_883, n_884, n_885, n_886, n_887, n_888;
  wire n_889, n_890, n_891, n_892, n_895, n_896, n_897, n_898;
  wire n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_907;
  wire n_908, n_911, n_912, n_913, n_914, n_915, n_916, n_921;
  wire n_922, n_923, n_924, n_925, n_926, n_927, n_929, n_930;
  wire n_931, n_932, n_933, n_934, n_935, n_936, n_939, n_940;
  wire n_942, n_943, n_944, n_945, n_948, n_950, n_951, n_952;
  wire n_955, n_958, n_959, n_963, n_964, n_968, n_969, n_971;
  wire n_972, n_975, n_978, n_979, n_980, n_981, n_982, n_983;
  wire n_984, n_985, n_986, n_987, n_988, n_990, n_991, n_992;
  wire n_993, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003;
  wire n_1004, n_1006, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013;
  wire n_1014, n_1016, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023;
  wire n_1024, n_1025, n_1028, n_1030, n_1031, n_1032, n_1033, n_1034;
  wire n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1044;
  wire n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055;
  wire n_1056, n_1057, n_1058, n_1059, n_1062, n_1063, n_1064, n_1066;
  wire n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074;
  wire n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1082, n_1083;
  wire n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092;
  wire n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100;
  wire n_1101, n_1102, n_1103, n_1105, n_1106, n_1108, n_1109, n_1110;
  wire n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118;
  wire n_1119, n_1120, n_1121, n_1122, n_1125, n_1126, n_1127, n_1128;
  wire n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137;
  wire n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145;
  wire n_1146, n_1147, n_1148, n_1154, n_1155, n_1158, n_1159, n_1160;
  wire n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168;
  wire n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1177;
  wire n_1178, n_1180, n_1181, n_1184, n_1185, n_1186, n_1187, n_1188;
  wire n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196;
  wire n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204;
  wire n_1208, n_1209, n_1210, n_1211, n_1212, n_1214, n_1215, n_1216;
  wire n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224;
  wire n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1242, n_1243, n_1244;
  wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253;
  wire n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261;
  wire n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269;
  wire n_1274, n_1276, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283;
  wire n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291;
  wire n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299;
  wire n_1300, n_1301, n_1304, n_1305, n_1306, n_1307, n_1308, n_1310;
  wire n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318;
  wire n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326;
  wire n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1336;
  wire n_1338, n_1339, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347;
  wire n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355;
  wire n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363;
  wire n_1364, n_1365, n_1368, n_1370, n_1371, n_1374, n_1375, n_1376;
  wire n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384;
  wire n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392;
  wire n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1400, n_1402;
  wire n_1403, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412;
  wire n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420;
  wire n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428;
  wire n_1429, n_1432, n_1434, n_1435, n_1438, n_1439, n_1440, n_1441;
  wire n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449;
  wire n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457;
  wire n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1466;
  wire n_1467, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476;
  wire n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484;
  wire n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492;
  wire n_1493, n_1496, n_1498, n_1499, n_1502, n_1503, n_1504, n_1505;
  wire n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513;
  wire n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521;
  wire n_1522, n_1523, n_1524, n_1525, n_1526, n_1528, n_1530, n_1531;
  wire n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541;
  wire n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557;
  wire n_1560, n_1562, n_1563, n_1566, n_1567, n_1568, n_1569, n_1570;
  wire n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578;
  wire n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586;
  wire n_1587, n_1588, n_1589, n_1590, n_1592, n_1594, n_1595, n_1598;
  wire n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606;
  wire n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614;
  wire n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1624;
  wire n_1626, n_1627, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635;
  wire n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643;
  wire n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651;
  wire n_1652, n_1653, n_1654, n_1655, n_1656, n_1658, n_1659, n_1662;
  wire n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670;
  wire n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678;
  wire n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1688;
  wire n_1690, n_1691, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699;
  wire n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707;
  wire n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715;
  wire n_1716, n_1717, n_1720, n_1722, n_1723, n_1726, n_1727, n_1728;
  wire n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736;
  wire n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744;
  wire n_1745, n_1746, n_1747, n_1748, n_1749, n_1752, n_1754, n_1755;
  wire n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765;
  wire n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773;
  wire n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781;
  wire n_1784, n_1786, n_1787, n_1790, n_1791, n_1792, n_1793, n_1794;
  wire n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802;
  wire n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810;
  wire n_1811, n_1812, n_1813, n_1816, n_1818, n_1819, n_1822, n_1823;
  wire n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831;
  wire n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839;
  wire n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1848, n_1850;
  wire n_1851, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860;
  wire n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868;
  wire n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876;
  wire n_1877, n_1880, n_1882, n_1883, n_1886, n_1887, n_1888, n_1889;
  wire n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897;
  wire n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905;
  wire n_1906, n_1907, n_1908, n_1909, n_1912, n_1914, n_1915, n_1918;
  wire n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926;
  wire n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934;
  wire n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1944;
  wire n_1946, n_1947, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955;
  wire n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963;
  wire n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971;
  wire n_1972, n_1973, n_1976, n_1978, n_1979, n_1982, n_1983, n_1984;
  wire n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992;
  wire n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000;
  wire n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008;
  wire n_2010, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019;
  wire n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027;
  wire n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035;
  wire n_2036, n_2037, n_2038, n_2039, n_2040, n_2042, n_2045, n_2046;
  wire n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054;
  wire n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062;
  wire n_2063, n_2064, n_2065, n_2069, n_2070, n_2072, n_2076, n_2077;
  wire n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085;
  wire n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093;
  wire n_2094, n_2095, n_2096, n_2097, n_2101, n_2102, n_2104, n_2108;
  wire n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116;
  wire n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124;
  wire n_2125, n_2126, n_2127, n_2128, n_2129, n_2133, n_2138, n_2139;
  wire n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147;
  wire n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155;
  wire n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2165, n_2170;
  wire n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178;
  wire n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186;
  wire n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194;
  wire n_2198, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208;
  wire n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216;
  wire n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224;
  wire n_2225, n_2226, n_2230, n_2234, n_2235, n_2236, n_2237, n_2238;
  wire n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246;
  wire n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254;
  wire n_2255, n_2256, n_2257, n_2258, n_2259, n_2261, n_2262, n_2266;
  wire n_2267, n_2268, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275;
  wire n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283;
  wire n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2292;
  wire n_2293, n_2294, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307;
  wire n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315;
  wire n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323;
  wire n_2325, n_2326, n_2327, n_2329, n_2334, n_2335, n_2336, n_2337;
  wire n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345;
  wire n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353;
  wire n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2369, n_2370;
  wire n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378;
  wire n_2379, n_2380, n_2381, n_2386, n_2387, n_2389, n_2390, n_2392;
  wire n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400;
  wire n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408;
  wire n_2409, n_2412, n_2413, n_2414, n_2417, n_2418, n_2419, n_2420;
  wire n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428;
  wire n_2429, n_2430, n_2431, n_2432, n_2433, n_2442, n_2444, n_2445;
  wire n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453;
  wire n_2454, n_2455, n_2456, n_2457, n_2458, n_2461, n_2462, n_2465;
  wire n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475;
  wire n_2476, n_2477, n_2480, n_2481, n_2482, n_2486, n_2487, n_2488;
  wire n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496;
  wire n_2497, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510;
  wire n_2511, n_2512, n_2513, n_2514, n_2517, n_2522, n_2523, n_2524;
  wire n_2525, n_2526, n_2527, n_2528, n_2529, n_2534, n_2535, n_2536;
  wire n_2537, n_2538, n_2539, n_2540, n_2541, n_2546, n_2547, n_2548;
  wire n_2549, n_2550, n_2551, n_2552, n_2553, n_2556, n_2557, n_2558;
  wire n_2559, n_2560, n_2561, n_2565, n_2566, n_2567, n_2568, n_2569;
  wire n_2570, n_2571, n_2572, n_2573, n_2576, n_2577, n_2589, n_2591;
  wire n_2593, n_2594, n_2595, n_2596, n_2597, n_2599, n_2600, n_2601;
  wire n_2602, n_2603, n_2605, n_2606, n_2607, n_2608, n_2609, n_2611;
  wire n_2612, n_2613, n_2614, n_2615, n_2617, n_2618, n_2619, n_2620;
  wire n_2621, n_2623, n_2624, n_2625, n_2626, n_2627, n_2629, n_2630;
  wire n_2631, n_2632, n_2633, n_2635, n_2636, n_2637, n_2638, n_2639;
  wire n_2641, n_2642, n_2643, n_2644, n_2645, n_2647, n_2648, n_2649;
  wire n_2650, n_2651, n_2653, n_2654, n_2655, n_2656, n_2657, n_2659;
  wire n_2660, n_2661, n_2662, n_2663, n_2665, n_2666, n_2667, n_2668;
  wire n_2669, n_2671, n_2672, n_2673, n_2674, n_2675, n_2677, n_2678;
  wire n_2679, n_2680, n_2681, n_2683, n_2684, n_2685, n_2686, n_2687;
  wire n_2689, n_2690, n_2691, n_2692, n_2693, n_2695, n_2696, n_2697;
  wire n_2698, n_2699, n_2701, n_2702, n_2703, n_2704, n_2705, n_2707;
  wire n_2708, n_2709, n_2710, n_2711, n_2713, n_2714, n_2715, n_2716;
  wire n_2717, n_2719, n_2720, n_2721, n_2722, n_2723, n_2725, n_2726;
  wire n_2727, n_2728, n_2729, n_2731, n_2732, n_2733, n_2734, n_2735;
  wire n_2737, n_2738, n_2739, n_2740, n_2741, n_2743, n_2744, n_2745;
  wire n_2746, n_2747, n_2749, n_2750, n_2751, n_2752, n_2753, n_2755;
  wire n_2756, n_2757, n_2758, n_2759, n_2761, n_2762, n_2763, n_2764;
  wire n_2765, n_2767, n_2768, n_2769, n_2770, n_2771, n_2773, n_2774;
  wire n_2775, n_2776, n_2777, n_2779, n_2780, n_2781, n_2782, n_2783;
  wire n_2785, n_2786, n_2787, n_2788, n_2789, n_2791, n_2792, n_2795;
  wire n_2798, n_2800, n_2801, n_2803, n_2804, n_2806, n_2807, n_2808;
  wire n_2810, n_2811, n_2813, n_2814, n_2815, n_2817, n_2818, n_2820;
  wire n_2821, n_2822, n_2824, n_2825, n_2827, n_2828, n_2829, n_2831;
  wire n_2832, n_2834, n_2835, n_2836, n_2838, n_2839, n_2841, n_2842;
  wire n_2843, n_2845, n_2846, n_2848, n_2849, n_2850, n_2852, n_2853;
  wire n_2855, n_2856, n_2857, n_2859, n_2860, n_2862, n_2863, n_2864;
  wire n_2866, n_2867, n_2869, n_2870, n_2871, n_2873, n_2874, n_2876;
  wire n_2877, n_2878, n_2880, n_2881, n_2883, n_2884, n_2885, n_2887;
  wire n_2888, n_2890, n_2891, n_2892, n_2894, n_2895, n_2897, n_2898;
  wire n_2899, n_2901, n_2902, n_2904, n_2905, n_2906, n_2908, n_2909;
  wire n_2911, n_2912, n_2913, n_2914, n_2917, n_2918, n_2919, n_2920;
  wire n_2921, n_2922, n_2924, n_2925, n_2926, n_2927, n_2928, n_2930;
  wire n_2931, n_2932, n_2933, n_2934, n_2936, n_2937, n_2938, n_2939;
  wire n_2940, n_2942, n_2943, n_2944, n_2945, n_2946, n_2948, n_2949;
  wire n_2950, n_2951, n_2952, n_2954, n_2955, n_2956, n_2957, n_2958;
  wire n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967;
  wire n_2968, n_2970, n_2971, n_2973, n_2974, n_2975, n_2977, n_2978;
  wire n_2980, n_2981, n_2982, n_2984, n_2985, n_2987, n_2988, n_2989;
  wire n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2998, n_2999;
  wire n_3000, n_3001, n_3002, n_3004, n_3005, n_3006, n_3007, n_3008;
  wire n_3009, n_3011, n_3013, n_3014, n_3016, n_3018, n_3019, n_3021;
  wire n_3023, n_3024, n_3026, n_3028, n_3029, n_3030, n_3031, n_3032;
  wire n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040;
  wire n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048;
  wire n_3049, n_3050, n_3051, n_3052, n_3053, n_3057, n_3058, n_3060;
  wire n_3062, n_3063, n_3065, n_3067, n_3068, n_3070, n_3072, n_3073;
  wire n_3075, n_3077, n_3078, n_3080, n_3082, n_3083, n_3085, n_3087;
  wire n_3088, n_3090, n_3092, n_3093, n_3095, n_3097, n_3098, n_3100;
  wire n_3102, n_3103, n_3105, n_3107, n_3108, n_3110, n_3112, n_3113;
  wire n_3115, n_3117, n_3118, n_3120, n_3122, n_3123, n_3125, n_3127;
  wire n_3128, n_3130, n_3132, n_3133, n_3135, n_3137, n_3138, n_3140;
  wire n_3142, n_3145, n_3146, n_3148, n_3149, n_3150, n_3152, n_3153;
  wire n_3154, n_3156, n_3157, n_3158, n_3160, n_3161, n_3162, n_3164;
  wire n_3165, n_3166, n_3168, n_3169, n_3170, n_3172, n_3173, n_3174;
  wire n_3176, n_3177, n_3178, n_3180, n_3181, n_3182, n_3184, n_3185;
  wire n_3186, n_3188, n_3189, n_3190, n_3192, n_3193, n_3194, n_3196;
  wire n_3197, n_3198, n_3200, n_3201, n_3202, n_3204, n_3205, n_3206;
  wire n_3208, n_3209, n_3210, n_3212, n_3213, n_3214, n_3216, n_3217;
  wire n_3218, n_3220, n_3221, n_3222, n_3224, n_3225, n_3226, n_3228;
  wire n_3229, n_3230, n_3232, n_3233, n_3234, n_3236, n_3237, n_3238;
  wire n_3240, n_3241, n_3242, n_3244, n_3245, n_3246, n_3248, n_3249;
  wire n_3250, n_3252, n_3253, n_3254, n_3256, n_3257, n_3258, n_3260;
  wire n_3261, n_3262, n_3264, n_3265, n_3266, n_3268, n_3269, n_3270;
  wire n_3272, n_3273, n_3274, n_3276, n_3277, n_3278, n_3280;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g420 (n_193, A[4], A[0]);
  and g2 (n_120, A[4], A[0]);
  xor g421 (n_978, A[1], A[3]);
  xor g422 (n_192, n_978, A[5]);
  nand g3 (n_979, A[1], A[3]);
  nand g423 (n_980, A[5], A[3]);
  nand g424 (n_981, A[1], A[5]);
  nand g425 (n_119, n_979, n_980, n_981);
  xor g426 (n_271, A[6], A[4]);
  and g427 (n_272, A[6], A[4]);
  xor g428 (n_982, A[0], A[2]);
  xor g429 (n_191, n_982, n_271);
  nand g430 (n_983, A[0], A[2]);
  nand g4 (n_984, n_271, A[2]);
  nand g5 (n_985, A[0], n_271);
  nand g431 (n_118, n_983, n_984, n_985);
  xor g432 (n_986, A[1], A[7]);
  xor g433 (n_273, n_986, A[5]);
  nand g434 (n_987, A[1], A[7]);
  nand g435 (n_988, A[5], A[7]);
  nand g6 (n_275, n_987, n_988, n_981);
  xor g437 (n_990, A[3], n_272);
  xor g438 (n_190, n_990, n_273);
  nand g439 (n_991, A[3], n_272);
  nand g440 (n_992, n_273, n_272);
  nand g441 (n_993, A[3], n_273);
  nand g442 (n_117, n_991, n_992, n_993);
  xor g443 (n_274, A[8], A[6]);
  and g444 (n_277, A[8], A[6]);
  xor g446 (n_276, n_982, A[4]);
  nand g449 (n_997, A[2], A[4]);
  xor g451 (n_998, n_274, n_275);
  xor g452 (n_189, n_998, n_276);
  nand g453 (n_999, n_274, n_275);
  nand g454 (n_1000, n_276, n_275);
  nand g455 (n_1001, n_274, n_276);
  nand g456 (n_116, n_999, n_1000, n_1001);
  xor g457 (n_1002, A[1], A[9]);
  xor g458 (n_279, n_1002, A[3]);
  nand g459 (n_1003, A[1], A[9]);
  nand g460 (n_1004, A[3], A[9]);
  nand g462 (n_282, n_1003, n_1004, n_979);
  xor g463 (n_1006, A[7], A[5]);
  xor g464 (n_280, n_1006, n_277);
  nand g466 (n_1008, n_277, A[5]);
  nand g467 (n_1009, A[7], n_277);
  nand g468 (n_284, n_988, n_1008, n_1009);
  xor g469 (n_1010, n_278, n_279);
  xor g470 (n_188, n_1010, n_280);
  nand g471 (n_1011, n_278, n_279);
  nand g472 (n_1012, n_280, n_279);
  nand g473 (n_1013, n_278, n_280);
  nand g474 (n_115, n_1011, n_1012, n_1013);
  xor g475 (n_281, A[10], A[8]);
  and g476 (n_286, A[10], A[8]);
  xor g477 (n_1014, A[4], A[2]);
  xor g478 (n_283, n_1014, A[6]);
  nand g480 (n_1016, A[6], A[2]);
  xor g483 (n_1018, A[0], n_281);
  xor g484 (n_285, n_1018, n_282);
  nand g485 (n_1019, A[0], n_281);
  nand g486 (n_1020, n_282, n_281);
  nand g487 (n_1021, A[0], n_282);
  nand g488 (n_290, n_1019, n_1020, n_1021);
  xor g489 (n_1022, n_283, n_284);
  xor g490 (n_187, n_1022, n_285);
  nand g491 (n_1023, n_283, n_284);
  nand g492 (n_1024, n_285, n_284);
  nand g493 (n_1025, n_283, n_285);
  nand g494 (n_114, n_1023, n_1024, n_1025);
  xor g496 (n_288, n_1002, A[5]);
  nand g498 (n_1028, A[5], A[9]);
  nand g500 (n_293, n_1003, n_1028, n_981);
  xor g501 (n_1030, A[3], A[11]);
  xor g502 (n_289, n_1030, A[7]);
  nand g503 (n_1031, A[3], A[11]);
  nand g504 (n_1032, A[7], A[11]);
  nand g505 (n_1033, A[3], A[7]);
  nand g506 (n_294, n_1031, n_1032, n_1033);
  xor g507 (n_1034, n_286, n_287);
  xor g508 (n_291, n_1034, n_288);
  nand g509 (n_1035, n_286, n_287);
  nand g510 (n_1036, n_288, n_287);
  nand g511 (n_1037, n_286, n_288);
  nand g512 (n_298, n_1035, n_1036, n_1037);
  xor g513 (n_1038, n_289, n_290);
  xor g514 (n_186, n_1038, n_291);
  nand g515 (n_1039, n_289, n_290);
  nand g516 (n_1040, n_291, n_290);
  nand g517 (n_1041, n_289, n_291);
  nand g518 (n_113, n_1039, n_1040, n_1041);
  xor g519 (n_292, A[12], A[10]);
  and g520 (n_299, A[12], A[10]);
  xor g522 (n_295, n_271, A[8]);
  nand g524 (n_1044, A[8], A[4]);
  xor g528 (n_296, n_982, n_292);
  nand g530 (n_1048, n_292, A[0]);
  nand g531 (n_1049, A[2], n_292);
  nand g532 (n_303, n_983, n_1048, n_1049);
  xor g533 (n_1050, n_293, n_294);
  xor g534 (n_297, n_1050, n_295);
  nand g535 (n_1051, n_293, n_294);
  nand g536 (n_1052, n_295, n_294);
  nand g537 (n_1053, n_293, n_295);
  nand g538 (n_305, n_1051, n_1052, n_1053);
  xor g539 (n_1054, n_296, n_297);
  xor g540 (n_185, n_1054, n_298);
  nand g541 (n_1055, n_296, n_297);
  nand g542 (n_1056, n_298, n_297);
  nand g543 (n_1057, n_296, n_298);
  nand g544 (n_112, n_1055, n_1056, n_1057);
  xor g545 (n_1058, A[1], A[11]);
  xor g546 (n_302, n_1058, A[7]);
  nand g547 (n_1059, A[1], A[11]);
  nand g550 (n_308, n_1059, n_1032, n_987);
  xor g551 (n_1062, A[5], A[13]);
  xor g552 (n_301, n_1062, A[3]);
  nand g553 (n_1063, A[5], A[13]);
  nand g554 (n_1064, A[3], A[13]);
  nand g556 (n_309, n_1063, n_1064, n_980);
  xor g557 (n_1066, A[9], n_299);
  xor g558 (n_304, n_1066, n_300);
  nand g559 (n_1067, A[9], n_299);
  nand g560 (n_1068, n_300, n_299);
  nand g561 (n_1069, A[9], n_300);
  nand g562 (n_312, n_1067, n_1068, n_1069);
  xor g563 (n_1070, n_301, n_302);
  xor g564 (n_306, n_1070, n_303);
  nand g565 (n_1071, n_301, n_302);
  nand g566 (n_1072, n_303, n_302);
  nand g567 (n_1073, n_301, n_303);
  nand g568 (n_314, n_1071, n_1072, n_1073);
  xor g569 (n_1074, n_304, n_305);
  xor g570 (n_184, n_1074, n_306);
  nand g571 (n_1075, n_304, n_305);
  nand g572 (n_1076, n_306, n_305);
  nand g573 (n_1077, n_304, n_306);
  nand g574 (n_111, n_1075, n_1076, n_1077);
  xor g575 (n_307, A[14], A[12]);
  and g576 (n_316, A[14], A[12]);
  xor g577 (n_1078, A[8], A[0]);
  xor g578 (n_311, n_1078, A[6]);
  nand g579 (n_1079, A[8], A[0]);
  nand g580 (n_1080, A[6], A[0]);
  xor g583 (n_1082, A[10], A[4]);
  xor g584 (n_310, n_1082, A[2]);
  nand g585 (n_1083, A[10], A[4]);
  nand g587 (n_1085, A[10], A[2]);
  nand g588 (n_318, n_1083, n_997, n_1085);
  xor g589 (n_1086, n_307, n_308);
  xor g590 (n_313, n_1086, n_309);
  nand g591 (n_1087, n_307, n_308);
  nand g592 (n_1088, n_309, n_308);
  nand g593 (n_1089, n_307, n_309);
  nand g594 (n_322, n_1087, n_1088, n_1089);
  xor g595 (n_1090, n_310, n_311);
  xor g596 (n_315, n_1090, n_312);
  nand g597 (n_1091, n_310, n_311);
  nand g598 (n_1092, n_312, n_311);
  nand g599 (n_1093, n_310, n_312);
  nand g600 (n_325, n_1091, n_1092, n_1093);
  xor g601 (n_1094, n_313, n_314);
  xor g602 (n_183, n_1094, n_315);
  nand g603 (n_1095, n_313, n_314);
  nand g604 (n_1096, n_315, n_314);
  nand g605 (n_1097, n_313, n_315);
  nand g606 (n_110, n_1095, n_1096, n_1097);
  xor g607 (n_1098, A[1], A[15]);
  xor g608 (n_319, n_1098, A[13]);
  nand g609 (n_1099, A[1], A[15]);
  nand g610 (n_1100, A[13], A[15]);
  nand g611 (n_1101, A[1], A[13]);
  nand g612 (n_327, n_1099, n_1100, n_1101);
  xor g613 (n_1102, A[9], A[7]);
  xor g614 (n_320, n_1102, A[11]);
  nand g615 (n_1103, A[9], A[7]);
  nand g617 (n_1105, A[9], A[11]);
  nand g618 (n_328, n_1103, n_1032, n_1105);
  xor g619 (n_1106, A[5], A[3]);
  xor g620 (n_321, n_1106, n_316);
  nand g622 (n_1108, n_316, A[3]);
  nand g623 (n_1109, A[5], n_316);
  nand g624 (n_331, n_980, n_1108, n_1109);
  xor g625 (n_1110, n_317, n_318);
  xor g626 (n_323, n_1110, n_319);
  nand g627 (n_1111, n_317, n_318);
  nand g628 (n_1112, n_319, n_318);
  nand g629 (n_1113, n_317, n_319);
  nand g630 (n_333, n_1111, n_1112, n_1113);
  xor g631 (n_1114, n_320, n_321);
  xor g632 (n_324, n_1114, n_322);
  nand g633 (n_1115, n_320, n_321);
  nand g634 (n_1116, n_322, n_321);
  nand g635 (n_1117, n_320, n_322);
  nand g636 (n_335, n_1115, n_1116, n_1117);
  xor g637 (n_1118, n_323, n_324);
  xor g638 (n_182, n_1118, n_325);
  nand g639 (n_1119, n_323, n_324);
  nand g640 (n_1120, n_325, n_324);
  nand g641 (n_1121, n_323, n_325);
  nand g642 (n_109, n_1119, n_1120, n_1121);
  xor g643 (n_326, A[16], A[14]);
  and g644 (n_337, A[16], A[14]);
  xor g645 (n_1122, A[10], A[2]);
  xor g646 (n_330, n_1122, A[0]);
  nand g649 (n_1125, A[10], A[0]);
  nand g650 (n_338, n_1085, n_983, n_1125);
  xor g651 (n_1126, A[8], A[12]);
  xor g652 (n_329, n_1126, A[6]);
  nand g653 (n_1127, A[8], A[12]);
  nand g654 (n_1128, A[6], A[12]);
  xor g657 (n_1130, A[4], n_326);
  xor g658 (n_332, n_1130, n_327);
  nand g659 (n_1131, A[4], n_326);
  nand g660 (n_1132, n_327, n_326);
  nand g661 (n_1133, A[4], n_327);
  nand g662 (n_343, n_1131, n_1132, n_1133);
  xor g663 (n_1134, n_328, n_329);
  xor g664 (n_334, n_1134, n_330);
  nand g665 (n_1135, n_328, n_329);
  nand g666 (n_1136, n_330, n_329);
  nand g667 (n_1137, n_328, n_330);
  nand g668 (n_345, n_1135, n_1136, n_1137);
  xor g669 (n_1138, n_331, n_332);
  xor g670 (n_336, n_1138, n_333);
  nand g671 (n_1139, n_331, n_332);
  nand g672 (n_1140, n_333, n_332);
  nand g673 (n_1141, n_331, n_333);
  nand g674 (n_347, n_1139, n_1140, n_1141);
  xor g675 (n_1142, n_334, n_335);
  xor g676 (n_181, n_1142, n_336);
  nand g677 (n_1143, n_334, n_335);
  nand g678 (n_1144, n_336, n_335);
  nand g679 (n_1145, n_334, n_336);
  nand g680 (n_108, n_1143, n_1144, n_1145);
  xor g681 (n_1146, A[1], A[17]);
  xor g682 (n_341, n_1146, A[15]);
  nand g683 (n_1147, A[1], A[17]);
  nand g684 (n_1148, A[15], A[17]);
  nand g686 (n_350, n_1147, n_1148, n_1099);
  xor g688 (n_342, n_1030, A[9]);
  nand g692 (n_352, n_1031, n_1105, n_1004);
  xor g693 (n_1154, A[13], A[7]);
  xor g694 (n_340, n_1154, A[5]);
  nand g695 (n_1155, A[13], A[7]);
  nand g698 (n_351, n_1155, n_988, n_1063);
  xor g699 (n_1158, n_337, n_338);
  xor g700 (n_344, n_1158, n_339);
  nand g701 (n_1159, n_337, n_338);
  nand g702 (n_1160, n_339, n_338);
  nand g703 (n_1161, n_337, n_339);
  nand g704 (n_356, n_1159, n_1160, n_1161);
  xor g705 (n_1162, n_340, n_341);
  xor g706 (n_346, n_1162, n_342);
  nand g707 (n_1163, n_340, n_341);
  nand g708 (n_1164, n_342, n_341);
  nand g709 (n_1165, n_340, n_342);
  nand g710 (n_358, n_1163, n_1164, n_1165);
  xor g711 (n_1166, n_343, n_344);
  xor g712 (n_348, n_1166, n_345);
  nand g713 (n_1167, n_343, n_344);
  nand g714 (n_1168, n_345, n_344);
  nand g715 (n_1169, n_343, n_345);
  nand g716 (n_360, n_1167, n_1168, n_1169);
  xor g717 (n_1170, n_346, n_347);
  xor g718 (n_180, n_1170, n_348);
  nand g719 (n_1171, n_346, n_347);
  nand g720 (n_1172, n_348, n_347);
  nand g721 (n_1173, n_346, n_348);
  nand g722 (n_107, n_1171, n_1172, n_1173);
  xor g723 (n_349, A[18], A[16]);
  and g724 (n_362, A[18], A[16]);
  xor g725 (n_1174, A[12], A[4]);
  xor g726 (n_353, n_1174, A[2]);
  nand g727 (n_1175, A[12], A[4]);
  nand g729 (n_1177, A[12], A[2]);
  nand g730 (n_363, n_1175, n_997, n_1177);
  xor g731 (n_1178, A[10], A[0]);
  xor g732 (n_354, n_1178, A[14]);
  nand g734 (n_1180, A[14], A[0]);
  nand g735 (n_1181, A[10], A[14]);
  nand g736 (n_364, n_1125, n_1180, n_1181);
  xor g738 (n_355, n_274, n_349);
  nand g740 (n_1184, n_349, A[6]);
  nand g741 (n_1185, A[8], n_349);
  xor g743 (n_1186, n_350, n_351);
  xor g744 (n_357, n_1186, n_352);
  nand g745 (n_1187, n_350, n_351);
  nand g746 (n_1188, n_352, n_351);
  nand g747 (n_1189, n_350, n_352);
  nand g748 (n_121, n_1187, n_1188, n_1189);
  xor g749 (n_1190, n_353, n_354);
  xor g750 (n_359, n_1190, n_355);
  nand g751 (n_1191, n_353, n_354);
  nand g752 (n_1192, n_355, n_354);
  nand g753 (n_1193, n_353, n_355);
  nand g754 (n_122, n_1191, n_1192, n_1193);
  xor g755 (n_1194, n_356, n_357);
  xor g756 (n_361, n_1194, n_358);
  nand g757 (n_1195, n_356, n_357);
  nand g758 (n_1196, n_358, n_357);
  nand g759 (n_1197, n_356, n_358);
  nand g760 (n_125, n_1195, n_1196, n_1197);
  xor g761 (n_1198, n_359, n_360);
  xor g762 (n_179, n_1198, n_361);
  nand g763 (n_1199, n_359, n_360);
  nand g764 (n_1200, n_361, n_360);
  nand g765 (n_1201, n_359, n_361);
  nand g766 (n_106, n_1199, n_1200, n_1201);
  xor g767 (n_1202, A[1], A[19]);
  xor g768 (n_366, n_1202, A[13]);
  nand g769 (n_1203, A[1], A[19]);
  nand g770 (n_1204, A[13], A[19]);
  nand g772 (n_371, n_1203, n_1204, n_1101);
  xor g774 (n_367, n_1106, A[17]);
  nand g776 (n_1208, A[17], A[3]);
  nand g777 (n_1209, A[5], A[17]);
  nand g778 (n_372, n_980, n_1208, n_1209);
  xor g779 (n_1210, A[11], A[15]);
  xor g780 (n_365, n_1210, A[9]);
  nand g781 (n_1211, A[11], A[15]);
  nand g782 (n_1212, A[9], A[15]);
  nand g784 (n_373, n_1211, n_1212, n_1105);
  xor g785 (n_1214, A[7], n_362);
  xor g786 (n_369, n_1214, n_363);
  nand g787 (n_1215, A[7], n_362);
  nand g788 (n_1216, n_363, n_362);
  nand g789 (n_1217, A[7], n_363);
  nand g790 (n_377, n_1215, n_1216, n_1217);
  xor g791 (n_1218, n_364, n_365);
  xor g792 (n_123, n_1218, n_366);
  nand g793 (n_1219, n_364, n_365);
  nand g794 (n_1220, n_366, n_365);
  nand g795 (n_1221, n_364, n_366);
  nand g796 (n_379, n_1219, n_1220, n_1221);
  xor g797 (n_1222, n_367, n_368);
  xor g798 (n_124, n_1222, n_369);
  nand g799 (n_1223, n_367, n_368);
  nand g800 (n_1224, n_369, n_368);
  nand g801 (n_1225, n_367, n_369);
  nand g802 (n_381, n_1223, n_1224, n_1225);
  xor g803 (n_1226, n_121, n_122);
  xor g804 (n_370, n_1226, n_123);
  nand g805 (n_1227, n_121, n_122);
  nand g806 (n_1228, n_123, n_122);
  nand g807 (n_1229, n_121, n_123);
  nand g808 (n_383, n_1227, n_1228, n_1229);
  xor g809 (n_1230, n_124, n_125);
  xor g810 (n_178, n_1230, n_370);
  nand g811 (n_1231, n_124, n_125);
  nand g812 (n_1232, n_370, n_125);
  nand g813 (n_1233, n_124, n_370);
  nand g814 (n_105, n_1231, n_1232, n_1233);
  xor g815 (n_1234, A[20], A[18]);
  xor g816 (n_375, n_1234, A[14]);
  nand g817 (n_1235, A[20], A[18]);
  nand g818 (n_1236, A[14], A[18]);
  nand g819 (n_1237, A[20], A[14]);
  nand g820 (n_385, n_1235, n_1236, n_1237);
  xor g822 (n_376, n_271, A[12]);
  xor g827 (n_1242, A[2], A[16]);
  xor g828 (n_374, n_1242, A[10]);
  nand g829 (n_1243, A[2], A[16]);
  nand g830 (n_1244, A[10], A[16]);
  nand g832 (n_387, n_1243, n_1244, n_1085);
  xor g833 (n_1246, A[8], n_371);
  xor g834 (n_378, n_1246, n_372);
  nand g835 (n_1247, A[8], n_371);
  nand g836 (n_1248, n_372, n_371);
  nand g837 (n_1249, A[8], n_372);
  nand g838 (n_391, n_1247, n_1248, n_1249);
  xor g839 (n_1250, n_373, n_374);
  xor g840 (n_380, n_1250, n_375);
  nand g841 (n_1251, n_373, n_374);
  nand g842 (n_1252, n_375, n_374);
  nand g843 (n_1253, n_373, n_375);
  nand g844 (n_393, n_1251, n_1252, n_1253);
  xor g845 (n_1254, n_376, n_377);
  xor g846 (n_382, n_1254, n_378);
  nand g847 (n_1255, n_376, n_377);
  nand g848 (n_1256, n_378, n_377);
  nand g849 (n_1257, n_376, n_378);
  nand g850 (n_395, n_1255, n_1256, n_1257);
  xor g851 (n_1258, n_379, n_380);
  xor g852 (n_384, n_1258, n_381);
  nand g853 (n_1259, n_379, n_380);
  nand g854 (n_1260, n_381, n_380);
  nand g855 (n_1261, n_379, n_381);
  nand g856 (n_397, n_1259, n_1260, n_1261);
  xor g857 (n_1262, n_382, n_383);
  xor g858 (n_177, n_1262, n_384);
  nand g859 (n_1263, n_382, n_383);
  nand g860 (n_1264, n_384, n_383);
  nand g861 (n_1265, n_382, n_384);
  nand g862 (n_104, n_1263, n_1264, n_1265);
  xor g863 (n_1266, A[21], A[19]);
  xor g864 (n_389, n_1266, A[15]);
  nand g865 (n_1267, A[21], A[19]);
  nand g866 (n_1268, A[15], A[19]);
  nand g867 (n_1269, A[21], A[15]);
  nand g868 (n_399, n_1267, n_1268, n_1269);
  xor g870 (n_390, n_1006, A[13]);
  xor g875 (n_1274, A[3], A[17]);
  xor g876 (n_388, n_1274, A[11]);
  nand g878 (n_1276, A[11], A[17]);
  nand g880 (n_401, n_1208, n_1276, n_1031);
  xor g881 (n_1278, A[9], n_385);
  xor g882 (n_392, n_1278, n_386);
  nand g883 (n_1279, A[9], n_385);
  nand g884 (n_1280, n_386, n_385);
  nand g885 (n_1281, A[9], n_386);
  nand g886 (n_405, n_1279, n_1280, n_1281);
  xor g887 (n_1282, n_387, n_388);
  xor g888 (n_394, n_1282, n_389);
  nand g889 (n_1283, n_387, n_388);
  nand g890 (n_1284, n_389, n_388);
  nand g891 (n_1285, n_387, n_389);
  nand g892 (n_407, n_1283, n_1284, n_1285);
  xor g893 (n_1286, n_390, n_391);
  xor g894 (n_396, n_1286, n_392);
  nand g895 (n_1287, n_390, n_391);
  nand g896 (n_1288, n_392, n_391);
  nand g897 (n_1289, n_390, n_392);
  nand g898 (n_409, n_1287, n_1288, n_1289);
  xor g899 (n_1290, n_393, n_394);
  xor g900 (n_398, n_1290, n_395);
  nand g901 (n_1291, n_393, n_394);
  nand g902 (n_1292, n_395, n_394);
  nand g903 (n_1293, n_393, n_395);
  nand g904 (n_412, n_1291, n_1292, n_1293);
  xor g905 (n_1294, n_396, n_397);
  xor g906 (n_176, n_1294, n_398);
  nand g907 (n_1295, n_396, n_397);
  nand g908 (n_1296, n_398, n_397);
  nand g909 (n_1297, n_396, n_398);
  nand g910 (n_103, n_1295, n_1296, n_1297);
  xor g911 (n_1298, A[22], A[20]);
  xor g912 (n_403, n_1298, A[16]);
  nand g913 (n_1299, A[22], A[20]);
  nand g914 (n_1300, A[16], A[20]);
  nand g915 (n_1301, A[22], A[16]);
  nand g916 (n_413, n_1299, n_1300, n_1301);
  xor g918 (n_404, n_274, A[14]);
  nand g920 (n_1304, A[14], A[6]);
  nand g921 (n_1305, A[8], A[14]);
  xor g923 (n_1306, A[4], A[18]);
  xor g924 (n_402, n_1306, A[12]);
  nand g925 (n_1307, A[4], A[18]);
  nand g926 (n_1308, A[12], A[18]);
  nand g928 (n_415, n_1307, n_1308, n_1175);
  xor g929 (n_1310, A[10], n_399);
  xor g930 (n_406, n_1310, n_351);
  nand g931 (n_1311, A[10], n_399);
  nand g932 (n_1312, n_351, n_399);
  nand g933 (n_1313, A[10], n_351);
  nand g934 (n_419, n_1311, n_1312, n_1313);
  xor g935 (n_1314, n_401, n_402);
  xor g936 (n_408, n_1314, n_403);
  nand g937 (n_1315, n_401, n_402);
  nand g938 (n_1316, n_403, n_402);
  nand g939 (n_1317, n_401, n_403);
  nand g940 (n_421, n_1315, n_1316, n_1317);
  xor g941 (n_1318, n_404, n_405);
  xor g942 (n_410, n_1318, n_406);
  nand g943 (n_1319, n_404, n_405);
  nand g944 (n_1320, n_406, n_405);
  nand g945 (n_1321, n_404, n_406);
  nand g946 (n_423, n_1319, n_1320, n_1321);
  xor g947 (n_1322, n_407, n_408);
  xor g948 (n_411, n_1322, n_409);
  nand g949 (n_1323, n_407, n_408);
  nand g950 (n_1324, n_409, n_408);
  nand g951 (n_1325, n_407, n_409);
  nand g952 (n_426, n_1323, n_1324, n_1325);
  xor g953 (n_1326, n_410, n_411);
  xor g954 (n_175, n_1326, n_412);
  nand g955 (n_1327, n_410, n_411);
  nand g956 (n_1328, n_412, n_411);
  nand g957 (n_1329, n_410, n_412);
  nand g958 (n_102, n_1327, n_1328, n_1329);
  xor g959 (n_1330, A[23], A[21]);
  xor g960 (n_417, n_1330, A[17]);
  nand g961 (n_1331, A[23], A[21]);
  nand g962 (n_1332, A[17], A[21]);
  nand g963 (n_1333, A[23], A[17]);
  nand g964 (n_427, n_1331, n_1332, n_1333);
  xor g966 (n_418, n_1102, A[15]);
  nand g968 (n_1336, A[15], A[7]);
  nand g970 (n_428, n_1103, n_1336, n_1212);
  xor g971 (n_1338, A[5], A[19]);
  xor g972 (n_416, n_1338, A[13]);
  nand g973 (n_1339, A[5], A[19]);
  nand g976 (n_429, n_1339, n_1204, n_1063);
  xor g977 (n_1342, A[11], n_413);
  xor g978 (n_420, n_1342, n_414);
  nand g979 (n_1343, A[11], n_413);
  nand g980 (n_1344, n_414, n_413);
  nand g981 (n_1345, A[11], n_414);
  nand g982 (n_194, n_1343, n_1344, n_1345);
  xor g983 (n_1346, n_415, n_416);
  xor g984 (n_422, n_1346, n_417);
  nand g985 (n_1347, n_415, n_416);
  nand g986 (n_1348, n_417, n_416);
  nand g987 (n_1349, n_415, n_417);
  nand g988 (n_433, n_1347, n_1348, n_1349);
  xor g989 (n_1350, n_418, n_419);
  xor g990 (n_424, n_1350, n_420);
  nand g991 (n_1351, n_418, n_419);
  nand g992 (n_1352, n_420, n_419);
  nand g993 (n_1353, n_418, n_420);
  nand g994 (n_435, n_1351, n_1352, n_1353);
  xor g995 (n_1354, n_421, n_422);
  xor g996 (n_425, n_1354, n_423);
  nand g997 (n_1355, n_421, n_422);
  nand g998 (n_1356, n_423, n_422);
  nand g999 (n_1357, n_421, n_423);
  nand g1000 (n_438, n_1355, n_1356, n_1357);
  xor g1001 (n_1358, n_424, n_425);
  xor g1002 (n_174, n_1358, n_426);
  nand g1003 (n_1359, n_424, n_425);
  nand g1004 (n_1360, n_426, n_425);
  nand g1005 (n_1361, n_424, n_426);
  nand g1006 (n_101, n_1359, n_1360, n_1361);
  xor g1007 (n_1362, A[24], A[22]);
  xor g1008 (n_431, n_1362, A[18]);
  nand g1009 (n_1363, A[24], A[22]);
  nand g1010 (n_1364, A[18], A[22]);
  nand g1011 (n_1365, A[24], A[18]);
  nand g1012 (n_439, n_1363, n_1364, n_1365);
  xor g1014 (n_432, n_281, A[16]);
  nand g1016 (n_1368, A[16], A[8]);
  xor g1019 (n_1370, A[6], A[20]);
  xor g1020 (n_430, n_1370, A[14]);
  nand g1021 (n_1371, A[6], A[20]);
  nand g1024 (n_441, n_1371, n_1237, n_1304);
  xor g1025 (n_1374, A[12], n_427);
  xor g1026 (n_195, n_1374, n_428);
  nand g1027 (n_1375, A[12], n_427);
  nand g1028 (n_1376, n_428, n_427);
  nand g1029 (n_1377, A[12], n_428);
  nand g1030 (n_445, n_1375, n_1376, n_1377);
  xor g1031 (n_1378, n_429, n_430);
  xor g1032 (n_434, n_1378, n_431);
  nand g1033 (n_1379, n_429, n_430);
  nand g1034 (n_1380, n_431, n_430);
  nand g1035 (n_1381, n_429, n_431);
  nand g1036 (n_447, n_1379, n_1380, n_1381);
  xor g1037 (n_1382, n_432, n_194);
  xor g1038 (n_436, n_1382, n_195);
  nand g1039 (n_1383, n_432, n_194);
  nand g1040 (n_1384, n_195, n_194);
  nand g1041 (n_1385, n_432, n_195);
  nand g1042 (n_449, n_1383, n_1384, n_1385);
  xor g1043 (n_1386, n_433, n_434);
  xor g1044 (n_437, n_1386, n_435);
  nand g1045 (n_1387, n_433, n_434);
  nand g1046 (n_1388, n_435, n_434);
  nand g1047 (n_1389, n_433, n_435);
  nand g1048 (n_452, n_1387, n_1388, n_1389);
  xor g1049 (n_1390, n_436, n_437);
  xor g1050 (n_173, n_1390, n_438);
  nand g1051 (n_1391, n_436, n_437);
  nand g1052 (n_1392, n_438, n_437);
  nand g1053 (n_1393, n_436, n_438);
  nand g1054 (n_100, n_1391, n_1392, n_1393);
  xor g1055 (n_1394, A[25], A[23]);
  xor g1056 (n_443, n_1394, A[19]);
  nand g1057 (n_1395, A[25], A[23]);
  nand g1058 (n_1396, A[19], A[23]);
  nand g1059 (n_1397, A[25], A[19]);
  nand g1060 (n_453, n_1395, n_1396, n_1397);
  xor g1061 (n_1398, A[11], A[9]);
  xor g1062 (n_444, n_1398, A[17]);
  nand g1064 (n_1400, A[17], A[9]);
  nand g1066 (n_454, n_1105, n_1400, n_1276);
  xor g1067 (n_1402, A[7], A[21]);
  xor g1068 (n_442, n_1402, A[15]);
  nand g1069 (n_1403, A[7], A[21]);
  nand g1072 (n_455, n_1403, n_1269, n_1336);
  xor g1073 (n_1406, A[13], n_439);
  xor g1074 (n_446, n_1406, n_440);
  nand g1075 (n_1407, A[13], n_439);
  nand g1076 (n_1408, n_440, n_439);
  nand g1077 (n_1409, A[13], n_440);
  nand g1078 (n_459, n_1407, n_1408, n_1409);
  xor g1079 (n_1410, n_441, n_442);
  xor g1080 (n_448, n_1410, n_443);
  nand g1081 (n_1411, n_441, n_442);
  nand g1082 (n_1412, n_443, n_442);
  nand g1083 (n_1413, n_441, n_443);
  nand g1084 (n_461, n_1411, n_1412, n_1413);
  xor g1085 (n_1414, n_444, n_445);
  xor g1086 (n_450, n_1414, n_446);
  nand g1087 (n_1415, n_444, n_445);
  nand g1088 (n_1416, n_446, n_445);
  nand g1089 (n_1417, n_444, n_446);
  nand g1090 (n_463, n_1415, n_1416, n_1417);
  xor g1091 (n_1418, n_447, n_448);
  xor g1092 (n_451, n_1418, n_449);
  nand g1093 (n_1419, n_447, n_448);
  nand g1094 (n_1420, n_449, n_448);
  nand g1095 (n_1421, n_447, n_449);
  nand g1096 (n_466, n_1419, n_1420, n_1421);
  xor g1097 (n_1422, n_450, n_451);
  xor g1098 (n_172, n_1422, n_452);
  nand g1099 (n_1423, n_450, n_451);
  nand g1100 (n_1424, n_452, n_451);
  nand g1101 (n_1425, n_450, n_452);
  nand g1102 (n_99, n_1423, n_1424, n_1425);
  xor g1103 (n_1426, A[26], A[24]);
  xor g1104 (n_457, n_1426, A[20]);
  nand g1105 (n_1427, A[26], A[24]);
  nand g1106 (n_1428, A[20], A[24]);
  nand g1107 (n_1429, A[26], A[20]);
  nand g1108 (n_467, n_1427, n_1428, n_1429);
  xor g1110 (n_458, n_292, A[18]);
  nand g1112 (n_1432, A[18], A[10]);
  xor g1115 (n_1434, A[8], A[22]);
  xor g1116 (n_456, n_1434, A[16]);
  nand g1117 (n_1435, A[8], A[22]);
  nand g1120 (n_469, n_1435, n_1301, n_1368);
  xor g1121 (n_1438, A[14], n_453);
  xor g1122 (n_460, n_1438, n_454);
  nand g1123 (n_1439, A[14], n_453);
  nand g1124 (n_1440, n_454, n_453);
  nand g1125 (n_1441, A[14], n_454);
  nand g1126 (n_473, n_1439, n_1440, n_1441);
  xor g1127 (n_1442, n_455, n_456);
  xor g1128 (n_462, n_1442, n_457);
  nand g1129 (n_1443, n_455, n_456);
  nand g1130 (n_1444, n_457, n_456);
  nand g1131 (n_1445, n_455, n_457);
  nand g1132 (n_475, n_1443, n_1444, n_1445);
  xor g1133 (n_1446, n_458, n_459);
  xor g1134 (n_464, n_1446, n_460);
  nand g1135 (n_1447, n_458, n_459);
  nand g1136 (n_1448, n_460, n_459);
  nand g1137 (n_1449, n_458, n_460);
  nand g1138 (n_477, n_1447, n_1448, n_1449);
  xor g1139 (n_1450, n_461, n_462);
  xor g1140 (n_465, n_1450, n_463);
  nand g1141 (n_1451, n_461, n_462);
  nand g1142 (n_1452, n_463, n_462);
  nand g1143 (n_1453, n_461, n_463);
  nand g1144 (n_480, n_1451, n_1452, n_1453);
  xor g1145 (n_1454, n_464, n_465);
  xor g1146 (n_171, n_1454, n_466);
  nand g1147 (n_1455, n_464, n_465);
  nand g1148 (n_1456, n_466, n_465);
  nand g1149 (n_1457, n_464, n_466);
  nand g1150 (n_98, n_1455, n_1456, n_1457);
  xor g1151 (n_1458, A[27], A[25]);
  xor g1152 (n_471, n_1458, A[21]);
  nand g1153 (n_1459, A[27], A[25]);
  nand g1154 (n_1460, A[21], A[25]);
  nand g1155 (n_1461, A[27], A[21]);
  nand g1156 (n_481, n_1459, n_1460, n_1461);
  xor g1157 (n_1462, A[13], A[11]);
  xor g1158 (n_472, n_1462, A[19]);
  nand g1159 (n_1463, A[13], A[11]);
  nand g1160 (n_1464, A[19], A[11]);
  nand g1162 (n_482, n_1463, n_1464, n_1204);
  xor g1163 (n_1466, A[9], A[23]);
  xor g1164 (n_470, n_1466, A[17]);
  nand g1165 (n_1467, A[9], A[23]);
  nand g1168 (n_483, n_1467, n_1333, n_1400);
  xor g1169 (n_1470, A[15], n_467);
  xor g1170 (n_474, n_1470, n_468);
  nand g1171 (n_1471, A[15], n_467);
  nand g1172 (n_1472, n_468, n_467);
  nand g1173 (n_1473, A[15], n_468);
  nand g1174 (n_487, n_1471, n_1472, n_1473);
  xor g1175 (n_1474, n_469, n_470);
  xor g1176 (n_476, n_1474, n_471);
  nand g1177 (n_1475, n_469, n_470);
  nand g1178 (n_1476, n_471, n_470);
  nand g1179 (n_1477, n_469, n_471);
  nand g1180 (n_489, n_1475, n_1476, n_1477);
  xor g1181 (n_1478, n_472, n_473);
  xor g1182 (n_478, n_1478, n_474);
  nand g1183 (n_1479, n_472, n_473);
  nand g1184 (n_1480, n_474, n_473);
  nand g1185 (n_1481, n_472, n_474);
  nand g1186 (n_491, n_1479, n_1480, n_1481);
  xor g1187 (n_1482, n_475, n_476);
  xor g1188 (n_479, n_1482, n_477);
  nand g1189 (n_1483, n_475, n_476);
  nand g1190 (n_1484, n_477, n_476);
  nand g1191 (n_1485, n_475, n_477);
  nand g1192 (n_494, n_1483, n_1484, n_1485);
  xor g1193 (n_1486, n_478, n_479);
  xor g1194 (n_170, n_1486, n_480);
  nand g1195 (n_1487, n_478, n_479);
  nand g1196 (n_1488, n_480, n_479);
  nand g1197 (n_1489, n_478, n_480);
  nand g1198 (n_97, n_1487, n_1488, n_1489);
  xor g1199 (n_1490, A[28], A[26]);
  xor g1200 (n_485, n_1490, A[22]);
  nand g1201 (n_1491, A[28], A[26]);
  nand g1202 (n_1492, A[22], A[26]);
  nand g1203 (n_1493, A[28], A[22]);
  nand g1204 (n_495, n_1491, n_1492, n_1493);
  xor g1206 (n_486, n_307, A[20]);
  nand g1208 (n_1496, A[20], A[12]);
  xor g1211 (n_1498, A[10], A[24]);
  xor g1212 (n_484, n_1498, A[18]);
  nand g1213 (n_1499, A[10], A[24]);
  nand g1216 (n_497, n_1499, n_1365, n_1432);
  xor g1217 (n_1502, A[16], n_481);
  xor g1218 (n_488, n_1502, n_482);
  nand g1219 (n_1503, A[16], n_481);
  nand g1220 (n_1504, n_482, n_481);
  nand g1221 (n_1505, A[16], n_482);
  nand g1222 (n_501, n_1503, n_1504, n_1505);
  xor g1223 (n_1506, n_483, n_484);
  xor g1224 (n_490, n_1506, n_485);
  nand g1225 (n_1507, n_483, n_484);
  nand g1226 (n_1508, n_485, n_484);
  nand g1227 (n_1509, n_483, n_485);
  nand g1228 (n_503, n_1507, n_1508, n_1509);
  xor g1229 (n_1510, n_486, n_487);
  xor g1230 (n_492, n_1510, n_488);
  nand g1231 (n_1511, n_486, n_487);
  nand g1232 (n_1512, n_488, n_487);
  nand g1233 (n_1513, n_486, n_488);
  nand g1234 (n_505, n_1511, n_1512, n_1513);
  xor g1235 (n_1514, n_489, n_490);
  xor g1236 (n_493, n_1514, n_491);
  nand g1237 (n_1515, n_489, n_490);
  nand g1238 (n_1516, n_491, n_490);
  nand g1239 (n_1517, n_489, n_491);
  nand g1240 (n_508, n_1515, n_1516, n_1517);
  xor g1241 (n_1518, n_492, n_493);
  xor g1242 (n_169, n_1518, n_494);
  nand g1243 (n_1519, n_492, n_493);
  nand g1244 (n_1520, n_494, n_493);
  nand g1245 (n_1521, n_492, n_494);
  nand g1246 (n_96, n_1519, n_1520, n_1521);
  xor g1247 (n_1522, A[29], A[27]);
  xor g1248 (n_499, n_1522, A[23]);
  nand g1249 (n_1523, A[29], A[27]);
  nand g1250 (n_1524, A[23], A[27]);
  nand g1251 (n_1525, A[29], A[23]);
  nand g1252 (n_509, n_1523, n_1524, n_1525);
  xor g1253 (n_1526, A[15], A[13]);
  xor g1254 (n_500, n_1526, A[21]);
  nand g1256 (n_1528, A[21], A[13]);
  nand g1258 (n_510, n_1100, n_1528, n_1269);
  xor g1259 (n_1530, A[11], A[25]);
  xor g1260 (n_498, n_1530, A[19]);
  nand g1261 (n_1531, A[11], A[25]);
  nand g1264 (n_511, n_1531, n_1397, n_1464);
  xor g1265 (n_1534, A[17], n_495);
  xor g1266 (n_502, n_1534, n_496);
  nand g1267 (n_1535, A[17], n_495);
  nand g1268 (n_1536, n_496, n_495);
  nand g1269 (n_1537, A[17], n_496);
  nand g1270 (n_515, n_1535, n_1536, n_1537);
  xor g1271 (n_1538, n_497, n_498);
  xor g1272 (n_504, n_1538, n_499);
  nand g1273 (n_1539, n_497, n_498);
  nand g1274 (n_1540, n_499, n_498);
  nand g1275 (n_1541, n_497, n_499);
  nand g1276 (n_517, n_1539, n_1540, n_1541);
  xor g1277 (n_1542, n_500, n_501);
  xor g1278 (n_506, n_1542, n_502);
  nand g1279 (n_1543, n_500, n_501);
  nand g1280 (n_1544, n_502, n_501);
  nand g1281 (n_1545, n_500, n_502);
  nand g1282 (n_519, n_1543, n_1544, n_1545);
  xor g1283 (n_1546, n_503, n_504);
  xor g1284 (n_507, n_1546, n_505);
  nand g1285 (n_1547, n_503, n_504);
  nand g1286 (n_1548, n_505, n_504);
  nand g1287 (n_1549, n_503, n_505);
  nand g1288 (n_522, n_1547, n_1548, n_1549);
  xor g1289 (n_1550, n_506, n_507);
  xor g1290 (n_168, n_1550, n_508);
  nand g1291 (n_1551, n_506, n_507);
  nand g1292 (n_1552, n_508, n_507);
  nand g1293 (n_1553, n_506, n_508);
  nand g1294 (n_95, n_1551, n_1552, n_1553);
  xor g1295 (n_1554, A[30], A[28]);
  xor g1296 (n_513, n_1554, A[24]);
  nand g1297 (n_1555, A[30], A[28]);
  nand g1298 (n_1556, A[24], A[28]);
  nand g1299 (n_1557, A[30], A[24]);
  nand g1300 (n_523, n_1555, n_1556, n_1557);
  xor g1302 (n_514, n_326, A[22]);
  nand g1304 (n_1560, A[22], A[14]);
  xor g1307 (n_1562, A[12], A[26]);
  xor g1308 (n_512, n_1562, A[20]);
  nand g1309 (n_1563, A[12], A[26]);
  nand g1312 (n_525, n_1563, n_1429, n_1496);
  xor g1313 (n_1566, A[18], n_509);
  xor g1314 (n_516, n_1566, n_510);
  nand g1315 (n_1567, A[18], n_509);
  nand g1316 (n_1568, n_510, n_509);
  nand g1317 (n_1569, A[18], n_510);
  nand g1318 (n_529, n_1567, n_1568, n_1569);
  xor g1319 (n_1570, n_511, n_512);
  xor g1320 (n_518, n_1570, n_513);
  nand g1321 (n_1571, n_511, n_512);
  nand g1322 (n_1572, n_513, n_512);
  nand g1323 (n_1573, n_511, n_513);
  nand g1324 (n_531, n_1571, n_1572, n_1573);
  xor g1325 (n_1574, n_514, n_515);
  xor g1326 (n_520, n_1574, n_516);
  nand g1327 (n_1575, n_514, n_515);
  nand g1328 (n_1576, n_516, n_515);
  nand g1329 (n_1577, n_514, n_516);
  nand g1330 (n_533, n_1575, n_1576, n_1577);
  xor g1331 (n_1578, n_517, n_518);
  xor g1332 (n_521, n_1578, n_519);
  nand g1333 (n_1579, n_517, n_518);
  nand g1334 (n_1580, n_519, n_518);
  nand g1335 (n_1581, n_517, n_519);
  nand g1336 (n_536, n_1579, n_1580, n_1581);
  xor g1337 (n_1582, n_520, n_521);
  xor g1338 (n_167, n_1582, n_522);
  nand g1339 (n_1583, n_520, n_521);
  nand g1340 (n_1584, n_522, n_521);
  nand g1341 (n_1585, n_520, n_522);
  nand g1342 (n_94, n_1583, n_1584, n_1585);
  xor g1343 (n_1586, A[31], A[29]);
  xor g1344 (n_527, n_1586, A[25]);
  nand g1345 (n_1587, A[31], A[29]);
  nand g1346 (n_1588, A[25], A[29]);
  nand g1347 (n_1589, A[31], A[25]);
  nand g1348 (n_537, n_1587, n_1588, n_1589);
  xor g1349 (n_1590, A[17], A[15]);
  xor g1350 (n_528, n_1590, A[23]);
  nand g1352 (n_1592, A[23], A[15]);
  nand g1354 (n_538, n_1148, n_1592, n_1333);
  xor g1355 (n_1594, A[13], A[27]);
  xor g1356 (n_526, n_1594, A[21]);
  nand g1357 (n_1595, A[13], A[27]);
  nand g1360 (n_539, n_1595, n_1461, n_1528);
  xor g1361 (n_1598, A[19], n_523);
  xor g1362 (n_530, n_1598, n_524);
  nand g1363 (n_1599, A[19], n_523);
  nand g1364 (n_1600, n_524, n_523);
  nand g1365 (n_1601, A[19], n_524);
  nand g1366 (n_543, n_1599, n_1600, n_1601);
  xor g1367 (n_1602, n_525, n_526);
  xor g1368 (n_532, n_1602, n_527);
  nand g1369 (n_1603, n_525, n_526);
  nand g1370 (n_1604, n_527, n_526);
  nand g1371 (n_1605, n_525, n_527);
  nand g1372 (n_545, n_1603, n_1604, n_1605);
  xor g1373 (n_1606, n_528, n_529);
  xor g1374 (n_534, n_1606, n_530);
  nand g1375 (n_1607, n_528, n_529);
  nand g1376 (n_1608, n_530, n_529);
  nand g1377 (n_1609, n_528, n_530);
  nand g1378 (n_547, n_1607, n_1608, n_1609);
  xor g1379 (n_1610, n_531, n_532);
  xor g1380 (n_535, n_1610, n_533);
  nand g1381 (n_1611, n_531, n_532);
  nand g1382 (n_1612, n_533, n_532);
  nand g1383 (n_1613, n_531, n_533);
  nand g1384 (n_550, n_1611, n_1612, n_1613);
  xor g1385 (n_1614, n_534, n_535);
  xor g1386 (n_166, n_1614, n_536);
  nand g1387 (n_1615, n_534, n_535);
  nand g1388 (n_1616, n_536, n_535);
  nand g1389 (n_1617, n_534, n_536);
  nand g1390 (n_93, n_1615, n_1616, n_1617);
  xor g1391 (n_1618, A[32], A[30]);
  xor g1392 (n_541, n_1618, A[26]);
  nand g1393 (n_1619, A[32], A[30]);
  nand g1394 (n_1620, A[26], A[30]);
  nand g1395 (n_1621, A[32], A[26]);
  nand g1396 (n_551, n_1619, n_1620, n_1621);
  xor g1398 (n_542, n_349, A[24]);
  nand g1400 (n_1624, A[24], A[16]);
  xor g1403 (n_1626, A[14], A[28]);
  xor g1404 (n_540, n_1626, A[22]);
  nand g1405 (n_1627, A[14], A[28]);
  nand g1408 (n_553, n_1627, n_1493, n_1560);
  xor g1409 (n_1630, A[20], n_537);
  xor g1410 (n_544, n_1630, n_538);
  nand g1411 (n_1631, A[20], n_537);
  nand g1412 (n_1632, n_538, n_537);
  nand g1413 (n_1633, A[20], n_538);
  nand g1414 (n_557, n_1631, n_1632, n_1633);
  xor g1415 (n_1634, n_539, n_540);
  xor g1416 (n_546, n_1634, n_541);
  nand g1417 (n_1635, n_539, n_540);
  nand g1418 (n_1636, n_541, n_540);
  nand g1419 (n_1637, n_539, n_541);
  nand g1420 (n_559, n_1635, n_1636, n_1637);
  xor g1421 (n_1638, n_542, n_543);
  xor g1422 (n_548, n_1638, n_544);
  nand g1423 (n_1639, n_542, n_543);
  nand g1424 (n_1640, n_544, n_543);
  nand g1425 (n_1641, n_542, n_544);
  nand g1426 (n_561, n_1639, n_1640, n_1641);
  xor g1427 (n_1642, n_545, n_546);
  xor g1428 (n_549, n_1642, n_547);
  nand g1429 (n_1643, n_545, n_546);
  nand g1430 (n_1644, n_547, n_546);
  nand g1431 (n_1645, n_545, n_547);
  nand g1432 (n_564, n_1643, n_1644, n_1645);
  xor g1433 (n_1646, n_548, n_549);
  xor g1434 (n_165, n_1646, n_550);
  nand g1435 (n_1647, n_548, n_549);
  nand g1436 (n_1648, n_550, n_549);
  nand g1437 (n_1649, n_548, n_550);
  nand g1438 (n_92, n_1647, n_1648, n_1649);
  xor g1439 (n_1650, A[33], A[31]);
  xor g1440 (n_555, n_1650, A[27]);
  nand g1441 (n_1651, A[33], A[31]);
  nand g1442 (n_1652, A[27], A[31]);
  nand g1443 (n_1653, A[33], A[27]);
  nand g1444 (n_565, n_1651, n_1652, n_1653);
  xor g1445 (n_1654, A[19], A[17]);
  xor g1446 (n_556, n_1654, A[25]);
  nand g1447 (n_1655, A[19], A[17]);
  nand g1448 (n_1656, A[25], A[17]);
  nand g1450 (n_566, n_1655, n_1656, n_1397);
  xor g1451 (n_1658, A[15], A[29]);
  xor g1452 (n_554, n_1658, A[23]);
  nand g1453 (n_1659, A[15], A[29]);
  nand g1456 (n_567, n_1659, n_1525, n_1592);
  xor g1457 (n_1662, A[21], n_551);
  xor g1458 (n_558, n_1662, n_552);
  nand g1459 (n_1663, A[21], n_551);
  nand g1460 (n_1664, n_552, n_551);
  nand g1461 (n_1665, A[21], n_552);
  nand g1462 (n_571, n_1663, n_1664, n_1665);
  xor g1463 (n_1666, n_553, n_554);
  xor g1464 (n_560, n_1666, n_555);
  nand g1465 (n_1667, n_553, n_554);
  nand g1466 (n_1668, n_555, n_554);
  nand g1467 (n_1669, n_553, n_555);
  nand g1468 (n_573, n_1667, n_1668, n_1669);
  xor g1469 (n_1670, n_556, n_557);
  xor g1470 (n_562, n_1670, n_558);
  nand g1471 (n_1671, n_556, n_557);
  nand g1472 (n_1672, n_558, n_557);
  nand g1473 (n_1673, n_556, n_558);
  nand g1474 (n_575, n_1671, n_1672, n_1673);
  xor g1475 (n_1674, n_559, n_560);
  xor g1476 (n_563, n_1674, n_561);
  nand g1477 (n_1675, n_559, n_560);
  nand g1478 (n_1676, n_561, n_560);
  nand g1479 (n_1677, n_559, n_561);
  nand g1480 (n_578, n_1675, n_1676, n_1677);
  xor g1481 (n_1678, n_562, n_563);
  xor g1482 (n_164, n_1678, n_564);
  nand g1483 (n_1679, n_562, n_563);
  nand g1484 (n_1680, n_564, n_563);
  nand g1485 (n_1681, n_562, n_564);
  nand g1486 (n_91, n_1679, n_1680, n_1681);
  xor g1487 (n_1682, A[34], A[32]);
  xor g1488 (n_569, n_1682, A[28]);
  nand g1489 (n_1683, A[34], A[32]);
  nand g1490 (n_1684, A[28], A[32]);
  nand g1491 (n_1685, A[34], A[28]);
  nand g1492 (n_579, n_1683, n_1684, n_1685);
  xor g1494 (n_570, n_1234, A[26]);
  nand g1496 (n_1688, A[26], A[18]);
  nand g1498 (n_580, n_1235, n_1688, n_1429);
  xor g1499 (n_1690, A[16], A[30]);
  xor g1500 (n_568, n_1690, A[24]);
  nand g1501 (n_1691, A[16], A[30]);
  nand g1504 (n_581, n_1691, n_1557, n_1624);
  xor g1505 (n_1694, A[22], n_565);
  xor g1506 (n_572, n_1694, n_566);
  nand g1507 (n_1695, A[22], n_565);
  nand g1508 (n_1696, n_566, n_565);
  nand g1509 (n_1697, A[22], n_566);
  nand g1510 (n_585, n_1695, n_1696, n_1697);
  xor g1511 (n_1698, n_567, n_568);
  xor g1512 (n_574, n_1698, n_569);
  nand g1513 (n_1699, n_567, n_568);
  nand g1514 (n_1700, n_569, n_568);
  nand g1515 (n_1701, n_567, n_569);
  nand g1516 (n_587, n_1699, n_1700, n_1701);
  xor g1517 (n_1702, n_570, n_571);
  xor g1518 (n_576, n_1702, n_572);
  nand g1519 (n_1703, n_570, n_571);
  nand g1520 (n_1704, n_572, n_571);
  nand g1521 (n_1705, n_570, n_572);
  nand g1522 (n_589, n_1703, n_1704, n_1705);
  xor g1523 (n_1706, n_573, n_574);
  xor g1524 (n_577, n_1706, n_575);
  nand g1525 (n_1707, n_573, n_574);
  nand g1526 (n_1708, n_575, n_574);
  nand g1527 (n_1709, n_573, n_575);
  nand g1528 (n_592, n_1707, n_1708, n_1709);
  xor g1529 (n_1710, n_576, n_577);
  xor g1530 (n_163, n_1710, n_578);
  nand g1531 (n_1711, n_576, n_577);
  nand g1532 (n_1712, n_578, n_577);
  nand g1533 (n_1713, n_576, n_578);
  nand g1534 (n_90, n_1711, n_1712, n_1713);
  xor g1535 (n_1714, A[35], A[33]);
  xor g1536 (n_583, n_1714, A[29]);
  nand g1537 (n_1715, A[35], A[33]);
  nand g1538 (n_1716, A[29], A[33]);
  nand g1539 (n_1717, A[35], A[29]);
  nand g1540 (n_593, n_1715, n_1716, n_1717);
  xor g1542 (n_584, n_1266, A[27]);
  nand g1544 (n_1720, A[27], A[19]);
  nand g1546 (n_594, n_1267, n_1720, n_1461);
  xor g1547 (n_1722, A[17], A[31]);
  xor g1548 (n_582, n_1722, A[25]);
  nand g1549 (n_1723, A[17], A[31]);
  nand g1552 (n_595, n_1723, n_1589, n_1656);
  xor g1553 (n_1726, A[23], n_579);
  xor g1554 (n_586, n_1726, n_580);
  nand g1555 (n_1727, A[23], n_579);
  nand g1556 (n_1728, n_580, n_579);
  nand g1557 (n_1729, A[23], n_580);
  nand g1558 (n_599, n_1727, n_1728, n_1729);
  xor g1559 (n_1730, n_581, n_582);
  xor g1560 (n_588, n_1730, n_583);
  nand g1561 (n_1731, n_581, n_582);
  nand g1562 (n_1732, n_583, n_582);
  nand g1563 (n_1733, n_581, n_583);
  nand g1564 (n_601, n_1731, n_1732, n_1733);
  xor g1565 (n_1734, n_584, n_585);
  xor g1566 (n_590, n_1734, n_586);
  nand g1567 (n_1735, n_584, n_585);
  nand g1568 (n_1736, n_586, n_585);
  nand g1569 (n_1737, n_584, n_586);
  nand g1570 (n_603, n_1735, n_1736, n_1737);
  xor g1571 (n_1738, n_587, n_588);
  xor g1572 (n_591, n_1738, n_589);
  nand g1573 (n_1739, n_587, n_588);
  nand g1574 (n_1740, n_589, n_588);
  nand g1575 (n_1741, n_587, n_589);
  nand g1576 (n_606, n_1739, n_1740, n_1741);
  xor g1577 (n_1742, n_590, n_591);
  xor g1578 (n_162, n_1742, n_592);
  nand g1579 (n_1743, n_590, n_591);
  nand g1580 (n_1744, n_592, n_591);
  nand g1581 (n_1745, n_590, n_592);
  nand g1582 (n_89, n_1743, n_1744, n_1745);
  xor g1583 (n_1746, A[36], A[34]);
  xor g1584 (n_597, n_1746, A[30]);
  nand g1585 (n_1747, A[36], A[34]);
  nand g1586 (n_1748, A[30], A[34]);
  nand g1587 (n_1749, A[36], A[30]);
  nand g1588 (n_607, n_1747, n_1748, n_1749);
  xor g1590 (n_598, n_1298, A[28]);
  nand g1592 (n_1752, A[28], A[20]);
  nand g1594 (n_608, n_1299, n_1752, n_1493);
  xor g1595 (n_1754, A[18], A[32]);
  xor g1596 (n_596, n_1754, A[26]);
  nand g1597 (n_1755, A[18], A[32]);
  nand g1600 (n_609, n_1755, n_1621, n_1688);
  xor g1601 (n_1758, A[24], n_593);
  xor g1602 (n_600, n_1758, n_594);
  nand g1603 (n_1759, A[24], n_593);
  nand g1604 (n_1760, n_594, n_593);
  nand g1605 (n_1761, A[24], n_594);
  nand g1606 (n_613, n_1759, n_1760, n_1761);
  xor g1607 (n_1762, n_595, n_596);
  xor g1608 (n_602, n_1762, n_597);
  nand g1609 (n_1763, n_595, n_596);
  nand g1610 (n_1764, n_597, n_596);
  nand g1611 (n_1765, n_595, n_597);
  nand g1612 (n_615, n_1763, n_1764, n_1765);
  xor g1613 (n_1766, n_598, n_599);
  xor g1614 (n_604, n_1766, n_600);
  nand g1615 (n_1767, n_598, n_599);
  nand g1616 (n_1768, n_600, n_599);
  nand g1617 (n_1769, n_598, n_600);
  nand g1618 (n_617, n_1767, n_1768, n_1769);
  xor g1619 (n_1770, n_601, n_602);
  xor g1620 (n_605, n_1770, n_603);
  nand g1621 (n_1771, n_601, n_602);
  nand g1622 (n_1772, n_603, n_602);
  nand g1623 (n_1773, n_601, n_603);
  nand g1624 (n_620, n_1771, n_1772, n_1773);
  xor g1625 (n_1774, n_604, n_605);
  xor g1626 (n_161, n_1774, n_606);
  nand g1627 (n_1775, n_604, n_605);
  nand g1628 (n_1776, n_606, n_605);
  nand g1629 (n_1777, n_604, n_606);
  nand g1630 (n_88, n_1775, n_1776, n_1777);
  xor g1631 (n_1778, A[37], A[35]);
  xor g1632 (n_611, n_1778, A[31]);
  nand g1633 (n_1779, A[37], A[35]);
  nand g1634 (n_1780, A[31], A[35]);
  nand g1635 (n_1781, A[37], A[31]);
  nand g1636 (n_621, n_1779, n_1780, n_1781);
  xor g1638 (n_612, n_1330, A[29]);
  nand g1640 (n_1784, A[29], A[21]);
  nand g1642 (n_622, n_1331, n_1784, n_1525);
  xor g1643 (n_1786, A[19], A[33]);
  xor g1644 (n_610, n_1786, A[27]);
  nand g1645 (n_1787, A[19], A[33]);
  nand g1648 (n_623, n_1787, n_1653, n_1720);
  xor g1649 (n_1790, A[25], n_607);
  xor g1650 (n_614, n_1790, n_608);
  nand g1651 (n_1791, A[25], n_607);
  nand g1652 (n_1792, n_608, n_607);
  nand g1653 (n_1793, A[25], n_608);
  nand g1654 (n_627, n_1791, n_1792, n_1793);
  xor g1655 (n_1794, n_609, n_610);
  xor g1656 (n_616, n_1794, n_611);
  nand g1657 (n_1795, n_609, n_610);
  nand g1658 (n_1796, n_611, n_610);
  nand g1659 (n_1797, n_609, n_611);
  nand g1660 (n_629, n_1795, n_1796, n_1797);
  xor g1661 (n_1798, n_612, n_613);
  xor g1662 (n_618, n_1798, n_614);
  nand g1663 (n_1799, n_612, n_613);
  nand g1664 (n_1800, n_614, n_613);
  nand g1665 (n_1801, n_612, n_614);
  nand g1666 (n_631, n_1799, n_1800, n_1801);
  xor g1667 (n_1802, n_615, n_616);
  xor g1668 (n_619, n_1802, n_617);
  nand g1669 (n_1803, n_615, n_616);
  nand g1670 (n_1804, n_617, n_616);
  nand g1671 (n_1805, n_615, n_617);
  nand g1672 (n_634, n_1803, n_1804, n_1805);
  xor g1673 (n_1806, n_618, n_619);
  xor g1674 (n_160, n_1806, n_620);
  nand g1675 (n_1807, n_618, n_619);
  nand g1676 (n_1808, n_620, n_619);
  nand g1677 (n_1809, n_618, n_620);
  nand g1678 (n_87, n_1807, n_1808, n_1809);
  xor g1679 (n_1810, A[38], A[36]);
  xor g1680 (n_625, n_1810, A[32]);
  nand g1681 (n_1811, A[38], A[36]);
  nand g1682 (n_1812, A[32], A[36]);
  nand g1683 (n_1813, A[38], A[32]);
  nand g1684 (n_635, n_1811, n_1812, n_1813);
  xor g1686 (n_626, n_1362, A[30]);
  nand g1688 (n_1816, A[30], A[22]);
  nand g1690 (n_636, n_1363, n_1816, n_1557);
  xor g1691 (n_1818, A[20], A[34]);
  xor g1692 (n_624, n_1818, A[28]);
  nand g1693 (n_1819, A[20], A[34]);
  nand g1696 (n_637, n_1819, n_1685, n_1752);
  xor g1697 (n_1822, A[26], n_621);
  xor g1698 (n_628, n_1822, n_622);
  nand g1699 (n_1823, A[26], n_621);
  nand g1700 (n_1824, n_622, n_621);
  nand g1701 (n_1825, A[26], n_622);
  nand g1702 (n_641, n_1823, n_1824, n_1825);
  xor g1703 (n_1826, n_623, n_624);
  xor g1704 (n_630, n_1826, n_625);
  nand g1705 (n_1827, n_623, n_624);
  nand g1706 (n_1828, n_625, n_624);
  nand g1707 (n_1829, n_623, n_625);
  nand g1708 (n_643, n_1827, n_1828, n_1829);
  xor g1709 (n_1830, n_626, n_627);
  xor g1710 (n_632, n_1830, n_628);
  nand g1711 (n_1831, n_626, n_627);
  nand g1712 (n_1832, n_628, n_627);
  nand g1713 (n_1833, n_626, n_628);
  nand g1714 (n_645, n_1831, n_1832, n_1833);
  xor g1715 (n_1834, n_629, n_630);
  xor g1716 (n_633, n_1834, n_631);
  nand g1717 (n_1835, n_629, n_630);
  nand g1718 (n_1836, n_631, n_630);
  nand g1719 (n_1837, n_629, n_631);
  nand g1720 (n_648, n_1835, n_1836, n_1837);
  xor g1721 (n_1838, n_632, n_633);
  xor g1722 (n_159, n_1838, n_634);
  nand g1723 (n_1839, n_632, n_633);
  nand g1724 (n_1840, n_634, n_633);
  nand g1725 (n_1841, n_632, n_634);
  nand g1726 (n_86, n_1839, n_1840, n_1841);
  xor g1727 (n_1842, A[39], A[37]);
  xor g1728 (n_639, n_1842, A[33]);
  nand g1729 (n_1843, A[39], A[37]);
  nand g1730 (n_1844, A[33], A[37]);
  nand g1731 (n_1845, A[39], A[33]);
  nand g1732 (n_649, n_1843, n_1844, n_1845);
  xor g1734 (n_640, n_1394, A[31]);
  nand g1736 (n_1848, A[31], A[23]);
  nand g1738 (n_650, n_1395, n_1848, n_1589);
  xor g1739 (n_1850, A[21], A[35]);
  xor g1740 (n_638, n_1850, A[29]);
  nand g1741 (n_1851, A[21], A[35]);
  nand g1744 (n_651, n_1851, n_1717, n_1784);
  xor g1745 (n_1854, A[27], n_635);
  xor g1746 (n_642, n_1854, n_636);
  nand g1747 (n_1855, A[27], n_635);
  nand g1748 (n_1856, n_636, n_635);
  nand g1749 (n_1857, A[27], n_636);
  nand g1750 (n_655, n_1855, n_1856, n_1857);
  xor g1751 (n_1858, n_637, n_638);
  xor g1752 (n_644, n_1858, n_639);
  nand g1753 (n_1859, n_637, n_638);
  nand g1754 (n_1860, n_639, n_638);
  nand g1755 (n_1861, n_637, n_639);
  nand g1756 (n_657, n_1859, n_1860, n_1861);
  xor g1757 (n_1862, n_640, n_641);
  xor g1758 (n_646, n_1862, n_642);
  nand g1759 (n_1863, n_640, n_641);
  nand g1760 (n_1864, n_642, n_641);
  nand g1761 (n_1865, n_640, n_642);
  nand g1762 (n_659, n_1863, n_1864, n_1865);
  xor g1763 (n_1866, n_643, n_644);
  xor g1764 (n_647, n_1866, n_645);
  nand g1765 (n_1867, n_643, n_644);
  nand g1766 (n_1868, n_645, n_644);
  nand g1767 (n_1869, n_643, n_645);
  nand g1768 (n_662, n_1867, n_1868, n_1869);
  xor g1769 (n_1870, n_646, n_647);
  xor g1770 (n_158, n_1870, n_648);
  nand g1771 (n_1871, n_646, n_647);
  nand g1772 (n_1872, n_648, n_647);
  nand g1773 (n_1873, n_646, n_648);
  nand g1774 (n_85, n_1871, n_1872, n_1873);
  xor g1775 (n_1874, A[40], A[38]);
  xor g1776 (n_653, n_1874, A[34]);
  nand g1777 (n_1875, A[40], A[38]);
  nand g1778 (n_1876, A[34], A[38]);
  nand g1779 (n_1877, A[40], A[34]);
  nand g1780 (n_663, n_1875, n_1876, n_1877);
  xor g1782 (n_654, n_1426, A[32]);
  nand g1784 (n_1880, A[32], A[24]);
  nand g1786 (n_664, n_1427, n_1880, n_1621);
  xor g1787 (n_1882, A[22], A[36]);
  xor g1788 (n_652, n_1882, A[30]);
  nand g1789 (n_1883, A[22], A[36]);
  nand g1792 (n_665, n_1883, n_1749, n_1816);
  xor g1793 (n_1886, A[28], n_649);
  xor g1794 (n_656, n_1886, n_650);
  nand g1795 (n_1887, A[28], n_649);
  nand g1796 (n_1888, n_650, n_649);
  nand g1797 (n_1889, A[28], n_650);
  nand g1798 (n_669, n_1887, n_1888, n_1889);
  xor g1799 (n_1890, n_651, n_652);
  xor g1800 (n_658, n_1890, n_653);
  nand g1801 (n_1891, n_651, n_652);
  nand g1802 (n_1892, n_653, n_652);
  nand g1803 (n_1893, n_651, n_653);
  nand g1804 (n_671, n_1891, n_1892, n_1893);
  xor g1805 (n_1894, n_654, n_655);
  xor g1806 (n_660, n_1894, n_656);
  nand g1807 (n_1895, n_654, n_655);
  nand g1808 (n_1896, n_656, n_655);
  nand g1809 (n_1897, n_654, n_656);
  nand g1810 (n_673, n_1895, n_1896, n_1897);
  xor g1811 (n_1898, n_657, n_658);
  xor g1812 (n_661, n_1898, n_659);
  nand g1813 (n_1899, n_657, n_658);
  nand g1814 (n_1900, n_659, n_658);
  nand g1815 (n_1901, n_657, n_659);
  nand g1816 (n_676, n_1899, n_1900, n_1901);
  xor g1817 (n_1902, n_660, n_661);
  xor g1818 (n_157, n_1902, n_662);
  nand g1819 (n_1903, n_660, n_661);
  nand g1820 (n_1904, n_662, n_661);
  nand g1821 (n_1905, n_660, n_662);
  nand g1822 (n_84, n_1903, n_1904, n_1905);
  xor g1823 (n_1906, A[41], A[39]);
  xor g1824 (n_667, n_1906, A[35]);
  nand g1825 (n_1907, A[41], A[39]);
  nand g1826 (n_1908, A[35], A[39]);
  nand g1827 (n_1909, A[41], A[35]);
  nand g1828 (n_677, n_1907, n_1908, n_1909);
  xor g1830 (n_668, n_1458, A[33]);
  nand g1832 (n_1912, A[33], A[25]);
  nand g1834 (n_678, n_1459, n_1912, n_1653);
  xor g1835 (n_1914, A[23], A[37]);
  xor g1836 (n_666, n_1914, A[31]);
  nand g1837 (n_1915, A[23], A[37]);
  nand g1840 (n_679, n_1915, n_1781, n_1848);
  xor g1841 (n_1918, A[29], n_663);
  xor g1842 (n_670, n_1918, n_664);
  nand g1843 (n_1919, A[29], n_663);
  nand g1844 (n_1920, n_664, n_663);
  nand g1845 (n_1921, A[29], n_664);
  nand g1846 (n_683, n_1919, n_1920, n_1921);
  xor g1847 (n_1922, n_665, n_666);
  xor g1848 (n_672, n_1922, n_667);
  nand g1849 (n_1923, n_665, n_666);
  nand g1850 (n_1924, n_667, n_666);
  nand g1851 (n_1925, n_665, n_667);
  nand g1852 (n_685, n_1923, n_1924, n_1925);
  xor g1853 (n_1926, n_668, n_669);
  xor g1854 (n_674, n_1926, n_670);
  nand g1855 (n_1927, n_668, n_669);
  nand g1856 (n_1928, n_670, n_669);
  nand g1857 (n_1929, n_668, n_670);
  nand g1858 (n_687, n_1927, n_1928, n_1929);
  xor g1859 (n_1930, n_671, n_672);
  xor g1860 (n_675, n_1930, n_673);
  nand g1861 (n_1931, n_671, n_672);
  nand g1862 (n_1932, n_673, n_672);
  nand g1863 (n_1933, n_671, n_673);
  nand g1864 (n_690, n_1931, n_1932, n_1933);
  xor g1865 (n_1934, n_674, n_675);
  xor g1866 (n_156, n_1934, n_676);
  nand g1867 (n_1935, n_674, n_675);
  nand g1868 (n_1936, n_676, n_675);
  nand g1869 (n_1937, n_674, n_676);
  nand g1870 (n_83, n_1935, n_1936, n_1937);
  xor g1871 (n_1938, A[42], A[40]);
  xor g1872 (n_681, n_1938, A[36]);
  nand g1873 (n_1939, A[42], A[40]);
  nand g1874 (n_1940, A[36], A[40]);
  nand g1875 (n_1941, A[42], A[36]);
  nand g1876 (n_691, n_1939, n_1940, n_1941);
  xor g1878 (n_682, n_1490, A[34]);
  nand g1880 (n_1944, A[34], A[26]);
  nand g1882 (n_692, n_1491, n_1944, n_1685);
  xor g1883 (n_1946, A[24], A[38]);
  xor g1884 (n_680, n_1946, A[32]);
  nand g1885 (n_1947, A[24], A[38]);
  nand g1888 (n_693, n_1947, n_1813, n_1880);
  xor g1889 (n_1950, A[30], n_677);
  xor g1890 (n_684, n_1950, n_678);
  nand g1891 (n_1951, A[30], n_677);
  nand g1892 (n_1952, n_678, n_677);
  nand g1893 (n_1953, A[30], n_678);
  nand g1894 (n_697, n_1951, n_1952, n_1953);
  xor g1895 (n_1954, n_679, n_680);
  xor g1896 (n_686, n_1954, n_681);
  nand g1897 (n_1955, n_679, n_680);
  nand g1898 (n_1956, n_681, n_680);
  nand g1899 (n_1957, n_679, n_681);
  nand g1900 (n_699, n_1955, n_1956, n_1957);
  xor g1901 (n_1958, n_682, n_683);
  xor g1902 (n_688, n_1958, n_684);
  nand g1903 (n_1959, n_682, n_683);
  nand g1904 (n_1960, n_684, n_683);
  nand g1905 (n_1961, n_682, n_684);
  nand g1906 (n_701, n_1959, n_1960, n_1961);
  xor g1907 (n_1962, n_685, n_686);
  xor g1908 (n_689, n_1962, n_687);
  nand g1909 (n_1963, n_685, n_686);
  nand g1910 (n_1964, n_687, n_686);
  nand g1911 (n_1965, n_685, n_687);
  nand g1912 (n_704, n_1963, n_1964, n_1965);
  xor g1913 (n_1966, n_688, n_689);
  xor g1914 (n_155, n_1966, n_690);
  nand g1915 (n_1967, n_688, n_689);
  nand g1916 (n_1968, n_690, n_689);
  nand g1917 (n_1969, n_688, n_690);
  nand g1918 (n_82, n_1967, n_1968, n_1969);
  xor g1919 (n_1970, A[43], A[41]);
  xor g1920 (n_695, n_1970, A[37]);
  nand g1921 (n_1971, A[43], A[41]);
  nand g1922 (n_1972, A[37], A[41]);
  nand g1923 (n_1973, A[43], A[37]);
  nand g1924 (n_705, n_1971, n_1972, n_1973);
  xor g1926 (n_696, n_1522, A[35]);
  nand g1928 (n_1976, A[35], A[27]);
  nand g1930 (n_707, n_1523, n_1976, n_1717);
  xor g1931 (n_1978, A[25], A[39]);
  xor g1932 (n_694, n_1978, A[33]);
  nand g1933 (n_1979, A[25], A[39]);
  nand g1936 (n_706, n_1979, n_1845, n_1912);
  xor g1937 (n_1982, A[31], n_691);
  xor g1938 (n_698, n_1982, n_692);
  nand g1939 (n_1983, A[31], n_691);
  nand g1940 (n_1984, n_692, n_691);
  nand g1941 (n_1985, A[31], n_692);
  nand g1942 (n_711, n_1983, n_1984, n_1985);
  xor g1943 (n_1986, n_693, n_694);
  xor g1944 (n_700, n_1986, n_695);
  nand g1945 (n_1987, n_693, n_694);
  nand g1946 (n_1988, n_695, n_694);
  nand g1947 (n_1989, n_693, n_695);
  nand g1948 (n_713, n_1987, n_1988, n_1989);
  xor g1949 (n_1990, n_696, n_697);
  xor g1950 (n_702, n_1990, n_698);
  nand g1951 (n_1991, n_696, n_697);
  nand g1952 (n_1992, n_698, n_697);
  nand g1953 (n_1993, n_696, n_698);
  nand g1954 (n_716, n_1991, n_1992, n_1993);
  xor g1955 (n_1994, n_699, n_700);
  xor g1956 (n_703, n_1994, n_701);
  nand g1957 (n_1995, n_699, n_700);
  nand g1958 (n_1996, n_701, n_700);
  nand g1959 (n_1997, n_699, n_701);
  nand g1960 (n_718, n_1995, n_1996, n_1997);
  xor g1961 (n_1998, n_702, n_703);
  xor g1962 (n_154, n_1998, n_704);
  nand g1963 (n_1999, n_702, n_703);
  nand g1964 (n_2000, n_704, n_703);
  nand g1965 (n_2001, n_702, n_704);
  nand g1966 (n_81, n_1999, n_2000, n_2001);
  xor g1967 (n_2002, A[42], A[38]);
  xor g1968 (n_709, n_2002, A[30]);
  nand g1969 (n_2003, A[42], A[38]);
  nand g1970 (n_2004, A[30], A[38]);
  nand g1971 (n_2005, A[42], A[30]);
  nand g1972 (n_719, n_2003, n_2004, n_2005);
  xor g1973 (n_2006, A[28], A[36]);
  xor g1974 (n_710, n_2006, A[26]);
  nand g1975 (n_2007, A[28], A[36]);
  nand g1976 (n_2008, A[26], A[36]);
  nand g1978 (n_721, n_2007, n_2008, n_1491);
  xor g1979 (n_2010, A[40], A[34]);
  xor g1980 (n_708, n_2010, A[32]);
  nand g1983 (n_2013, A[40], A[32]);
  nand g1984 (n_720, n_1877, n_1683, n_2013);
  xor g1985 (n_2014, A[44], n_705);
  xor g1986 (n_712, n_2014, n_706);
  nand g1987 (n_2015, A[44], n_705);
  nand g1988 (n_2016, n_706, n_705);
  nand g1989 (n_2017, A[44], n_706);
  nand g1990 (n_725, n_2015, n_2016, n_2017);
  xor g1991 (n_2018, n_707, n_708);
  xor g1992 (n_714, n_2018, n_709);
  nand g1993 (n_2019, n_707, n_708);
  nand g1994 (n_2020, n_709, n_708);
  nand g1995 (n_2021, n_707, n_709);
  nand g1996 (n_727, n_2019, n_2020, n_2021);
  xor g1997 (n_2022, n_710, n_711);
  xor g1998 (n_715, n_2022, n_712);
  nand g1999 (n_2023, n_710, n_711);
  nand g2000 (n_2024, n_712, n_711);
  nand g2001 (n_2025, n_710, n_712);
  nand g2002 (n_730, n_2023, n_2024, n_2025);
  xor g2003 (n_2026, n_713, n_714);
  xor g2004 (n_717, n_2026, n_715);
  nand g2005 (n_2027, n_713, n_714);
  nand g2006 (n_2028, n_715, n_714);
  nand g2007 (n_2029, n_713, n_715);
  nand g2008 (n_732, n_2027, n_2028, n_2029);
  xor g2009 (n_2030, n_716, n_717);
  xor g2010 (n_153, n_2030, n_718);
  nand g2011 (n_2031, n_716, n_717);
  nand g2012 (n_2032, n_718, n_717);
  nand g2013 (n_2033, n_716, n_718);
  nand g2014 (n_80, n_2031, n_2032, n_2033);
  xor g2015 (n_2034, A[43], A[39]);
  xor g2016 (n_723, n_2034, A[31]);
  nand g2017 (n_2035, A[43], A[39]);
  nand g2018 (n_2036, A[31], A[39]);
  nand g2019 (n_2037, A[43], A[31]);
  nand g2020 (n_734, n_2035, n_2036, n_2037);
  xor g2021 (n_2038, A[29], A[37]);
  xor g2022 (n_724, n_2038, A[27]);
  nand g2023 (n_2039, A[29], A[37]);
  nand g2024 (n_2040, A[27], A[37]);
  nand g2026 (n_735, n_2039, n_2040, n_1523);
  xor g2027 (n_2042, A[41], A[35]);
  xor g2028 (n_722, n_2042, A[33]);
  nand g2031 (n_2045, A[41], A[33]);
  nand g2032 (n_733, n_1909, n_1715, n_2045);
  xor g2033 (n_2046, A[45], n_719);
  xor g2034 (n_726, n_2046, n_720);
  nand g2035 (n_2047, A[45], n_719);
  nand g2036 (n_2048, n_720, n_719);
  nand g2037 (n_2049, A[45], n_720);
  nand g2038 (n_739, n_2047, n_2048, n_2049);
  xor g2039 (n_2050, n_721, n_722);
  xor g2040 (n_728, n_2050, n_723);
  nand g2041 (n_2051, n_721, n_722);
  nand g2042 (n_2052, n_723, n_722);
  nand g2043 (n_2053, n_721, n_723);
  nand g2044 (n_740, n_2051, n_2052, n_2053);
  xor g2045 (n_2054, n_724, n_725);
  xor g2046 (n_729, n_2054, n_726);
  nand g2047 (n_2055, n_724, n_725);
  nand g2048 (n_2056, n_726, n_725);
  nand g2049 (n_2057, n_724, n_726);
  nand g2050 (n_744, n_2055, n_2056, n_2057);
  xor g2051 (n_2058, n_727, n_728);
  xor g2052 (n_731, n_2058, n_729);
  nand g2053 (n_2059, n_727, n_728);
  nand g2054 (n_2060, n_729, n_728);
  nand g2055 (n_2061, n_727, n_729);
  nand g2056 (n_746, n_2059, n_2060, n_2061);
  xor g2057 (n_2062, n_730, n_731);
  xor g2058 (n_152, n_2062, n_732);
  nand g2059 (n_2063, n_730, n_731);
  nand g2060 (n_2064, n_732, n_731);
  nand g2061 (n_2065, n_730, n_732);
  nand g2062 (n_79, n_2063, n_2064, n_2065);
  xor g2064 (n_736, n_1938, A[32]);
  nand g2067 (n_2069, A[42], A[32]);
  nand g2068 (n_747, n_1939, n_2013, n_2069);
  xor g2069 (n_2070, A[30], A[38]);
  xor g2070 (n_738, n_2070, A[28]);
  nand g2072 (n_2072, A[28], A[38]);
  nand g2074 (n_748, n_2004, n_2072, n_1555);
  xor g2076 (n_737, n_1746, A[44]);
  nand g2078 (n_2076, A[44], A[34]);
  nand g2079 (n_2077, A[36], A[44]);
  nand g2080 (n_750, n_1747, n_2076, n_2077);
  xor g2081 (n_2078, A[46], n_733);
  xor g2082 (n_741, n_2078, n_734);
  nand g2083 (n_2079, A[46], n_733);
  nand g2084 (n_2080, n_734, n_733);
  nand g2085 (n_2081, A[46], n_734);
  nand g2086 (n_753, n_2079, n_2080, n_2081);
  xor g2087 (n_2082, n_735, n_736);
  xor g2088 (n_742, n_2082, n_737);
  nand g2089 (n_2083, n_735, n_736);
  nand g2090 (n_2084, n_737, n_736);
  nand g2091 (n_2085, n_735, n_737);
  nand g2092 (n_754, n_2083, n_2084, n_2085);
  xor g2093 (n_2086, n_738, n_739);
  xor g2094 (n_743, n_2086, n_740);
  nand g2095 (n_2087, n_738, n_739);
  nand g2096 (n_2088, n_740, n_739);
  nand g2097 (n_2089, n_738, n_740);
  nand g2098 (n_758, n_2087, n_2088, n_2089);
  xor g2099 (n_2090, n_741, n_742);
  xor g2100 (n_745, n_2090, n_743);
  nand g2101 (n_2091, n_741, n_742);
  nand g2102 (n_2092, n_743, n_742);
  nand g2103 (n_2093, n_741, n_743);
  nand g2104 (n_760, n_2091, n_2092, n_2093);
  xor g2105 (n_2094, n_744, n_745);
  xor g2106 (n_151, n_2094, n_746);
  nand g2107 (n_2095, n_744, n_745);
  nand g2108 (n_2096, n_746, n_745);
  nand g2109 (n_2097, n_744, n_746);
  nand g2110 (n_78, n_2095, n_2096, n_2097);
  xor g2112 (n_749, n_1970, A[33]);
  nand g2115 (n_2101, A[43], A[33]);
  nand g2116 (n_761, n_1971, n_2045, n_2101);
  xor g2117 (n_2102, A[31], A[39]);
  xor g2118 (n_752, n_2102, A[29]);
  nand g2120 (n_2104, A[29], A[39]);
  nand g2122 (n_762, n_2036, n_2104, n_1587);
  xor g2124 (n_751, n_1778, A[45]);
  nand g2126 (n_2108, A[45], A[35]);
  nand g2127 (n_2109, A[37], A[45]);
  nand g2128 (n_764, n_1779, n_2108, n_2109);
  xor g2129 (n_2110, A[47], n_747);
  xor g2130 (n_755, n_2110, n_748);
  nand g2131 (n_2111, A[47], n_747);
  nand g2132 (n_2112, n_748, n_747);
  nand g2133 (n_2113, A[47], n_748);
  nand g2134 (n_767, n_2111, n_2112, n_2113);
  xor g2135 (n_2114, n_749, n_750);
  xor g2136 (n_756, n_2114, n_751);
  nand g2137 (n_2115, n_749, n_750);
  nand g2138 (n_2116, n_751, n_750);
  nand g2139 (n_2117, n_749, n_751);
  nand g2140 (n_768, n_2115, n_2116, n_2117);
  xor g2141 (n_2118, n_752, n_753);
  xor g2142 (n_757, n_2118, n_754);
  nand g2143 (n_2119, n_752, n_753);
  nand g2144 (n_2120, n_754, n_753);
  nand g2145 (n_2121, n_752, n_754);
  nand g2146 (n_772, n_2119, n_2120, n_2121);
  xor g2147 (n_2122, n_755, n_756);
  xor g2148 (n_759, n_2122, n_757);
  nand g2149 (n_2123, n_755, n_756);
  nand g2150 (n_2124, n_757, n_756);
  nand g2151 (n_2125, n_755, n_757);
  nand g2152 (n_774, n_2123, n_2124, n_2125);
  xor g2153 (n_2126, n_758, n_759);
  xor g2154 (n_150, n_2126, n_760);
  nand g2155 (n_2127, n_758, n_759);
  nand g2156 (n_2128, n_760, n_759);
  nand g2157 (n_2129, n_758, n_760);
  nand g2158 (n_77, n_2127, n_2128, n_2129);
  xor g2160 (n_763, n_1938, A[34]);
  nand g2163 (n_2133, A[42], A[34]);
  nand g2164 (n_775, n_1939, n_1877, n_2133);
  xor g2166 (n_765, n_1618, A[38]);
  nand g2170 (n_776, n_1619, n_2004, n_1813);
  xor g2171 (n_2138, A[36], A[46]);
  xor g2172 (n_766, n_2138, A[48]);
  nand g2173 (n_2139, A[36], A[46]);
  nand g2174 (n_2140, A[48], A[46]);
  nand g2175 (n_2141, A[36], A[48]);
  nand g2176 (n_778, n_2139, n_2140, n_2141);
  xor g2177 (n_2142, A[44], n_761);
  xor g2178 (n_769, n_2142, n_762);
  nand g2179 (n_2143, A[44], n_761);
  nand g2180 (n_2144, n_762, n_761);
  nand g2181 (n_2145, A[44], n_762);
  nand g2182 (n_781, n_2143, n_2144, n_2145);
  xor g2183 (n_2146, n_763, n_764);
  xor g2184 (n_770, n_2146, n_765);
  nand g2185 (n_2147, n_763, n_764);
  nand g2186 (n_2148, n_765, n_764);
  nand g2187 (n_2149, n_763, n_765);
  nand g2188 (n_782, n_2147, n_2148, n_2149);
  xor g2189 (n_2150, n_766, n_767);
  xor g2190 (n_771, n_2150, n_768);
  nand g2191 (n_2151, n_766, n_767);
  nand g2192 (n_2152, n_768, n_767);
  nand g2193 (n_2153, n_766, n_768);
  nand g2194 (n_786, n_2151, n_2152, n_2153);
  xor g2195 (n_2154, n_769, n_770);
  xor g2196 (n_773, n_2154, n_771);
  nand g2197 (n_2155, n_769, n_770);
  nand g2198 (n_2156, n_771, n_770);
  nand g2199 (n_2157, n_769, n_771);
  nand g2200 (n_788, n_2155, n_2156, n_2157);
  xor g2201 (n_2158, n_772, n_773);
  xor g2202 (n_149, n_2158, n_774);
  nand g2203 (n_2159, n_772, n_773);
  nand g2204 (n_2160, n_774, n_773);
  nand g2205 (n_2161, n_772, n_774);
  nand g2206 (n_76, n_2159, n_2160, n_2161);
  xor g2208 (n_777, n_1970, A[35]);
  nand g2211 (n_2165, A[43], A[35]);
  nand g2212 (n_789, n_1971, n_1909, n_2165);
  xor g2214 (n_779, n_1650, A[39]);
  nand g2218 (n_790, n_1651, n_2036, n_1845);
  xor g2219 (n_2170, A[37], A[47]);
  xor g2220 (n_780, n_2170, A[49]);
  nand g2221 (n_2171, A[37], A[47]);
  nand g2222 (n_2172, A[49], A[47]);
  nand g2223 (n_2173, A[37], A[49]);
  nand g2224 (n_792, n_2171, n_2172, n_2173);
  xor g2225 (n_2174, A[45], n_775);
  xor g2226 (n_783, n_2174, n_776);
  nand g2227 (n_2175, A[45], n_775);
  nand g2228 (n_2176, n_776, n_775);
  nand g2229 (n_2177, A[45], n_776);
  nand g2230 (n_795, n_2175, n_2176, n_2177);
  xor g2231 (n_2178, n_777, n_778);
  xor g2232 (n_784, n_2178, n_779);
  nand g2233 (n_2179, n_777, n_778);
  nand g2234 (n_2180, n_779, n_778);
  nand g2235 (n_2181, n_777, n_779);
  nand g2236 (n_796, n_2179, n_2180, n_2181);
  xor g2237 (n_2182, n_780, n_781);
  xor g2238 (n_785, n_2182, n_782);
  nand g2239 (n_2183, n_780, n_781);
  nand g2240 (n_2184, n_782, n_781);
  nand g2241 (n_2185, n_780, n_782);
  nand g2242 (n_800, n_2183, n_2184, n_2185);
  xor g2243 (n_2186, n_783, n_784);
  xor g2244 (n_787, n_2186, n_785);
  nand g2245 (n_2187, n_783, n_784);
  nand g2246 (n_2188, n_785, n_784);
  nand g2247 (n_2189, n_783, n_785);
  nand g2248 (n_802, n_2187, n_2188, n_2189);
  xor g2249 (n_2190, n_786, n_787);
  xor g2250 (n_148, n_2190, n_788);
  nand g2251 (n_2191, n_786, n_787);
  nand g2252 (n_2192, n_788, n_787);
  nand g2253 (n_2193, n_786, n_788);
  nand g2254 (n_75, n_2191, n_2192, n_2193);
  xor g2255 (n_2194, A[42], A[36]);
  xor g2256 (n_791, n_2194, A[34]);
  nand g2260 (n_803, n_1941, n_1747, n_2133);
  xor g2261 (n_2198, A[32], A[40]);
  xor g2262 (n_793, n_2198, A[38]);
  nand g2266 (n_804, n_2013, n_1875, n_1813);
  xor g2267 (n_2202, A[44], A[50]);
  xor g2268 (n_794, n_2202, A[48]);
  nand g2269 (n_2203, A[44], A[50]);
  nand g2270 (n_2204, A[48], A[50]);
  nand g2271 (n_2205, A[44], A[48]);
  nand g2272 (n_806, n_2203, n_2204, n_2205);
  xor g2273 (n_2206, A[46], n_789);
  xor g2274 (n_797, n_2206, n_790);
  nand g2275 (n_2207, A[46], n_789);
  nand g2276 (n_2208, n_790, n_789);
  nand g2277 (n_2209, A[46], n_790);
  nand g2278 (n_809, n_2207, n_2208, n_2209);
  xor g2279 (n_2210, n_791, n_792);
  xor g2280 (n_798, n_2210, n_793);
  nand g2281 (n_2211, n_791, n_792);
  nand g2282 (n_2212, n_793, n_792);
  nand g2283 (n_2213, n_791, n_793);
  nand g2284 (n_810, n_2211, n_2212, n_2213);
  xor g2285 (n_2214, n_794, n_795);
  xor g2286 (n_799, n_2214, n_796);
  nand g2287 (n_2215, n_794, n_795);
  nand g2288 (n_2216, n_796, n_795);
  nand g2289 (n_2217, n_794, n_796);
  nand g2290 (n_814, n_2215, n_2216, n_2217);
  xor g2291 (n_2218, n_797, n_798);
  xor g2292 (n_801, n_2218, n_799);
  nand g2293 (n_2219, n_797, n_798);
  nand g2294 (n_2220, n_799, n_798);
  nand g2295 (n_2221, n_797, n_799);
  nand g2296 (n_816, n_2219, n_2220, n_2221);
  xor g2297 (n_2222, n_800, n_801);
  xor g2298 (n_147, n_2222, n_802);
  nand g2299 (n_2223, n_800, n_801);
  nand g2300 (n_2224, n_802, n_801);
  nand g2301 (n_2225, n_800, n_802);
  nand g2302 (n_74, n_2223, n_2224, n_2225);
  xor g2303 (n_2226, A[43], A[37]);
  xor g2304 (n_805, n_2226, A[35]);
  nand g2308 (n_820, n_1973, n_1779, n_2165);
  xor g2309 (n_2230, A[33], A[41]);
  xor g2310 (n_807, n_2230, A[39]);
  nand g2314 (n_819, n_2045, n_1907, n_1845);
  xor g2315 (n_2234, A[45], A[51]);
  xor g2316 (n_808, n_2234, A[49]);
  nand g2317 (n_2235, A[45], A[51]);
  nand g2318 (n_2236, A[49], A[51]);
  nand g2319 (n_2237, A[45], A[49]);
  nand g2320 (n_823, n_2235, n_2236, n_2237);
  xor g2321 (n_2238, A[47], n_803);
  xor g2322 (n_811, n_2238, n_804);
  nand g2323 (n_2239, A[47], n_803);
  nand g2324 (n_2240, n_804, n_803);
  nand g2325 (n_2241, A[47], n_804);
  nand g2326 (n_825, n_2239, n_2240, n_2241);
  xor g2327 (n_2242, n_805, n_806);
  xor g2328 (n_812, n_2242, n_807);
  nand g2329 (n_2243, n_805, n_806);
  nand g2330 (n_2244, n_807, n_806);
  nand g2331 (n_2245, n_805, n_807);
  nand g2332 (n_826, n_2243, n_2244, n_2245);
  xor g2333 (n_2246, n_808, n_809);
  xor g2334 (n_813, n_2246, n_810);
  nand g2335 (n_2247, n_808, n_809);
  nand g2336 (n_2248, n_810, n_809);
  nand g2337 (n_2249, n_808, n_810);
  nand g2338 (n_830, n_2247, n_2248, n_2249);
  xor g2339 (n_2250, n_811, n_812);
  xor g2340 (n_815, n_2250, n_813);
  nand g2341 (n_2251, n_811, n_812);
  nand g2342 (n_2252, n_813, n_812);
  nand g2343 (n_2253, n_811, n_813);
  nand g2344 (n_832, n_2251, n_2252, n_2253);
  xor g2345 (n_2254, n_814, n_815);
  xor g2346 (n_146, n_2254, n_816);
  nand g2347 (n_2255, n_814, n_815);
  nand g2348 (n_2256, n_816, n_815);
  nand g2349 (n_2257, n_814, n_816);
  nand g2350 (n_73, n_2255, n_2256, n_2257);
  xor g2353 (n_2258, A[52], A[36]);
  xor g2354 (n_821, n_2258, A[38]);
  nand g2355 (n_2259, A[52], A[36]);
  nand g2357 (n_2261, A[52], A[38]);
  nand g2358 (n_837, n_2259, n_1811, n_2261);
  xor g2359 (n_2262, A[34], A[42]);
  xor g2360 (n_822, n_2262, A[40]);
  xor g2365 (n_2266, A[50], A[46]);
  xor g2366 (n_824, n_2266, A[44]);
  nand g2367 (n_2267, A[50], A[46]);
  nand g2368 (n_2268, A[44], A[46]);
  nand g2370 (n_840, n_2267, n_2268, n_2203);
  xor g2371 (n_2270, A[48], n_819);
  xor g2372 (n_827, n_2270, n_820);
  nand g2373 (n_2271, A[48], n_819);
  nand g2374 (n_2272, n_820, n_819);
  nand g2375 (n_2273, A[48], n_820);
  nand g2376 (n_842, n_2271, n_2272, n_2273);
  xor g2377 (n_2274, n_821, n_822);
  xor g2378 (n_828, n_2274, n_823);
  nand g2379 (n_2275, n_821, n_822);
  nand g2380 (n_2276, n_823, n_822);
  nand g2381 (n_2277, n_821, n_823);
  nand g2382 (n_843, n_2275, n_2276, n_2277);
  xor g2383 (n_2278, n_824, n_825);
  xor g2384 (n_829, n_2278, n_826);
  nand g2385 (n_2279, n_824, n_825);
  nand g2386 (n_2280, n_826, n_825);
  nand g2387 (n_2281, n_824, n_826);
  nand g2388 (n_847, n_2279, n_2280, n_2281);
  xor g2389 (n_2282, n_827, n_828);
  xor g2390 (n_831, n_2282, n_829);
  nand g2391 (n_2283, n_827, n_828);
  nand g2392 (n_2284, n_829, n_828);
  nand g2393 (n_2285, n_827, n_829);
  nand g2394 (n_849, n_2283, n_2284, n_2285);
  xor g2395 (n_2286, n_830, n_831);
  xor g2396 (n_145, n_2286, n_832);
  nand g2397 (n_2287, n_830, n_831);
  nand g2398 (n_2288, n_832, n_831);
  nand g2399 (n_2289, n_830, n_832);
  nand g2400 (n_72, n_2287, n_2288, n_2289);
  xor g2403 (n_2290, A[35], A[43]);
  xor g2404 (n_838, n_2290, A[52]);
  nand g2406 (n_2292, A[52], A[43]);
  nand g2407 (n_2293, A[35], A[52]);
  nand g2408 (n_851, n_2165, n_2292, n_2293);
  xor g2409 (n_2294, A[37], A[41]);
  xor g2410 (n_839, n_2294, A[39]);
  nand g2414 (n_852, n_1972, n_1907, n_1843);
  xor g2421 (n_2302, A[47], n_775);
  xor g2422 (n_844, n_2302, n_837);
  nand g2423 (n_2303, A[47], n_775);
  nand g2424 (n_2304, n_837, n_775);
  nand g2425 (n_2305, A[47], n_837);
  nand g2426 (n_857, n_2303, n_2304, n_2305);
  xor g2427 (n_2306, n_838, n_839);
  xor g2428 (n_845, n_2306, n_840);
  nand g2429 (n_2307, n_838, n_839);
  nand g2430 (n_2308, n_840, n_839);
  nand g2431 (n_2309, n_838, n_840);
  nand g2432 (n_858, n_2307, n_2308, n_2309);
  xor g2433 (n_2310, n_808, n_842);
  xor g2434 (n_846, n_2310, n_843);
  nand g2435 (n_2311, n_808, n_842);
  nand g2436 (n_2312, n_843, n_842);
  nand g2437 (n_2313, n_808, n_843);
  nand g2438 (n_862, n_2311, n_2312, n_2313);
  xor g2439 (n_2314, n_844, n_845);
  xor g2440 (n_848, n_2314, n_846);
  nand g2441 (n_2315, n_844, n_845);
  nand g2442 (n_2316, n_846, n_845);
  nand g2443 (n_2317, n_844, n_846);
  nand g2444 (n_864, n_2315, n_2316, n_2317);
  xor g2445 (n_2318, n_847, n_848);
  xor g2446 (n_144, n_2318, n_849);
  nand g2447 (n_2319, n_847, n_848);
  nand g2448 (n_2320, n_849, n_848);
  nand g2449 (n_2321, n_847, n_849);
  nand g2450 (n_71, n_2319, n_2320, n_2321);
  xor g2452 (n_853, n_2322, A[36]);
  nand g2456 (n_867, n_2323, n_1811, n_2325);
  xor g2469 (n_2334, A[48], n_851);
  xor g2470 (n_859, n_2334, n_852);
  nand g2471 (n_2335, A[48], n_851);
  nand g2472 (n_2336, n_852, n_851);
  nand g2473 (n_2337, A[48], n_852);
  nand g2474 (n_872, n_2335, n_2336, n_2337);
  xor g2475 (n_2338, n_853, n_823);
  xor g2476 (n_860, n_2338, n_855);
  nand g2477 (n_2339, n_853, n_823);
  nand g2478 (n_2340, n_855, n_823);
  nand g2479 (n_2341, n_853, n_855);
  nand g2480 (n_874, n_2339, n_2340, n_2341);
  xor g2481 (n_2342, n_824, n_857);
  xor g2482 (n_861, n_2342, n_858);
  nand g2483 (n_2343, n_824, n_857);
  nand g2484 (n_2344, n_858, n_857);
  nand g2485 (n_2345, n_824, n_858);
  nand g2486 (n_876, n_2343, n_2344, n_2345);
  xor g2487 (n_2346, n_859, n_860);
  xor g2488 (n_863, n_2346, n_861);
  nand g2489 (n_2347, n_859, n_860);
  nand g2490 (n_2348, n_861, n_860);
  nand g2491 (n_2349, n_859, n_861);
  nand g2492 (n_879, n_2347, n_2348, n_2349);
  xor g2493 (n_2350, n_862, n_863);
  xor g2494 (n_143, n_2350, n_864);
  nand g2495 (n_2351, n_862, n_863);
  nand g2496 (n_2352, n_864, n_863);
  nand g2497 (n_2353, n_862, n_864);
  nand g2498 (n_70, n_2351, n_2352, n_2353);
  xor g2514 (n_873, n_2362, n_867);
  nand g2517 (n_2365, A[47], n_867);
  nand g2518 (n_886, n_2363, n_2364, n_2365);
  xor g2520 (n_875, n_2366, n_839);
  nand g2523 (n_2369, n_868, n_839);
  nand g2524 (n_887, n_2367, n_2308, n_2369);
  xor g2525 (n_2370, n_808, n_872);
  xor g2526 (n_877, n_2370, n_873);
  nand g2527 (n_2371, n_808, n_872);
  nand g2528 (n_2372, n_873, n_872);
  nand g2529 (n_2373, n_808, n_873);
  nand g2530 (n_890, n_2371, n_2372, n_2373);
  xor g2531 (n_2374, n_874, n_875);
  xor g2532 (n_878, n_2374, n_876);
  nand g2533 (n_2375, n_874, n_875);
  nand g2534 (n_2376, n_876, n_875);
  nand g2535 (n_2377, n_874, n_876);
  nand g2536 (n_892, n_2375, n_2376, n_2377);
  xor g2537 (n_2378, n_877, n_878);
  xor g2538 (n_142, n_2378, n_879);
  nand g2539 (n_2379, n_877, n_878);
  nand g2540 (n_2380, n_879, n_878);
  nand g2541 (n_2381, n_877, n_879);
  nand g2542 (n_69, n_2379, n_2380, n_2381);
  xor g2544 (n_883, n_2322, A[42]);
  nand g2548 (n_895, n_2323, n_2003, n_2327);
  xor g2549 (n_2386, A[40], A[50]);
  xor g2550 (n_885, n_2386, A[46]);
  nand g2551 (n_2387, A[40], A[50]);
  nand g2553 (n_2389, A[40], A[46]);
  nand g2554 (n_896, n_2387, n_2267, n_2389);
  xor g2555 (n_2390, A[44], A[48]);
  xor g2556 (n_884, n_2390, A[43]);
  nand g2558 (n_2392, A[43], A[48]);
  nand g2559 (n_2393, A[44], A[43]);
  nand g2560 (n_899, n_2205, n_2392, n_2393);
  xor g2561 (n_2394, n_852, n_823);
  xor g2562 (n_888, n_2394, n_883);
  nand g2563 (n_2395, n_852, n_823);
  nand g2564 (n_2396, n_883, n_823);
  nand g2565 (n_2397, n_852, n_883);
  nand g2566 (n_901, n_2395, n_2396, n_2397);
  xor g2567 (n_2398, n_884, n_885);
  xor g2568 (n_889, n_2398, n_886);
  nand g2569 (n_2399, n_884, n_885);
  nand g2570 (n_2400, n_886, n_885);
  nand g2571 (n_2401, n_884, n_886);
  nand g2572 (n_902, n_2399, n_2400, n_2401);
  xor g2573 (n_2402, n_887, n_888);
  xor g2574 (n_891, n_2402, n_889);
  nand g2575 (n_2403, n_887, n_888);
  nand g2576 (n_2404, n_889, n_888);
  nand g2577 (n_2405, n_887, n_889);
  nand g2578 (n_905, n_2403, n_2404, n_2405);
  xor g2579 (n_2406, n_890, n_891);
  xor g2580 (n_141, n_2406, n_892);
  nand g2581 (n_2407, n_890, n_891);
  nand g2582 (n_2408, n_892, n_891);
  nand g2583 (n_2409, n_890, n_892);
  nand g2584 (n_68, n_2407, n_2408, n_2409);
  xor g2588 (n_897, n_1906, A[51]);
  nand g2590 (n_2412, A[51], A[39]);
  nand g2591 (n_2413, A[41], A[51]);
  nand g2592 (n_907, n_1907, n_2412, n_2413);
  xor g2593 (n_2414, A[45], A[49]);
  xor g2594 (n_898, n_2414, A[47]);
  nand g2597 (n_2417, A[45], A[47]);
  nand g2598 (n_908, n_2237, n_2172, n_2417);
  xor g2600 (n_900, n_2418, n_896);
  nand g2602 (n_2420, n_896, n_895);
  nand g2604 (n_912, n_2419, n_2420, n_2421);
  xor g2605 (n_2422, n_897, n_898);
  xor g2606 (n_903, n_2422, n_899);
  nand g2607 (n_2423, n_897, n_898);
  nand g2608 (n_2424, n_899, n_898);
  nand g2609 (n_2425, n_897, n_899);
  nand g2610 (n_914, n_2423, n_2424, n_2425);
  xor g2611 (n_2426, n_900, n_901);
  xor g2612 (n_904, n_2426, n_902);
  nand g2613 (n_2427, n_900, n_901);
  nand g2614 (n_2428, n_902, n_901);
  nand g2615 (n_2429, n_900, n_902);
  nand g2616 (n_916, n_2427, n_2428, n_2429);
  xor g2617 (n_2430, n_903, n_904);
  xor g2618 (n_140, n_2430, n_905);
  nand g2619 (n_2431, n_903, n_904);
  nand g2620 (n_2432, n_905, n_904);
  nand g2621 (n_2433, n_903, n_905);
  nand g2622 (n_67, n_2431, n_2432, n_2433);
  xor g2624 (n_855, n_2326, A[40]);
  nand g2628 (n_868, n_2327, n_1939, n_2329);
  xor g2635 (n_2442, A[48], A[43]);
  xor g2636 (n_911, n_2442, n_907);
  nand g2638 (n_2444, n_907, A[43]);
  nand g2639 (n_2445, A[48], n_907);
  nand g2640 (n_923, n_2392, n_2444, n_2445);
  xor g2641 (n_2446, n_908, n_855);
  xor g2642 (n_913, n_2446, n_824);
  nand g2643 (n_2447, n_908, n_855);
  nand g2644 (n_2448, n_824, n_855);
  nand g2645 (n_2449, n_908, n_824);
  nand g2646 (n_924, n_2447, n_2448, n_2449);
  xor g2647 (n_2450, n_911, n_912);
  xor g2648 (n_915, n_2450, n_913);
  nand g2649 (n_2451, n_911, n_912);
  nand g2650 (n_2452, n_913, n_912);
  nand g2651 (n_2453, n_911, n_913);
  nand g2652 (n_927, n_2451, n_2452, n_2453);
  xor g2653 (n_2454, n_914, n_915);
  xor g2654 (n_139, n_2454, n_916);
  nand g2655 (n_2455, n_914, n_915);
  nand g2656 (n_2456, n_916, n_915);
  nand g2657 (n_2457, n_914, n_916);
  nand g2658 (n_66, n_2455, n_2456, n_2457);
  xor g2661 (n_2458, A[41], A[51]);
  xor g2662 (n_922, n_2458, A[45]);
  nand g2665 (n_2461, A[41], A[45]);
  nand g2666 (n_929, n_2413, n_2235, n_2461);
  xor g2667 (n_2462, A[49], A[47]);
  nand g2672 (n_931, n_2172, n_2363, n_2465);
  xor g2673 (n_2366, n_868, n_840);
  xor g2674 (n_925, n_2366, n_921);
  nand g2675 (n_2367, n_868, n_840);
  nand g2676 (n_2468, n_921, n_840);
  nand g2677 (n_2469, n_868, n_921);
  nand g2678 (n_934, n_2367, n_2468, n_2469);
  xor g2679 (n_2470, n_922, n_923);
  xor g2680 (n_926, n_2470, n_924);
  nand g2681 (n_2471, n_922, n_923);
  nand g2682 (n_2472, n_924, n_923);
  nand g2683 (n_2473, n_922, n_924);
  nand g2684 (n_936, n_2471, n_2472, n_2473);
  xor g2685 (n_2474, n_925, n_926);
  xor g2686 (n_138, n_2474, n_927);
  nand g2687 (n_2475, n_925, n_926);
  nand g2688 (n_2476, n_927, n_926);
  nand g2689 (n_2477, n_925, n_927);
  nand g2690 (n_65, n_2475, n_2476, n_2477);
  xor g2692 (n_930, n_2326, A[50]);
  nand g2694 (n_2480, A[50], A[42]);
  nand g2696 (n_940, n_2327, n_2480, n_2481);
  xor g2697 (n_2482, A[46], A[44]);
  xor g2698 (n_932, n_2482, A[48]);
  nand g2702 (n_939, n_2268, n_2205, n_2140);
  xor g2703 (n_2486, A[43], n_929);
  xor g2704 (n_933, n_2486, n_930);
  nand g2705 (n_2487, A[43], n_929);
  nand g2706 (n_2488, n_930, n_929);
  nand g2707 (n_2489, A[43], n_930);
  nand g2708 (n_942, n_2487, n_2488, n_2489);
  xor g2709 (n_2490, n_931, n_932);
  xor g2710 (n_935, n_2490, n_933);
  nand g2711 (n_2491, n_931, n_932);
  nand g2712 (n_2492, n_933, n_932);
  nand g2713 (n_2493, n_931, n_933);
  nand g2714 (n_945, n_2491, n_2492, n_2493);
  xor g2715 (n_2494, n_934, n_935);
  xor g2716 (n_137, n_2494, n_936);
  nand g2717 (n_2495, n_934, n_935);
  nand g2718 (n_2496, n_936, n_935);
  nand g2719 (n_2497, n_934, n_936);
  nand g2720 (n_64, n_2495, n_2496, n_2497);
  xor g2730 (n_943, n_2362, n_939);
  nand g2733 (n_2505, A[47], n_939);
  nand g2734 (n_950, n_2363, n_2504, n_2505);
  xor g2735 (n_2506, n_940, n_808);
  xor g2736 (n_944, n_2506, n_942);
  nand g2737 (n_2507, n_940, n_808);
  nand g2738 (n_2508, n_942, n_808);
  nand g2739 (n_2509, n_940, n_942);
  nand g2740 (n_952, n_2507, n_2508, n_2509);
  xor g2741 (n_2510, n_943, n_944);
  xor g2742 (n_136, n_2510, n_945);
  nand g2743 (n_2511, n_943, n_944);
  nand g2744 (n_2512, n_945, n_944);
  nand g2745 (n_2513, n_943, n_945);
  nand g2746 (n_135, n_2511, n_2512, n_2513);
  xor g2748 (n_948, n_2514, A[46]);
  nand g2752 (n_955, n_2481, n_2267, n_2517);
  xor g2759 (n_2522, n_823, n_948);
  xor g2760 (n_951, n_2522, n_884);
  nand g2761 (n_2523, n_823, n_948);
  nand g2762 (n_2524, n_884, n_948);
  nand g2763 (n_2525, n_823, n_884);
  nand g2764 (n_959, n_2523, n_2524, n_2525);
  xor g2765 (n_2526, n_950, n_951);
  xor g2766 (n_63, n_2526, n_952);
  nand g2767 (n_2527, n_950, n_951);
  nand g2768 (n_2528, n_952, n_951);
  nand g2769 (n_2529, n_950, n_952);
  nand g2770 (n_134, n_2527, n_2528, n_2529);
  xor g2780 (n_958, n_2534, n_899);
  nand g2782 (n_2536, n_899, n_955);
  nand g2784 (n_964, n_2535, n_2536, n_2537);
  xor g2785 (n_2538, n_898, n_958);
  xor g2786 (n_62, n_2538, n_959);
  nand g2787 (n_2539, n_898, n_958);
  nand g2788 (n_2540, n_959, n_958);
  nand g2789 (n_2541, n_898, n_959);
  nand g2790 (n_61, n_2539, n_2540, n_2541);
  xor g2797 (n_2546, A[48], A[51]);
  xor g2798 (n_963, n_2546, n_908);
  nand g2799 (n_2547, A[48], A[51]);
  nand g2800 (n_2548, n_908, A[51]);
  nand g2801 (n_2549, A[48], n_908);
  nand g2802 (n_969, n_2547, n_2548, n_2549);
  xor g2803 (n_2550, n_948, n_963);
  xor g2804 (n_133, n_2550, n_964);
  nand g2805 (n_2551, n_948, n_963);
  nand g2806 (n_2552, n_964, n_963);
  nand g2807 (n_2553, n_948, n_964);
  nand g2808 (n_132, n_2551, n_2552, n_2553);
  nand g2816 (n_972, n_2172, n_2556, n_2557);
  xor g2817 (n_2558, n_955, n_968);
  xor g2818 (n_60, n_2558, n_969);
  nand g2819 (n_2559, n_955, n_968);
  nand g2820 (n_2560, n_969, n_968);
  nand g2821 (n_2561, n_955, n_969);
  nand g2822 (n_131, n_2559, n_2560, n_2561);
  xor g2824 (n_971, n_2514, A[48]);
  nand g2828 (n_975, n_2481, n_2204, n_2565);
  xor g2829 (n_2566, A[51], n_971);
  xor g2830 (n_59, n_2566, n_972);
  nand g2831 (n_2567, A[51], n_971);
  nand g2832 (n_2568, n_972, n_971);
  nand g2833 (n_2569, A[51], n_972);
  nand g2834 (n_130, n_2567, n_2568, n_2569);
  xor g2838 (n_58, n_2570, n_975);
  nand g2841 (n_2573, A[51], n_975);
  nand g2842 (n_129, n_2571, n_2572, n_2573);
  xor g2844 (n_57, n_2514, A[49]);
  nand g2846 (n_2576, A[49], A[50]);
  nand g2848 (n_128, n_2481, n_2576, n_2577);
  nor g11 (n_2593, A[2], A[0]);
  nor g13 (n_2589, A[1], A[3]);
  nor g15 (n_2599, A[2], n_193);
  nand g16 (n_2594, A[2], n_193);
  nor g17 (n_2595, n_120, n_192);
  nand g18 (n_2596, n_120, n_192);
  nor g19 (n_2605, n_119, n_191);
  nand g20 (n_2600, n_119, n_191);
  nor g21 (n_2601, n_118, n_190);
  nand g22 (n_2602, n_118, n_190);
  nor g23 (n_2611, n_117, n_189);
  nand g24 (n_2606, n_117, n_189);
  nor g25 (n_2607, n_116, n_188);
  nand g26 (n_2608, n_116, n_188);
  nor g27 (n_2617, n_115, n_187);
  nand g28 (n_2612, n_115, n_187);
  nor g29 (n_2613, n_114, n_186);
  nand g30 (n_2614, n_114, n_186);
  nor g31 (n_2623, n_113, n_185);
  nand g32 (n_2618, n_113, n_185);
  nor g33 (n_2619, n_112, n_184);
  nand g34 (n_2620, n_112, n_184);
  nor g35 (n_2629, n_111, n_183);
  nand g36 (n_2624, n_111, n_183);
  nor g37 (n_2625, n_110, n_182);
  nand g38 (n_2626, n_110, n_182);
  nor g39 (n_2635, n_109, n_181);
  nand g40 (n_2630, n_109, n_181);
  nor g41 (n_2631, n_108, n_180);
  nand g42 (n_2632, n_108, n_180);
  nor g43 (n_2641, n_107, n_179);
  nand g44 (n_2636, n_107, n_179);
  nor g45 (n_2637, n_106, n_178);
  nand g46 (n_2638, n_106, n_178);
  nor g47 (n_2647, n_105, n_177);
  nand g48 (n_2642, n_105, n_177);
  nor g49 (n_2643, n_104, n_176);
  nand g50 (n_2644, n_104, n_176);
  nor g51 (n_2653, n_103, n_175);
  nand g52 (n_2648, n_103, n_175);
  nor g53 (n_2649, n_102, n_174);
  nand g54 (n_2650, n_102, n_174);
  nor g55 (n_2659, n_101, n_173);
  nand g56 (n_2654, n_101, n_173);
  nor g57 (n_2655, n_100, n_172);
  nand g58 (n_2656, n_100, n_172);
  nor g59 (n_2665, n_99, n_171);
  nand g60 (n_2660, n_99, n_171);
  nor g61 (n_2661, n_98, n_170);
  nand g62 (n_2662, n_98, n_170);
  nor g63 (n_2671, n_97, n_169);
  nand g64 (n_2666, n_97, n_169);
  nor g65 (n_2667, n_96, n_168);
  nand g66 (n_2668, n_96, n_168);
  nor g67 (n_2677, n_95, n_167);
  nand g68 (n_2672, n_95, n_167);
  nor g69 (n_2673, n_94, n_166);
  nand g70 (n_2674, n_94, n_166);
  nor g71 (n_2683, n_93, n_165);
  nand g72 (n_2678, n_93, n_165);
  nor g73 (n_2679, n_92, n_164);
  nand g74 (n_2680, n_92, n_164);
  nor g75 (n_2689, n_91, n_163);
  nand g76 (n_2684, n_91, n_163);
  nor g77 (n_2685, n_90, n_162);
  nand g78 (n_2686, n_90, n_162);
  nor g79 (n_2695, n_89, n_161);
  nand g80 (n_2690, n_89, n_161);
  nor g81 (n_2691, n_88, n_160);
  nand g82 (n_2692, n_88, n_160);
  nor g83 (n_2701, n_87, n_159);
  nand g84 (n_2696, n_87, n_159);
  nor g85 (n_2697, n_86, n_158);
  nand g86 (n_2698, n_86, n_158);
  nor g87 (n_2707, n_85, n_157);
  nand g88 (n_2702, n_85, n_157);
  nor g89 (n_2703, n_84, n_156);
  nand g90 (n_2704, n_84, n_156);
  nor g91 (n_2713, n_83, n_155);
  nand g92 (n_2708, n_83, n_155);
  nor g93 (n_2709, n_82, n_154);
  nand g94 (n_2710, n_82, n_154);
  nor g95 (n_2719, n_81, n_153);
  nand g96 (n_2714, n_81, n_153);
  nor g97 (n_2715, n_80, n_152);
  nand g98 (n_2716, n_80, n_152);
  nor g99 (n_2725, n_79, n_151);
  nand g100 (n_2720, n_79, n_151);
  nor g101 (n_2721, n_78, n_150);
  nand g102 (n_2722, n_78, n_150);
  nor g103 (n_2731, n_77, n_149);
  nand g104 (n_2726, n_77, n_149);
  nor g105 (n_2727, n_76, n_148);
  nand g106 (n_2728, n_76, n_148);
  nor g107 (n_2737, n_75, n_147);
  nand g108 (n_2732, n_75, n_147);
  nor g109 (n_2733, n_74, n_146);
  nand g110 (n_2734, n_74, n_146);
  nor g111 (n_2743, n_73, n_145);
  nand g112 (n_2738, n_73, n_145);
  nor g113 (n_2739, n_72, n_144);
  nand g114 (n_2740, n_72, n_144);
  nor g115 (n_2749, n_71, n_143);
  nand g116 (n_2744, n_71, n_143);
  nor g117 (n_2745, n_70, n_142);
  nand g118 (n_2746, n_70, n_142);
  nor g119 (n_2755, n_69, n_141);
  nand g120 (n_2750, n_69, n_141);
  nor g121 (n_2751, n_68, n_140);
  nand g122 (n_2752, n_68, n_140);
  nor g123 (n_2761, n_67, n_139);
  nand g124 (n_2756, n_67, n_139);
  nor g125 (n_2757, n_66, n_138);
  nand g126 (n_2758, n_66, n_138);
  nor g127 (n_2767, n_65, n_137);
  nand g128 (n_2762, n_65, n_137);
  nor g129 (n_2763, n_64, n_136);
  nand g130 (n_2764, n_64, n_136);
  nor g131 (n_2773, n_63, n_135);
  nand g132 (n_2768, n_63, n_135);
  nor g133 (n_2769, n_62, n_134);
  nand g134 (n_2770, n_62, n_134);
  nor g135 (n_2779, n_61, n_133);
  nand g136 (n_2774, n_61, n_133);
  nor g137 (n_2775, n_60, n_132);
  nand g138 (n_2776, n_60, n_132);
  nor g139 (n_2785, n_59, n_131);
  nand g140 (n_2780, n_59, n_131);
  nor g141 (n_2781, n_58, n_130);
  nand g142 (n_2782, n_58, n_130);
  nor g143 (n_2791, n_57, n_129);
  nand g144 (n_2786, n_57, n_129);
  nor g154 (n_2591, n_983, n_2589);
  nor g158 (n_2597, n_2594, n_2595);
  nor g161 (n_2806, n_2599, n_2595);
  nor g162 (n_2603, n_2600, n_2601);
  nor g165 (n_2800, n_2605, n_2601);
  nor g166 (n_2609, n_2606, n_2607);
  nor g169 (n_2813, n_2611, n_2607);
  nor g170 (n_2615, n_2612, n_2613);
  nor g173 (n_2807, n_2617, n_2613);
  nor g174 (n_2621, n_2618, n_2619);
  nor g177 (n_2820, n_2623, n_2619);
  nor g178 (n_2627, n_2624, n_2625);
  nor g181 (n_2814, n_2629, n_2625);
  nor g182 (n_2633, n_2630, n_2631);
  nor g185 (n_2827, n_2635, n_2631);
  nor g186 (n_2639, n_2636, n_2637);
  nor g189 (n_2821, n_2641, n_2637);
  nor g190 (n_2645, n_2642, n_2643);
  nor g193 (n_2834, n_2647, n_2643);
  nor g194 (n_2651, n_2648, n_2649);
  nor g197 (n_2828, n_2653, n_2649);
  nor g198 (n_2657, n_2654, n_2655);
  nor g201 (n_2841, n_2659, n_2655);
  nor g202 (n_2663, n_2660, n_2661);
  nor g205 (n_2835, n_2665, n_2661);
  nor g206 (n_2669, n_2666, n_2667);
  nor g209 (n_2848, n_2671, n_2667);
  nor g210 (n_2675, n_2672, n_2673);
  nor g213 (n_2842, n_2677, n_2673);
  nor g214 (n_2681, n_2678, n_2679);
  nor g217 (n_2855, n_2683, n_2679);
  nor g218 (n_2687, n_2684, n_2685);
  nor g221 (n_2849, n_2689, n_2685);
  nor g222 (n_2693, n_2690, n_2691);
  nor g225 (n_2862, n_2695, n_2691);
  nor g226 (n_2699, n_2696, n_2697);
  nor g229 (n_2856, n_2701, n_2697);
  nor g230 (n_2705, n_2702, n_2703);
  nor g233 (n_2869, n_2707, n_2703);
  nor g234 (n_2711, n_2708, n_2709);
  nor g237 (n_2863, n_2713, n_2709);
  nor g238 (n_2717, n_2714, n_2715);
  nor g241 (n_2876, n_2719, n_2715);
  nor g242 (n_2723, n_2720, n_2721);
  nor g245 (n_2870, n_2725, n_2721);
  nor g246 (n_2729, n_2726, n_2727);
  nor g249 (n_2883, n_2731, n_2727);
  nor g250 (n_2735, n_2732, n_2733);
  nor g253 (n_2877, n_2737, n_2733);
  nor g254 (n_2741, n_2738, n_2739);
  nor g257 (n_2890, n_2743, n_2739);
  nor g258 (n_2747, n_2744, n_2745);
  nor g261 (n_2884, n_2749, n_2745);
  nor g262 (n_2753, n_2750, n_2751);
  nor g265 (n_2897, n_2755, n_2751);
  nor g266 (n_2759, n_2756, n_2757);
  nor g269 (n_2891, n_2761, n_2757);
  nor g270 (n_2765, n_2762, n_2763);
  nor g273 (n_2904, n_2767, n_2763);
  nor g274 (n_2771, n_2768, n_2769);
  nor g277 (n_2898, n_2773, n_2769);
  nor g278 (n_2777, n_2774, n_2775);
  nor g281 (n_2911, n_2779, n_2775);
  nor g282 (n_2783, n_2780, n_2781);
  nor g285 (n_2905, n_2785, n_2781);
  nor g286 (n_2789, n_2786, n_2787);
  nor g289 (n_2913, n_2791, n_2787);
  nand g300 (n_2914, n_2806, n_2800);
  nand g305 (n_2924, n_2813, n_2807);
  nand g310 (n_2919, n_2820, n_2814);
  nand g315 (n_2930, n_2827, n_2821);
  nand g320 (n_2925, n_2834, n_2828);
  nand g325 (n_2936, n_2841, n_2835);
  nand g330 (n_2931, n_2848, n_2842);
  nand g335 (n_2942, n_2855, n_2849);
  nand g340 (n_2937, n_2862, n_2856);
  nand g345 (n_2948, n_2869, n_2863);
  nand g350 (n_2943, n_2876, n_2870);
  nand g355 (n_2954, n_2883, n_2877);
  nand g360 (n_2949, n_2890, n_2884);
  nand g365 (n_2960, n_2897, n_2891);
  nand g370 (n_2955, n_2904, n_2898);
  nand g375 (n_2962, n_2911, n_2905);
  nand g383 (n_2964, n_2917, n_2918);
  nor g384 (n_2922, n_2919, n_2920);
  nor g387 (n_2963, n_2924, n_2919);
  nor g388 (n_2928, n_2925, n_2926);
  nor g391 (n_2973, n_2930, n_2925);
  nor g392 (n_2934, n_2931, n_2932);
  nor g395 (n_2967, n_2936, n_2931);
  nor g396 (n_2940, n_2937, n_2938);
  nor g399 (n_2980, n_2942, n_2937);
  nor g400 (n_2946, n_2943, n_2944);
  nor g403 (n_2974, n_2948, n_2943);
  nor g404 (n_2952, n_2949, n_2950);
  nor g407 (n_2987, n_2954, n_2949);
  nor g408 (n_2958, n_2955, n_2956);
  nor g411 (n_2981, n_2960, n_2955);
  nand g416 (n_2966, n_2963, n_2964);
  nand g417 (n_2989, n_2965, n_2966);
  nand g2858 (n_2988, n_2973, n_2967);
  nand g2863 (n_2998, n_2980, n_2974);
  nand g2868 (n_2993, n_2987, n_2981);
  nand g2871 (n_3000, n_2991, n_2992);
  nor g2872 (n_2996, n_2993, n_2994);
  nor g2875 (n_2999, n_2998, n_2993);
  nand g2876 (n_3002, n_2999, n_3000);
  nand g2877 (n_3009, n_3001, n_3002);
  nand g2880 (n_3007, n_2994, n_3004);
  nand g2881 (n_3005, n_2973, n_2989);
  nand g2882 (n_3014, n_2968, n_3005);
  nand g2883 (n_3006, n_2980, n_3000);
  nand g2884 (n_3019, n_2975, n_3006);
  nand g2885 (n_3008, n_2987, n_3007);
  nand g2886 (n_3024, n_2982, n_3008);
  nand g2889 (n_3031, n_2920, n_3011);
  nand g2892 (n_3034, n_2926, n_3013);
  nand g2895 (n_3037, n_2932, n_3016);
  nand g2898 (n_3040, n_2938, n_3018);
  nand g2901 (n_3043, n_2944, n_3021);
  nand g2904 (n_3046, n_2950, n_3023);
  nand g2907 (n_3049, n_2956, n_3026);
  nand g2910 (n_3052, n_2961, n_3028);
  nand g2912 (n_3058, n_2801, n_3029);
  nand g2913 (n_3030, n_2813, n_2964);
  nand g2914 (n_3063, n_2808, n_3030);
  nand g2915 (n_3032, n_2820, n_3031);
  nand g2916 (n_3068, n_2815, n_3032);
  nand g2917 (n_3033, n_2827, n_2989);
  nand g2918 (n_3073, n_2822, n_3033);
  nand g2919 (n_3035, n_2834, n_3034);
  nand g2920 (n_3078, n_2829, n_3035);
  nand g2921 (n_3036, n_2841, n_3014);
  nand g2922 (n_3083, n_2836, n_3036);
  nand g2923 (n_3038, n_2848, n_3037);
  nand g2924 (n_3088, n_2843, n_3038);
  nand g2925 (n_3039, n_2855, n_3000);
  nand g2926 (n_3093, n_2850, n_3039);
  nand g2927 (n_3041, n_2862, n_3040);
  nand g2928 (n_3098, n_2857, n_3041);
  nand g2929 (n_3042, n_2869, n_3019);
  nand g2930 (n_3103, n_2864, n_3042);
  nand g2931 (n_3044, n_2876, n_3043);
  nand g2932 (n_3108, n_2871, n_3044);
  nand g2933 (n_3045, n_2883, n_3007);
  nand g2934 (n_3113, n_2878, n_3045);
  nand g2935 (n_3047, n_2890, n_3046);
  nand g2936 (n_3118, n_2885, n_3047);
  nand g2937 (n_3048, n_2897, n_3024);
  nand g2938 (n_3123, n_2892, n_3048);
  nand g2939 (n_3050, n_2904, n_3049);
  nand g2940 (n_3128, n_2899, n_3050);
  nand g2941 (n_3051, n_2911, n_3009);
  nand g2942 (n_3133, n_2906, n_3051);
  nand g2943 (n_3053, n_2913, n_3052);
  nand g2944 (n_3138, n_2912, n_3053);
  nand g2950 (n_3148, n_2594, n_3057);
  nand g2953 (n_3152, n_2600, n_3060);
  nand g2956 (n_3156, n_2606, n_3062);
  nand g2959 (n_3160, n_2612, n_3065);
  nand g2962 (n_3164, n_2618, n_3067);
  nand g2965 (n_3168, n_2624, n_3070);
  nand g2968 (n_3172, n_2630, n_3072);
  nand g2971 (n_3176, n_2636, n_3075);
  nand g2974 (n_3180, n_2642, n_3077);
  nand g2977 (n_3184, n_2648, n_3080);
  nand g2980 (n_3188, n_2654, n_3082);
  nand g2983 (n_3192, n_2660, n_3085);
  nand g2986 (n_3196, n_2666, n_3087);
  nand g2989 (n_3200, n_2672, n_3090);
  nand g2992 (n_3204, n_2678, n_3092);
  nand g2995 (n_3208, n_2684, n_3095);
  nand g2998 (n_3212, n_2690, n_3097);
  nand g3001 (n_3216, n_2696, n_3100);
  nand g3004 (n_3220, n_2702, n_3102);
  nand g3007 (n_3224, n_2708, n_3105);
  nand g3010 (n_3228, n_2714, n_3107);
  nand g3013 (n_3232, n_2720, n_3110);
  nand g3016 (n_3236, n_2726, n_3112);
  nand g3019 (n_3240, n_2732, n_3115);
  nand g3022 (n_3244, n_2738, n_3117);
  nand g3025 (n_3248, n_2744, n_3120);
  nand g3028 (n_3252, n_2750, n_3122);
  nand g3031 (n_3256, n_2756, n_3125);
  nand g3034 (n_3260, n_2762, n_3127);
  nand g3037 (n_3264, n_2768, n_3130);
  nand g3040 (n_3268, n_2774, n_3132);
  nand g3043 (n_3272, n_2780, n_3135);
  nand g3046 (n_3276, n_2786, n_3137);
  nand g3049 (n_3280, n_2792, n_3140);
  xnor g3061 (Z[5], n_3148, n_3149);
  xnor g3063 (Z[6], n_3058, n_3150);
  xnor g3066 (Z[7], n_3152, n_3153);
  xnor g3068 (Z[8], n_2964, n_3154);
  xnor g3071 (Z[9], n_3156, n_3157);
  xnor g3073 (Z[10], n_3063, n_3158);
  xnor g3076 (Z[11], n_3160, n_3161);
  xnor g3078 (Z[12], n_3031, n_3162);
  xnor g3081 (Z[13], n_3164, n_3165);
  xnor g3083 (Z[14], n_3068, n_3166);
  xnor g3086 (Z[15], n_3168, n_3169);
  xnor g3088 (Z[16], n_2989, n_3170);
  xnor g3091 (Z[17], n_3172, n_3173);
  xnor g3093 (Z[18], n_3073, n_3174);
  xnor g3096 (Z[19], n_3176, n_3177);
  xnor g3098 (Z[20], n_3034, n_3178);
  xnor g3101 (Z[21], n_3180, n_3181);
  xnor g3103 (Z[22], n_3078, n_3182);
  xnor g3106 (Z[23], n_3184, n_3185);
  xnor g3108 (Z[24], n_3014, n_3186);
  xnor g3111 (Z[25], n_3188, n_3189);
  xnor g3113 (Z[26], n_3083, n_3190);
  xnor g3116 (Z[27], n_3192, n_3193);
  xnor g3118 (Z[28], n_3037, n_3194);
  xnor g3121 (Z[29], n_3196, n_3197);
  xnor g3123 (Z[30], n_3088, n_3198);
  xnor g3126 (Z[31], n_3200, n_3201);
  xnor g3128 (Z[32], n_3000, n_3202);
  xnor g3131 (Z[33], n_3204, n_3205);
  xnor g3133 (Z[34], n_3093, n_3206);
  xnor g3136 (Z[35], n_3208, n_3209);
  xnor g3138 (Z[36], n_3040, n_3210);
  xnor g3141 (Z[37], n_3212, n_3213);
  xnor g3143 (Z[38], n_3098, n_3214);
  xnor g3146 (Z[39], n_3216, n_3217);
  xnor g3148 (Z[40], n_3019, n_3218);
  xnor g3151 (Z[41], n_3220, n_3221);
  xnor g3153 (Z[42], n_3103, n_3222);
  xnor g3156 (Z[43], n_3224, n_3225);
  xnor g3158 (Z[44], n_3043, n_3226);
  xnor g3161 (Z[45], n_3228, n_3229);
  xnor g3163 (Z[46], n_3108, n_3230);
  xnor g3166 (Z[47], n_3232, n_3233);
  xnor g3168 (Z[48], n_3007, n_3234);
  xnor g3171 (Z[49], n_3236, n_3237);
  xnor g3173 (Z[50], n_3113, n_3238);
  xnor g3176 (Z[51], n_3240, n_3241);
  xnor g3178 (Z[52], n_3046, n_3242);
  xnor g3181 (Z[53], n_3244, n_3245);
  xnor g3183 (Z[54], n_3118, n_3246);
  xnor g3186 (Z[55], n_3248, n_3249);
  xnor g3188 (Z[56], n_3024, n_3250);
  xnor g3191 (Z[57], n_3252, n_3253);
  xnor g3193 (Z[58], n_3123, n_3254);
  xnor g3196 (Z[59], n_3256, n_3257);
  xnor g3198 (Z[60], n_3049, n_3258);
  xnor g3201 (Z[61], n_3260, n_3261);
  xnor g3203 (Z[62], n_3128, n_3262);
  xnor g3206 (Z[63], n_3264, n_3265);
  xnor g3208 (Z[64], n_3009, n_3266);
  xnor g3211 (Z[65], n_3268, n_3269);
  xnor g3213 (Z[66], n_3133, n_3270);
  xnor g3216 (Z[67], n_3272, n_3273);
  xnor g3218 (Z[68], n_3052, n_3274);
  xnor g3221 (Z[69], n_3276, n_3277);
  xnor g3223 (Z[70], n_3138, n_3278);
  or g3240 (n_278, wc, wc0, n_120);
  not gc0 (wc0, n_983);
  not gc (wc, n_997);
  or g3241 (n_287, wc1, wc2, n_272);
  not gc2 (wc2, n_997);
  not gc1 (wc1, n_1016);
  or g3242 (n_300, wc3, n_277, n_272);
  not gc3 (wc3, n_1044);
  or g3243 (n_317, wc4, wc5, n_277);
  not gc5 (wc5, n_1079);
  not gc4 (wc4, n_1080);
  or g3244 (n_339, wc6, wc7, n_277);
  not gc7 (wc7, n_1127);
  not gc6 (wc6, n_1128);
  or g3245 (n_386, wc8, wc9, n_272);
  not gc9 (wc9, n_1128);
  not gc8 (wc8, n_1175);
  or g3246 (n_414, wc10, wc11, n_277);
  not gc11 (wc11, n_1304);
  not gc10 (wc10, n_1305);
  or g3247 (n_440, wc12, wc13, n_286);
  not gc13 (wc13, n_1244);
  not gc12 (wc12, n_1368);
  or g3248 (n_468, wc14, wc15, n_299);
  not gc15 (wc15, n_1308);
  not gc14 (wc14, n_1432);
  or g3249 (n_496, wc16, wc17, n_316);
  not gc17 (wc17, n_1237);
  not gc16 (wc16, n_1496);
  or g3250 (n_524, wc18, wc19, n_337);
  not gc19 (wc19, n_1301);
  not gc18 (wc18, n_1560);
  or g3251 (n_552, wc20, wc21, n_362);
  not gc21 (wc21, n_1365);
  not gc20 (wc20, n_1624);
  xnor g3252 (n_2322, A[52], A[38]);
  or g3253 (n_2323, wc22, A[52]);
  not gc22 (wc22, A[38]);
  or g3254 (n_2325, wc23, A[52]);
  not gc23 (wc23, A[36]);
  xnor g3255 (n_2362, A[47], A[43]);
  or g3256 (n_2363, A[43], wc24);
  not gc24 (wc24, A[47]);
  or g3257 (n_2327, wc25, A[52]);
  not gc25 (wc25, A[42]);
  xnor g3258 (n_2326, A[52], A[42]);
  or g3259 (n_2329, wc26, A[52]);
  not gc26 (wc26, A[40]);
  xnor g3260 (n_921, n_2462, A[43]);
  or g3261 (n_2465, A[43], wc27);
  not gc27 (wc27, A[49]);
  or g3262 (n_2481, wc28, A[52]);
  not gc28 (wc28, A[50]);
  xnor g3263 (n_2514, A[52], A[50]);
  or g3264 (n_2517, wc29, A[52]);
  not gc29 (wc29, A[46]);
  xnor g3265 (n_968, n_2462, A[51]);
  or g3266 (n_2556, wc30, A[51]);
  not gc30 (wc30, A[47]);
  or g3267 (n_2557, wc31, A[51]);
  not gc31 (wc31, A[49]);
  or g3268 (n_2565, wc32, A[52]);
  not gc32 (wc32, A[48]);
  xnor g3269 (n_2570, A[51], A[49]);
  or g3270 (n_2571, A[49], wc33);
  not gc33 (wc33, A[51]);
  or g3271 (n_2577, wc34, A[52]);
  not gc34 (wc34, A[49]);
  and g3272 (n_2795, wc35, A[52]);
  not gc35 (wc35, A[51]);
  or g3273 (n_2792, wc36, A[52]);
  not gc36 (wc36, A[51]);
  or g3274 (n_368, wc37, wc38, n_277);
  not gc38 (wc38, n_1184);
  not gc37 (wc37, n_1185);
  or g3275 (n_2421, A[43], wc39);
  not gc39 (wc39, n_896);
  or g3276 (n_2504, A[43], wc40);
  not gc40 (wc40, n_939);
  and g3277 (n_2798, wc41, n_979);
  not gc41 (wc41, n_2591);
  or g3279 (n_3142, n_2593, wc42);
  not gc42 (wc42, n_983);
  or g3280 (n_3145, n_2589, wc43);
  not gc43 (wc43, n_979);
  or g3281 (n_2364, A[43], wc44);
  not gc44 (wc44, n_867);
  xnor g3282 (n_2418, n_895, A[43]);
  or g3283 (n_2419, A[43], wc45);
  not gc45 (wc45, n_895);
  xnor g3284 (n_2534, n_955, A[51]);
  or g3285 (n_2535, A[51], wc46);
  not gc46 (wc46, n_955);
  or g3286 (n_2537, A[51], wc47);
  not gc47 (wc47, n_899);
  or g3287 (n_2572, A[49], wc48);
  not gc48 (wc48, n_975);
  and g3288 (n_2787, A[51], wc49);
  not gc49 (wc49, n_128);
  or g3289 (n_2788, A[51], wc50);
  not gc50 (wc50, n_128);
  or g3290 (n_3146, wc51, n_2599);
  not gc51 (wc51, n_2594);
  or g3291 (n_3278, wc52, n_2795);
  not gc52 (wc52, n_2792);
  and g3292 (n_2801, wc53, n_2596);
  not gc53 (wc53, n_2597);
  not g3293 (Z[2], n_3142);
  or g3294 (n_3149, wc54, n_2595);
  not gc54 (wc54, n_2596);
  or g3295 (n_3150, wc55, n_2605);
  not gc55 (wc55, n_2600);
  and g3296 (n_2803, wc56, n_2602);
  not gc56 (wc56, n_2603);
  or g3299 (n_3153, wc57, n_2601);
  not gc57 (wc57, n_2602);
  or g3300 (n_3277, wc58, n_2787);
  not gc58 (wc58, n_2788);
  and g3301 (n_2808, wc59, n_2608);
  not gc59 (wc59, n_2609);
  and g3302 (n_2804, wc60, n_2800);
  not gc60 (wc60, n_2801);
  or g3303 (n_3029, n_2798, wc61);
  not gc61 (wc61, n_2806);
  or g3304 (n_3057, n_2599, n_2798);
  xor g3305 (Z[3], n_983, n_3145);
  xor g3306 (Z[4], n_2798, n_3146);
  or g3307 (n_3154, wc62, n_2611);
  not gc62 (wc62, n_2606);
  or g3308 (n_3157, wc63, n_2607);
  not gc63 (wc63, n_2608);
  and g3309 (n_2912, n_2788, wc64);
  not gc64 (wc64, n_2789);
  and g3310 (n_2917, wc65, n_2803);
  not gc65 (wc65, n_2804);
  or g3311 (n_2918, n_2914, n_2798);
  or g3312 (n_3158, wc66, n_2617);
  not gc66 (wc66, n_2612);
  or g3313 (n_3273, wc67, n_2781);
  not gc67 (wc67, n_2782);
  or g3314 (n_3274, wc68, n_2791);
  not gc68 (wc68, n_2786);
  and g3315 (n_2810, wc69, n_2614);
  not gc69 (wc69, n_2615);
  and g3316 (n_2815, wc70, n_2620);
  not gc70 (wc70, n_2621);
  and g3317 (n_2908, wc71, n_2782);
  not gc71 (wc71, n_2783);
  or g3318 (n_3060, wc72, n_2605);
  not gc72 (wc72, n_3058);
  or g3319 (n_3161, wc73, n_2613);
  not gc73 (wc73, n_2614);
  or g3320 (n_3162, wc74, n_2623);
  not gc74 (wc74, n_2618);
  or g3321 (n_3165, wc75, n_2619);
  not gc75 (wc75, n_2620);
  or g3322 (n_3270, wc76, n_2785);
  not gc76 (wc76, n_2780);
  and g3323 (n_2817, wc77, n_2626);
  not gc77 (wc77, n_2627);
  and g3324 (n_2906, wc78, n_2776);
  not gc78 (wc78, n_2777);
  and g3325 (n_2811, wc79, n_2807);
  not gc79 (wc79, n_2808);
  or g3326 (n_3062, wc80, n_2611);
  not gc80 (wc80, n_2964);
  or g3327 (n_3166, wc81, n_2629);
  not gc81 (wc81, n_2624);
  or g3328 (n_3169, wc82, n_2625);
  not gc82 (wc82, n_2626);
  or g3329 (n_3266, wc83, n_2779);
  not gc83 (wc83, n_2774);
  or g3330 (n_3269, wc84, n_2775);
  not gc84 (wc84, n_2776);
  and g3331 (n_2822, wc85, n_2632);
  not gc85 (wc85, n_2633);
  and g3332 (n_2824, wc86, n_2638);
  not gc86 (wc86, n_2639);
  and g3333 (n_2920, wc87, n_2810);
  not gc87 (wc87, n_2811);
  and g3334 (n_2818, wc88, n_2814);
  not gc88 (wc88, n_2815);
  and g3335 (n_2909, wc89, n_2905);
  not gc89 (wc89, n_2906);
  or g3336 (n_3011, wc90, n_2924);
  not gc90 (wc90, n_2964);
  or g3337 (n_3170, wc91, n_2635);
  not gc91 (wc91, n_2630);
  or g3338 (n_3173, wc92, n_2631);
  not gc92 (wc92, n_2632);
  or g3339 (n_3174, wc93, n_2641);
  not gc93 (wc93, n_2636);
  or g3340 (n_3177, wc94, n_2637);
  not gc94 (wc94, n_2638);
  or g3341 (n_3178, wc95, n_2647);
  not gc95 (wc95, n_2642);
  or g3342 (n_3262, wc96, n_2773);
  not gc96 (wc96, n_2768);
  and g3343 (n_2829, wc97, n_2644);
  not gc97 (wc97, n_2645);
  and g3344 (n_2899, wc98, n_2764);
  not gc98 (wc98, n_2765);
  and g3345 (n_2901, wc99, n_2770);
  not gc99 (wc99, n_2771);
  and g3346 (n_2921, wc100, n_2817);
  not gc100 (wc100, n_2818);
  and g3347 (n_2825, wc101, n_2821);
  not gc101 (wc101, n_2822);
  and g3348 (n_2961, wc102, n_2908);
  not gc102 (wc102, n_2909);
  or g3349 (n_3065, wc103, n_2617);
  not gc103 (wc103, n_3063);
  or g3350 (n_3181, wc104, n_2643);
  not gc104 (wc104, n_2644);
  or g3351 (n_3182, wc105, n_2653);
  not gc105 (wc105, n_2648);
  or g3352 (n_3258, wc106, n_2767);
  not gc106 (wc106, n_2762);
  or g3353 (n_3261, wc107, n_2763);
  not gc107 (wc107, n_2764);
  or g3354 (n_3265, wc108, n_2769);
  not gc108 (wc108, n_2770);
  and g3355 (n_2831, wc109, n_2650);
  not gc109 (wc109, n_2651);
  and g3356 (n_2836, wc110, n_2656);
  not gc110 (wc110, n_2657);
  and g3357 (n_2838, wc111, n_2662);
  not gc111 (wc111, n_2663);
  and g3358 (n_2843, wc112, n_2668);
  not gc112 (wc112, n_2669);
  and g3359 (n_2845, wc113, n_2674);
  not gc113 (wc113, n_2675);
  and g3360 (n_2850, wc114, n_2680);
  not gc114 (wc114, n_2681);
  and g3361 (n_2852, wc115, n_2686);
  not gc115 (wc115, n_2687);
  and g3362 (n_2857, wc116, n_2692);
  not gc116 (wc116, n_2693);
  and g3363 (n_2859, wc117, n_2698);
  not gc117 (wc117, n_2699);
  and g3364 (n_2864, wc118, n_2704);
  not gc118 (wc118, n_2705);
  and g3365 (n_2866, wc119, n_2710);
  not gc119 (wc119, n_2711);
  and g3366 (n_2871, wc120, n_2716);
  not gc120 (wc120, n_2717);
  and g3367 (n_2873, wc121, n_2722);
  not gc121 (wc121, n_2723);
  and g3368 (n_2878, wc122, n_2728);
  not gc122 (wc122, n_2729);
  and g3369 (n_2880, wc123, n_2734);
  not gc123 (wc123, n_2735);
  and g3370 (n_2885, wc124, n_2740);
  not gc124 (wc124, n_2741);
  and g3371 (n_2926, wc125, n_2824);
  not gc125 (wc125, n_2825);
  and g3372 (n_2902, wc126, n_2898);
  not gc126 (wc126, n_2899);
  or g3373 (n_3067, wc127, n_2623);
  not gc127 (wc127, n_3031);
  or g3374 (n_3185, wc128, n_2649);
  not gc128 (wc128, n_2650);
  or g3375 (n_3186, wc129, n_2659);
  not gc129 (wc129, n_2654);
  or g3376 (n_3189, wc130, n_2655);
  not gc130 (wc130, n_2656);
  or g3377 (n_3190, wc131, n_2665);
  not gc131 (wc131, n_2660);
  or g3378 (n_3193, wc132, n_2661);
  not gc132 (wc132, n_2662);
  or g3379 (n_3194, wc133, n_2671);
  not gc133 (wc133, n_2666);
  or g3380 (n_3197, wc134, n_2667);
  not gc134 (wc134, n_2668);
  or g3381 (n_3198, wc135, n_2677);
  not gc135 (wc135, n_2672);
  or g3382 (n_3201, wc136, n_2673);
  not gc136 (wc136, n_2674);
  or g3383 (n_3202, wc137, n_2683);
  not gc137 (wc137, n_2678);
  or g3384 (n_3205, wc138, n_2679);
  not gc138 (wc138, n_2680);
  or g3385 (n_3206, wc139, n_2689);
  not gc139 (wc139, n_2684);
  or g3386 (n_3209, wc140, n_2685);
  not gc140 (wc140, n_2686);
  or g3387 (n_3210, wc141, n_2695);
  not gc141 (wc141, n_2690);
  or g3388 (n_3213, wc142, n_2691);
  not gc142 (wc142, n_2692);
  or g3389 (n_3214, wc143, n_2701);
  not gc143 (wc143, n_2696);
  or g3390 (n_3217, wc144, n_2697);
  not gc144 (wc144, n_2698);
  or g3391 (n_3218, wc145, n_2707);
  not gc145 (wc145, n_2702);
  or g3392 (n_3221, wc146, n_2703);
  not gc146 (wc146, n_2704);
  or g3393 (n_3222, wc147, n_2713);
  not gc147 (wc147, n_2708);
  or g3394 (n_3225, wc148, n_2709);
  not gc148 (wc148, n_2710);
  or g3395 (n_3226, wc149, n_2719);
  not gc149 (wc149, n_2714);
  or g3396 (n_3229, wc150, n_2715);
  not gc150 (wc150, n_2716);
  or g3397 (n_3230, wc151, n_2725);
  not gc151 (wc151, n_2720);
  or g3398 (n_3233, wc152, n_2721);
  not gc152 (wc152, n_2722);
  or g3399 (n_3234, wc153, n_2731);
  not gc153 (wc153, n_2726);
  or g3400 (n_3237, wc154, n_2727);
  not gc154 (wc154, n_2728);
  or g3401 (n_3238, wc155, n_2737);
  not gc155 (wc155, n_2732);
  or g3402 (n_3241, wc156, n_2733);
  not gc156 (wc156, n_2734);
  or g3403 (n_3242, wc157, n_2743);
  not gc157 (wc157, n_2738);
  or g3404 (n_3245, wc158, n_2739);
  not gc158 (wc158, n_2740);
  and g3405 (n_2887, wc159, n_2746);
  not gc159 (wc159, n_2747);
  and g3406 (n_2894, wc160, n_2758);
  not gc160 (wc160, n_2759);
  and g3407 (n_2832, wc161, n_2828);
  not gc161 (wc161, n_2829);
  and g3408 (n_2839, wc162, n_2835);
  not gc162 (wc162, n_2836);
  and g3409 (n_2846, wc163, n_2842);
  not gc163 (wc163, n_2843);
  and g3410 (n_2853, wc164, n_2849);
  not gc164 (wc164, n_2850);
  and g3411 (n_2860, wc165, n_2856);
  not gc165 (wc165, n_2857);
  and g3412 (n_2867, wc166, n_2863);
  not gc166 (wc166, n_2864);
  and g3413 (n_2874, wc167, n_2870);
  not gc167 (wc167, n_2871);
  and g3414 (n_2881, wc168, n_2877);
  not gc168 (wc168, n_2878);
  and g3415 (n_2957, wc169, n_2901);
  not gc169 (wc169, n_2902);
  and g3416 (n_2965, n_2921, wc170);
  not gc170 (wc170, n_2922);
  or g3417 (n_3246, wc171, n_2749);
  not gc171 (wc171, n_2744);
  or g3418 (n_3249, wc172, n_2745);
  not gc172 (wc172, n_2746);
  or g3419 (n_3254, wc173, n_2761);
  not gc173 (wc173, n_2756);
  or g3420 (n_3257, wc174, n_2757);
  not gc174 (wc174, n_2758);
  and g3421 (n_2892, wc175, n_2752);
  not gc175 (wc175, n_2753);
  and g3422 (n_2927, wc176, n_2831);
  not gc176 (wc176, n_2832);
  and g3423 (n_2932, wc177, n_2838);
  not gc177 (wc177, n_2839);
  and g3424 (n_2933, wc178, n_2845);
  not gc178 (wc178, n_2846);
  and g3425 (n_2938, wc179, n_2852);
  not gc179 (wc179, n_2853);
  and g3426 (n_2939, wc180, n_2859);
  not gc180 (wc180, n_2860);
  and g3427 (n_2944, wc181, n_2866);
  not gc181 (wc181, n_2867);
  and g3428 (n_2945, wc182, n_2873);
  not gc182 (wc182, n_2874);
  and g3429 (n_2950, wc183, n_2880);
  not gc183 (wc183, n_2881);
  and g3430 (n_2888, wc184, n_2884);
  not gc184 (wc184, n_2885);
  or g3431 (n_3070, wc185, n_2629);
  not gc185 (wc185, n_3068);
  or g3432 (n_3250, wc186, n_2755);
  not gc186 (wc186, n_2750);
  or g3433 (n_3253, wc187, n_2751);
  not gc187 (wc187, n_2752);
  and g3434 (n_2951, wc188, n_2887);
  not gc188 (wc188, n_2888);
  and g3435 (n_2895, wc189, n_2891);
  not gc189 (wc189, n_2892);
  or g3436 (n_3013, wc190, n_2930);
  not gc190 (wc190, n_2989);
  or g3437 (n_3072, wc191, n_2635);
  not gc191 (wc191, n_2989);
  and g3438 (n_2956, wc192, n_2894);
  not gc192 (wc192, n_2895);
  and g3439 (n_2968, n_2927, wc193);
  not gc193 (wc193, n_2928);
  and g3440 (n_2970, n_2933, wc194);
  not gc194 (wc194, n_2934);
  and g3441 (n_2975, n_2939, wc195);
  not gc195 (wc195, n_2940);
  and g3442 (n_2977, n_2945, wc196);
  not gc196 (wc196, n_2946);
  or g3443 (n_2992, n_2988, wc197);
  not gc197 (wc197, n_2989);
  and g3444 (n_2982, n_2951, wc198);
  not gc198 (wc198, n_2952);
  and g3445 (n_2971, wc199, n_2967);
  not gc199 (wc199, n_2968);
  and g3446 (n_2978, wc200, n_2974);
  not gc200 (wc200, n_2975);
  or g3447 (n_3075, wc201, n_2641);
  not gc201 (wc201, n_3073);
  or g3448 (n_3077, wc202, n_2647);
  not gc202 (wc202, n_3034);
  and g3449 (n_2984, n_2957, wc203);
  not gc203 (wc203, n_2958);
  and g3450 (n_2991, wc204, n_2970);
  not gc204 (wc204, n_2971);
  and g3451 (n_2994, wc205, n_2977);
  not gc205 (wc205, n_2978);
  and g3452 (n_2985, wc206, n_2981);
  not gc206 (wc206, n_2982);
  or g3453 (n_3016, wc207, n_2936);
  not gc207 (wc207, n_3014);
  or g3454 (n_3082, wc208, n_2659);
  not gc208 (wc208, n_3014);
  or g3455 (n_3080, wc209, n_2653);
  not gc209 (wc209, n_3078);
  and g3456 (n_2995, wc210, n_2984);
  not gc210 (wc210, n_2985);
  or g3457 (n_3004, wc211, n_2998);
  not gc211 (wc211, n_3000);
  or g3458 (n_3018, wc212, n_2942);
  not gc212 (wc212, n_3000);
  or g3459 (n_3085, wc213, n_2665);
  not gc213 (wc213, n_3083);
  or g3460 (n_3087, wc214, n_2671);
  not gc214 (wc214, n_3037);
  or g3461 (n_3092, wc215, n_2683);
  not gc215 (wc215, n_3000);
  and g3462 (n_3001, n_2995, wc216);
  not gc216 (wc216, n_2996);
  or g3463 (n_3021, wc217, n_2948);
  not gc217 (wc217, n_3019);
  or g3464 (n_3023, wc218, n_2954);
  not gc218 (wc218, n_3007);
  or g3465 (n_3090, wc219, n_2677);
  not gc219 (wc219, n_3088);
  or g3466 (n_3095, wc220, n_2689);
  not gc220 (wc220, n_3093);
  or g3467 (n_3097, wc221, n_2695);
  not gc221 (wc221, n_3040);
  or g3468 (n_3102, wc222, n_2707);
  not gc222 (wc222, n_3019);
  or g3469 (n_3112, wc223, n_2731);
  not gc223 (wc223, n_3007);
  or g3470 (n_3026, wc224, n_2960);
  not gc224 (wc224, n_3024);
  or g3471 (n_3028, wc225, n_2962);
  not gc225 (wc225, n_3009);
  or g3472 (n_3100, wc226, n_2701);
  not gc226 (wc226, n_3098);
  or g3473 (n_3105, wc227, n_2713);
  not gc227 (wc227, n_3103);
  or g3474 (n_3107, wc228, n_2719);
  not gc228 (wc228, n_3043);
  or g3475 (n_3115, wc229, n_2737);
  not gc229 (wc229, n_3113);
  or g3476 (n_3117, wc230, n_2743);
  not gc230 (wc230, n_3046);
  or g3477 (n_3122, wc231, n_2755);
  not gc231 (wc231, n_3024);
  or g3478 (n_3132, wc232, n_2779);
  not gc232 (wc232, n_3009);
  or g3479 (n_3110, wc233, n_2725);
  not gc233 (wc233, n_3108);
  or g3480 (n_3120, wc234, n_2749);
  not gc234 (wc234, n_3118);
  or g3481 (n_3125, wc235, n_2761);
  not gc235 (wc235, n_3123);
  or g3482 (n_3127, wc236, n_2767);
  not gc236 (wc236, n_3049);
  or g3483 (n_3135, wc237, n_2785);
  not gc237 (wc237, n_3133);
  or g3484 (n_3137, wc238, n_2791);
  not gc238 (wc238, n_3052);
  or g3485 (n_3130, wc239, n_2773);
  not gc239 (wc239, n_3128);
  or g3486 (n_3140, n_2795, wc240);
  not gc240 (wc240, n_3138);
  not g3487 (Z[71], n_3280);
endmodule

module mult_signed_const_11946_GENERIC(A, Z);
  input [52:0] A;
  output [71:0] Z;
  wire [52:0] A;
  wire [71:0] Z;
  mult_signed_const_11946_GENERIC_REAL g1(.A ({A[52:2], A[0], A[0]}),
       .Z (Z));
endmodule

module mult_signed_const_12373_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [53:0] A;
  output [72:0] Z;
  wire [53:0] A;
  wire [72:0] Z;
  wire n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_275, n_276, n_277, n_278, n_279, n_280;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593;
  wire n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601;
  wire n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609;
  wire n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617;
  wire n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681;
  wire n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697;
  wire n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705;
  wire n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721;
  wire n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729;
  wire n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737;
  wire n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745;
  wire n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753;
  wire n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761;
  wire n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769;
  wire n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777;
  wire n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785;
  wire n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793;
  wire n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801;
  wire n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809;
  wire n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817;
  wire n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825;
  wire n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833;
  wire n_834, n_835, n_838, n_839, n_840, n_841, n_842, n_843;
  wire n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851;
  wire n_855, n_856, n_858, n_859, n_860, n_861, n_862, n_863;
  wire n_864, n_865, n_866, n_867, n_868, n_870, n_871, n_872;
  wire n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882;
  wire n_883, n_886, n_887, n_890, n_891, n_892, n_893, n_894;
  wire n_895, n_896, n_897, n_898, n_900, n_902, n_904, n_905;
  wire n_906, n_907, n_908, n_909, n_910, n_911, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_926, n_928, n_929, n_930, n_931, n_932, n_933, n_934;
  wire n_935, n_938, n_940, n_941, n_942, n_943, n_944, n_945;
  wire n_946, n_948, n_950, n_951, n_952, n_953, n_954, n_955;
  wire n_959, n_960, n_961, n_962, n_963, n_964, n_967, n_968;
  wire n_969, n_970, n_971, n_975, n_976, n_977, n_978, n_980;
  wire n_981, n_982, n_983, n_986, n_987, n_988, n_990, n_991;
  wire n_994, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003;
  wire n_1004, n_1005, n_1006, n_1008, n_1009, n_1010, n_1011, n_1012;
  wire n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023;
  wire n_1024, n_1025, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1035, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042;
  wire n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1053;
  wire n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1063;
  wire n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074;
  wire n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1085;
  wire n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093;
  wire n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1101, n_1102;
  wire n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111;
  wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119;
  wire n_1120, n_1121, n_1124, n_1127, n_1128, n_1129, n_1130, n_1131;
  wire n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139;
  wire n_1140, n_1141, n_1144, n_1145, n_1146, n_1147, n_1149, n_1150;
  wire n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158;
  wire n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166;
  wire n_1167, n_1168, n_1169, n_1171, n_1173, n_1176, n_1177, n_1178;
  wire n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186;
  wire n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194;
  wire n_1196, n_1197, n_1199, n_1200, n_1203, n_1204, n_1205, n_1206;
  wire n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214;
  wire n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222;
  wire n_1223, n_1224, n_1227, n_1229, n_1230, n_1233, n_1234, n_1235;
  wire n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243;
  wire n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251;
  wire n_1252, n_1253, n_1254, n_1255, n_1256, n_1261, n_1262, n_1263;
  wire n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272;
  wire n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280;
  wire n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288;
  wire n_1293, n_1294, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302;
  wire n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310;
  wire n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318;
  wire n_1319, n_1320, n_1323, n_1324, n_1325, n_1326, n_1327, n_1329;
  wire n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337;
  wire n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345;
  wire n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1355;
  wire n_1357, n_1358, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366;
  wire n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374;
  wire n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382;
  wire n_1383, n_1384, n_1387, n_1389, n_1390, n_1393, n_1394, n_1395;
  wire n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403;
  wire n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411;
  wire n_1412, n_1413, n_1414, n_1415, n_1416, n_1419, n_1421, n_1422;
  wire n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432;
  wire n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440;
  wire n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448;
  wire n_1451, n_1453, n_1454, n_1457, n_1458, n_1459, n_1460, n_1461;
  wire n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469;
  wire n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477;
  wire n_1478, n_1479, n_1480, n_1483, n_1485, n_1486, n_1489, n_1490;
  wire n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498;
  wire n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506;
  wire n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1515, n_1517;
  wire n_1518, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527;
  wire n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535;
  wire n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543;
  wire n_1544, n_1547, n_1549, n_1550, n_1553, n_1554, n_1555, n_1556;
  wire n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564;
  wire n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572;
  wire n_1573, n_1574, n_1575, n_1576, n_1579, n_1581, n_1582, n_1585;
  wire n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593;
  wire n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601;
  wire n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1611;
  wire n_1613, n_1614, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622;
  wire n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630;
  wire n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638;
  wire n_1639, n_1640, n_1643, n_1645, n_1646, n_1649, n_1650, n_1651;
  wire n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659;
  wire n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667;
  wire n_1668, n_1669, n_1670, n_1671, n_1672, n_1675, n_1677, n_1678;
  wire n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688;
  wire n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696;
  wire n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704;
  wire n_1707, n_1709, n_1710, n_1713, n_1714, n_1715, n_1716, n_1717;
  wire n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725;
  wire n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733;
  wire n_1734, n_1735, n_1736, n_1739, n_1741, n_1742, n_1745, n_1746;
  wire n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754;
  wire n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762;
  wire n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1771, n_1773;
  wire n_1774, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
  wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1803, n_1805, n_1806, n_1809, n_1810, n_1811, n_1812;
  wire n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820;
  wire n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
  wire n_1829, n_1830, n_1831, n_1832, n_1835, n_1837, n_1838, n_1841;
  wire n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849;
  wire n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857;
  wire n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1867;
  wire n_1869, n_1870, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878;
  wire n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886;
  wire n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894;
  wire n_1895, n_1896, n_1899, n_1901, n_1902, n_1905, n_1906, n_1907;
  wire n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915;
  wire n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923;
  wire n_1924, n_1925, n_1926, n_1927, n_1928, n_1931, n_1933, n_1934;
  wire n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944;
  wire n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952;
  wire n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960;
  wire n_1963, n_1965, n_1966, n_1969, n_1970, n_1971, n_1972, n_1973;
  wire n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981;
  wire n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989;
  wire n_1990, n_1991, n_1992, n_1995, n_1997, n_1998, n_2001, n_2002;
  wire n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010;
  wire n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018;
  wire n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2027, n_2029;
  wire n_2030, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039;
  wire n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047;
  wire n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055;
  wire n_2056, n_2059, n_2061, n_2062, n_2065, n_2066, n_2067, n_2068;
  wire n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076;
  wire n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084;
  wire n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2093;
  wire n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103;
  wire n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111;
  wire n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119;
  wire n_2120, n_2121, n_2122, n_2123, n_2125, n_2128, n_2129, n_2130;
  wire n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138;
  wire n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146;
  wire n_2147, n_2148, n_2152, n_2153, n_2155, n_2159, n_2160, n_2161;
  wire n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169;
  wire n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177;
  wire n_2178, n_2179, n_2180, n_2184, n_2185, n_2187, n_2191, n_2192;
  wire n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200;
  wire n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208;
  wire n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216;
  wire n_2217, n_2219, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228;
  wire n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236;
  wire n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244;
  wire n_2245, n_2246, n_2247, n_2248, n_2249, n_2251, n_2255, n_2256;
  wire n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264;
  wire n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272;
  wire n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280;
  wire n_2281, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293;
  wire n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301;
  wire n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309;
  wire n_2310, n_2312, n_2313, n_2314, n_2319, n_2320, n_2321, n_2322;
  wire n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330;
  wire n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338;
  wire n_2339, n_2340, n_2343, n_2344, n_2345, n_2346, n_2353, n_2354;
  wire n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362;
  wire n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370;
  wire n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2379;
  wire n_2380, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391;
  wire n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399;
  wire n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2413, n_2414;
  wire n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422;
  wire n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430;
  wire n_2431, n_2432, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446;
  wire n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454;
  wire n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2464, n_2465;
  wire n_2467, n_2469, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476;
  wire n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484;
  wire n_2493, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501;
  wire n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2511;
  wire n_2513, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521;
  wire n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2533;
  wire n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543;
  wire n_2544, n_2545, n_2546, n_2547, n_2548, n_2551, n_2552, n_2555;
  wire n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563;
  wire n_2564, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577;
  wire n_2578, n_2579, n_2580, n_2581, n_2582, n_2584, n_2585, n_2586;
  wire n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2595, n_2596;
  wire n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2608;
  wire n_2609, n_2610, n_2611, n_2612, n_2615, n_2616, n_2617, n_2618;
  wire n_2619, n_2620, n_2622, n_2623, n_2624, n_2627, n_2628, n_2640;
  wire n_2642, n_2644, n_2645, n_2646, n_2647, n_2648, n_2650, n_2651;
  wire n_2652, n_2653, n_2654, n_2656, n_2657, n_2658, n_2659, n_2660;
  wire n_2662, n_2663, n_2664, n_2665, n_2666, n_2668, n_2669, n_2670;
  wire n_2671, n_2672, n_2674, n_2675, n_2676, n_2677, n_2678, n_2680;
  wire n_2681, n_2682, n_2683, n_2684, n_2686, n_2687, n_2688, n_2689;
  wire n_2690, n_2692, n_2693, n_2694, n_2695, n_2696, n_2698, n_2699;
  wire n_2700, n_2701, n_2702, n_2704, n_2705, n_2706, n_2707, n_2708;
  wire n_2710, n_2711, n_2712, n_2713, n_2714, n_2716, n_2717, n_2718;
  wire n_2719, n_2720, n_2722, n_2723, n_2724, n_2725, n_2726, n_2728;
  wire n_2729, n_2730, n_2731, n_2732, n_2734, n_2735, n_2736, n_2737;
  wire n_2738, n_2740, n_2741, n_2742, n_2743, n_2744, n_2746, n_2747;
  wire n_2748, n_2749, n_2750, n_2752, n_2753, n_2754, n_2755, n_2756;
  wire n_2758, n_2759, n_2760, n_2761, n_2762, n_2764, n_2765, n_2766;
  wire n_2767, n_2768, n_2770, n_2771, n_2772, n_2773, n_2774, n_2776;
  wire n_2777, n_2778, n_2779, n_2780, n_2782, n_2783, n_2784, n_2785;
  wire n_2786, n_2788, n_2789, n_2790, n_2791, n_2792, n_2794, n_2795;
  wire n_2796, n_2797, n_2798, n_2800, n_2801, n_2802, n_2803, n_2804;
  wire n_2806, n_2807, n_2808, n_2809, n_2810, n_2812, n_2813, n_2814;
  wire n_2815, n_2816, n_2818, n_2819, n_2820, n_2821, n_2822, n_2824;
  wire n_2825, n_2826, n_2827, n_2828, n_2830, n_2831, n_2832, n_2833;
  wire n_2834, n_2836, n_2837, n_2838, n_2839, n_2840, n_2842, n_2843;
  wire n_2844, n_2845, n_2846, n_2848, n_2851, n_2853, n_2854, n_2856;
  wire n_2857, n_2859, n_2860, n_2861, n_2863, n_2864, n_2866, n_2867;
  wire n_2868, n_2870, n_2871, n_2873, n_2874, n_2875, n_2877, n_2878;
  wire n_2880, n_2881, n_2882, n_2884, n_2885, n_2887, n_2888, n_2889;
  wire n_2891, n_2892, n_2894, n_2895, n_2896, n_2898, n_2899, n_2901;
  wire n_2902, n_2903, n_2905, n_2906, n_2908, n_2909, n_2910, n_2912;
  wire n_2913, n_2915, n_2916, n_2917, n_2919, n_2920, n_2922, n_2923;
  wire n_2924, n_2926, n_2927, n_2929, n_2930, n_2931, n_2933, n_2934;
  wire n_2936, n_2937, n_2938, n_2940, n_2941, n_2943, n_2944, n_2945;
  wire n_2947, n_2948, n_2950, n_2951, n_2952, n_2954, n_2955, n_2957;
  wire n_2958, n_2959, n_2961, n_2962, n_2964, n_2965, n_2966, n_2968;
  wire n_2969, n_2971, n_2972, n_2975, n_2976, n_2977, n_2978, n_2979;
  wire n_2980, n_2982, n_2983, n_2984, n_2985, n_2986, n_2988, n_2989;
  wire n_2990, n_2991, n_2992, n_2994, n_2995, n_2996, n_2997, n_2998;
  wire n_3000, n_3001, n_3002, n_3003, n_3004, n_3006, n_3007, n_3008;
  wire n_3009, n_3010, n_3012, n_3013, n_3014, n_3015, n_3016, n_3018;
  wire n_3019, n_3020, n_3021, n_3022, n_3024, n_3025, n_3026, n_3027;
  wire n_3028, n_3029, n_3030, n_3032, n_3033, n_3035, n_3036, n_3037;
  wire n_3039, n_3040, n_3042, n_3043, n_3044, n_3046, n_3047, n_3049;
  wire n_3050, n_3051, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058;
  wire n_3060, n_3061, n_3062, n_3063, n_3064, n_3066, n_3067, n_3068;
  wire n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3076, n_3078;
  wire n_3079, n_3081, n_3083, n_3084, n_3086, n_3088, n_3089, n_3091;
  wire n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100;
  wire n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108;
  wire n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116;
  wire n_3117, n_3118, n_3122, n_3123, n_3125, n_3127, n_3128, n_3130;
  wire n_3132, n_3133, n_3135, n_3137, n_3138, n_3140, n_3142, n_3143;
  wire n_3145, n_3147, n_3148, n_3150, n_3152, n_3153, n_3155, n_3157;
  wire n_3158, n_3160, n_3162, n_3163, n_3165, n_3167, n_3168, n_3170;
  wire n_3172, n_3173, n_3175, n_3177, n_3178, n_3180, n_3182, n_3183;
  wire n_3185, n_3187, n_3188, n_3190, n_3192, n_3193, n_3195, n_3197;
  wire n_3198, n_3200, n_3202, n_3203, n_3205, n_3207, n_3211, n_3214;
  wire n_3215, n_3217, n_3218, n_3219, n_3221, n_3222, n_3223, n_3225;
  wire n_3226, n_3227, n_3229, n_3230, n_3231, n_3233, n_3234, n_3235;
  wire n_3237, n_3238, n_3239, n_3241, n_3242, n_3243, n_3245, n_3246;
  wire n_3247, n_3249, n_3250, n_3251, n_3253, n_3254, n_3255, n_3257;
  wire n_3258, n_3259, n_3261, n_3262, n_3263, n_3265, n_3266, n_3267;
  wire n_3269, n_3270, n_3271, n_3273, n_3274, n_3275, n_3277, n_3278;
  wire n_3279, n_3281, n_3282, n_3283, n_3285, n_3286, n_3287, n_3289;
  wire n_3290, n_3291, n_3293, n_3294, n_3295, n_3297, n_3298, n_3299;
  wire n_3301, n_3302, n_3303, n_3305, n_3306, n_3307, n_3309, n_3310;
  wire n_3311, n_3313, n_3314, n_3315, n_3317, n_3318, n_3319, n_3321;
  wire n_3322, n_3323, n_3325, n_3326, n_3327, n_3329, n_3330, n_3331;
  wire n_3333, n_3334, n_3335, n_3337, n_3338, n_3339, n_3341, n_3342;
  wire n_3343, n_3345, n_3346, n_3347, n_3349, n_3350;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g428 (n_196, A[4], A[0]);
  and g2 (n_122, A[4], A[0]);
  xor g429 (n_997, A[5], A[3]);
  xor g430 (n_195, n_997, A[1]);
  nand g3 (n_998, A[5], A[3]);
  nand g431 (n_999, A[1], A[3]);
  nand g432 (n_1000, A[5], A[1]);
  nand g433 (n_121, n_998, n_999, n_1000);
  xor g434 (n_275, A[6], A[4]);
  and g435 (n_276, A[6], A[4]);
  xor g436 (n_1001, A[0], A[2]);
  xor g437 (n_194, n_1001, n_275);
  nand g438 (n_1002, A[0], A[2]);
  nand g4 (n_1003, n_275, A[2]);
  nand g5 (n_1004, A[0], n_275);
  nand g439 (n_120, n_1002, n_1003, n_1004);
  xor g440 (n_1005, A[7], A[5]);
  xor g441 (n_277, n_1005, A[1]);
  nand g442 (n_1006, A[7], A[5]);
  nand g444 (n_1008, A[7], A[1]);
  nand g6 (n_279, n_1006, n_1000, n_1008);
  xor g445 (n_1009, A[3], n_276);
  xor g446 (n_193, n_1009, n_277);
  nand g447 (n_1010, A[3], n_276);
  nand g448 (n_1011, n_277, n_276);
  nand g449 (n_1012, A[3], n_277);
  nand g450 (n_119, n_1010, n_1011, n_1012);
  xor g451 (n_278, A[8], A[6]);
  and g452 (n_281, A[8], A[6]);
  xor g454 (n_280, n_1001, A[4]);
  nand g457 (n_1016, A[2], A[4]);
  xor g459 (n_1017, n_278, n_279);
  xor g460 (n_192, n_1017, n_280);
  nand g461 (n_1018, n_278, n_279);
  nand g462 (n_1019, n_280, n_279);
  nand g463 (n_1020, n_278, n_280);
  nand g464 (n_118, n_1018, n_1019, n_1020);
  xor g465 (n_1021, A[9], A[7]);
  xor g466 (n_283, n_1021, A[3]);
  nand g467 (n_1022, A[9], A[7]);
  nand g468 (n_1023, A[3], A[7]);
  nand g469 (n_1024, A[9], A[3]);
  nand g470 (n_286, n_1022, n_1023, n_1024);
  xor g471 (n_1025, A[1], A[5]);
  xor g472 (n_284, n_1025, n_281);
  nand g474 (n_1027, n_281, A[5]);
  nand g475 (n_1028, A[1], n_281);
  nand g476 (n_288, n_1000, n_1027, n_1028);
  xor g477 (n_1029, n_282, n_283);
  xor g478 (n_191, n_1029, n_284);
  nand g479 (n_1030, n_282, n_283);
  nand g480 (n_1031, n_284, n_283);
  nand g481 (n_1032, n_282, n_284);
  nand g482 (n_117, n_1030, n_1031, n_1032);
  xor g483 (n_285, A[10], A[8]);
  and g484 (n_290, A[10], A[8]);
  xor g485 (n_1033, A[4], A[2]);
  xor g486 (n_287, n_1033, A[6]);
  nand g488 (n_1035, A[6], A[2]);
  xor g491 (n_1037, A[0], n_285);
  xor g492 (n_289, n_1037, n_286);
  nand g493 (n_1038, A[0], n_285);
  nand g494 (n_1039, n_286, n_285);
  nand g495 (n_1040, A[0], n_286);
  nand g496 (n_294, n_1038, n_1039, n_1040);
  xor g497 (n_1041, n_287, n_288);
  xor g498 (n_190, n_1041, n_289);
  nand g499 (n_1042, n_287, n_288);
  nand g500 (n_1043, n_289, n_288);
  nand g501 (n_1044, n_287, n_289);
  nand g502 (n_116, n_1042, n_1043, n_1044);
  xor g503 (n_1045, A[11], A[9]);
  xor g504 (n_292, n_1045, A[5]);
  nand g505 (n_1046, A[11], A[9]);
  nand g506 (n_1047, A[5], A[9]);
  nand g507 (n_1048, A[11], A[5]);
  nand g508 (n_297, n_1046, n_1047, n_1048);
  xor g509 (n_1049, A[3], A[7]);
  xor g510 (n_293, n_1049, A[1]);
  nand g514 (n_298, n_1023, n_1008, n_999);
  xor g515 (n_1053, n_290, n_291);
  xor g516 (n_295, n_1053, n_292);
  nand g517 (n_1054, n_290, n_291);
  nand g518 (n_1055, n_292, n_291);
  nand g519 (n_1056, n_290, n_292);
  nand g520 (n_302, n_1054, n_1055, n_1056);
  xor g521 (n_1057, n_293, n_294);
  xor g522 (n_189, n_1057, n_295);
  nand g523 (n_1058, n_293, n_294);
  nand g524 (n_1059, n_295, n_294);
  nand g525 (n_1060, n_293, n_295);
  nand g526 (n_115, n_1058, n_1059, n_1060);
  xor g527 (n_296, A[12], A[10]);
  and g528 (n_303, A[12], A[10]);
  xor g530 (n_299, n_275, A[8]);
  nand g532 (n_1063, A[8], A[4]);
  xor g536 (n_300, n_1001, n_296);
  nand g538 (n_1067, n_296, A[0]);
  nand g539 (n_1068, A[2], n_296);
  nand g540 (n_307, n_1002, n_1067, n_1068);
  xor g541 (n_1069, n_297, n_298);
  xor g542 (n_301, n_1069, n_299);
  nand g543 (n_1070, n_297, n_298);
  nand g544 (n_1071, n_299, n_298);
  nand g545 (n_1072, n_297, n_299);
  nand g546 (n_309, n_1070, n_1071, n_1072);
  xor g547 (n_1073, n_300, n_301);
  xor g548 (n_188, n_1073, n_302);
  nand g549 (n_1074, n_300, n_301);
  nand g550 (n_1075, n_302, n_301);
  nand g551 (n_1076, n_300, n_302);
  nand g552 (n_114, n_1074, n_1075, n_1076);
  xor g553 (n_1077, A[13], A[11]);
  xor g554 (n_306, n_1077, A[7]);
  nand g555 (n_1078, A[13], A[11]);
  nand g556 (n_1079, A[7], A[11]);
  nand g557 (n_1080, A[13], A[7]);
  nand g558 (n_312, n_1078, n_1079, n_1080);
  xor g559 (n_1081, A[5], A[9]);
  xor g560 (n_305, n_1081, A[3]);
  nand g564 (n_313, n_1047, n_1024, n_998);
  xor g565 (n_1085, A[1], n_303);
  xor g566 (n_308, n_1085, n_304);
  nand g567 (n_1086, A[1], n_303);
  nand g568 (n_1087, n_304, n_303);
  nand g569 (n_1088, A[1], n_304);
  nand g570 (n_316, n_1086, n_1087, n_1088);
  xor g571 (n_1089, n_305, n_306);
  xor g572 (n_310, n_1089, n_307);
  nand g573 (n_1090, n_305, n_306);
  nand g574 (n_1091, n_307, n_306);
  nand g575 (n_1092, n_305, n_307);
  nand g576 (n_318, n_1090, n_1091, n_1092);
  xor g577 (n_1093, n_308, n_309);
  xor g578 (n_187, n_1093, n_310);
  nand g579 (n_1094, n_308, n_309);
  nand g580 (n_1095, n_310, n_309);
  nand g581 (n_1096, n_308, n_310);
  nand g582 (n_113, n_1094, n_1095, n_1096);
  xor g583 (n_311, A[14], A[12]);
  and g584 (n_320, A[14], A[12]);
  xor g585 (n_1097, A[8], A[0]);
  xor g586 (n_315, n_1097, A[6]);
  nand g587 (n_1098, A[8], A[0]);
  nand g588 (n_1099, A[6], A[0]);
  xor g591 (n_1101, A[10], A[4]);
  xor g592 (n_314, n_1101, A[2]);
  nand g593 (n_1102, A[10], A[4]);
  nand g595 (n_1104, A[10], A[2]);
  nand g596 (n_322, n_1102, n_1016, n_1104);
  xor g597 (n_1105, n_311, n_312);
  xor g598 (n_317, n_1105, n_313);
  nand g599 (n_1106, n_311, n_312);
  nand g600 (n_1107, n_313, n_312);
  nand g601 (n_1108, n_311, n_313);
  nand g602 (n_326, n_1106, n_1107, n_1108);
  xor g603 (n_1109, n_314, n_315);
  xor g604 (n_319, n_1109, n_316);
  nand g605 (n_1110, n_314, n_315);
  nand g606 (n_1111, n_316, n_315);
  nand g607 (n_1112, n_314, n_316);
  nand g608 (n_329, n_1110, n_1111, n_1112);
  xor g609 (n_1113, n_317, n_318);
  xor g610 (n_186, n_1113, n_319);
  nand g611 (n_1114, n_317, n_318);
  nand g612 (n_1115, n_319, n_318);
  nand g613 (n_1116, n_317, n_319);
  nand g614 (n_112, n_1114, n_1115, n_1116);
  xor g615 (n_1117, A[15], A[13]);
  xor g616 (n_323, n_1117, A[9]);
  nand g617 (n_1118, A[15], A[13]);
  nand g618 (n_1119, A[9], A[13]);
  nand g619 (n_1120, A[15], A[9]);
  nand g620 (n_331, n_1118, n_1119, n_1120);
  xor g621 (n_1121, A[1], A[7]);
  xor g622 (n_324, n_1121, A[11]);
  nand g625 (n_1124, A[1], A[11]);
  nand g626 (n_332, n_1008, n_1079, n_1124);
  xor g628 (n_325, n_997, n_320);
  nand g630 (n_1127, n_320, A[3]);
  nand g631 (n_1128, A[5], n_320);
  nand g632 (n_335, n_998, n_1127, n_1128);
  xor g633 (n_1129, n_321, n_322);
  xor g634 (n_327, n_1129, n_323);
  nand g635 (n_1130, n_321, n_322);
  nand g636 (n_1131, n_323, n_322);
  nand g637 (n_1132, n_321, n_323);
  nand g638 (n_337, n_1130, n_1131, n_1132);
  xor g639 (n_1133, n_324, n_325);
  xor g640 (n_328, n_1133, n_326);
  nand g641 (n_1134, n_324, n_325);
  nand g642 (n_1135, n_326, n_325);
  nand g643 (n_1136, n_324, n_326);
  nand g644 (n_339, n_1134, n_1135, n_1136);
  xor g645 (n_1137, n_327, n_328);
  xor g646 (n_185, n_1137, n_329);
  nand g647 (n_1138, n_327, n_328);
  nand g648 (n_1139, n_329, n_328);
  nand g649 (n_1140, n_327, n_329);
  nand g650 (n_111, n_1138, n_1139, n_1140);
  xor g651 (n_330, A[16], A[14]);
  and g652 (n_341, A[16], A[14]);
  xor g653 (n_1141, A[10], A[2]);
  xor g654 (n_334, n_1141, A[0]);
  nand g657 (n_1144, A[10], A[0]);
  nand g658 (n_342, n_1104, n_1002, n_1144);
  xor g659 (n_1145, A[8], A[12]);
  xor g660 (n_333, n_1145, A[6]);
  nand g661 (n_1146, A[8], A[12]);
  nand g662 (n_1147, A[6], A[12]);
  xor g665 (n_1149, A[4], n_330);
  xor g666 (n_336, n_1149, n_331);
  nand g667 (n_1150, A[4], n_330);
  nand g668 (n_1151, n_331, n_330);
  nand g669 (n_1152, A[4], n_331);
  nand g670 (n_347, n_1150, n_1151, n_1152);
  xor g671 (n_1153, n_332, n_333);
  xor g672 (n_338, n_1153, n_334);
  nand g673 (n_1154, n_332, n_333);
  nand g674 (n_1155, n_334, n_333);
  nand g675 (n_1156, n_332, n_334);
  nand g676 (n_349, n_1154, n_1155, n_1156);
  xor g677 (n_1157, n_335, n_336);
  xor g678 (n_340, n_1157, n_337);
  nand g679 (n_1158, n_335, n_336);
  nand g680 (n_1159, n_337, n_336);
  nand g681 (n_1160, n_335, n_337);
  nand g682 (n_351, n_1158, n_1159, n_1160);
  xor g683 (n_1161, n_338, n_339);
  xor g684 (n_184, n_1161, n_340);
  nand g685 (n_1162, n_338, n_339);
  nand g686 (n_1163, n_340, n_339);
  nand g687 (n_1164, n_338, n_340);
  nand g688 (n_110, n_1162, n_1163, n_1164);
  xor g689 (n_1165, A[17], A[15]);
  xor g690 (n_345, n_1165, A[11]);
  nand g691 (n_1166, A[17], A[15]);
  nand g692 (n_1167, A[11], A[15]);
  nand g693 (n_1168, A[17], A[11]);
  nand g694 (n_354, n_1166, n_1167, n_1168);
  xor g695 (n_1169, A[3], A[1]);
  xor g696 (n_346, n_1169, A[9]);
  nand g698 (n_1171, A[9], A[1]);
  nand g700 (n_356, n_999, n_1171, n_1024);
  xor g701 (n_1173, A[13], A[7]);
  xor g702 (n_344, n_1173, A[5]);
  nand g705 (n_1176, A[13], A[5]);
  nand g706 (n_355, n_1080, n_1006, n_1176);
  xor g707 (n_1177, n_341, n_342);
  xor g708 (n_348, n_1177, n_343);
  nand g709 (n_1178, n_341, n_342);
  nand g710 (n_1179, n_343, n_342);
  nand g711 (n_1180, n_341, n_343);
  nand g712 (n_360, n_1178, n_1179, n_1180);
  xor g713 (n_1181, n_344, n_345);
  xor g714 (n_350, n_1181, n_346);
  nand g715 (n_1182, n_344, n_345);
  nand g716 (n_1183, n_346, n_345);
  nand g717 (n_1184, n_344, n_346);
  nand g718 (n_362, n_1182, n_1183, n_1184);
  xor g719 (n_1185, n_347, n_348);
  xor g720 (n_352, n_1185, n_349);
  nand g721 (n_1186, n_347, n_348);
  nand g722 (n_1187, n_349, n_348);
  nand g723 (n_1188, n_347, n_349);
  nand g724 (n_364, n_1186, n_1187, n_1188);
  xor g725 (n_1189, n_350, n_351);
  xor g726 (n_183, n_1189, n_352);
  nand g727 (n_1190, n_350, n_351);
  nand g728 (n_1191, n_352, n_351);
  nand g729 (n_1192, n_350, n_352);
  nand g730 (n_109, n_1190, n_1191, n_1192);
  xor g731 (n_353, A[18], A[16]);
  and g732 (n_366, A[18], A[16]);
  xor g733 (n_1193, A[12], A[4]);
  xor g734 (n_357, n_1193, A[2]);
  nand g735 (n_1194, A[12], A[4]);
  nand g737 (n_1196, A[12], A[2]);
  nand g738 (n_367, n_1194, n_1016, n_1196);
  xor g739 (n_1197, A[10], A[0]);
  xor g740 (n_358, n_1197, A[14]);
  nand g742 (n_1199, A[14], A[0]);
  nand g743 (n_1200, A[10], A[14]);
  nand g744 (n_368, n_1144, n_1199, n_1200);
  xor g746 (n_359, n_278, n_353);
  nand g748 (n_1203, n_353, A[6]);
  nand g749 (n_1204, A[8], n_353);
  xor g751 (n_1205, n_354, n_355);
  xor g752 (n_361, n_1205, n_356);
  nand g753 (n_1206, n_354, n_355);
  nand g754 (n_1207, n_356, n_355);
  nand g755 (n_1208, n_354, n_356);
  nand g756 (n_374, n_1206, n_1207, n_1208);
  xor g757 (n_1209, n_357, n_358);
  xor g758 (n_363, n_1209, n_359);
  nand g759 (n_1210, n_357, n_358);
  nand g760 (n_1211, n_359, n_358);
  nand g761 (n_1212, n_357, n_359);
  nand g762 (n_375, n_1210, n_1211, n_1212);
  xor g763 (n_1213, n_360, n_361);
  xor g764 (n_365, n_1213, n_362);
  nand g765 (n_1214, n_360, n_361);
  nand g766 (n_1215, n_362, n_361);
  nand g767 (n_1216, n_360, n_362);
  nand g768 (n_125, n_1214, n_1215, n_1216);
  xor g769 (n_1217, n_363, n_364);
  xor g770 (n_182, n_1217, n_365);
  nand g771 (n_1218, n_363, n_364);
  nand g772 (n_1219, n_365, n_364);
  nand g773 (n_1220, n_363, n_365);
  nand g774 (n_108, n_1218, n_1219, n_1220);
  xor g775 (n_1221, A[19], A[17]);
  xor g776 (n_370, n_1221, A[13]);
  nand g777 (n_1222, A[19], A[17]);
  nand g778 (n_1223, A[13], A[17]);
  nand g779 (n_1224, A[19], A[13]);
  nand g780 (n_376, n_1222, n_1223, n_1224);
  xor g782 (n_371, n_997, A[11]);
  nand g784 (n_1227, A[11], A[3]);
  nand g786 (n_377, n_998, n_1227, n_1048);
  xor g787 (n_1229, A[1], A[15]);
  xor g788 (n_369, n_1229, A[9]);
  nand g789 (n_1230, A[1], A[15]);
  nand g792 (n_378, n_1230, n_1120, n_1171);
  xor g793 (n_1233, A[7], n_366);
  xor g794 (n_373, n_1233, n_367);
  nand g795 (n_1234, A[7], n_366);
  nand g796 (n_1235, n_367, n_366);
  nand g797 (n_1236, A[7], n_367);
  nand g798 (n_382, n_1234, n_1235, n_1236);
  xor g799 (n_1237, n_368, n_369);
  xor g800 (n_123, n_1237, n_370);
  nand g801 (n_1238, n_368, n_369);
  nand g802 (n_1239, n_370, n_369);
  nand g803 (n_1240, n_368, n_370);
  nand g804 (n_384, n_1238, n_1239, n_1240);
  xor g805 (n_1241, n_371, n_372);
  xor g806 (n_124, n_1241, n_373);
  nand g807 (n_1242, n_371, n_372);
  nand g808 (n_1243, n_373, n_372);
  nand g809 (n_1244, n_371, n_373);
  nand g810 (n_386, n_1242, n_1243, n_1244);
  xor g811 (n_1245, n_374, n_375);
  xor g812 (n_126, n_1245, n_123);
  nand g813 (n_1246, n_374, n_375);
  nand g814 (n_1247, n_123, n_375);
  nand g815 (n_1248, n_374, n_123);
  nand g816 (n_388, n_1246, n_1247, n_1248);
  xor g817 (n_1249, n_124, n_125);
  xor g818 (n_181, n_1249, n_126);
  nand g819 (n_1250, n_124, n_125);
  nand g820 (n_1251, n_126, n_125);
  nand g821 (n_1252, n_124, n_126);
  nand g822 (n_107, n_1250, n_1251, n_1252);
  xor g823 (n_1253, A[20], A[18]);
  xor g824 (n_380, n_1253, A[14]);
  nand g825 (n_1254, A[20], A[18]);
  nand g826 (n_1255, A[14], A[18]);
  nand g827 (n_1256, A[20], A[14]);
  nand g828 (n_390, n_1254, n_1255, n_1256);
  xor g830 (n_381, n_275, A[12]);
  xor g835 (n_1261, A[2], A[16]);
  xor g836 (n_379, n_1261, A[10]);
  nand g837 (n_1262, A[2], A[16]);
  nand g838 (n_1263, A[10], A[16]);
  nand g840 (n_392, n_1262, n_1263, n_1104);
  xor g841 (n_1265, A[8], n_376);
  xor g842 (n_383, n_1265, n_377);
  nand g843 (n_1266, A[8], n_376);
  nand g844 (n_1267, n_377, n_376);
  nand g845 (n_1268, A[8], n_377);
  nand g846 (n_396, n_1266, n_1267, n_1268);
  xor g847 (n_1269, n_378, n_379);
  xor g848 (n_385, n_1269, n_380);
  nand g849 (n_1270, n_378, n_379);
  nand g850 (n_1271, n_380, n_379);
  nand g851 (n_1272, n_378, n_380);
  nand g852 (n_398, n_1270, n_1271, n_1272);
  xor g853 (n_1273, n_381, n_382);
  xor g854 (n_387, n_1273, n_383);
  nand g855 (n_1274, n_381, n_382);
  nand g856 (n_1275, n_383, n_382);
  nand g857 (n_1276, n_381, n_383);
  nand g858 (n_400, n_1274, n_1275, n_1276);
  xor g859 (n_1277, n_384, n_385);
  xor g860 (n_389, n_1277, n_386);
  nand g861 (n_1278, n_384, n_385);
  nand g862 (n_1279, n_386, n_385);
  nand g863 (n_1280, n_384, n_386);
  nand g864 (n_402, n_1278, n_1279, n_1280);
  xor g865 (n_1281, n_387, n_388);
  xor g866 (n_180, n_1281, n_389);
  nand g867 (n_1282, n_387, n_388);
  nand g868 (n_1283, n_389, n_388);
  nand g869 (n_1284, n_387, n_389);
  nand g870 (n_106, n_1282, n_1283, n_1284);
  xor g871 (n_1285, A[21], A[19]);
  xor g872 (n_394, n_1285, A[15]);
  nand g873 (n_1286, A[21], A[19]);
  nand g874 (n_1287, A[15], A[19]);
  nand g875 (n_1288, A[21], A[15]);
  nand g876 (n_404, n_1286, n_1287, n_1288);
  xor g878 (n_395, n_1005, A[13]);
  xor g883 (n_1293, A[3], A[17]);
  xor g884 (n_393, n_1293, A[11]);
  nand g885 (n_1294, A[3], A[17]);
  nand g888 (n_406, n_1294, n_1168, n_1227);
  xor g889 (n_1297, A[9], n_390);
  xor g890 (n_397, n_1297, n_391);
  nand g891 (n_1298, A[9], n_390);
  nand g892 (n_1299, n_391, n_390);
  nand g893 (n_1300, A[9], n_391);
  nand g894 (n_410, n_1298, n_1299, n_1300);
  xor g895 (n_1301, n_392, n_393);
  xor g896 (n_399, n_1301, n_394);
  nand g897 (n_1302, n_392, n_393);
  nand g898 (n_1303, n_394, n_393);
  nand g899 (n_1304, n_392, n_394);
  nand g900 (n_412, n_1302, n_1303, n_1304);
  xor g901 (n_1305, n_395, n_396);
  xor g902 (n_401, n_1305, n_397);
  nand g903 (n_1306, n_395, n_396);
  nand g904 (n_1307, n_397, n_396);
  nand g905 (n_1308, n_395, n_397);
  nand g906 (n_414, n_1306, n_1307, n_1308);
  xor g907 (n_1309, n_398, n_399);
  xor g908 (n_403, n_1309, n_400);
  nand g909 (n_1310, n_398, n_399);
  nand g910 (n_1311, n_400, n_399);
  nand g911 (n_1312, n_398, n_400);
  nand g912 (n_417, n_1310, n_1311, n_1312);
  xor g913 (n_1313, n_401, n_402);
  xor g914 (n_179, n_1313, n_403);
  nand g915 (n_1314, n_401, n_402);
  nand g916 (n_1315, n_403, n_402);
  nand g917 (n_1316, n_401, n_403);
  nand g918 (n_105, n_1314, n_1315, n_1316);
  xor g919 (n_1317, A[22], A[20]);
  xor g920 (n_408, n_1317, A[16]);
  nand g921 (n_1318, A[22], A[20]);
  nand g922 (n_1319, A[16], A[20]);
  nand g923 (n_1320, A[22], A[16]);
  nand g924 (n_418, n_1318, n_1319, n_1320);
  xor g926 (n_409, n_278, A[14]);
  nand g928 (n_1323, A[14], A[6]);
  nand g929 (n_1324, A[8], A[14]);
  xor g931 (n_1325, A[4], A[18]);
  xor g932 (n_407, n_1325, A[12]);
  nand g933 (n_1326, A[4], A[18]);
  nand g934 (n_1327, A[12], A[18]);
  nand g936 (n_420, n_1326, n_1327, n_1194);
  xor g937 (n_1329, A[10], n_404);
  xor g938 (n_411, n_1329, n_355);
  nand g939 (n_1330, A[10], n_404);
  nand g940 (n_1331, n_355, n_404);
  nand g941 (n_1332, A[10], n_355);
  nand g942 (n_424, n_1330, n_1331, n_1332);
  xor g943 (n_1333, n_406, n_407);
  xor g944 (n_413, n_1333, n_408);
  nand g945 (n_1334, n_406, n_407);
  nand g946 (n_1335, n_408, n_407);
  nand g947 (n_1336, n_406, n_408);
  nand g948 (n_426, n_1334, n_1335, n_1336);
  xor g949 (n_1337, n_409, n_410);
  xor g950 (n_415, n_1337, n_411);
  nand g951 (n_1338, n_409, n_410);
  nand g952 (n_1339, n_411, n_410);
  nand g953 (n_1340, n_409, n_411);
  nand g954 (n_428, n_1338, n_1339, n_1340);
  xor g955 (n_1341, n_412, n_413);
  xor g956 (n_416, n_1341, n_414);
  nand g957 (n_1342, n_412, n_413);
  nand g958 (n_1343, n_414, n_413);
  nand g959 (n_1344, n_412, n_414);
  nand g960 (n_431, n_1342, n_1343, n_1344);
  xor g961 (n_1345, n_415, n_416);
  xor g962 (n_178, n_1345, n_417);
  nand g963 (n_1346, n_415, n_416);
  nand g964 (n_1347, n_417, n_416);
  nand g965 (n_1348, n_415, n_417);
  nand g966 (n_104, n_1346, n_1347, n_1348);
  xor g967 (n_1349, A[23], A[21]);
  xor g968 (n_422, n_1349, A[17]);
  nand g969 (n_1350, A[23], A[21]);
  nand g970 (n_1351, A[17], A[21]);
  nand g971 (n_1352, A[23], A[17]);
  nand g972 (n_432, n_1350, n_1351, n_1352);
  xor g974 (n_423, n_1021, A[15]);
  nand g976 (n_1355, A[15], A[7]);
  nand g978 (n_433, n_1022, n_1355, n_1120);
  xor g979 (n_1357, A[5], A[19]);
  xor g980 (n_421, n_1357, A[13]);
  nand g981 (n_1358, A[5], A[19]);
  nand g984 (n_434, n_1358, n_1224, n_1176);
  xor g985 (n_1361, A[11], n_418);
  xor g986 (n_425, n_1361, n_419);
  nand g987 (n_1362, A[11], n_418);
  nand g988 (n_1363, n_419, n_418);
  nand g989 (n_1364, A[11], n_419);
  nand g990 (n_438, n_1362, n_1363, n_1364);
  xor g991 (n_1365, n_420, n_421);
  xor g992 (n_427, n_1365, n_422);
  nand g993 (n_1366, n_420, n_421);
  nand g994 (n_1367, n_422, n_421);
  nand g995 (n_1368, n_420, n_422);
  nand g996 (n_440, n_1366, n_1367, n_1368);
  xor g997 (n_1369, n_423, n_424);
  xor g998 (n_429, n_1369, n_425);
  nand g999 (n_1370, n_423, n_424);
  nand g1000 (n_1371, n_425, n_424);
  nand g1001 (n_1372, n_423, n_425);
  nand g1002 (n_198, n_1370, n_1371, n_1372);
  xor g1003 (n_1373, n_426, n_427);
  xor g1004 (n_430, n_1373, n_428);
  nand g1005 (n_1374, n_426, n_427);
  nand g1006 (n_1375, n_428, n_427);
  nand g1007 (n_1376, n_426, n_428);
  nand g1008 (n_443, n_1374, n_1375, n_1376);
  xor g1009 (n_1377, n_429, n_430);
  xor g1010 (n_177, n_1377, n_431);
  nand g1011 (n_1378, n_429, n_430);
  nand g1012 (n_1379, n_431, n_430);
  nand g1013 (n_1380, n_429, n_431);
  nand g1014 (n_103, n_1378, n_1379, n_1380);
  xor g1015 (n_1381, A[24], A[22]);
  xor g1016 (n_436, n_1381, A[18]);
  nand g1017 (n_1382, A[24], A[22]);
  nand g1018 (n_1383, A[18], A[22]);
  nand g1019 (n_1384, A[24], A[18]);
  nand g1020 (n_444, n_1382, n_1383, n_1384);
  xor g1022 (n_437, n_285, A[16]);
  nand g1024 (n_1387, A[16], A[8]);
  xor g1027 (n_1389, A[6], A[20]);
  xor g1028 (n_435, n_1389, A[14]);
  nand g1029 (n_1390, A[6], A[20]);
  nand g1032 (n_446, n_1390, n_1256, n_1323);
  xor g1033 (n_1393, A[12], n_432);
  xor g1034 (n_439, n_1393, n_433);
  nand g1035 (n_1394, A[12], n_432);
  nand g1036 (n_1395, n_433, n_432);
  nand g1037 (n_1396, A[12], n_433);
  nand g1038 (n_450, n_1394, n_1395, n_1396);
  xor g1039 (n_1397, n_434, n_435);
  xor g1040 (n_197, n_1397, n_436);
  nand g1041 (n_1398, n_434, n_435);
  nand g1042 (n_1399, n_436, n_435);
  nand g1043 (n_1400, n_434, n_436);
  nand g1044 (n_452, n_1398, n_1399, n_1400);
  xor g1045 (n_1401, n_437, n_438);
  xor g1046 (n_441, n_1401, n_439);
  nand g1047 (n_1402, n_437, n_438);
  nand g1048 (n_1403, n_439, n_438);
  nand g1049 (n_1404, n_437, n_439);
  nand g1050 (n_454, n_1402, n_1403, n_1404);
  xor g1051 (n_1405, n_440, n_197);
  xor g1052 (n_442, n_1405, n_198);
  nand g1053 (n_1406, n_440, n_197);
  nand g1054 (n_1407, n_198, n_197);
  nand g1055 (n_1408, n_440, n_198);
  nand g1056 (n_457, n_1406, n_1407, n_1408);
  xor g1057 (n_1409, n_441, n_442);
  xor g1058 (n_176, n_1409, n_443);
  nand g1059 (n_1410, n_441, n_442);
  nand g1060 (n_1411, n_443, n_442);
  nand g1061 (n_1412, n_441, n_443);
  nand g1062 (n_102, n_1410, n_1411, n_1412);
  xor g1063 (n_1413, A[25], A[23]);
  xor g1064 (n_448, n_1413, A[19]);
  nand g1065 (n_1414, A[25], A[23]);
  nand g1066 (n_1415, A[19], A[23]);
  nand g1067 (n_1416, A[25], A[19]);
  nand g1068 (n_458, n_1414, n_1415, n_1416);
  xor g1070 (n_449, n_1045, A[17]);
  nand g1072 (n_1419, A[17], A[9]);
  nand g1074 (n_459, n_1046, n_1419, n_1168);
  xor g1075 (n_1421, A[7], A[21]);
  xor g1076 (n_447, n_1421, A[15]);
  nand g1077 (n_1422, A[7], A[21]);
  nand g1080 (n_460, n_1422, n_1288, n_1355);
  xor g1081 (n_1425, A[13], n_444);
  xor g1082 (n_451, n_1425, n_445);
  nand g1083 (n_1426, A[13], n_444);
  nand g1084 (n_1427, n_445, n_444);
  nand g1085 (n_1428, A[13], n_445);
  nand g1086 (n_464, n_1426, n_1427, n_1428);
  xor g1087 (n_1429, n_446, n_447);
  xor g1088 (n_453, n_1429, n_448);
  nand g1089 (n_1430, n_446, n_447);
  nand g1090 (n_1431, n_448, n_447);
  nand g1091 (n_1432, n_446, n_448);
  nand g1092 (n_466, n_1430, n_1431, n_1432);
  xor g1093 (n_1433, n_449, n_450);
  xor g1094 (n_455, n_1433, n_451);
  nand g1095 (n_1434, n_449, n_450);
  nand g1096 (n_1435, n_451, n_450);
  nand g1097 (n_1436, n_449, n_451);
  nand g1098 (n_468, n_1434, n_1435, n_1436);
  xor g1099 (n_1437, n_452, n_453);
  xor g1100 (n_456, n_1437, n_454);
  nand g1101 (n_1438, n_452, n_453);
  nand g1102 (n_1439, n_454, n_453);
  nand g1103 (n_1440, n_452, n_454);
  nand g1104 (n_471, n_1438, n_1439, n_1440);
  xor g1105 (n_1441, n_455, n_456);
  xor g1106 (n_175, n_1441, n_457);
  nand g1107 (n_1442, n_455, n_456);
  nand g1108 (n_1443, n_457, n_456);
  nand g1109 (n_1444, n_455, n_457);
  nand g1110 (n_101, n_1442, n_1443, n_1444);
  xor g1111 (n_1445, A[26], A[24]);
  xor g1112 (n_462, n_1445, A[20]);
  nand g1113 (n_1446, A[26], A[24]);
  nand g1114 (n_1447, A[20], A[24]);
  nand g1115 (n_1448, A[26], A[20]);
  nand g1116 (n_472, n_1446, n_1447, n_1448);
  xor g1118 (n_463, n_296, A[18]);
  nand g1120 (n_1451, A[18], A[10]);
  xor g1123 (n_1453, A[8], A[22]);
  xor g1124 (n_461, n_1453, A[16]);
  nand g1125 (n_1454, A[8], A[22]);
  nand g1128 (n_474, n_1454, n_1320, n_1387);
  xor g1129 (n_1457, A[14], n_458);
  xor g1130 (n_465, n_1457, n_459);
  nand g1131 (n_1458, A[14], n_458);
  nand g1132 (n_1459, n_459, n_458);
  nand g1133 (n_1460, A[14], n_459);
  nand g1134 (n_478, n_1458, n_1459, n_1460);
  xor g1135 (n_1461, n_460, n_461);
  xor g1136 (n_467, n_1461, n_462);
  nand g1137 (n_1462, n_460, n_461);
  nand g1138 (n_1463, n_462, n_461);
  nand g1139 (n_1464, n_460, n_462);
  nand g1140 (n_480, n_1462, n_1463, n_1464);
  xor g1141 (n_1465, n_463, n_464);
  xor g1142 (n_469, n_1465, n_465);
  nand g1143 (n_1466, n_463, n_464);
  nand g1144 (n_1467, n_465, n_464);
  nand g1145 (n_1468, n_463, n_465);
  nand g1146 (n_482, n_1466, n_1467, n_1468);
  xor g1147 (n_1469, n_466, n_467);
  xor g1148 (n_470, n_1469, n_468);
  nand g1149 (n_1470, n_466, n_467);
  nand g1150 (n_1471, n_468, n_467);
  nand g1151 (n_1472, n_466, n_468);
  nand g1152 (n_485, n_1470, n_1471, n_1472);
  xor g1153 (n_1473, n_469, n_470);
  xor g1154 (n_174, n_1473, n_471);
  nand g1155 (n_1474, n_469, n_470);
  nand g1156 (n_1475, n_471, n_470);
  nand g1157 (n_1476, n_469, n_471);
  nand g1158 (n_100, n_1474, n_1475, n_1476);
  xor g1159 (n_1477, A[27], A[25]);
  xor g1160 (n_476, n_1477, A[21]);
  nand g1161 (n_1478, A[27], A[25]);
  nand g1162 (n_1479, A[21], A[25]);
  nand g1163 (n_1480, A[27], A[21]);
  nand g1164 (n_486, n_1478, n_1479, n_1480);
  xor g1166 (n_477, n_1077, A[19]);
  nand g1168 (n_1483, A[19], A[11]);
  nand g1170 (n_487, n_1078, n_1483, n_1224);
  xor g1171 (n_1485, A[9], A[23]);
  xor g1172 (n_475, n_1485, A[17]);
  nand g1173 (n_1486, A[9], A[23]);
  nand g1176 (n_488, n_1486, n_1352, n_1419);
  xor g1177 (n_1489, A[15], n_472);
  xor g1178 (n_479, n_1489, n_473);
  nand g1179 (n_1490, A[15], n_472);
  nand g1180 (n_1491, n_473, n_472);
  nand g1181 (n_1492, A[15], n_473);
  nand g1182 (n_492, n_1490, n_1491, n_1492);
  xor g1183 (n_1493, n_474, n_475);
  xor g1184 (n_481, n_1493, n_476);
  nand g1185 (n_1494, n_474, n_475);
  nand g1186 (n_1495, n_476, n_475);
  nand g1187 (n_1496, n_474, n_476);
  nand g1188 (n_494, n_1494, n_1495, n_1496);
  xor g1189 (n_1497, n_477, n_478);
  xor g1190 (n_483, n_1497, n_479);
  nand g1191 (n_1498, n_477, n_478);
  nand g1192 (n_1499, n_479, n_478);
  nand g1193 (n_1500, n_477, n_479);
  nand g1194 (n_496, n_1498, n_1499, n_1500);
  xor g1195 (n_1501, n_480, n_481);
  xor g1196 (n_484, n_1501, n_482);
  nand g1197 (n_1502, n_480, n_481);
  nand g1198 (n_1503, n_482, n_481);
  nand g1199 (n_1504, n_480, n_482);
  nand g1200 (n_499, n_1502, n_1503, n_1504);
  xor g1201 (n_1505, n_483, n_484);
  xor g1202 (n_173, n_1505, n_485);
  nand g1203 (n_1506, n_483, n_484);
  nand g1204 (n_1507, n_485, n_484);
  nand g1205 (n_1508, n_483, n_485);
  nand g1206 (n_99, n_1506, n_1507, n_1508);
  xor g1207 (n_1509, A[28], A[26]);
  xor g1208 (n_490, n_1509, A[22]);
  nand g1209 (n_1510, A[28], A[26]);
  nand g1210 (n_1511, A[22], A[26]);
  nand g1211 (n_1512, A[28], A[22]);
  nand g1212 (n_500, n_1510, n_1511, n_1512);
  xor g1214 (n_491, n_311, A[20]);
  nand g1216 (n_1515, A[20], A[12]);
  xor g1219 (n_1517, A[10], A[24]);
  xor g1220 (n_489, n_1517, A[18]);
  nand g1221 (n_1518, A[10], A[24]);
  nand g1224 (n_502, n_1518, n_1384, n_1451);
  xor g1225 (n_1521, A[16], n_486);
  xor g1226 (n_493, n_1521, n_487);
  nand g1227 (n_1522, A[16], n_486);
  nand g1228 (n_1523, n_487, n_486);
  nand g1229 (n_1524, A[16], n_487);
  nand g1230 (n_506, n_1522, n_1523, n_1524);
  xor g1231 (n_1525, n_488, n_489);
  xor g1232 (n_495, n_1525, n_490);
  nand g1233 (n_1526, n_488, n_489);
  nand g1234 (n_1527, n_490, n_489);
  nand g1235 (n_1528, n_488, n_490);
  nand g1236 (n_508, n_1526, n_1527, n_1528);
  xor g1237 (n_1529, n_491, n_492);
  xor g1238 (n_497, n_1529, n_493);
  nand g1239 (n_1530, n_491, n_492);
  nand g1240 (n_1531, n_493, n_492);
  nand g1241 (n_1532, n_491, n_493);
  nand g1242 (n_510, n_1530, n_1531, n_1532);
  xor g1243 (n_1533, n_494, n_495);
  xor g1244 (n_498, n_1533, n_496);
  nand g1245 (n_1534, n_494, n_495);
  nand g1246 (n_1535, n_496, n_495);
  nand g1247 (n_1536, n_494, n_496);
  nand g1248 (n_513, n_1534, n_1535, n_1536);
  xor g1249 (n_1537, n_497, n_498);
  xor g1250 (n_172, n_1537, n_499);
  nand g1251 (n_1538, n_497, n_498);
  nand g1252 (n_1539, n_499, n_498);
  nand g1253 (n_1540, n_497, n_499);
  nand g1254 (n_98, n_1538, n_1539, n_1540);
  xor g1255 (n_1541, A[29], A[27]);
  xor g1256 (n_504, n_1541, A[23]);
  nand g1257 (n_1542, A[29], A[27]);
  nand g1258 (n_1543, A[23], A[27]);
  nand g1259 (n_1544, A[29], A[23]);
  nand g1260 (n_514, n_1542, n_1543, n_1544);
  xor g1262 (n_505, n_1117, A[21]);
  nand g1264 (n_1547, A[21], A[13]);
  nand g1266 (n_515, n_1118, n_1547, n_1288);
  xor g1267 (n_1549, A[11], A[25]);
  xor g1268 (n_503, n_1549, A[19]);
  nand g1269 (n_1550, A[11], A[25]);
  nand g1272 (n_516, n_1550, n_1416, n_1483);
  xor g1273 (n_1553, A[17], n_500);
  xor g1274 (n_507, n_1553, n_501);
  nand g1275 (n_1554, A[17], n_500);
  nand g1276 (n_1555, n_501, n_500);
  nand g1277 (n_1556, A[17], n_501);
  nand g1278 (n_520, n_1554, n_1555, n_1556);
  xor g1279 (n_1557, n_502, n_503);
  xor g1280 (n_509, n_1557, n_504);
  nand g1281 (n_1558, n_502, n_503);
  nand g1282 (n_1559, n_504, n_503);
  nand g1283 (n_1560, n_502, n_504);
  nand g1284 (n_522, n_1558, n_1559, n_1560);
  xor g1285 (n_1561, n_505, n_506);
  xor g1286 (n_511, n_1561, n_507);
  nand g1287 (n_1562, n_505, n_506);
  nand g1288 (n_1563, n_507, n_506);
  nand g1289 (n_1564, n_505, n_507);
  nand g1290 (n_524, n_1562, n_1563, n_1564);
  xor g1291 (n_1565, n_508, n_509);
  xor g1292 (n_512, n_1565, n_510);
  nand g1293 (n_1566, n_508, n_509);
  nand g1294 (n_1567, n_510, n_509);
  nand g1295 (n_1568, n_508, n_510);
  nand g1296 (n_527, n_1566, n_1567, n_1568);
  xor g1297 (n_1569, n_511, n_512);
  xor g1298 (n_171, n_1569, n_513);
  nand g1299 (n_1570, n_511, n_512);
  nand g1300 (n_1571, n_513, n_512);
  nand g1301 (n_1572, n_511, n_513);
  nand g1302 (n_97, n_1570, n_1571, n_1572);
  xor g1303 (n_1573, A[30], A[28]);
  xor g1304 (n_518, n_1573, A[24]);
  nand g1305 (n_1574, A[30], A[28]);
  nand g1306 (n_1575, A[24], A[28]);
  nand g1307 (n_1576, A[30], A[24]);
  nand g1308 (n_528, n_1574, n_1575, n_1576);
  xor g1310 (n_519, n_330, A[22]);
  nand g1312 (n_1579, A[22], A[14]);
  xor g1315 (n_1581, A[12], A[26]);
  xor g1316 (n_517, n_1581, A[20]);
  nand g1317 (n_1582, A[12], A[26]);
  nand g1320 (n_530, n_1582, n_1448, n_1515);
  xor g1321 (n_1585, A[18], n_514);
  xor g1322 (n_521, n_1585, n_515);
  nand g1323 (n_1586, A[18], n_514);
  nand g1324 (n_1587, n_515, n_514);
  nand g1325 (n_1588, A[18], n_515);
  nand g1326 (n_534, n_1586, n_1587, n_1588);
  xor g1327 (n_1589, n_516, n_517);
  xor g1328 (n_523, n_1589, n_518);
  nand g1329 (n_1590, n_516, n_517);
  nand g1330 (n_1591, n_518, n_517);
  nand g1331 (n_1592, n_516, n_518);
  nand g1332 (n_536, n_1590, n_1591, n_1592);
  xor g1333 (n_1593, n_519, n_520);
  xor g1334 (n_525, n_1593, n_521);
  nand g1335 (n_1594, n_519, n_520);
  nand g1336 (n_1595, n_521, n_520);
  nand g1337 (n_1596, n_519, n_521);
  nand g1338 (n_538, n_1594, n_1595, n_1596);
  xor g1339 (n_1597, n_522, n_523);
  xor g1340 (n_526, n_1597, n_524);
  nand g1341 (n_1598, n_522, n_523);
  nand g1342 (n_1599, n_524, n_523);
  nand g1343 (n_1600, n_522, n_524);
  nand g1344 (n_541, n_1598, n_1599, n_1600);
  xor g1345 (n_1601, n_525, n_526);
  xor g1346 (n_170, n_1601, n_527);
  nand g1347 (n_1602, n_525, n_526);
  nand g1348 (n_1603, n_527, n_526);
  nand g1349 (n_1604, n_525, n_527);
  nand g1350 (n_96, n_1602, n_1603, n_1604);
  xor g1351 (n_1605, A[31], A[29]);
  xor g1352 (n_532, n_1605, A[25]);
  nand g1353 (n_1606, A[31], A[29]);
  nand g1354 (n_1607, A[25], A[29]);
  nand g1355 (n_1608, A[31], A[25]);
  nand g1356 (n_542, n_1606, n_1607, n_1608);
  xor g1358 (n_533, n_1165, A[23]);
  nand g1360 (n_1611, A[23], A[15]);
  nand g1362 (n_543, n_1166, n_1611, n_1352);
  xor g1363 (n_1613, A[13], A[27]);
  xor g1364 (n_531, n_1613, A[21]);
  nand g1365 (n_1614, A[13], A[27]);
  nand g1368 (n_544, n_1614, n_1480, n_1547);
  xor g1369 (n_1617, A[19], n_528);
  xor g1370 (n_535, n_1617, n_529);
  nand g1371 (n_1618, A[19], n_528);
  nand g1372 (n_1619, n_529, n_528);
  nand g1373 (n_1620, A[19], n_529);
  nand g1374 (n_548, n_1618, n_1619, n_1620);
  xor g1375 (n_1621, n_530, n_531);
  xor g1376 (n_537, n_1621, n_532);
  nand g1377 (n_1622, n_530, n_531);
  nand g1378 (n_1623, n_532, n_531);
  nand g1379 (n_1624, n_530, n_532);
  nand g1380 (n_550, n_1622, n_1623, n_1624);
  xor g1381 (n_1625, n_533, n_534);
  xor g1382 (n_539, n_1625, n_535);
  nand g1383 (n_1626, n_533, n_534);
  nand g1384 (n_1627, n_535, n_534);
  nand g1385 (n_1628, n_533, n_535);
  nand g1386 (n_552, n_1626, n_1627, n_1628);
  xor g1387 (n_1629, n_536, n_537);
  xor g1388 (n_540, n_1629, n_538);
  nand g1389 (n_1630, n_536, n_537);
  nand g1390 (n_1631, n_538, n_537);
  nand g1391 (n_1632, n_536, n_538);
  nand g1392 (n_555, n_1630, n_1631, n_1632);
  xor g1393 (n_1633, n_539, n_540);
  xor g1394 (n_169, n_1633, n_541);
  nand g1395 (n_1634, n_539, n_540);
  nand g1396 (n_1635, n_541, n_540);
  nand g1397 (n_1636, n_539, n_541);
  nand g1398 (n_95, n_1634, n_1635, n_1636);
  xor g1399 (n_1637, A[32], A[30]);
  xor g1400 (n_546, n_1637, A[26]);
  nand g1401 (n_1638, A[32], A[30]);
  nand g1402 (n_1639, A[26], A[30]);
  nand g1403 (n_1640, A[32], A[26]);
  nand g1404 (n_556, n_1638, n_1639, n_1640);
  xor g1406 (n_547, n_353, A[24]);
  nand g1408 (n_1643, A[24], A[16]);
  xor g1411 (n_1645, A[14], A[28]);
  xor g1412 (n_545, n_1645, A[22]);
  nand g1413 (n_1646, A[14], A[28]);
  nand g1416 (n_558, n_1646, n_1512, n_1579);
  xor g1417 (n_1649, A[20], n_542);
  xor g1418 (n_549, n_1649, n_543);
  nand g1419 (n_1650, A[20], n_542);
  nand g1420 (n_1651, n_543, n_542);
  nand g1421 (n_1652, A[20], n_543);
  nand g1422 (n_562, n_1650, n_1651, n_1652);
  xor g1423 (n_1653, n_544, n_545);
  xor g1424 (n_551, n_1653, n_546);
  nand g1425 (n_1654, n_544, n_545);
  nand g1426 (n_1655, n_546, n_545);
  nand g1427 (n_1656, n_544, n_546);
  nand g1428 (n_564, n_1654, n_1655, n_1656);
  xor g1429 (n_1657, n_547, n_548);
  xor g1430 (n_553, n_1657, n_549);
  nand g1431 (n_1658, n_547, n_548);
  nand g1432 (n_1659, n_549, n_548);
  nand g1433 (n_1660, n_547, n_549);
  nand g1434 (n_566, n_1658, n_1659, n_1660);
  xor g1435 (n_1661, n_550, n_551);
  xor g1436 (n_554, n_1661, n_552);
  nand g1437 (n_1662, n_550, n_551);
  nand g1438 (n_1663, n_552, n_551);
  nand g1439 (n_1664, n_550, n_552);
  nand g1440 (n_569, n_1662, n_1663, n_1664);
  xor g1441 (n_1665, n_553, n_554);
  xor g1442 (n_168, n_1665, n_555);
  nand g1443 (n_1666, n_553, n_554);
  nand g1444 (n_1667, n_555, n_554);
  nand g1445 (n_1668, n_553, n_555);
  nand g1446 (n_94, n_1666, n_1667, n_1668);
  xor g1447 (n_1669, A[33], A[31]);
  xor g1448 (n_560, n_1669, A[27]);
  nand g1449 (n_1670, A[33], A[31]);
  nand g1450 (n_1671, A[27], A[31]);
  nand g1451 (n_1672, A[33], A[27]);
  nand g1452 (n_570, n_1670, n_1671, n_1672);
  xor g1454 (n_561, n_1221, A[25]);
  nand g1456 (n_1675, A[25], A[17]);
  nand g1458 (n_571, n_1222, n_1675, n_1416);
  xor g1459 (n_1677, A[15], A[29]);
  xor g1460 (n_559, n_1677, A[23]);
  nand g1461 (n_1678, A[15], A[29]);
  nand g1464 (n_572, n_1678, n_1544, n_1611);
  xor g1465 (n_1681, A[21], n_556);
  xor g1466 (n_563, n_1681, n_557);
  nand g1467 (n_1682, A[21], n_556);
  nand g1468 (n_1683, n_557, n_556);
  nand g1469 (n_1684, A[21], n_557);
  nand g1470 (n_576, n_1682, n_1683, n_1684);
  xor g1471 (n_1685, n_558, n_559);
  xor g1472 (n_565, n_1685, n_560);
  nand g1473 (n_1686, n_558, n_559);
  nand g1474 (n_1687, n_560, n_559);
  nand g1475 (n_1688, n_558, n_560);
  nand g1476 (n_578, n_1686, n_1687, n_1688);
  xor g1477 (n_1689, n_561, n_562);
  xor g1478 (n_567, n_1689, n_563);
  nand g1479 (n_1690, n_561, n_562);
  nand g1480 (n_1691, n_563, n_562);
  nand g1481 (n_1692, n_561, n_563);
  nand g1482 (n_580, n_1690, n_1691, n_1692);
  xor g1483 (n_1693, n_564, n_565);
  xor g1484 (n_568, n_1693, n_566);
  nand g1485 (n_1694, n_564, n_565);
  nand g1486 (n_1695, n_566, n_565);
  nand g1487 (n_1696, n_564, n_566);
  nand g1488 (n_583, n_1694, n_1695, n_1696);
  xor g1489 (n_1697, n_567, n_568);
  xor g1490 (n_167, n_1697, n_569);
  nand g1491 (n_1698, n_567, n_568);
  nand g1492 (n_1699, n_569, n_568);
  nand g1493 (n_1700, n_567, n_569);
  nand g1494 (n_93, n_1698, n_1699, n_1700);
  xor g1495 (n_1701, A[34], A[32]);
  xor g1496 (n_574, n_1701, A[28]);
  nand g1497 (n_1702, A[34], A[32]);
  nand g1498 (n_1703, A[28], A[32]);
  nand g1499 (n_1704, A[34], A[28]);
  nand g1500 (n_584, n_1702, n_1703, n_1704);
  xor g1502 (n_575, n_1253, A[26]);
  nand g1504 (n_1707, A[26], A[18]);
  nand g1506 (n_585, n_1254, n_1707, n_1448);
  xor g1507 (n_1709, A[16], A[30]);
  xor g1508 (n_573, n_1709, A[24]);
  nand g1509 (n_1710, A[16], A[30]);
  nand g1512 (n_586, n_1710, n_1576, n_1643);
  xor g1513 (n_1713, A[22], n_570);
  xor g1514 (n_577, n_1713, n_571);
  nand g1515 (n_1714, A[22], n_570);
  nand g1516 (n_1715, n_571, n_570);
  nand g1517 (n_1716, A[22], n_571);
  nand g1518 (n_590, n_1714, n_1715, n_1716);
  xor g1519 (n_1717, n_572, n_573);
  xor g1520 (n_579, n_1717, n_574);
  nand g1521 (n_1718, n_572, n_573);
  nand g1522 (n_1719, n_574, n_573);
  nand g1523 (n_1720, n_572, n_574);
  nand g1524 (n_592, n_1718, n_1719, n_1720);
  xor g1525 (n_1721, n_575, n_576);
  xor g1526 (n_581, n_1721, n_577);
  nand g1527 (n_1722, n_575, n_576);
  nand g1528 (n_1723, n_577, n_576);
  nand g1529 (n_1724, n_575, n_577);
  nand g1530 (n_594, n_1722, n_1723, n_1724);
  xor g1531 (n_1725, n_578, n_579);
  xor g1532 (n_582, n_1725, n_580);
  nand g1533 (n_1726, n_578, n_579);
  nand g1534 (n_1727, n_580, n_579);
  nand g1535 (n_1728, n_578, n_580);
  nand g1536 (n_597, n_1726, n_1727, n_1728);
  xor g1537 (n_1729, n_581, n_582);
  xor g1538 (n_166, n_1729, n_583);
  nand g1539 (n_1730, n_581, n_582);
  nand g1540 (n_1731, n_583, n_582);
  nand g1541 (n_1732, n_581, n_583);
  nand g1542 (n_92, n_1730, n_1731, n_1732);
  xor g1543 (n_1733, A[35], A[33]);
  xor g1544 (n_588, n_1733, A[29]);
  nand g1545 (n_1734, A[35], A[33]);
  nand g1546 (n_1735, A[29], A[33]);
  nand g1547 (n_1736, A[35], A[29]);
  nand g1548 (n_598, n_1734, n_1735, n_1736);
  xor g1550 (n_589, n_1285, A[27]);
  nand g1552 (n_1739, A[27], A[19]);
  nand g1554 (n_599, n_1286, n_1739, n_1480);
  xor g1555 (n_1741, A[17], A[31]);
  xor g1556 (n_587, n_1741, A[25]);
  nand g1557 (n_1742, A[17], A[31]);
  nand g1560 (n_600, n_1742, n_1608, n_1675);
  xor g1561 (n_1745, A[23], n_584);
  xor g1562 (n_591, n_1745, n_585);
  nand g1563 (n_1746, A[23], n_584);
  nand g1564 (n_1747, n_585, n_584);
  nand g1565 (n_1748, A[23], n_585);
  nand g1566 (n_604, n_1746, n_1747, n_1748);
  xor g1567 (n_1749, n_586, n_587);
  xor g1568 (n_593, n_1749, n_588);
  nand g1569 (n_1750, n_586, n_587);
  nand g1570 (n_1751, n_588, n_587);
  nand g1571 (n_1752, n_586, n_588);
  nand g1572 (n_606, n_1750, n_1751, n_1752);
  xor g1573 (n_1753, n_589, n_590);
  xor g1574 (n_595, n_1753, n_591);
  nand g1575 (n_1754, n_589, n_590);
  nand g1576 (n_1755, n_591, n_590);
  nand g1577 (n_1756, n_589, n_591);
  nand g1578 (n_608, n_1754, n_1755, n_1756);
  xor g1579 (n_1757, n_592, n_593);
  xor g1580 (n_596, n_1757, n_594);
  nand g1581 (n_1758, n_592, n_593);
  nand g1582 (n_1759, n_594, n_593);
  nand g1583 (n_1760, n_592, n_594);
  nand g1584 (n_611, n_1758, n_1759, n_1760);
  xor g1585 (n_1761, n_595, n_596);
  xor g1586 (n_165, n_1761, n_597);
  nand g1587 (n_1762, n_595, n_596);
  nand g1588 (n_1763, n_597, n_596);
  nand g1589 (n_1764, n_595, n_597);
  nand g1590 (n_91, n_1762, n_1763, n_1764);
  xor g1591 (n_1765, A[36], A[34]);
  xor g1592 (n_602, n_1765, A[30]);
  nand g1593 (n_1766, A[36], A[34]);
  nand g1594 (n_1767, A[30], A[34]);
  nand g1595 (n_1768, A[36], A[30]);
  nand g1596 (n_612, n_1766, n_1767, n_1768);
  xor g1598 (n_603, n_1317, A[28]);
  nand g1600 (n_1771, A[28], A[20]);
  nand g1602 (n_613, n_1318, n_1771, n_1512);
  xor g1603 (n_1773, A[18], A[32]);
  xor g1604 (n_601, n_1773, A[26]);
  nand g1605 (n_1774, A[18], A[32]);
  nand g1608 (n_614, n_1774, n_1640, n_1707);
  xor g1609 (n_1777, A[24], n_598);
  xor g1610 (n_605, n_1777, n_599);
  nand g1611 (n_1778, A[24], n_598);
  nand g1612 (n_1779, n_599, n_598);
  nand g1613 (n_1780, A[24], n_599);
  nand g1614 (n_618, n_1778, n_1779, n_1780);
  xor g1615 (n_1781, n_600, n_601);
  xor g1616 (n_607, n_1781, n_602);
  nand g1617 (n_1782, n_600, n_601);
  nand g1618 (n_1783, n_602, n_601);
  nand g1619 (n_1784, n_600, n_602);
  nand g1620 (n_620, n_1782, n_1783, n_1784);
  xor g1621 (n_1785, n_603, n_604);
  xor g1622 (n_609, n_1785, n_605);
  nand g1623 (n_1786, n_603, n_604);
  nand g1624 (n_1787, n_605, n_604);
  nand g1625 (n_1788, n_603, n_605);
  nand g1626 (n_622, n_1786, n_1787, n_1788);
  xor g1627 (n_1789, n_606, n_607);
  xor g1628 (n_610, n_1789, n_608);
  nand g1629 (n_1790, n_606, n_607);
  nand g1630 (n_1791, n_608, n_607);
  nand g1631 (n_1792, n_606, n_608);
  nand g1632 (n_625, n_1790, n_1791, n_1792);
  xor g1633 (n_1793, n_609, n_610);
  xor g1634 (n_164, n_1793, n_611);
  nand g1635 (n_1794, n_609, n_610);
  nand g1636 (n_1795, n_611, n_610);
  nand g1637 (n_1796, n_609, n_611);
  nand g1638 (n_90, n_1794, n_1795, n_1796);
  xor g1639 (n_1797, A[37], A[35]);
  xor g1640 (n_616, n_1797, A[31]);
  nand g1641 (n_1798, A[37], A[35]);
  nand g1642 (n_1799, A[31], A[35]);
  nand g1643 (n_1800, A[37], A[31]);
  nand g1644 (n_626, n_1798, n_1799, n_1800);
  xor g1646 (n_617, n_1349, A[29]);
  nand g1648 (n_1803, A[29], A[21]);
  nand g1650 (n_627, n_1350, n_1803, n_1544);
  xor g1651 (n_1805, A[19], A[33]);
  xor g1652 (n_615, n_1805, A[27]);
  nand g1653 (n_1806, A[19], A[33]);
  nand g1656 (n_628, n_1806, n_1672, n_1739);
  xor g1657 (n_1809, A[25], n_612);
  xor g1658 (n_619, n_1809, n_613);
  nand g1659 (n_1810, A[25], n_612);
  nand g1660 (n_1811, n_613, n_612);
  nand g1661 (n_1812, A[25], n_613);
  nand g1662 (n_632, n_1810, n_1811, n_1812);
  xor g1663 (n_1813, n_614, n_615);
  xor g1664 (n_621, n_1813, n_616);
  nand g1665 (n_1814, n_614, n_615);
  nand g1666 (n_1815, n_616, n_615);
  nand g1667 (n_1816, n_614, n_616);
  nand g1668 (n_634, n_1814, n_1815, n_1816);
  xor g1669 (n_1817, n_617, n_618);
  xor g1670 (n_623, n_1817, n_619);
  nand g1671 (n_1818, n_617, n_618);
  nand g1672 (n_1819, n_619, n_618);
  nand g1673 (n_1820, n_617, n_619);
  nand g1674 (n_636, n_1818, n_1819, n_1820);
  xor g1675 (n_1821, n_620, n_621);
  xor g1676 (n_624, n_1821, n_622);
  nand g1677 (n_1822, n_620, n_621);
  nand g1678 (n_1823, n_622, n_621);
  nand g1679 (n_1824, n_620, n_622);
  nand g1680 (n_639, n_1822, n_1823, n_1824);
  xor g1681 (n_1825, n_623, n_624);
  xor g1682 (n_163, n_1825, n_625);
  nand g1683 (n_1826, n_623, n_624);
  nand g1684 (n_1827, n_625, n_624);
  nand g1685 (n_1828, n_623, n_625);
  nand g1686 (n_89, n_1826, n_1827, n_1828);
  xor g1687 (n_1829, A[38], A[36]);
  xor g1688 (n_630, n_1829, A[32]);
  nand g1689 (n_1830, A[38], A[36]);
  nand g1690 (n_1831, A[32], A[36]);
  nand g1691 (n_1832, A[38], A[32]);
  nand g1692 (n_640, n_1830, n_1831, n_1832);
  xor g1694 (n_631, n_1381, A[30]);
  nand g1696 (n_1835, A[30], A[22]);
  nand g1698 (n_641, n_1382, n_1835, n_1576);
  xor g1699 (n_1837, A[20], A[34]);
  xor g1700 (n_629, n_1837, A[28]);
  nand g1701 (n_1838, A[20], A[34]);
  nand g1704 (n_642, n_1838, n_1704, n_1771);
  xor g1705 (n_1841, A[26], n_626);
  xor g1706 (n_633, n_1841, n_627);
  nand g1707 (n_1842, A[26], n_626);
  nand g1708 (n_1843, n_627, n_626);
  nand g1709 (n_1844, A[26], n_627);
  nand g1710 (n_646, n_1842, n_1843, n_1844);
  xor g1711 (n_1845, n_628, n_629);
  xor g1712 (n_635, n_1845, n_630);
  nand g1713 (n_1846, n_628, n_629);
  nand g1714 (n_1847, n_630, n_629);
  nand g1715 (n_1848, n_628, n_630);
  nand g1716 (n_648, n_1846, n_1847, n_1848);
  xor g1717 (n_1849, n_631, n_632);
  xor g1718 (n_637, n_1849, n_633);
  nand g1719 (n_1850, n_631, n_632);
  nand g1720 (n_1851, n_633, n_632);
  nand g1721 (n_1852, n_631, n_633);
  nand g1722 (n_650, n_1850, n_1851, n_1852);
  xor g1723 (n_1853, n_634, n_635);
  xor g1724 (n_638, n_1853, n_636);
  nand g1725 (n_1854, n_634, n_635);
  nand g1726 (n_1855, n_636, n_635);
  nand g1727 (n_1856, n_634, n_636);
  nand g1728 (n_653, n_1854, n_1855, n_1856);
  xor g1729 (n_1857, n_637, n_638);
  xor g1730 (n_162, n_1857, n_639);
  nand g1731 (n_1858, n_637, n_638);
  nand g1732 (n_1859, n_639, n_638);
  nand g1733 (n_1860, n_637, n_639);
  nand g1734 (n_88, n_1858, n_1859, n_1860);
  xor g1735 (n_1861, A[39], A[37]);
  xor g1736 (n_644, n_1861, A[33]);
  nand g1737 (n_1862, A[39], A[37]);
  nand g1738 (n_1863, A[33], A[37]);
  nand g1739 (n_1864, A[39], A[33]);
  nand g1740 (n_654, n_1862, n_1863, n_1864);
  xor g1742 (n_645, n_1413, A[31]);
  nand g1744 (n_1867, A[31], A[23]);
  nand g1746 (n_655, n_1414, n_1867, n_1608);
  xor g1747 (n_1869, A[21], A[35]);
  xor g1748 (n_643, n_1869, A[29]);
  nand g1749 (n_1870, A[21], A[35]);
  nand g1752 (n_656, n_1870, n_1736, n_1803);
  xor g1753 (n_1873, A[27], n_640);
  xor g1754 (n_647, n_1873, n_641);
  nand g1755 (n_1874, A[27], n_640);
  nand g1756 (n_1875, n_641, n_640);
  nand g1757 (n_1876, A[27], n_641);
  nand g1758 (n_660, n_1874, n_1875, n_1876);
  xor g1759 (n_1877, n_642, n_643);
  xor g1760 (n_649, n_1877, n_644);
  nand g1761 (n_1878, n_642, n_643);
  nand g1762 (n_1879, n_644, n_643);
  nand g1763 (n_1880, n_642, n_644);
  nand g1764 (n_662, n_1878, n_1879, n_1880);
  xor g1765 (n_1881, n_645, n_646);
  xor g1766 (n_651, n_1881, n_647);
  nand g1767 (n_1882, n_645, n_646);
  nand g1768 (n_1883, n_647, n_646);
  nand g1769 (n_1884, n_645, n_647);
  nand g1770 (n_664, n_1882, n_1883, n_1884);
  xor g1771 (n_1885, n_648, n_649);
  xor g1772 (n_652, n_1885, n_650);
  nand g1773 (n_1886, n_648, n_649);
  nand g1774 (n_1887, n_650, n_649);
  nand g1775 (n_1888, n_648, n_650);
  nand g1776 (n_667, n_1886, n_1887, n_1888);
  xor g1777 (n_1889, n_651, n_652);
  xor g1778 (n_161, n_1889, n_653);
  nand g1779 (n_1890, n_651, n_652);
  nand g1780 (n_1891, n_653, n_652);
  nand g1781 (n_1892, n_651, n_653);
  nand g1782 (n_87, n_1890, n_1891, n_1892);
  xor g1783 (n_1893, A[40], A[38]);
  xor g1784 (n_658, n_1893, A[34]);
  nand g1785 (n_1894, A[40], A[38]);
  nand g1786 (n_1895, A[34], A[38]);
  nand g1787 (n_1896, A[40], A[34]);
  nand g1788 (n_668, n_1894, n_1895, n_1896);
  xor g1790 (n_659, n_1445, A[32]);
  nand g1792 (n_1899, A[32], A[24]);
  nand g1794 (n_669, n_1446, n_1899, n_1640);
  xor g1795 (n_1901, A[22], A[36]);
  xor g1796 (n_657, n_1901, A[30]);
  nand g1797 (n_1902, A[22], A[36]);
  nand g1800 (n_670, n_1902, n_1768, n_1835);
  xor g1801 (n_1905, A[28], n_654);
  xor g1802 (n_661, n_1905, n_655);
  nand g1803 (n_1906, A[28], n_654);
  nand g1804 (n_1907, n_655, n_654);
  nand g1805 (n_1908, A[28], n_655);
  nand g1806 (n_674, n_1906, n_1907, n_1908);
  xor g1807 (n_1909, n_656, n_657);
  xor g1808 (n_663, n_1909, n_658);
  nand g1809 (n_1910, n_656, n_657);
  nand g1810 (n_1911, n_658, n_657);
  nand g1811 (n_1912, n_656, n_658);
  nand g1812 (n_676, n_1910, n_1911, n_1912);
  xor g1813 (n_1913, n_659, n_660);
  xor g1814 (n_665, n_1913, n_661);
  nand g1815 (n_1914, n_659, n_660);
  nand g1816 (n_1915, n_661, n_660);
  nand g1817 (n_1916, n_659, n_661);
  nand g1818 (n_678, n_1914, n_1915, n_1916);
  xor g1819 (n_1917, n_662, n_663);
  xor g1820 (n_666, n_1917, n_664);
  nand g1821 (n_1918, n_662, n_663);
  nand g1822 (n_1919, n_664, n_663);
  nand g1823 (n_1920, n_662, n_664);
  nand g1824 (n_681, n_1918, n_1919, n_1920);
  xor g1825 (n_1921, n_665, n_666);
  xor g1826 (n_160, n_1921, n_667);
  nand g1827 (n_1922, n_665, n_666);
  nand g1828 (n_1923, n_667, n_666);
  nand g1829 (n_1924, n_665, n_667);
  nand g1830 (n_86, n_1922, n_1923, n_1924);
  xor g1831 (n_1925, A[41], A[39]);
  xor g1832 (n_672, n_1925, A[35]);
  nand g1833 (n_1926, A[41], A[39]);
  nand g1834 (n_1927, A[35], A[39]);
  nand g1835 (n_1928, A[41], A[35]);
  nand g1836 (n_682, n_1926, n_1927, n_1928);
  xor g1838 (n_673, n_1477, A[33]);
  nand g1840 (n_1931, A[33], A[25]);
  nand g1842 (n_683, n_1478, n_1931, n_1672);
  xor g1843 (n_1933, A[23], A[37]);
  xor g1844 (n_671, n_1933, A[31]);
  nand g1845 (n_1934, A[23], A[37]);
  nand g1848 (n_684, n_1934, n_1800, n_1867);
  xor g1849 (n_1937, A[29], n_668);
  xor g1850 (n_675, n_1937, n_669);
  nand g1851 (n_1938, A[29], n_668);
  nand g1852 (n_1939, n_669, n_668);
  nand g1853 (n_1940, A[29], n_669);
  nand g1854 (n_688, n_1938, n_1939, n_1940);
  xor g1855 (n_1941, n_670, n_671);
  xor g1856 (n_677, n_1941, n_672);
  nand g1857 (n_1942, n_670, n_671);
  nand g1858 (n_1943, n_672, n_671);
  nand g1859 (n_1944, n_670, n_672);
  nand g1860 (n_690, n_1942, n_1943, n_1944);
  xor g1861 (n_1945, n_673, n_674);
  xor g1862 (n_679, n_1945, n_675);
  nand g1863 (n_1946, n_673, n_674);
  nand g1864 (n_1947, n_675, n_674);
  nand g1865 (n_1948, n_673, n_675);
  nand g1866 (n_692, n_1946, n_1947, n_1948);
  xor g1867 (n_1949, n_676, n_677);
  xor g1868 (n_680, n_1949, n_678);
  nand g1869 (n_1950, n_676, n_677);
  nand g1870 (n_1951, n_678, n_677);
  nand g1871 (n_1952, n_676, n_678);
  nand g1872 (n_695, n_1950, n_1951, n_1952);
  xor g1873 (n_1953, n_679, n_680);
  xor g1874 (n_159, n_1953, n_681);
  nand g1875 (n_1954, n_679, n_680);
  nand g1876 (n_1955, n_681, n_680);
  nand g1877 (n_1956, n_679, n_681);
  nand g1878 (n_85, n_1954, n_1955, n_1956);
  xor g1879 (n_1957, A[42], A[40]);
  xor g1880 (n_686, n_1957, A[36]);
  nand g1881 (n_1958, A[42], A[40]);
  nand g1882 (n_1959, A[36], A[40]);
  nand g1883 (n_1960, A[42], A[36]);
  nand g1884 (n_696, n_1958, n_1959, n_1960);
  xor g1886 (n_687, n_1509, A[34]);
  nand g1888 (n_1963, A[34], A[26]);
  nand g1890 (n_697, n_1510, n_1963, n_1704);
  xor g1891 (n_1965, A[24], A[38]);
  xor g1892 (n_685, n_1965, A[32]);
  nand g1893 (n_1966, A[24], A[38]);
  nand g1896 (n_698, n_1966, n_1832, n_1899);
  xor g1897 (n_1969, A[30], n_682);
  xor g1898 (n_689, n_1969, n_683);
  nand g1899 (n_1970, A[30], n_682);
  nand g1900 (n_1971, n_683, n_682);
  nand g1901 (n_1972, A[30], n_683);
  nand g1902 (n_702, n_1970, n_1971, n_1972);
  xor g1903 (n_1973, n_684, n_685);
  xor g1904 (n_691, n_1973, n_686);
  nand g1905 (n_1974, n_684, n_685);
  nand g1906 (n_1975, n_686, n_685);
  nand g1907 (n_1976, n_684, n_686);
  nand g1908 (n_704, n_1974, n_1975, n_1976);
  xor g1909 (n_1977, n_687, n_688);
  xor g1910 (n_693, n_1977, n_689);
  nand g1911 (n_1978, n_687, n_688);
  nand g1912 (n_1979, n_689, n_688);
  nand g1913 (n_1980, n_687, n_689);
  nand g1914 (n_706, n_1978, n_1979, n_1980);
  xor g1915 (n_1981, n_690, n_691);
  xor g1916 (n_694, n_1981, n_692);
  nand g1917 (n_1982, n_690, n_691);
  nand g1918 (n_1983, n_692, n_691);
  nand g1919 (n_1984, n_690, n_692);
  nand g1920 (n_709, n_1982, n_1983, n_1984);
  xor g1921 (n_1985, n_693, n_694);
  xor g1922 (n_158, n_1985, n_695);
  nand g1923 (n_1986, n_693, n_694);
  nand g1924 (n_1987, n_695, n_694);
  nand g1925 (n_1988, n_693, n_695);
  nand g1926 (n_84, n_1986, n_1987, n_1988);
  xor g1927 (n_1989, A[43], A[41]);
  xor g1928 (n_700, n_1989, A[37]);
  nand g1929 (n_1990, A[43], A[41]);
  nand g1930 (n_1991, A[37], A[41]);
  nand g1931 (n_1992, A[43], A[37]);
  nand g1932 (n_710, n_1990, n_1991, n_1992);
  xor g1934 (n_701, n_1541, A[35]);
  nand g1936 (n_1995, A[35], A[27]);
  nand g1938 (n_711, n_1542, n_1995, n_1736);
  xor g1939 (n_1997, A[25], A[39]);
  xor g1940 (n_699, n_1997, A[33]);
  nand g1941 (n_1998, A[25], A[39]);
  nand g1944 (n_712, n_1998, n_1864, n_1931);
  xor g1945 (n_2001, A[31], n_696);
  xor g1946 (n_703, n_2001, n_697);
  nand g1947 (n_2002, A[31], n_696);
  nand g1948 (n_2003, n_697, n_696);
  nand g1949 (n_2004, A[31], n_697);
  nand g1950 (n_716, n_2002, n_2003, n_2004);
  xor g1951 (n_2005, n_698, n_699);
  xor g1952 (n_705, n_2005, n_700);
  nand g1953 (n_2006, n_698, n_699);
  nand g1954 (n_2007, n_700, n_699);
  nand g1955 (n_2008, n_698, n_700);
  nand g1956 (n_718, n_2006, n_2007, n_2008);
  xor g1957 (n_2009, n_701, n_702);
  xor g1958 (n_707, n_2009, n_703);
  nand g1959 (n_2010, n_701, n_702);
  nand g1960 (n_2011, n_703, n_702);
  nand g1961 (n_2012, n_701, n_703);
  nand g1962 (n_720, n_2010, n_2011, n_2012);
  xor g1963 (n_2013, n_704, n_705);
  xor g1964 (n_708, n_2013, n_706);
  nand g1965 (n_2014, n_704, n_705);
  nand g1966 (n_2015, n_706, n_705);
  nand g1967 (n_2016, n_704, n_706);
  nand g1968 (n_723, n_2014, n_2015, n_2016);
  xor g1969 (n_2017, n_707, n_708);
  xor g1970 (n_157, n_2017, n_709);
  nand g1971 (n_2018, n_707, n_708);
  nand g1972 (n_2019, n_709, n_708);
  nand g1973 (n_2020, n_707, n_709);
  nand g1974 (n_83, n_2018, n_2019, n_2020);
  xor g1975 (n_2021, A[44], A[42]);
  xor g1976 (n_714, n_2021, A[38]);
  nand g1977 (n_2022, A[44], A[42]);
  nand g1978 (n_2023, A[38], A[42]);
  nand g1979 (n_2024, A[44], A[38]);
  nand g1980 (n_724, n_2022, n_2023, n_2024);
  xor g1982 (n_715, n_1573, A[36]);
  nand g1984 (n_2027, A[36], A[28]);
  nand g1986 (n_725, n_1574, n_2027, n_1768);
  xor g1987 (n_2029, A[26], A[40]);
  xor g1988 (n_713, n_2029, A[34]);
  nand g1989 (n_2030, A[26], A[40]);
  nand g1992 (n_726, n_2030, n_1896, n_1963);
  xor g1993 (n_2033, A[32], n_710);
  xor g1994 (n_717, n_2033, n_711);
  nand g1995 (n_2034, A[32], n_710);
  nand g1996 (n_2035, n_711, n_710);
  nand g1997 (n_2036, A[32], n_711);
  nand g1998 (n_730, n_2034, n_2035, n_2036);
  xor g1999 (n_2037, n_712, n_713);
  xor g2000 (n_719, n_2037, n_714);
  nand g2001 (n_2038, n_712, n_713);
  nand g2002 (n_2039, n_714, n_713);
  nand g2003 (n_2040, n_712, n_714);
  nand g2004 (n_732, n_2038, n_2039, n_2040);
  xor g2005 (n_2041, n_715, n_716);
  xor g2006 (n_721, n_2041, n_717);
  nand g2007 (n_2042, n_715, n_716);
  nand g2008 (n_2043, n_717, n_716);
  nand g2009 (n_2044, n_715, n_717);
  nand g2010 (n_734, n_2042, n_2043, n_2044);
  xor g2011 (n_2045, n_718, n_719);
  xor g2012 (n_722, n_2045, n_720);
  nand g2013 (n_2046, n_718, n_719);
  nand g2014 (n_2047, n_720, n_719);
  nand g2015 (n_2048, n_718, n_720);
  nand g2016 (n_737, n_2046, n_2047, n_2048);
  xor g2017 (n_2049, n_721, n_722);
  xor g2018 (n_156, n_2049, n_723);
  nand g2019 (n_2050, n_721, n_722);
  nand g2020 (n_2051, n_723, n_722);
  nand g2021 (n_2052, n_721, n_723);
  nand g2022 (n_82, n_2050, n_2051, n_2052);
  xor g2023 (n_2053, A[45], A[43]);
  xor g2024 (n_728, n_2053, A[39]);
  nand g2025 (n_2054, A[45], A[43]);
  nand g2026 (n_2055, A[39], A[43]);
  nand g2027 (n_2056, A[45], A[39]);
  nand g2028 (n_738, n_2054, n_2055, n_2056);
  xor g2030 (n_729, n_1605, A[37]);
  nand g2032 (n_2059, A[37], A[29]);
  nand g2034 (n_740, n_1606, n_2059, n_1800);
  xor g2035 (n_2061, A[27], A[41]);
  xor g2036 (n_727, n_2061, A[35]);
  nand g2037 (n_2062, A[27], A[41]);
  nand g2040 (n_739, n_2062, n_1928, n_1995);
  xor g2041 (n_2065, A[33], n_724);
  xor g2042 (n_731, n_2065, n_725);
  nand g2043 (n_2066, A[33], n_724);
  nand g2044 (n_2067, n_725, n_724);
  nand g2045 (n_2068, A[33], n_725);
  nand g2046 (n_744, n_2066, n_2067, n_2068);
  xor g2047 (n_2069, n_726, n_727);
  xor g2048 (n_733, n_2069, n_728);
  nand g2049 (n_2070, n_726, n_727);
  nand g2050 (n_2071, n_728, n_727);
  nand g2051 (n_2072, n_726, n_728);
  nand g2052 (n_746, n_2070, n_2071, n_2072);
  xor g2053 (n_2073, n_729, n_730);
  xor g2054 (n_735, n_2073, n_731);
  nand g2055 (n_2074, n_729, n_730);
  nand g2056 (n_2075, n_731, n_730);
  nand g2057 (n_2076, n_729, n_731);
  nand g2058 (n_749, n_2074, n_2075, n_2076);
  xor g2059 (n_2077, n_732, n_733);
  xor g2060 (n_736, n_2077, n_734);
  nand g2061 (n_2078, n_732, n_733);
  nand g2062 (n_2079, n_734, n_733);
  nand g2063 (n_2080, n_732, n_734);
  nand g2064 (n_751, n_2078, n_2079, n_2080);
  xor g2065 (n_2081, n_735, n_736);
  xor g2066 (n_155, n_2081, n_737);
  nand g2067 (n_2082, n_735, n_736);
  nand g2068 (n_2083, n_737, n_736);
  nand g2069 (n_2084, n_735, n_737);
  nand g2070 (n_81, n_2082, n_2083, n_2084);
  xor g2071 (n_2085, A[44], A[40]);
  xor g2072 (n_742, n_2085, A[32]);
  nand g2073 (n_2086, A[44], A[40]);
  nand g2074 (n_2087, A[32], A[40]);
  nand g2075 (n_2088, A[44], A[32]);
  nand g2076 (n_752, n_2086, n_2087, n_2088);
  xor g2077 (n_2089, A[30], A[38]);
  xor g2078 (n_743, n_2089, A[28]);
  nand g2079 (n_2090, A[30], A[38]);
  nand g2080 (n_2091, A[28], A[38]);
  nand g2082 (n_754, n_2090, n_2091, n_1574);
  xor g2083 (n_2093, A[42], A[36]);
  xor g2084 (n_741, n_2093, A[34]);
  nand g2087 (n_2096, A[42], A[34]);
  nand g2088 (n_753, n_1960, n_1766, n_2096);
  xor g2089 (n_2097, A[46], n_738);
  xor g2090 (n_745, n_2097, n_739);
  nand g2091 (n_2098, A[46], n_738);
  nand g2092 (n_2099, n_739, n_738);
  nand g2093 (n_2100, A[46], n_739);
  nand g2094 (n_758, n_2098, n_2099, n_2100);
  xor g2095 (n_2101, n_740, n_741);
  xor g2096 (n_747, n_2101, n_742);
  nand g2097 (n_2102, n_740, n_741);
  nand g2098 (n_2103, n_742, n_741);
  nand g2099 (n_2104, n_740, n_742);
  nand g2100 (n_760, n_2102, n_2103, n_2104);
  xor g2101 (n_2105, n_743, n_744);
  xor g2102 (n_748, n_2105, n_745);
  nand g2103 (n_2106, n_743, n_744);
  nand g2104 (n_2107, n_745, n_744);
  nand g2105 (n_2108, n_743, n_745);
  nand g2106 (n_763, n_2106, n_2107, n_2108);
  xor g2107 (n_2109, n_746, n_747);
  xor g2108 (n_750, n_2109, n_748);
  nand g2109 (n_2110, n_746, n_747);
  nand g2110 (n_2111, n_748, n_747);
  nand g2111 (n_2112, n_746, n_748);
  nand g2112 (n_765, n_2110, n_2111, n_2112);
  xor g2113 (n_2113, n_749, n_750);
  xor g2114 (n_154, n_2113, n_751);
  nand g2115 (n_2114, n_749, n_750);
  nand g2116 (n_2115, n_751, n_750);
  nand g2117 (n_2116, n_749, n_751);
  nand g2118 (n_80, n_2114, n_2115, n_2116);
  xor g2119 (n_2117, A[45], A[41]);
  xor g2120 (n_756, n_2117, A[33]);
  nand g2121 (n_2118, A[45], A[41]);
  nand g2122 (n_2119, A[33], A[41]);
  nand g2123 (n_2120, A[45], A[33]);
  nand g2124 (n_767, n_2118, n_2119, n_2120);
  xor g2125 (n_2121, A[31], A[39]);
  xor g2126 (n_757, n_2121, A[29]);
  nand g2127 (n_2122, A[31], A[39]);
  nand g2128 (n_2123, A[29], A[39]);
  nand g2130 (n_768, n_2122, n_2123, n_1606);
  xor g2131 (n_2125, A[43], A[37]);
  xor g2132 (n_755, n_2125, A[35]);
  nand g2135 (n_2128, A[43], A[35]);
  nand g2136 (n_766, n_1992, n_1798, n_2128);
  xor g2137 (n_2129, A[47], n_752);
  xor g2138 (n_759, n_2129, n_753);
  nand g2139 (n_2130, A[47], n_752);
  nand g2140 (n_2131, n_753, n_752);
  nand g2141 (n_2132, A[47], n_753);
  nand g2142 (n_772, n_2130, n_2131, n_2132);
  xor g2143 (n_2133, n_754, n_755);
  xor g2144 (n_761, n_2133, n_756);
  nand g2145 (n_2134, n_754, n_755);
  nand g2146 (n_2135, n_756, n_755);
  nand g2147 (n_2136, n_754, n_756);
  nand g2148 (n_773, n_2134, n_2135, n_2136);
  xor g2149 (n_2137, n_757, n_758);
  xor g2150 (n_762, n_2137, n_759);
  nand g2151 (n_2138, n_757, n_758);
  nand g2152 (n_2139, n_759, n_758);
  nand g2153 (n_2140, n_757, n_759);
  nand g2154 (n_777, n_2138, n_2139, n_2140);
  xor g2155 (n_2141, n_760, n_761);
  xor g2156 (n_764, n_2141, n_762);
  nand g2157 (n_2142, n_760, n_761);
  nand g2158 (n_2143, n_762, n_761);
  nand g2159 (n_2144, n_760, n_762);
  nand g2160 (n_779, n_2142, n_2143, n_2144);
  xor g2161 (n_2145, n_763, n_764);
  xor g2162 (n_153, n_2145, n_765);
  nand g2163 (n_2146, n_763, n_764);
  nand g2164 (n_2147, n_765, n_764);
  nand g2165 (n_2148, n_763, n_765);
  nand g2166 (n_79, n_2146, n_2147, n_2148);
  xor g2168 (n_769, n_2021, A[34]);
  nand g2171 (n_2152, A[44], A[34]);
  nand g2172 (n_780, n_2022, n_2096, n_2152);
  xor g2173 (n_2153, A[32], A[40]);
  xor g2174 (n_771, n_2153, A[30]);
  nand g2176 (n_2155, A[30], A[40]);
  nand g2178 (n_781, n_2087, n_2155, n_1638);
  xor g2180 (n_770, n_1829, A[46]);
  nand g2182 (n_2159, A[46], A[36]);
  nand g2183 (n_2160, A[38], A[46]);
  nand g2184 (n_783, n_1830, n_2159, n_2160);
  xor g2185 (n_2161, A[48], n_766);
  xor g2186 (n_774, n_2161, n_767);
  nand g2187 (n_2162, A[48], n_766);
  nand g2188 (n_2163, n_767, n_766);
  nand g2189 (n_2164, A[48], n_767);
  nand g2190 (n_786, n_2162, n_2163, n_2164);
  xor g2191 (n_2165, n_768, n_769);
  xor g2192 (n_775, n_2165, n_770);
  nand g2193 (n_2166, n_768, n_769);
  nand g2194 (n_2167, n_770, n_769);
  nand g2195 (n_2168, n_768, n_770);
  nand g2196 (n_787, n_2166, n_2167, n_2168);
  xor g2197 (n_2169, n_771, n_772);
  xor g2198 (n_776, n_2169, n_773);
  nand g2199 (n_2170, n_771, n_772);
  nand g2200 (n_2171, n_773, n_772);
  nand g2201 (n_2172, n_771, n_773);
  nand g2202 (n_791, n_2170, n_2171, n_2172);
  xor g2203 (n_2173, n_774, n_775);
  xor g2204 (n_778, n_2173, n_776);
  nand g2205 (n_2174, n_774, n_775);
  nand g2206 (n_2175, n_776, n_775);
  nand g2207 (n_2176, n_774, n_776);
  nand g2208 (n_793, n_2174, n_2175, n_2176);
  xor g2209 (n_2177, n_777, n_778);
  xor g2210 (n_152, n_2177, n_779);
  nand g2211 (n_2178, n_777, n_778);
  nand g2212 (n_2179, n_779, n_778);
  nand g2213 (n_2180, n_777, n_779);
  nand g2214 (n_78, n_2178, n_2179, n_2180);
  xor g2216 (n_782, n_2053, A[35]);
  nand g2219 (n_2184, A[45], A[35]);
  nand g2220 (n_794, n_2054, n_2128, n_2184);
  xor g2221 (n_2185, A[33], A[41]);
  xor g2222 (n_785, n_2185, A[31]);
  nand g2224 (n_2187, A[31], A[41]);
  nand g2226 (n_795, n_2119, n_2187, n_1670);
  xor g2228 (n_784, n_1861, A[47]);
  nand g2230 (n_2191, A[47], A[37]);
  nand g2231 (n_2192, A[39], A[47]);
  nand g2232 (n_797, n_1862, n_2191, n_2192);
  xor g2233 (n_2193, A[49], n_780);
  xor g2234 (n_788, n_2193, n_781);
  nand g2235 (n_2194, A[49], n_780);
  nand g2236 (n_2195, n_781, n_780);
  nand g2237 (n_2196, A[49], n_781);
  nand g2238 (n_800, n_2194, n_2195, n_2196);
  xor g2239 (n_2197, n_782, n_783);
  xor g2240 (n_789, n_2197, n_784);
  nand g2241 (n_2198, n_782, n_783);
  nand g2242 (n_2199, n_784, n_783);
  nand g2243 (n_2200, n_782, n_784);
  nand g2244 (n_801, n_2198, n_2199, n_2200);
  xor g2245 (n_2201, n_785, n_786);
  xor g2246 (n_790, n_2201, n_787);
  nand g2247 (n_2202, n_785, n_786);
  nand g2248 (n_2203, n_787, n_786);
  nand g2249 (n_2204, n_785, n_787);
  nand g2250 (n_805, n_2202, n_2203, n_2204);
  xor g2251 (n_2205, n_788, n_789);
  xor g2252 (n_792, n_2205, n_790);
  nand g2253 (n_2206, n_788, n_789);
  nand g2254 (n_2207, n_790, n_789);
  nand g2255 (n_2208, n_788, n_790);
  nand g2256 (n_807, n_2206, n_2207, n_2208);
  xor g2257 (n_2209, n_791, n_792);
  xor g2258 (n_151, n_2209, n_793);
  nand g2259 (n_2210, n_791, n_792);
  nand g2260 (n_2211, n_793, n_792);
  nand g2261 (n_2212, n_791, n_793);
  nand g2262 (n_77, n_2210, n_2211, n_2212);
  xor g2263 (n_2213, A[50], A[44]);
  xor g2264 (n_796, n_2213, A[36]);
  nand g2265 (n_2214, A[50], A[44]);
  nand g2266 (n_2215, A[36], A[44]);
  nand g2267 (n_2216, A[50], A[36]);
  nand g2268 (n_808, n_2214, n_2215, n_2216);
  xor g2269 (n_2217, A[34], A[42]);
  xor g2270 (n_799, n_2217, A[32]);
  nand g2272 (n_2219, A[32], A[42]);
  nand g2274 (n_809, n_2096, n_2219, n_1702);
  xor g2276 (n_798, n_1893, A[48]);
  nand g2278 (n_2223, A[48], A[38]);
  nand g2279 (n_2224, A[40], A[48]);
  nand g2280 (n_811, n_1894, n_2223, n_2224);
  xor g2281 (n_2225, A[46], n_794);
  xor g2282 (n_802, n_2225, n_795);
  nand g2283 (n_2226, A[46], n_794);
  nand g2284 (n_2227, n_795, n_794);
  nand g2285 (n_2228, A[46], n_795);
  nand g2286 (n_814, n_2226, n_2227, n_2228);
  xor g2287 (n_2229, n_796, n_797);
  xor g2288 (n_803, n_2229, n_798);
  nand g2289 (n_2230, n_796, n_797);
  nand g2290 (n_2231, n_798, n_797);
  nand g2291 (n_2232, n_796, n_798);
  nand g2292 (n_815, n_2230, n_2231, n_2232);
  xor g2293 (n_2233, n_799, n_800);
  xor g2294 (n_804, n_2233, n_801);
  nand g2295 (n_2234, n_799, n_800);
  nand g2296 (n_2235, n_801, n_800);
  nand g2297 (n_2236, n_799, n_801);
  nand g2298 (n_819, n_2234, n_2235, n_2236);
  xor g2299 (n_2237, n_802, n_803);
  xor g2300 (n_806, n_2237, n_804);
  nand g2301 (n_2238, n_802, n_803);
  nand g2302 (n_2239, n_804, n_803);
  nand g2303 (n_2240, n_802, n_804);
  nand g2304 (n_821, n_2238, n_2239, n_2240);
  xor g2305 (n_2241, n_805, n_806);
  xor g2306 (n_150, n_2241, n_807);
  nand g2307 (n_2242, n_805, n_806);
  nand g2308 (n_2243, n_807, n_806);
  nand g2309 (n_2244, n_805, n_807);
  nand g2310 (n_76, n_2242, n_2243, n_2244);
  xor g2311 (n_2245, A[51], A[45]);
  xor g2312 (n_810, n_2245, A[37]);
  nand g2313 (n_2246, A[51], A[45]);
  nand g2314 (n_2247, A[37], A[45]);
  nand g2315 (n_2248, A[51], A[37]);
  nand g2316 (n_822, n_2246, n_2247, n_2248);
  xor g2317 (n_2249, A[35], A[43]);
  xor g2318 (n_813, n_2249, A[33]);
  nand g2320 (n_2251, A[33], A[43]);
  nand g2322 (n_823, n_2128, n_2251, n_1734);
  xor g2324 (n_812, n_1925, A[49]);
  nand g2326 (n_2255, A[49], A[39]);
  nand g2327 (n_2256, A[41], A[49]);
  nand g2328 (n_825, n_1926, n_2255, n_2256);
  xor g2329 (n_2257, A[47], n_808);
  xor g2330 (n_816, n_2257, n_809);
  nand g2331 (n_2258, A[47], n_808);
  nand g2332 (n_2259, n_809, n_808);
  nand g2333 (n_2260, A[47], n_809);
  nand g2334 (n_828, n_2258, n_2259, n_2260);
  xor g2335 (n_2261, n_810, n_811);
  xor g2336 (n_817, n_2261, n_812);
  nand g2337 (n_2262, n_810, n_811);
  nand g2338 (n_2263, n_812, n_811);
  nand g2339 (n_2264, n_810, n_812);
  nand g2340 (n_829, n_2262, n_2263, n_2264);
  xor g2341 (n_2265, n_813, n_814);
  xor g2342 (n_818, n_2265, n_815);
  nand g2343 (n_2266, n_813, n_814);
  nand g2344 (n_2267, n_815, n_814);
  nand g2345 (n_2268, n_813, n_815);
  nand g2346 (n_833, n_2266, n_2267, n_2268);
  xor g2347 (n_2269, n_816, n_817);
  xor g2348 (n_820, n_2269, n_818);
  nand g2349 (n_2270, n_816, n_817);
  nand g2350 (n_2271, n_818, n_817);
  nand g2351 (n_2272, n_816, n_818);
  nand g2352 (n_835, n_2270, n_2271, n_2272);
  xor g2353 (n_2273, n_819, n_820);
  xor g2354 (n_149, n_2273, n_821);
  nand g2355 (n_2274, n_819, n_820);
  nand g2356 (n_2275, n_821, n_820);
  nand g2357 (n_2276, n_819, n_821);
  nand g2358 (n_75, n_2274, n_2275, n_2276);
  xor g2359 (n_2277, A[52], A[50]);
  xor g2360 (n_824, n_2277, A[38]);
  nand g2361 (n_2278, A[52], A[50]);
  nand g2362 (n_2279, A[38], A[50]);
  nand g2363 (n_2280, A[52], A[38]);
  nand g2364 (n_839, n_2278, n_2279, n_2280);
  xor g2365 (n_2281, A[36], A[44]);
  xor g2366 (n_827, n_2281, A[34]);
  nand g2370 (n_838, n_2215, n_2152, n_1766);
  xor g2372 (n_826, n_1957, A[46]);
  nand g2374 (n_2287, A[46], A[40]);
  nand g2375 (n_2288, A[42], A[46]);
  nand g2376 (n_843, n_1958, n_2287, n_2288);
  xor g2377 (n_2289, A[48], n_822);
  xor g2378 (n_830, n_2289, n_823);
  nand g2379 (n_2290, A[48], n_822);
  nand g2380 (n_2291, n_823, n_822);
  nand g2381 (n_2292, A[48], n_823);
  nand g2382 (n_844, n_2290, n_2291, n_2292);
  xor g2383 (n_2293, n_824, n_825);
  xor g2384 (n_831, n_2293, n_826);
  nand g2385 (n_2294, n_824, n_825);
  nand g2386 (n_2295, n_826, n_825);
  nand g2387 (n_2296, n_824, n_826);
  nand g2388 (n_846, n_2294, n_2295, n_2296);
  xor g2389 (n_2297, n_827, n_828);
  xor g2390 (n_832, n_2297, n_829);
  nand g2391 (n_2298, n_827, n_828);
  nand g2392 (n_2299, n_829, n_828);
  nand g2393 (n_2300, n_827, n_829);
  nand g2394 (n_849, n_2298, n_2299, n_2300);
  xor g2395 (n_2301, n_830, n_831);
  xor g2396 (n_834, n_2301, n_832);
  nand g2397 (n_2302, n_830, n_831);
  nand g2398 (n_2303, n_832, n_831);
  nand g2399 (n_2304, n_830, n_832);
  nand g2400 (n_851, n_2302, n_2303, n_2304);
  xor g2401 (n_2305, n_833, n_834);
  xor g2402 (n_148, n_2305, n_835);
  nand g2403 (n_2306, n_833, n_834);
  nand g2404 (n_2307, n_835, n_834);
  nand g2405 (n_2308, n_833, n_835);
  nand g2406 (n_74, n_2306, n_2307, n_2308);
  xor g2409 (n_2309, A[53], A[39]);
  xor g2410 (n_841, n_2309, A[37]);
  nand g2411 (n_2310, A[53], A[39]);
  nand g2413 (n_2312, A[53], A[37]);
  nand g2414 (n_856, n_2310, n_1862, n_2312);
  xor g2415 (n_2313, A[51], A[35]);
  xor g2416 (n_842, n_2313, A[45]);
  nand g2417 (n_2314, A[51], A[35]);
  nand g2420 (n_855, n_2314, n_2184, n_2246);
  xor g2422 (n_840, n_1989, A[47]);
  nand g2424 (n_2319, A[47], A[41]);
  nand g2425 (n_2320, A[43], A[47]);
  nand g2426 (n_860, n_1990, n_2319, n_2320);
  xor g2427 (n_2321, A[49], n_838);
  xor g2428 (n_845, n_2321, n_839);
  nand g2429 (n_2322, A[49], n_838);
  nand g2430 (n_2323, n_839, n_838);
  nand g2431 (n_2324, A[49], n_839);
  nand g2432 (n_861, n_2322, n_2323, n_2324);
  xor g2433 (n_2325, n_840, n_841);
  xor g2434 (n_847, n_2325, n_842);
  nand g2435 (n_2326, n_840, n_841);
  nand g2436 (n_2327, n_842, n_841);
  nand g2437 (n_2328, n_840, n_842);
  nand g2438 (n_863, n_2326, n_2327, n_2328);
  xor g2439 (n_2329, n_843, n_844);
  xor g2440 (n_848, n_2329, n_845);
  nand g2441 (n_2330, n_843, n_844);
  nand g2442 (n_2331, n_845, n_844);
  nand g2443 (n_2332, n_843, n_845);
  nand g2444 (n_866, n_2330, n_2331, n_2332);
  xor g2445 (n_2333, n_846, n_847);
  xor g2446 (n_850, n_2333, n_848);
  nand g2447 (n_2334, n_846, n_847);
  nand g2448 (n_2335, n_848, n_847);
  nand g2449 (n_2336, n_846, n_848);
  nand g2450 (n_868, n_2334, n_2335, n_2336);
  xor g2451 (n_2337, n_849, n_850);
  xor g2452 (n_147, n_2337, n_851);
  nand g2453 (n_2338, n_849, n_850);
  nand g2454 (n_2339, n_851, n_850);
  nand g2455 (n_2340, n_849, n_851);
  nand g2456 (n_73, n_2338, n_2339, n_2340);
  xor g2460 (n_858, n_1829, A[53]);
  nand g2462 (n_2343, A[53], A[36]);
  nand g2463 (n_2344, A[38], A[53]);
  nand g2464 (n_870, n_1830, n_2343, n_2344);
  xor g2465 (n_2345, A[52], A[44]);
  xor g2466 (n_859, n_2345, A[50]);
  nand g2467 (n_2346, A[52], A[44]);
  nand g2470 (n_871, n_2346, n_2214, n_2278);
  xor g2477 (n_2353, A[48], n_855);
  xor g2478 (n_862, n_2353, n_856);
  nand g2479 (n_2354, A[48], n_855);
  nand g2480 (n_2355, n_856, n_855);
  nand g2481 (n_2356, A[48], n_856);
  nand g2482 (n_876, n_2354, n_2355, n_2356);
  xor g2483 (n_2357, n_826, n_858);
  xor g2484 (n_864, n_2357, n_859);
  nand g2485 (n_2358, n_826, n_858);
  nand g2486 (n_2359, n_859, n_858);
  nand g2487 (n_2360, n_826, n_859);
  nand g2488 (n_877, n_2358, n_2359, n_2360);
  xor g2489 (n_2361, n_860, n_861);
  xor g2490 (n_865, n_2361, n_862);
  nand g2491 (n_2362, n_860, n_861);
  nand g2492 (n_2363, n_862, n_861);
  nand g2493 (n_2364, n_860, n_862);
  nand g2494 (n_881, n_2362, n_2363, n_2364);
  xor g2495 (n_2365, n_863, n_864);
  xor g2496 (n_867, n_2365, n_865);
  nand g2497 (n_2366, n_863, n_864);
  nand g2498 (n_2367, n_865, n_864);
  nand g2499 (n_2368, n_863, n_865);
  nand g2500 (n_883, n_2366, n_2367, n_2368);
  xor g2501 (n_2369, n_866, n_867);
  xor g2502 (n_146, n_2369, n_868);
  nand g2503 (n_2370, n_866, n_867);
  nand g2504 (n_2371, n_868, n_867);
  nand g2505 (n_2372, n_866, n_868);
  nand g2506 (n_72, n_2370, n_2371, n_2372);
  xor g2508 (n_872, n_2373, A[39]);
  nand g2510 (n_2375, A[39], A[51]);
  nand g2512 (n_886, n_2374, n_2375, n_2376);
  xor g2513 (n_2377, A[37], A[45]);
  nand g2518 (n_887, n_2247, n_2379, n_2380);
  xor g2525 (n_2385, A[49], n_870);
  xor g2526 (n_878, n_2385, n_871);
  nand g2527 (n_2386, A[49], n_870);
  nand g2528 (n_2387, n_871, n_870);
  nand g2529 (n_2388, A[49], n_871);
  nand g2530 (n_891, n_2386, n_2387, n_2388);
  xor g2531 (n_2389, n_872, n_843);
  xor g2532 (n_879, n_2389, n_840);
  nand g2533 (n_2390, n_872, n_843);
  nand g2534 (n_2391, n_840, n_843);
  nand g2535 (n_2392, n_872, n_840);
  nand g2536 (n_893, n_2390, n_2391, n_2392);
  xor g2537 (n_2393, n_875, n_876);
  xor g2538 (n_880, n_2393, n_877);
  nand g2539 (n_2394, n_875, n_876);
  nand g2540 (n_2395, n_877, n_876);
  nand g2541 (n_2396, n_875, n_877);
  nand g2542 (n_895, n_2394, n_2395, n_2396);
  xor g2543 (n_2397, n_878, n_879);
  xor g2544 (n_882, n_2397, n_880);
  nand g2545 (n_2398, n_878, n_879);
  nand g2546 (n_2399, n_880, n_879);
  nand g2547 (n_2400, n_878, n_880);
  nand g2548 (n_898, n_2398, n_2399, n_2400);
  xor g2549 (n_2401, n_881, n_882);
  xor g2550 (n_145, n_2401, n_883);
  nand g2551 (n_2402, n_881, n_882);
  nand g2552 (n_2403, n_883, n_882);
  nand g2553 (n_2404, n_881, n_883);
  nand g2554 (n_71, n_2402, n_2403, n_2404);
  xor g2557 (n_2405, A[50], A[38]);
  xor g2558 (n_890, n_2405, A[44]);
  nand g2562 (n_900, n_2279, n_2024, n_2214);
  xor g2570 (n_892, n_2413, n_886);
  nand g2573 (n_2416, A[48], n_886);
  nand g2574 (n_905, n_2414, n_2415, n_2416);
  xor g2575 (n_2417, n_887, n_860);
  xor g2576 (n_894, n_2417, n_826);
  nand g2577 (n_2418, n_887, n_860);
  nand g2578 (n_2419, n_826, n_860);
  nand g2579 (n_2420, n_887, n_826);
  nand g2580 (n_906, n_2418, n_2419, n_2420);
  xor g2581 (n_2421, n_890, n_891);
  xor g2582 (n_896, n_2421, n_892);
  nand g2583 (n_2422, n_890, n_891);
  nand g2584 (n_2423, n_892, n_891);
  nand g2585 (n_2424, n_890, n_892);
  nand g2586 (n_909, n_2422, n_2423, n_2424);
  xor g2587 (n_2425, n_893, n_894);
  xor g2588 (n_897, n_2425, n_895);
  nand g2589 (n_2426, n_893, n_894);
  nand g2590 (n_2427, n_895, n_894);
  nand g2591 (n_2428, n_893, n_895);
  nand g2592 (n_911, n_2426, n_2427, n_2428);
  xor g2593 (n_2429, n_896, n_897);
  xor g2594 (n_144, n_2429, n_898);
  nand g2595 (n_2430, n_896, n_897);
  nand g2596 (n_2431, n_898, n_897);
  nand g2597 (n_2432, n_896, n_898);
  nand g2598 (n_70, n_2430, n_2431, n_2432);
  xor g2606 (n_902, n_2053, A[41]);
  nand g2610 (n_915, n_2054, n_1990, n_2118);
  xor g2611 (n_2441, A[47], A[49]);
  xor g2612 (n_904, n_2441, A[52]);
  nand g2613 (n_2442, A[47], A[49]);
  nand g2614 (n_2443, A[52], A[49]);
  nand g2615 (n_2444, A[47], A[52]);
  nand g2616 (n_918, n_2442, n_2443, n_2444);
  xor g2617 (n_2445, n_900, n_843);
  xor g2618 (n_907, n_2445, n_902);
  nand g2619 (n_2446, n_900, n_843);
  nand g2620 (n_2447, n_902, n_843);
  nand g2621 (n_2448, n_900, n_902);
  nand g2622 (n_920, n_2446, n_2447, n_2448);
  xor g2623 (n_2449, n_872, n_904);
  xor g2624 (n_908, n_2449, n_905);
  nand g2625 (n_2450, n_872, n_904);
  nand g2626 (n_2451, n_905, n_904);
  nand g2627 (n_2452, n_872, n_905);
  nand g2628 (n_922, n_2450, n_2451, n_2452);
  xor g2629 (n_2453, n_906, n_907);
  xor g2630 (n_910, n_2453, n_908);
  nand g2631 (n_2454, n_906, n_907);
  nand g2632 (n_2455, n_908, n_907);
  nand g2633 (n_2456, n_906, n_908);
  nand g2634 (n_924, n_2454, n_2455, n_2456);
  xor g2635 (n_2457, n_909, n_910);
  xor g2636 (n_143, n_2457, n_911);
  nand g2637 (n_2458, n_909, n_910);
  nand g2638 (n_2459, n_911, n_910);
  nand g2639 (n_2460, n_909, n_911);
  nand g2640 (n_69, n_2458, n_2459, n_2460);
  xor g2644 (n_916, n_2213, A[42]);
  nand g2647 (n_2464, A[50], A[42]);
  nand g2648 (n_926, n_2214, n_2022, n_2464);
  xor g2649 (n_2465, A[40], A[46]);
  xor g2650 (n_917, n_2465, A[48]);
  nand g2652 (n_2467, A[48], A[46]);
  nand g2654 (n_928, n_2287, n_2467, n_2224);
  xor g2656 (n_919, n_2469, n_915);
  nand g2658 (n_2471, n_915, n_886);
  nand g2660 (n_931, n_2415, n_2471, n_2472);
  xor g2661 (n_2473, n_916, n_917);
  xor g2662 (n_921, n_2473, n_918);
  nand g2663 (n_2474, n_916, n_917);
  nand g2664 (n_2475, n_918, n_917);
  nand g2665 (n_2476, n_916, n_918);
  nand g2666 (n_933, n_2474, n_2475, n_2476);
  xor g2667 (n_2477, n_919, n_920);
  xor g2668 (n_923, n_2477, n_921);
  nand g2669 (n_2478, n_919, n_920);
  nand g2670 (n_2479, n_921, n_920);
  nand g2671 (n_2480, n_919, n_921);
  nand g2672 (n_935, n_2478, n_2479, n_2480);
  xor g2673 (n_2481, n_922, n_923);
  xor g2674 (n_142, n_2481, n_924);
  nand g2675 (n_2482, n_922, n_923);
  nand g2676 (n_2483, n_924, n_923);
  nand g2677 (n_2484, n_922, n_924);
  nand g2678 (n_68, n_2482, n_2483, n_2484);
  xor g2680 (n_929, n_2373, A[45]);
  nand g2684 (n_938, n_2374, n_2246, n_2379);
  xor g2691 (n_2493, A[49], A[52]);
  xor g2692 (n_930, n_2493, n_926);
  nand g2694 (n_2495, n_926, A[52]);
  nand g2695 (n_2496, A[49], n_926);
  nand g2696 (n_942, n_2443, n_2495, n_2496);
  xor g2697 (n_2497, n_840, n_928);
  xor g2698 (n_932, n_2497, n_929);
  nand g2699 (n_2498, n_840, n_928);
  nand g2700 (n_2499, n_929, n_928);
  nand g2701 (n_2500, n_840, n_929);
  nand g2702 (n_943, n_2498, n_2499, n_2500);
  xor g2703 (n_2501, n_930, n_931);
  xor g2704 (n_934, n_2501, n_932);
  nand g2705 (n_2502, n_930, n_931);
  nand g2706 (n_2503, n_932, n_931);
  nand g2707 (n_2504, n_930, n_932);
  nand g2708 (n_946, n_2502, n_2503, n_2504);
  xor g2709 (n_2505, n_933, n_934);
  xor g2710 (n_141, n_2505, n_935);
  nand g2711 (n_2506, n_933, n_934);
  nand g2712 (n_2507, n_935, n_934);
  nand g2713 (n_2508, n_933, n_935);
  nand g2714 (n_140, n_2506, n_2507, n_2508);
  xor g2718 (n_940, n_2345, A[42]);
  nand g2720 (n_2511, A[42], A[52]);
  nand g2722 (n_948, n_2346, n_2511, n_2022);
  xor g2723 (n_2513, A[46], A[48]);
  nand g2728 (n_950, n_2467, n_2515, n_2516);
  xor g2729 (n_2517, n_938, n_860);
  xor g2730 (n_944, n_2517, n_940);
  nand g2731 (n_2518, n_938, n_860);
  nand g2732 (n_2519, n_940, n_860);
  nand g2733 (n_2520, n_938, n_940);
  nand g2734 (n_953, n_2518, n_2519, n_2520);
  xor g2735 (n_2521, n_941, n_942);
  xor g2736 (n_945, n_2521, n_943);
  nand g2737 (n_2522, n_941, n_942);
  nand g2738 (n_2523, n_943, n_942);
  nand g2739 (n_2524, n_941, n_943);
  nand g2740 (n_955, n_2522, n_2523, n_2524);
  xor g2741 (n_2525, n_944, n_945);
  xor g2742 (n_67, n_2525, n_946);
  nand g2743 (n_2526, n_944, n_945);
  nand g2744 (n_2527, n_946, n_945);
  nand g2745 (n_2528, n_944, n_946);
  nand g2746 (n_66, n_2526, n_2527, n_2528);
  xor g2753 (n_2533, A[43], A[47]);
  xor g2754 (n_951, n_2533, A[49]);
  nand g2757 (n_2536, A[43], A[49]);
  nand g2758 (n_960, n_2320, n_2442, n_2536);
  xor g2759 (n_2537, A[50], n_948);
  xor g2760 (n_952, n_2537, n_929);
  nand g2761 (n_2538, A[50], n_948);
  nand g2762 (n_2539, n_929, n_948);
  nand g2763 (n_2540, A[50], n_929);
  nand g2764 (n_962, n_2538, n_2539, n_2540);
  xor g2765 (n_2541, n_950, n_951);
  xor g2766 (n_954, n_2541, n_952);
  nand g2767 (n_2542, n_950, n_951);
  nand g2768 (n_2543, n_952, n_951);
  nand g2769 (n_2544, n_950, n_952);
  nand g2770 (n_964, n_2542, n_2543, n_2544);
  xor g2771 (n_2545, n_953, n_954);
  xor g2772 (n_139, n_2545, n_955);
  nand g2773 (n_2546, n_953, n_954);
  nand g2774 (n_2547, n_955, n_954);
  nand g2775 (n_2548, n_953, n_955);
  nand g2776 (n_65, n_2546, n_2547, n_2548);
  xor g2780 (n_959, n_2345, A[46]);
  nand g2782 (n_2551, A[46], A[52]);
  nand g2783 (n_2552, A[44], A[46]);
  nand g2784 (n_967, n_2346, n_2551, n_2552);
  nand g2789 (n_2556, A[48], n_938);
  nand g2790 (n_969, n_2515, n_2555, n_2556);
  xor g2791 (n_2557, n_959, n_960);
  xor g2792 (n_963, n_2557, n_961);
  nand g2793 (n_2558, n_959, n_960);
  nand g2794 (n_2559, n_961, n_960);
  nand g2795 (n_2560, n_959, n_961);
  nand g2796 (n_971, n_2558, n_2559, n_2560);
  xor g2797 (n_2561, n_962, n_963);
  xor g2798 (n_138, n_2561, n_964);
  nand g2799 (n_2562, n_962, n_963);
  nand g2800 (n_2563, n_964, n_963);
  nand g2801 (n_2564, n_962, n_964);
  nand g2802 (n_137, n_2562, n_2563, n_2564);
  xor g2810 (n_968, n_2441, A[50]);
  nand g2812 (n_2571, A[50], A[49]);
  nand g2813 (n_2572, A[47], A[50]);
  nand g2814 (n_975, n_2442, n_2571, n_2572);
  xor g2815 (n_2573, n_929, n_967);
  xor g2816 (n_970, n_2573, n_968);
  nand g2817 (n_2574, n_929, n_967);
  nand g2818 (n_2575, n_968, n_967);
  nand g2819 (n_2576, n_929, n_968);
  nand g2820 (n_978, n_2574, n_2575, n_2576);
  xor g2821 (n_2577, n_969, n_970);
  xor g2822 (n_64, n_2577, n_971);
  nand g2823 (n_2578, n_969, n_970);
  nand g2824 (n_2579, n_971, n_970);
  nand g2825 (n_2580, n_969, n_971);
  nand g2826 (n_63, n_2578, n_2579, n_2580);
  xor g2829 (n_2581, A[50], A[46]);
  xor g2830 (n_976, n_2581, A[48]);
  nand g2831 (n_2582, A[50], A[46]);
  nand g2833 (n_2584, A[50], A[48]);
  nand g2834 (n_981, n_2582, n_2467, n_2584);
  xor g2836 (n_977, n_2585, n_975);
  nand g2838 (n_2587, n_975, n_938);
  nand g2840 (n_983, n_2586, n_2587, n_2588);
  xor g2841 (n_2589, n_976, n_977);
  xor g2842 (n_136, n_2589, n_978);
  nand g2843 (n_2590, n_976, n_977);
  nand g2844 (n_2591, n_978, n_977);
  nand g2845 (n_2592, n_976, n_978);
  nand g2846 (n_62, n_2590, n_2591, n_2592);
  xor g2848 (n_980, n_2373, A[47]);
  nand g2850 (n_2595, A[47], A[51]);
  nand g2852 (n_986, n_2374, n_2595, n_2596);
  xor g2854 (n_982, n_2493, n_980);
  nand g2856 (n_2599, n_980, A[52]);
  nand g2857 (n_2600, A[49], n_980);
  nand g2858 (n_988, n_2443, n_2599, n_2600);
  xor g2859 (n_2601, n_981, n_982);
  xor g2860 (n_135, n_2601, n_983);
  nand g2861 (n_2602, n_981, n_982);
  nand g2862 (n_2603, n_983, n_982);
  nand g2863 (n_2604, n_981, n_983);
  nand g2864 (n_134, n_2602, n_2603, n_2604);
  xor g2867 (n_2605, A[50], A[48]);
  nand g2872 (n_991, n_2584, n_2414, n_2608);
  xor g2873 (n_2609, n_986, n_987);
  xor g2874 (n_61, n_2609, n_988);
  nand g2875 (n_2610, n_986, n_987);
  nand g2876 (n_2611, n_988, n_987);
  nand g2877 (n_2612, n_986, n_988);
  nand g2878 (n_133, n_2610, n_2611, n_2612);
  xor g2880 (n_990, n_2373, A[49]);
  nand g2882 (n_2615, A[49], A[51]);
  nand g2884 (n_994, n_2374, n_2615, n_2616);
  xor g2885 (n_2617, A[52], n_990);
  xor g2886 (n_60, n_2617, n_991);
  nand g2887 (n_2618, A[52], n_990);
  nand g2888 (n_2619, n_991, n_990);
  nand g2889 (n_2620, A[52], n_991);
  nand g2890 (n_132, n_2618, n_2619, n_2620);
  nand g2897 (n_2624, A[52], n_994);
  nand g2898 (n_131, n_2622, n_2623, n_2624);
  xor g2900 (n_58, n_2373, A[50]);
  nand g2902 (n_2627, A[50], A[51]);
  nand g2904 (n_130, n_2374, n_2627, n_2628);
  nor g11 (n_2644, A[2], A[0]);
  nor g13 (n_2640, A[3], A[1]);
  nor g15 (n_2650, A[2], n_196);
  nand g16 (n_2645, A[2], n_196);
  nor g17 (n_2646, n_122, n_195);
  nand g18 (n_2647, n_122, n_195);
  nor g19 (n_2656, n_121, n_194);
  nand g20 (n_2651, n_121, n_194);
  nor g21 (n_2652, n_120, n_193);
  nand g22 (n_2653, n_120, n_193);
  nor g23 (n_2662, n_119, n_192);
  nand g24 (n_2657, n_119, n_192);
  nor g25 (n_2658, n_118, n_191);
  nand g26 (n_2659, n_118, n_191);
  nor g27 (n_2668, n_117, n_190);
  nand g28 (n_2663, n_117, n_190);
  nor g29 (n_2664, n_116, n_189);
  nand g30 (n_2665, n_116, n_189);
  nor g31 (n_2674, n_115, n_188);
  nand g32 (n_2669, n_115, n_188);
  nor g33 (n_2670, n_114, n_187);
  nand g34 (n_2671, n_114, n_187);
  nor g35 (n_2680, n_113, n_186);
  nand g36 (n_2675, n_113, n_186);
  nor g37 (n_2676, n_112, n_185);
  nand g38 (n_2677, n_112, n_185);
  nor g39 (n_2686, n_111, n_184);
  nand g40 (n_2681, n_111, n_184);
  nor g41 (n_2682, n_110, n_183);
  nand g42 (n_2683, n_110, n_183);
  nor g43 (n_2692, n_109, n_182);
  nand g44 (n_2687, n_109, n_182);
  nor g45 (n_2688, n_108, n_181);
  nand g46 (n_2689, n_108, n_181);
  nor g47 (n_2698, n_107, n_180);
  nand g48 (n_2693, n_107, n_180);
  nor g49 (n_2694, n_106, n_179);
  nand g50 (n_2695, n_106, n_179);
  nor g51 (n_2704, n_105, n_178);
  nand g52 (n_2699, n_105, n_178);
  nor g53 (n_2700, n_104, n_177);
  nand g54 (n_2701, n_104, n_177);
  nor g55 (n_2710, n_103, n_176);
  nand g56 (n_2705, n_103, n_176);
  nor g57 (n_2706, n_102, n_175);
  nand g58 (n_2707, n_102, n_175);
  nor g59 (n_2716, n_101, n_174);
  nand g60 (n_2711, n_101, n_174);
  nor g61 (n_2712, n_100, n_173);
  nand g62 (n_2713, n_100, n_173);
  nor g63 (n_2722, n_99, n_172);
  nand g64 (n_2717, n_99, n_172);
  nor g65 (n_2718, n_98, n_171);
  nand g66 (n_2719, n_98, n_171);
  nor g67 (n_2728, n_97, n_170);
  nand g68 (n_2723, n_97, n_170);
  nor g69 (n_2724, n_96, n_169);
  nand g70 (n_2725, n_96, n_169);
  nor g71 (n_2734, n_95, n_168);
  nand g72 (n_2729, n_95, n_168);
  nor g73 (n_2730, n_94, n_167);
  nand g74 (n_2731, n_94, n_167);
  nor g75 (n_2740, n_93, n_166);
  nand g76 (n_2735, n_93, n_166);
  nor g77 (n_2736, n_92, n_165);
  nand g78 (n_2737, n_92, n_165);
  nor g79 (n_2746, n_91, n_164);
  nand g80 (n_2741, n_91, n_164);
  nor g81 (n_2742, n_90, n_163);
  nand g82 (n_2743, n_90, n_163);
  nor g83 (n_2752, n_89, n_162);
  nand g84 (n_2747, n_89, n_162);
  nor g85 (n_2748, n_88, n_161);
  nand g86 (n_2749, n_88, n_161);
  nor g87 (n_2758, n_87, n_160);
  nand g88 (n_2753, n_87, n_160);
  nor g89 (n_2754, n_86, n_159);
  nand g90 (n_2755, n_86, n_159);
  nor g91 (n_2764, n_85, n_158);
  nand g92 (n_2759, n_85, n_158);
  nor g93 (n_2760, n_84, n_157);
  nand g94 (n_2761, n_84, n_157);
  nor g95 (n_2770, n_83, n_156);
  nand g96 (n_2765, n_83, n_156);
  nor g97 (n_2766, n_82, n_155);
  nand g98 (n_2767, n_82, n_155);
  nor g99 (n_2776, n_81, n_154);
  nand g100 (n_2771, n_81, n_154);
  nor g101 (n_2772, n_80, n_153);
  nand g102 (n_2773, n_80, n_153);
  nor g103 (n_2782, n_79, n_152);
  nand g104 (n_2777, n_79, n_152);
  nor g105 (n_2778, n_78, n_151);
  nand g106 (n_2779, n_78, n_151);
  nor g107 (n_2788, n_77, n_150);
  nand g108 (n_2783, n_77, n_150);
  nor g109 (n_2784, n_76, n_149);
  nand g110 (n_2785, n_76, n_149);
  nor g111 (n_2794, n_75, n_148);
  nand g112 (n_2789, n_75, n_148);
  nor g113 (n_2790, n_74, n_147);
  nand g114 (n_2791, n_74, n_147);
  nor g115 (n_2800, n_73, n_146);
  nand g116 (n_2795, n_73, n_146);
  nor g117 (n_2796, n_72, n_145);
  nand g118 (n_2797, n_72, n_145);
  nor g119 (n_2806, n_71, n_144);
  nand g120 (n_2801, n_71, n_144);
  nor g121 (n_2802, n_70, n_143);
  nand g122 (n_2803, n_70, n_143);
  nor g123 (n_2812, n_69, n_142);
  nand g124 (n_2807, n_69, n_142);
  nor g125 (n_2808, n_68, n_141);
  nand g126 (n_2809, n_68, n_141);
  nor g127 (n_2818, n_67, n_140);
  nand g128 (n_2813, n_67, n_140);
  nor g129 (n_2814, n_66, n_139);
  nand g130 (n_2815, n_66, n_139);
  nor g131 (n_2824, n_65, n_138);
  nand g132 (n_2819, n_65, n_138);
  nor g133 (n_2820, n_64, n_137);
  nand g134 (n_2821, n_64, n_137);
  nor g135 (n_2830, n_63, n_136);
  nand g136 (n_2825, n_63, n_136);
  nor g137 (n_2826, n_62, n_135);
  nand g138 (n_2827, n_62, n_135);
  nor g139 (n_2836, n_61, n_134);
  nand g140 (n_2831, n_61, n_134);
  nor g141 (n_2832, n_60, n_133);
  nand g142 (n_2833, n_60, n_133);
  nor g143 (n_2842, n_59, n_132);
  nand g144 (n_2837, n_59, n_132);
  nor g145 (n_2838, n_58, n_131);
  nand g146 (n_2839, n_58, n_131);
  nor g156 (n_2642, n_1002, n_2640);
  nor g160 (n_2648, n_2645, n_2646);
  nor g163 (n_2859, n_2650, n_2646);
  nor g164 (n_2654, n_2651, n_2652);
  nor g167 (n_2853, n_2656, n_2652);
  nor g168 (n_2660, n_2657, n_2658);
  nor g171 (n_2866, n_2662, n_2658);
  nor g172 (n_2666, n_2663, n_2664);
  nor g175 (n_2860, n_2668, n_2664);
  nor g176 (n_2672, n_2669, n_2670);
  nor g179 (n_2873, n_2674, n_2670);
  nor g180 (n_2678, n_2675, n_2676);
  nor g183 (n_2867, n_2680, n_2676);
  nor g184 (n_2684, n_2681, n_2682);
  nor g187 (n_2880, n_2686, n_2682);
  nor g188 (n_2690, n_2687, n_2688);
  nor g191 (n_2874, n_2692, n_2688);
  nor g192 (n_2696, n_2693, n_2694);
  nor g195 (n_2887, n_2698, n_2694);
  nor g196 (n_2702, n_2699, n_2700);
  nor g199 (n_2881, n_2704, n_2700);
  nor g200 (n_2708, n_2705, n_2706);
  nor g203 (n_2894, n_2710, n_2706);
  nor g204 (n_2714, n_2711, n_2712);
  nor g207 (n_2888, n_2716, n_2712);
  nor g208 (n_2720, n_2717, n_2718);
  nor g211 (n_2901, n_2722, n_2718);
  nor g212 (n_2726, n_2723, n_2724);
  nor g215 (n_2895, n_2728, n_2724);
  nor g216 (n_2732, n_2729, n_2730);
  nor g219 (n_2908, n_2734, n_2730);
  nor g220 (n_2738, n_2735, n_2736);
  nor g223 (n_2902, n_2740, n_2736);
  nor g224 (n_2744, n_2741, n_2742);
  nor g227 (n_2915, n_2746, n_2742);
  nor g228 (n_2750, n_2747, n_2748);
  nor g231 (n_2909, n_2752, n_2748);
  nor g232 (n_2756, n_2753, n_2754);
  nor g235 (n_2922, n_2758, n_2754);
  nor g236 (n_2762, n_2759, n_2760);
  nor g239 (n_2916, n_2764, n_2760);
  nor g240 (n_2768, n_2765, n_2766);
  nor g243 (n_2929, n_2770, n_2766);
  nor g244 (n_2774, n_2771, n_2772);
  nor g247 (n_2923, n_2776, n_2772);
  nor g248 (n_2780, n_2777, n_2778);
  nor g251 (n_2936, n_2782, n_2778);
  nor g252 (n_2786, n_2783, n_2784);
  nor g255 (n_2930, n_2788, n_2784);
  nor g256 (n_2792, n_2789, n_2790);
  nor g259 (n_2943, n_2794, n_2790);
  nor g260 (n_2798, n_2795, n_2796);
  nor g263 (n_2937, n_2800, n_2796);
  nor g264 (n_2804, n_2801, n_2802);
  nor g267 (n_2950, n_2806, n_2802);
  nor g268 (n_2810, n_2807, n_2808);
  nor g271 (n_2944, n_2812, n_2808);
  nor g272 (n_2816, n_2813, n_2814);
  nor g275 (n_2957, n_2818, n_2814);
  nor g276 (n_2822, n_2819, n_2820);
  nor g279 (n_2951, n_2824, n_2820);
  nor g280 (n_2828, n_2825, n_2826);
  nor g283 (n_2964, n_2830, n_2826);
  nor g284 (n_2834, n_2831, n_2832);
  nor g287 (n_2958, n_2836, n_2832);
  nor g288 (n_2840, n_2837, n_2838);
  nor g291 (n_2971, n_2842, n_2838);
  nor g292 (n_2846, n_2843, n_2844);
  nor g295 (n_2965, n_2848, n_2844);
  nand g302 (n_2972, n_2859, n_2853);
  nand g307 (n_2982, n_2866, n_2860);
  nand g312 (n_2977, n_2873, n_2867);
  nand g317 (n_2988, n_2880, n_2874);
  nand g322 (n_2983, n_2887, n_2881);
  nand g327 (n_2994, n_2894, n_2888);
  nand g332 (n_2989, n_2901, n_2895);
  nand g337 (n_3000, n_2908, n_2902);
  nand g342 (n_2995, n_2915, n_2909);
  nand g347 (n_3006, n_2922, n_2916);
  nand g352 (n_3001, n_2929, n_2923);
  nand g357 (n_3012, n_2936, n_2930);
  nand g362 (n_3007, n_2943, n_2937);
  nand g367 (n_3018, n_2950, n_2944);
  nand g372 (n_3013, n_2957, n_2951);
  nand g377 (n_3024, n_2964, n_2958);
  nand g382 (n_3019, n_2971, n_2965);
  nand g385 (n_3026, n_2975, n_2976);
  nor g386 (n_2980, n_2977, n_2978);
  nor g389 (n_3025, n_2982, n_2977);
  nor g390 (n_2986, n_2983, n_2984);
  nor g393 (n_3035, n_2988, n_2983);
  nor g394 (n_2992, n_2989, n_2990);
  nor g397 (n_3029, n_2994, n_2989);
  nor g398 (n_2998, n_2995, n_2996);
  nor g401 (n_3042, n_3000, n_2995);
  nor g402 (n_3004, n_3001, n_3002);
  nor g405 (n_3036, n_3006, n_3001);
  nor g406 (n_3010, n_3007, n_3008);
  nor g409 (n_3049, n_3012, n_3007);
  nor g410 (n_3016, n_3013, n_3014);
  nor g413 (n_3043, n_3018, n_3013);
  nor g414 (n_3022, n_3019, n_3020);
  nor g417 (n_3071, n_3024, n_3019);
  nand g418 (n_3028, n_3025, n_3026);
  nand g419 (n_3051, n_3027, n_3028);
  nand g424 (n_3050, n_3035, n_3029);
  nand g2913 (n_3060, n_3042, n_3036);
  nand g2918 (n_3055, n_3049, n_3043);
  nand g2921 (n_3062, n_3053, n_3054);
  nor g2922 (n_3058, n_3055, n_3056);
  nor g2925 (n_3061, n_3060, n_3055);
  nand g2926 (n_3064, n_3061, n_3062);
  nand g2927 (n_3072, n_3063, n_3064);
  nand g2930 (n_3069, n_3056, n_3066);
  nand g2931 (n_3067, n_3035, n_3051);
  nand g2932 (n_3079, n_3030, n_3067);
  nand g2933 (n_3068, n_3042, n_3062);
  nand g2934 (n_3084, n_3037, n_3068);
  nand g2935 (n_3070, n_3049, n_3069);
  nand g2936 (n_3089, n_3044, n_3070);
  nand g2937 (n_3074, n_3071, n_3072);
  nand g2938 (n_3207, n_3073, n_3074);
  nand g2941 (n_3096, n_2978, n_3076);
  nand g2944 (n_3099, n_2984, n_3078);
  nand g2947 (n_3102, n_2990, n_3081);
  nand g2950 (n_3105, n_2996, n_3083);
  nand g2953 (n_3108, n_3002, n_3086);
  nand g2956 (n_3111, n_3008, n_3088);
  nand g2959 (n_3114, n_3014, n_3091);
  nand g2962 (n_3117, n_3020, n_3093);
  nand g2964 (n_3123, n_2854, n_3094);
  nand g2965 (n_3095, n_2866, n_3026);
  nand g2966 (n_3128, n_2861, n_3095);
  nand g2967 (n_3097, n_2873, n_3096);
  nand g2968 (n_3133, n_2868, n_3097);
  nand g2969 (n_3098, n_2880, n_3051);
  nand g2970 (n_3138, n_2875, n_3098);
  nand g2971 (n_3100, n_2887, n_3099);
  nand g2972 (n_3143, n_2882, n_3100);
  nand g2973 (n_3101, n_2894, n_3079);
  nand g2974 (n_3148, n_2889, n_3101);
  nand g2975 (n_3103, n_2901, n_3102);
  nand g2976 (n_3153, n_2896, n_3103);
  nand g2977 (n_3104, n_2908, n_3062);
  nand g2978 (n_3158, n_2903, n_3104);
  nand g2979 (n_3106, n_2915, n_3105);
  nand g2980 (n_3163, n_2910, n_3106);
  nand g2981 (n_3107, n_2922, n_3084);
  nand g2982 (n_3168, n_2917, n_3107);
  nand g2983 (n_3109, n_2929, n_3108);
  nand g2984 (n_3173, n_2924, n_3109);
  nand g2985 (n_3110, n_2936, n_3069);
  nand g2986 (n_3178, n_2931, n_3110);
  nand g2987 (n_3112, n_2943, n_3111);
  nand g2988 (n_3183, n_2938, n_3112);
  nand g2989 (n_3113, n_2950, n_3089);
  nand g2990 (n_3188, n_2945, n_3113);
  nand g2991 (n_3115, n_2957, n_3114);
  nand g2992 (n_3193, n_2952, n_3115);
  nand g2993 (n_3116, n_2964, n_3072);
  nand g2994 (n_3198, n_2959, n_3116);
  nand g2995 (n_3118, n_2971, n_3117);
  nand g2996 (n_3203, n_2966, n_3118);
  nand g3002 (n_3217, n_2645, n_3122);
  nand g3005 (n_3221, n_2651, n_3125);
  nand g3008 (n_3225, n_2657, n_3127);
  nand g3011 (n_3229, n_2663, n_3130);
  nand g3014 (n_3233, n_2669, n_3132);
  nand g3017 (n_3237, n_2675, n_3135);
  nand g3020 (n_3241, n_2681, n_3137);
  nand g3023 (n_3245, n_2687, n_3140);
  nand g3026 (n_3249, n_2693, n_3142);
  nand g3029 (n_3253, n_2699, n_3145);
  nand g3032 (n_3257, n_2705, n_3147);
  nand g3035 (n_3261, n_2711, n_3150);
  nand g3038 (n_3265, n_2717, n_3152);
  nand g3041 (n_3269, n_2723, n_3155);
  nand g3044 (n_3273, n_2729, n_3157);
  nand g3047 (n_3277, n_2735, n_3160);
  nand g3050 (n_3281, n_2741, n_3162);
  nand g3053 (n_3285, n_2747, n_3165);
  nand g3056 (n_3289, n_2753, n_3167);
  nand g3059 (n_3293, n_2759, n_3170);
  nand g3062 (n_3297, n_2765, n_3172);
  nand g3065 (n_3301, n_2771, n_3175);
  nand g3068 (n_3305, n_2777, n_3177);
  nand g3071 (n_3309, n_2783, n_3180);
  nand g3074 (n_3313, n_2789, n_3182);
  nand g3077 (n_3317, n_2795, n_3185);
  nand g3080 (n_3321, n_2801, n_3187);
  nand g3083 (n_3325, n_2807, n_3190);
  nand g3086 (n_3329, n_2813, n_3192);
  nand g3089 (n_3333, n_2819, n_3195);
  nand g3092 (n_3337, n_2825, n_3197);
  nand g3095 (n_3341, n_2831, n_3200);
  nand g3098 (n_3345, n_2837, n_3202);
  nand g3101 (n_3349, n_2843, n_3205);
  xnor g3114 (Z[5], n_3217, n_3218);
  xnor g3116 (Z[6], n_3123, n_3219);
  xnor g3119 (Z[7], n_3221, n_3222);
  xnor g3121 (Z[8], n_3026, n_3223);
  xnor g3124 (Z[9], n_3225, n_3226);
  xnor g3126 (Z[10], n_3128, n_3227);
  xnor g3129 (Z[11], n_3229, n_3230);
  xnor g3131 (Z[12], n_3096, n_3231);
  xnor g3134 (Z[13], n_3233, n_3234);
  xnor g3136 (Z[14], n_3133, n_3235);
  xnor g3139 (Z[15], n_3237, n_3238);
  xnor g3141 (Z[16], n_3051, n_3239);
  xnor g3144 (Z[17], n_3241, n_3242);
  xnor g3146 (Z[18], n_3138, n_3243);
  xnor g3149 (Z[19], n_3245, n_3246);
  xnor g3151 (Z[20], n_3099, n_3247);
  xnor g3154 (Z[21], n_3249, n_3250);
  xnor g3156 (Z[22], n_3143, n_3251);
  xnor g3159 (Z[23], n_3253, n_3254);
  xnor g3161 (Z[24], n_3079, n_3255);
  xnor g3164 (Z[25], n_3257, n_3258);
  xnor g3166 (Z[26], n_3148, n_3259);
  xnor g3169 (Z[27], n_3261, n_3262);
  xnor g3171 (Z[28], n_3102, n_3263);
  xnor g3174 (Z[29], n_3265, n_3266);
  xnor g3176 (Z[30], n_3153, n_3267);
  xnor g3179 (Z[31], n_3269, n_3270);
  xnor g3181 (Z[32], n_3062, n_3271);
  xnor g3184 (Z[33], n_3273, n_3274);
  xnor g3186 (Z[34], n_3158, n_3275);
  xnor g3189 (Z[35], n_3277, n_3278);
  xnor g3191 (Z[36], n_3105, n_3279);
  xnor g3194 (Z[37], n_3281, n_3282);
  xnor g3196 (Z[38], n_3163, n_3283);
  xnor g3199 (Z[39], n_3285, n_3286);
  xnor g3201 (Z[40], n_3084, n_3287);
  xnor g3204 (Z[41], n_3289, n_3290);
  xnor g3206 (Z[42], n_3168, n_3291);
  xnor g3209 (Z[43], n_3293, n_3294);
  xnor g3211 (Z[44], n_3108, n_3295);
  xnor g3214 (Z[45], n_3297, n_3298);
  xnor g3216 (Z[46], n_3173, n_3299);
  xnor g3219 (Z[47], n_3301, n_3302);
  xnor g3221 (Z[48], n_3069, n_3303);
  xnor g3224 (Z[49], n_3305, n_3306);
  xnor g3226 (Z[50], n_3178, n_3307);
  xnor g3229 (Z[51], n_3309, n_3310);
  xnor g3231 (Z[52], n_3111, n_3311);
  xnor g3234 (Z[53], n_3313, n_3314);
  xnor g3236 (Z[54], n_3183, n_3315);
  xnor g3239 (Z[55], n_3317, n_3318);
  xnor g3241 (Z[56], n_3089, n_3319);
  xnor g3244 (Z[57], n_3321, n_3322);
  xnor g3246 (Z[58], n_3188, n_3323);
  xnor g3249 (Z[59], n_3325, n_3326);
  xnor g3251 (Z[60], n_3114, n_3327);
  xnor g3254 (Z[61], n_3329, n_3330);
  xnor g3256 (Z[62], n_3193, n_3331);
  xnor g3259 (Z[63], n_3333, n_3334);
  xnor g3261 (Z[64], n_3072, n_3335);
  xnor g3264 (Z[65], n_3337, n_3338);
  xnor g3266 (Z[66], n_3198, n_3339);
  xnor g3269 (Z[67], n_3341, n_3342);
  xnor g3271 (Z[68], n_3117, n_3343);
  xnor g3274 (Z[69], n_3345, n_3346);
  xnor g3276 (Z[70], n_3203, n_3347);
  xnor g3279 (Z[71], n_3349, n_3350);
  or g3294 (n_282, wc, wc0, n_122);
  not gc0 (wc0, n_1002);
  not gc (wc, n_1016);
  or g3295 (n_291, wc1, wc2, n_276);
  not gc2 (wc2, n_1016);
  not gc1 (wc1, n_1035);
  or g3296 (n_304, wc3, n_281, n_276);
  not gc3 (wc3, n_1063);
  or g3297 (n_321, wc4, wc5, n_281);
  not gc5 (wc5, n_1098);
  not gc4 (wc4, n_1099);
  or g3298 (n_343, wc6, wc7, n_281);
  not gc7 (wc7, n_1146);
  not gc6 (wc6, n_1147);
  or g3299 (n_391, wc8, wc9, n_276);
  not gc9 (wc9, n_1147);
  not gc8 (wc8, n_1194);
  or g3300 (n_419, wc10, wc11, n_281);
  not gc11 (wc11, n_1323);
  not gc10 (wc10, n_1324);
  or g3301 (n_445, wc12, wc13, n_290);
  not gc13 (wc13, n_1263);
  not gc12 (wc12, n_1387);
  or g3302 (n_473, wc14, wc15, n_303);
  not gc15 (wc15, n_1327);
  not gc14 (wc14, n_1451);
  or g3303 (n_501, wc16, wc17, n_320);
  not gc17 (wc17, n_1256);
  not gc16 (wc16, n_1515);
  or g3304 (n_529, wc18, wc19, n_341);
  not gc19 (wc19, n_1320);
  not gc18 (wc18, n_1579);
  or g3305 (n_557, wc20, wc21, n_366);
  not gc21 (wc21, n_1384);
  not gc20 (wc20, n_1643);
  xnor g3306 (n_2373, A[53], A[51]);
  or g3307 (n_2374, wc22, A[53]);
  not gc22 (wc22, A[51]);
  or g3308 (n_2376, wc23, A[53]);
  not gc23 (wc23, A[39]);
  xnor g3309 (n_2413, A[52], A[48]);
  or g3310 (n_2414, wc24, A[52]);
  not gc24 (wc24, A[48]);
  or g3311 (n_2379, wc25, A[53]);
  not gc25 (wc25, A[45]);
  xnor g3312 (n_941, n_2513, A[50]);
  or g3313 (n_2515, wc26, A[50]);
  not gc26 (wc26, A[48]);
  or g3314 (n_2516, wc27, A[50]);
  not gc27 (wc27, A[46]);
  or g3316 (n_2596, wc28, A[53]);
  not gc28 (wc28, A[47]);
  xnor g3317 (n_987, n_2605, A[52]);
  or g3318 (n_2608, wc29, A[52]);
  not gc29 (wc29, A[50]);
  or g3319 (n_2616, wc30, A[53]);
  not gc30 (wc30, A[49]);
  or g3321 (n_2622, A[50], wc31);
  not gc31 (wc31, A[52]);
  or g3322 (n_2628, wc32, A[53]);
  not gc32 (wc32, A[50]);
  and g3323 (n_2844, wc33, A[53]);
  not gc33 (wc33, A[52]);
  or g3324 (n_2845, wc34, A[53]);
  not gc34 (wc34, A[52]);
  or g3325 (n_372, wc35, wc36, n_281);
  not gc36 (wc36, n_1203);
  not gc35 (wc35, n_1204);
  or g3326 (n_2472, A[52], wc37);
  not gc37 (wc37, n_915);
  and g3327 (n_2851, wc38, n_999);
  not gc38 (wc38, n_2642);
  or g3329 (n_3211, n_2644, wc39);
  not gc39 (wc39, n_1002);
  or g3330 (n_3214, n_2640, wc40);
  not gc40 (wc40, n_999);
  xnor g3331 (n_875, n_2377, A[53]);
  or g3332 (n_2380, wc41, A[53]);
  not gc41 (wc41, A[37]);
  or g3333 (n_2415, A[52], wc42);
  not gc42 (wc42, n_886);
  xnor g3334 (n_2469, n_886, A[52]);
  xnor g3335 (n_961, n_938, n_2605);
  or g3336 (n_2555, A[50], wc43);
  not gc43 (wc43, n_938);
  xnor g3337 (n_2585, n_938, A[52]);
  or g3338 (n_2586, A[52], wc44);
  not gc44 (wc44, n_938);
  or g3339 (n_2588, A[52], wc45);
  not gc45 (wc45, n_975);
  xnor g3340 (n_59, n_2277, n_994);
  or g3341 (n_2623, A[50], wc46);
  not gc46 (wc46, n_994);
  and g3342 (n_2848, A[52], wc47);
  not gc47 (wc47, n_130);
  or g3343 (n_2843, A[52], wc48);
  not gc48 (wc48, n_130);
  or g3344 (n_3215, wc49, n_2650);
  not gc49 (wc49, n_2645);
  or g3345 (n_3350, wc50, n_2844);
  not gc50 (wc50, n_2845);
  and g3346 (n_2854, wc51, n_2647);
  not gc51 (wc51, n_2648);
  not g3347 (Z[2], n_3211);
  or g3348 (n_3218, wc52, n_2646);
  not gc52 (wc52, n_2647);
  or g3349 (n_3219, wc53, n_2656);
  not gc53 (wc53, n_2651);
  and g3350 (n_2856, wc54, n_2653);
  not gc54 (wc54, n_2654);
  and g3351 (n_2968, n_2845, wc55);
  not gc55 (wc55, n_2846);
  or g3354 (n_3222, wc56, n_2652);
  not gc56 (wc56, n_2653);
  or g3355 (n_3347, wc57, n_2848);
  not gc57 (wc57, n_2843);
  and g3356 (n_2861, wc58, n_2659);
  not gc58 (wc58, n_2660);
  and g3357 (n_2857, wc59, n_2853);
  not gc59 (wc59, n_2854);
  or g3358 (n_3094, n_2851, wc60);
  not gc60 (wc60, n_2859);
  or g3359 (n_3122, n_2650, n_2851);
  xor g3360 (Z[3], n_1002, n_3214);
  xor g3361 (Z[4], n_2851, n_3215);
  or g3362 (n_3223, wc61, n_2662);
  not gc61 (wc61, n_2657);
  or g3363 (n_3226, wc62, n_2658);
  not gc62 (wc62, n_2659);
  and g3364 (n_2966, wc63, n_2839);
  not gc63 (wc63, n_2840);
  and g3365 (n_2975, wc64, n_2856);
  not gc64 (wc64, n_2857);
  or g3366 (n_2976, n_2972, n_2851);
  or g3367 (n_3227, wc65, n_2668);
  not gc65 (wc65, n_2663);
  or g3368 (n_3343, wc66, n_2842);
  not gc66 (wc66, n_2837);
  or g3369 (n_3346, wc67, n_2838);
  not gc67 (wc67, n_2839);
  and g3370 (n_2863, wc68, n_2665);
  not gc68 (wc68, n_2666);
  and g3371 (n_2868, wc69, n_2671);
  not gc69 (wc69, n_2672);
  and g3372 (n_2969, wc70, n_2965);
  not gc70 (wc70, n_2966);
  or g3373 (n_3125, wc71, n_2656);
  not gc71 (wc71, n_3123);
  or g3374 (n_3230, wc72, n_2664);
  not gc72 (wc72, n_2665);
  or g3375 (n_3231, wc73, n_2674);
  not gc73 (wc73, n_2669);
  or g3376 (n_3234, wc74, n_2670);
  not gc74 (wc74, n_2671);
  and g3377 (n_2870, wc75, n_2677);
  not gc75 (wc75, n_2678);
  and g3378 (n_2961, wc76, n_2833);
  not gc76 (wc76, n_2834);
  and g3379 (n_2864, wc77, n_2860);
  not gc77 (wc77, n_2861);
  and g3380 (n_3021, wc78, n_2968);
  not gc78 (wc78, n_2969);
  or g3381 (n_3127, wc79, n_2662);
  not gc79 (wc79, n_3026);
  or g3382 (n_3235, wc80, n_2680);
  not gc80 (wc80, n_2675);
  or g3383 (n_3238, wc81, n_2676);
  not gc81 (wc81, n_2677);
  or g3384 (n_3338, wc82, n_2826);
  not gc82 (wc82, n_2827);
  or g3385 (n_3339, wc83, n_2836);
  not gc83 (wc83, n_2831);
  or g3386 (n_3342, wc84, n_2832);
  not gc84 (wc84, n_2833);
  and g3387 (n_2875, wc85, n_2683);
  not gc85 (wc85, n_2684);
  and g3388 (n_2877, wc86, n_2689);
  not gc86 (wc86, n_2690);
  and g3389 (n_2959, wc87, n_2827);
  not gc87 (wc87, n_2828);
  and g3390 (n_2978, wc88, n_2863);
  not gc88 (wc88, n_2864);
  and g3391 (n_2871, wc89, n_2867);
  not gc89 (wc89, n_2868);
  or g3392 (n_3076, wc90, n_2982);
  not gc90 (wc90, n_3026);
  or g3393 (n_3239, wc91, n_2686);
  not gc91 (wc91, n_2681);
  or g3394 (n_3242, wc92, n_2682);
  not gc92 (wc92, n_2683);
  or g3395 (n_3243, wc93, n_2692);
  not gc93 (wc93, n_2687);
  or g3396 (n_3246, wc94, n_2688);
  not gc94 (wc94, n_2689);
  or g3397 (n_3247, wc95, n_2698);
  not gc95 (wc95, n_2693);
  or g3398 (n_3334, wc96, n_2820);
  not gc96 (wc96, n_2821);
  or g3399 (n_3335, wc97, n_2830);
  not gc97 (wc97, n_2825);
  and g3400 (n_2882, wc98, n_2695);
  not gc98 (wc98, n_2696);
  and g3401 (n_2952, wc99, n_2815);
  not gc99 (wc99, n_2816);
  and g3402 (n_2954, wc100, n_2821);
  not gc100 (wc100, n_2822);
  and g3403 (n_2979, wc101, n_2870);
  not gc101 (wc101, n_2871);
  and g3404 (n_2878, wc102, n_2874);
  not gc102 (wc102, n_2875);
  and g3405 (n_2962, wc103, n_2958);
  not gc103 (wc103, n_2959);
  or g3406 (n_3130, wc104, n_2668);
  not gc104 (wc104, n_3128);
  or g3407 (n_3250, wc105, n_2694);
  not gc105 (wc105, n_2695);
  or g3408 (n_3251, wc106, n_2704);
  not gc106 (wc106, n_2699);
  or g3409 (n_3327, wc107, n_2818);
  not gc107 (wc107, n_2813);
  or g3410 (n_3330, wc108, n_2814);
  not gc108 (wc108, n_2815);
  or g3411 (n_3331, wc109, n_2824);
  not gc109 (wc109, n_2819);
  and g3412 (n_2884, wc110, n_2701);
  not gc110 (wc110, n_2702);
  and g3413 (n_2889, wc111, n_2707);
  not gc111 (wc111, n_2708);
  and g3414 (n_2891, wc112, n_2713);
  not gc112 (wc112, n_2714);
  and g3415 (n_2896, wc113, n_2719);
  not gc113 (wc113, n_2720);
  and g3416 (n_2898, wc114, n_2725);
  not gc114 (wc114, n_2726);
  and g3417 (n_2903, wc115, n_2731);
  not gc115 (wc115, n_2732);
  and g3418 (n_2905, wc116, n_2737);
  not gc116 (wc116, n_2738);
  and g3419 (n_2910, wc117, n_2743);
  not gc117 (wc117, n_2744);
  and g3420 (n_2912, wc118, n_2749);
  not gc118 (wc118, n_2750);
  and g3421 (n_2917, wc119, n_2755);
  not gc119 (wc119, n_2756);
  and g3422 (n_2919, wc120, n_2761);
  not gc120 (wc120, n_2762);
  and g3423 (n_2924, wc121, n_2767);
  not gc121 (wc121, n_2768);
  and g3424 (n_2926, wc122, n_2773);
  not gc122 (wc122, n_2774);
  and g3425 (n_2931, wc123, n_2779);
  not gc123 (wc123, n_2780);
  and g3426 (n_2933, wc124, n_2785);
  not gc124 (wc124, n_2786);
  and g3427 (n_2938, wc125, n_2791);
  not gc125 (wc125, n_2792);
  and g3428 (n_2984, wc126, n_2877);
  not gc126 (wc126, n_2878);
  and g3429 (n_2955, wc127, n_2951);
  not gc127 (wc127, n_2952);
  and g3430 (n_3020, wc128, n_2961);
  not gc128 (wc128, n_2962);
  or g3431 (n_3132, wc129, n_2674);
  not gc129 (wc129, n_3096);
  or g3432 (n_3254, wc130, n_2700);
  not gc130 (wc130, n_2701);
  or g3433 (n_3255, wc131, n_2710);
  not gc131 (wc131, n_2705);
  or g3434 (n_3258, wc132, n_2706);
  not gc132 (wc132, n_2707);
  or g3435 (n_3259, wc133, n_2716);
  not gc133 (wc133, n_2711);
  or g3436 (n_3262, wc134, n_2712);
  not gc134 (wc134, n_2713);
  or g3437 (n_3263, wc135, n_2722);
  not gc135 (wc135, n_2717);
  or g3438 (n_3266, wc136, n_2718);
  not gc136 (wc136, n_2719);
  or g3439 (n_3267, wc137, n_2728);
  not gc137 (wc137, n_2723);
  or g3440 (n_3270, wc138, n_2724);
  not gc138 (wc138, n_2725);
  or g3441 (n_3271, wc139, n_2734);
  not gc139 (wc139, n_2729);
  or g3442 (n_3274, wc140, n_2730);
  not gc140 (wc140, n_2731);
  or g3443 (n_3275, wc141, n_2740);
  not gc141 (wc141, n_2735);
  or g3444 (n_3278, wc142, n_2736);
  not gc142 (wc142, n_2737);
  or g3445 (n_3279, wc143, n_2746);
  not gc143 (wc143, n_2741);
  or g3446 (n_3282, wc144, n_2742);
  not gc144 (wc144, n_2743);
  or g3447 (n_3283, wc145, n_2752);
  not gc145 (wc145, n_2747);
  or g3448 (n_3286, wc146, n_2748);
  not gc146 (wc146, n_2749);
  or g3449 (n_3287, wc147, n_2758);
  not gc147 (wc147, n_2753);
  or g3450 (n_3290, wc148, n_2754);
  not gc148 (wc148, n_2755);
  or g3451 (n_3291, wc149, n_2764);
  not gc149 (wc149, n_2759);
  or g3452 (n_3294, wc150, n_2760);
  not gc150 (wc150, n_2761);
  or g3453 (n_3295, wc151, n_2770);
  not gc151 (wc151, n_2765);
  or g3454 (n_3298, wc152, n_2766);
  not gc152 (wc152, n_2767);
  or g3455 (n_3299, wc153, n_2776);
  not gc153 (wc153, n_2771);
  or g3456 (n_3302, wc154, n_2772);
  not gc154 (wc154, n_2773);
  or g3457 (n_3303, wc155, n_2782);
  not gc155 (wc155, n_2777);
  or g3458 (n_3306, wc156, n_2778);
  not gc156 (wc156, n_2779);
  or g3459 (n_3307, wc157, n_2788);
  not gc157 (wc157, n_2783);
  or g3460 (n_3310, wc158, n_2784);
  not gc158 (wc158, n_2785);
  or g3461 (n_3311, wc159, n_2794);
  not gc159 (wc159, n_2789);
  or g3462 (n_3314, wc160, n_2790);
  not gc160 (wc160, n_2791);
  or g3463 (n_3315, wc161, n_2800);
  not gc161 (wc161, n_2795);
  and g3464 (n_2940, wc162, n_2797);
  not gc162 (wc162, n_2798);
  and g3465 (n_2885, wc163, n_2881);
  not gc163 (wc163, n_2882);
  and g3466 (n_2892, wc164, n_2888);
  not gc164 (wc164, n_2889);
  and g3467 (n_2899, wc165, n_2895);
  not gc165 (wc165, n_2896);
  and g3468 (n_2906, wc166, n_2902);
  not gc166 (wc166, n_2903);
  and g3469 (n_2913, wc167, n_2909);
  not gc167 (wc167, n_2910);
  and g3470 (n_2920, wc168, n_2916);
  not gc168 (wc168, n_2917);
  and g3471 (n_2927, wc169, n_2923);
  not gc169 (wc169, n_2924);
  and g3472 (n_2934, wc170, n_2930);
  not gc170 (wc170, n_2931);
  and g3473 (n_3015, wc171, n_2954);
  not gc171 (wc171, n_2955);
  and g3474 (n_3027, n_2979, wc172);
  not gc172 (wc172, n_2980);
  or g3475 (n_3318, wc173, n_2796);
  not gc173 (wc173, n_2797);
  or g3476 (n_3319, wc174, n_2806);
  not gc174 (wc174, n_2801);
  or g3477 (n_3326, wc175, n_2808);
  not gc175 (wc175, n_2809);
  and g3478 (n_2945, wc176, n_2803);
  not gc176 (wc176, n_2804);
  and g3479 (n_2947, wc177, n_2809);
  not gc177 (wc177, n_2810);
  and g3480 (n_2985, wc178, n_2884);
  not gc178 (wc178, n_2885);
  and g3481 (n_2990, wc179, n_2891);
  not gc179 (wc179, n_2892);
  and g3482 (n_2991, wc180, n_2898);
  not gc180 (wc180, n_2899);
  and g3483 (n_2996, wc181, n_2905);
  not gc181 (wc181, n_2906);
  and g3484 (n_2997, wc182, n_2912);
  not gc182 (wc182, n_2913);
  and g3485 (n_3002, wc183, n_2919);
  not gc183 (wc183, n_2920);
  and g3486 (n_3003, wc184, n_2926);
  not gc184 (wc184, n_2927);
  and g3487 (n_3008, wc185, n_2933);
  not gc185 (wc185, n_2934);
  and g3488 (n_2941, wc186, n_2937);
  not gc186 (wc186, n_2938);
  and g3489 (n_3073, n_3021, wc187);
  not gc187 (wc187, n_3022);
  or g3490 (n_3135, wc188, n_2680);
  not gc188 (wc188, n_3133);
  or g3491 (n_3322, wc189, n_2802);
  not gc189 (wc189, n_2803);
  or g3492 (n_3323, wc190, n_2812);
  not gc190 (wc190, n_2807);
  and g3493 (n_3009, wc191, n_2940);
  not gc191 (wc191, n_2941);
  and g3494 (n_2948, wc192, n_2944);
  not gc192 (wc192, n_2945);
  or g3495 (n_3078, wc193, n_2988);
  not gc193 (wc193, n_3051);
  or g3496 (n_3137, wc194, n_2686);
  not gc194 (wc194, n_3051);
  and g3497 (n_3014, wc195, n_2947);
  not gc195 (wc195, n_2948);
  and g3498 (n_3030, n_2985, wc196);
  not gc196 (wc196, n_2986);
  and g3499 (n_3032, n_2991, wc197);
  not gc197 (wc197, n_2992);
  and g3500 (n_3037, n_2997, wc198);
  not gc198 (wc198, n_2998);
  and g3501 (n_3039, n_3003, wc199);
  not gc199 (wc199, n_3004);
  or g3502 (n_3054, n_3050, wc200);
  not gc200 (wc200, n_3051);
  and g3503 (n_3044, n_3009, wc201);
  not gc201 (wc201, n_3010);
  and g3504 (n_3033, wc202, n_3029);
  not gc202 (wc202, n_3030);
  and g3505 (n_3040, wc203, n_3036);
  not gc203 (wc203, n_3037);
  or g3506 (n_3140, wc204, n_2692);
  not gc204 (wc204, n_3138);
  or g3507 (n_3142, wc205, n_2698);
  not gc205 (wc205, n_3099);
  and g3508 (n_3046, n_3015, wc206);
  not gc206 (wc206, n_3016);
  and g3509 (n_3053, wc207, n_3032);
  not gc207 (wc207, n_3033);
  and g3510 (n_3056, wc208, n_3039);
  not gc208 (wc208, n_3040);
  and g3511 (n_3047, wc209, n_3043);
  not gc209 (wc209, n_3044);
  or g3512 (n_3081, wc210, n_2994);
  not gc210 (wc210, n_3079);
  or g3513 (n_3147, wc211, n_2710);
  not gc211 (wc211, n_3079);
  or g3514 (n_3145, wc212, n_2704);
  not gc212 (wc212, n_3143);
  and g3515 (n_3057, wc213, n_3046);
  not gc213 (wc213, n_3047);
  or g3516 (n_3066, wc214, n_3060);
  not gc214 (wc214, n_3062);
  or g3517 (n_3083, wc215, n_3000);
  not gc215 (wc215, n_3062);
  or g3518 (n_3150, wc216, n_2716);
  not gc216 (wc216, n_3148);
  or g3519 (n_3152, wc217, n_2722);
  not gc217 (wc217, n_3102);
  or g3520 (n_3157, wc218, n_2734);
  not gc218 (wc218, n_3062);
  and g3521 (n_3063, n_3057, wc219);
  not gc219 (wc219, n_3058);
  or g3522 (n_3086, wc220, n_3006);
  not gc220 (wc220, n_3084);
  or g3523 (n_3088, wc221, n_3012);
  not gc221 (wc221, n_3069);
  or g3524 (n_3155, wc222, n_2728);
  not gc222 (wc222, n_3153);
  or g3525 (n_3160, wc223, n_2740);
  not gc223 (wc223, n_3158);
  or g3526 (n_3162, wc224, n_2746);
  not gc224 (wc224, n_3105);
  or g3527 (n_3167, wc225, n_2758);
  not gc225 (wc225, n_3084);
  or g3528 (n_3177, wc226, n_2782);
  not gc226 (wc226, n_3069);
  or g3529 (n_3091, wc227, n_3018);
  not gc227 (wc227, n_3089);
  or g3530 (n_3093, wc228, n_3024);
  not gc228 (wc228, n_3072);
  or g3531 (n_3165, wc229, n_2752);
  not gc229 (wc229, n_3163);
  or g3532 (n_3170, wc230, n_2764);
  not gc230 (wc230, n_3168);
  or g3533 (n_3172, wc231, n_2770);
  not gc231 (wc231, n_3108);
  or g3534 (n_3180, wc232, n_2788);
  not gc232 (wc232, n_3178);
  or g3535 (n_3182, wc233, n_2794);
  not gc233 (wc233, n_3111);
  or g3536 (n_3187, wc234, n_2806);
  not gc234 (wc234, n_3089);
  or g3537 (n_3197, wc235, n_2830);
  not gc235 (wc235, n_3072);
  or g3538 (n_3175, wc236, n_2776);
  not gc236 (wc236, n_3173);
  or g3539 (n_3185, wc237, n_2800);
  not gc237 (wc237, n_3183);
  or g3540 (n_3190, wc238, n_2812);
  not gc238 (wc238, n_3188);
  or g3541 (n_3192, wc239, n_2818);
  not gc239 (wc239, n_3114);
  or g3542 (n_3200, wc240, n_2836);
  not gc240 (wc240, n_3198);
  or g3543 (n_3202, wc241, n_2842);
  not gc241 (wc241, n_3117);
  not g3544 (Z[72], n_3207);
  or g3545 (n_3195, wc242, n_2824);
  not gc242 (wc242, n_3193);
  or g3546 (n_3205, n_2848, wc243);
  not gc243 (wc243, n_3203);
endmodule

module mult_signed_const_12373_GENERIC(A, Z);
  input [53:0] A;
  output [72:0] Z;
  wire [53:0] A;
  wire [72:0] Z;
  mult_signed_const_12373_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_12824_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [56:0] A;
  output [75:0] Z;
  wire [56:0] A;
  wire [75:0] Z;
  wire n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68;
  wire n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190;
  wire n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201, n_202, n_203, n_204, n_205, n_206;
  wire n_207, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_298, n_299, n_300, n_301, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_310, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371;
  wire n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395;
  wire n_396, n_397, n_398, n_399, n_400, n_401, n_403, n_404;
  wire n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412;
  wire n_413, n_414, n_415, n_417, n_418, n_419, n_420, n_421;
  wire n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429;
  wire n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437;
  wire n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445;
  wire n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453;
  wire n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461;
  wire n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477;
  wire n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485;
  wire n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501;
  wire n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509;
  wire n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517;
  wire n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_530, n_531, n_532, n_533;
  wire n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541;
  wire n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_555, n_556, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_566, n_567, n_568, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581;
  wire n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589;
  wire n_590, n_591, n_592, n_593, n_594, n_595, n_596, n_597;
  wire n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605;
  wire n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613;
  wire n_614, n_615, n_616, n_617, n_618, n_619, n_620, n_621;
  wire n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629;
  wire n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637;
  wire n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645;
  wire n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
  wire n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669;
  wire n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677;
  wire n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685;
  wire n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693;
  wire n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701;
  wire n_702, n_703, n_704, n_705, n_706, n_707, n_708, n_709;
  wire n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717;
  wire n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725;
  wire n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733;
  wire n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741;
  wire n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749;
  wire n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757;
  wire n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765;
  wire n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781;
  wire n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789;
  wire n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797;
  wire n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805;
  wire n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813;
  wire n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821;
  wire n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829;
  wire n_830, n_831, n_832, n_833, n_834, n_835, n_836, n_837;
  wire n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845;
  wire n_846, n_847, n_848, n_849, n_850, n_851, n_852, n_853;
  wire n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_861;
  wire n_862, n_863, n_864, n_865, n_866, n_867, n_868, n_869;
  wire n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877;
  wire n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885;
  wire n_886, n_887, n_888, n_891, n_892, n_893, n_894, n_895;
  wire n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903;
  wire n_904, n_908, n_909, n_910, n_911, n_912, n_913, n_914;
  wire n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_923;
  wire n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931;
  wire n_932, n_933, n_934, n_935, n_936, n_939, n_940, n_941;
  wire n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949;
  wire n_950, n_951, n_953, n_954, n_956, n_957, n_958, n_959;
  wire n_960, n_961, n_962, n_963, n_964, n_968, n_969, n_970;
  wire n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_979;
  wire n_980, n_983, n_984, n_985, n_986, n_987, n_988, n_993;
  wire n_994, n_995, n_996, n_997, n_998, n_999, n_1001, n_1004;
  wire n_1005, n_1006, n_1007, n_1008, n_1014, n_1015, n_1016, n_1017;
  wire n_1021, n_1022, n_1023, n_1024, n_1028, n_1029, n_1030, n_1031;
  wire n_1033, n_1035, n_1036, n_1040, n_1041, n_1043, n_1044, n_1047;
  wire n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057;
  wire n_1058, n_1059, n_1060, n_1062, n_1063, n_1064, n_1065, n_1066;
  wire n_1067, n_1068, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075;
  wire n_1076, n_1078, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085;
  wire n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095;
  wire n_1096, n_1097, n_1100, n_1102, n_1103, n_1104, n_1105, n_1106;
  wire n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114;
  wire n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123;
  wire n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131;
  wire n_1134, n_1135, n_1136, n_1138, n_1139, n_1140, n_1141, n_1142;
  wire n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150;
  wire n_1151, n_1152, n_1154, n_1158, n_1159, n_1160, n_1161, n_1162;
  wire n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170;
  wire n_1171, n_1172, n_1173, n_1174, n_1175, n_1177, n_1178, n_1180;
  wire n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188;
  wire n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1197;
  wire n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209;
  wire n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217;
  wire n_1218, n_1219, n_1220, n_1226, n_1227, n_1230, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240;
  wire n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1249, n_1250;
  wire n_1251, n_1253, n_1254, n_1256, n_1257, n_1258, n_1259, n_1260;
  wire n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268;
  wire n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276;
  wire n_1280, n_1281, n_1282, n_1283, n_1284, n_1286, n_1287, n_1288;
  wire n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304;
  wire n_1305, n_1306, n_1307, n_1308, n_1309, n_1314, n_1315, n_1318;
  wire n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326;
  wire n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334;
  wire n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1346;
  wire n_1348, n_1350, n_1351, n_1352, n_1354, n_1355, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373;
  wire n_1376, n_1377, n_1378, n_1379, n_1380, n_1382, n_1383, n_1384;
  wire n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392;
  wire n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400;
  wire n_1401, n_1402, n_1403, n_1404, n_1405, n_1408, n_1410, n_1411;
  wire n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421;
  wire n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429;
  wire n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437;
  wire n_1438, n_1439, n_1440, n_1442, n_1443, n_1446, n_1447, n_1448;
  wire n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456;
  wire n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464;
  wire n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1472, n_1474;
  wire n_1475, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484;
  wire n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492;
  wire n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500;
  wire n_1501, n_1502, n_1503, n_1504, n_1506, n_1507, n_1510, n_1511;
  wire n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519;
  wire n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527;
  wire n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535;
  wire n_1536, n_1538, n_1539, n_1542, n_1543, n_1544, n_1545, n_1546;
  wire n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554;
  wire n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562;
  wire n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1570, n_1571;
  wire n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581;
  wire n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589;
  wire n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597;
  wire n_1598, n_1600, n_1602, n_1603, n_1606, n_1607, n_1608, n_1609;
  wire n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617;
  wire n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625;
  wire n_1626, n_1627, n_1628, n_1629, n_1630, n_1632, n_1634, n_1635;
  wire n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645;
  wire n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653;
  wire n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661;
  wire n_1662, n_1664, n_1666, n_1667, n_1670, n_1671, n_1672, n_1673;
  wire n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681;
  wire n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689;
  wire n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1698;
  wire n_1699, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708;
  wire n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716;
  wire n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724;
  wire n_1725, n_1726, n_1727, n_1728, n_1730, n_1731, n_1734, n_1735;
  wire n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743;
  wire n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751;
  wire n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1760, n_1762;
  wire n_1763, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772;
  wire n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780;
  wire n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788;
  wire n_1789, n_1792, n_1794, n_1795, n_1798, n_1799, n_1800, n_1801;
  wire n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809;
  wire n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817;
  wire n_1818, n_1819, n_1820, n_1821, n_1824, n_1826, n_1827, n_1830;
  wire n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838;
  wire n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846;
  wire n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1856;
  wire n_1858, n_1859, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867;
  wire n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875;
  wire n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883;
  wire n_1884, n_1885, n_1888, n_1890, n_1891, n_1894, n_1895, n_1896;
  wire n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904;
  wire n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912;
  wire n_1913, n_1914, n_1915, n_1916, n_1917, n_1920, n_1922, n_1923;
  wire n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933;
  wire n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941;
  wire n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949;
  wire n_1952, n_1954, n_1955, n_1958, n_1959, n_1960, n_1961, n_1962;
  wire n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970;
  wire n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978;
  wire n_1979, n_1980, n_1981, n_1984, n_1986, n_1987, n_1990, n_1991;
  wire n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999;
  wire n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007;
  wire n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2016, n_2018;
  wire n_2019, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028;
  wire n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036;
  wire n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044;
  wire n_2045, n_2048, n_2050, n_2051, n_2054, n_2055, n_2056, n_2057;
  wire n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065;
  wire n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073;
  wire n_2074, n_2075, n_2076, n_2077, n_2080, n_2082, n_2083, n_2086;
  wire n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094;
  wire n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102;
  wire n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2112;
  wire n_2114, n_2115, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123;
  wire n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131;
  wire n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139;
  wire n_2140, n_2141, n_2144, n_2146, n_2147, n_2150, n_2151, n_2152;
  wire n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160;
  wire n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168;
  wire n_2169, n_2170, n_2171, n_2172, n_2173, n_2176, n_2178, n_2179;
  wire n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189;
  wire n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197;
  wire n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205;
  wire n_2208, n_2210, n_2211, n_2214, n_2215, n_2216, n_2217, n_2218;
  wire n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226;
  wire n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234;
  wire n_2235, n_2236, n_2237, n_2240, n_2242, n_2243, n_2246, n_2247;
  wire n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255;
  wire n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263;
  wire n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2272, n_2274;
  wire n_2275, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284;
  wire n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292;
  wire n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300;
  wire n_2301, n_2304, n_2306, n_2307, n_2310, n_2311, n_2312, n_2313;
  wire n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321;
  wire n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329;
  wire n_2330, n_2331, n_2332, n_2333, n_2336, n_2338, n_2339, n_2342;
  wire n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350;
  wire n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358;
  wire n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2368;
  wire n_2370, n_2371, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379;
  wire n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387;
  wire n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395;
  wire n_2396, n_2397, n_2400, n_2402, n_2403, n_2406, n_2407, n_2408;
  wire n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416;
  wire n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424;
  wire n_2425, n_2426, n_2427, n_2428, n_2429, n_2432, n_2434, n_2435;
  wire n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445;
  wire n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453;
  wire n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461;
  wire n_2462, n_2463, n_2464, n_2466, n_2470, n_2471, n_2472, n_2473;
  wire n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481;
  wire n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489;
  wire n_2490, n_2491, n_2493, n_2494, n_2495, n_2496, n_2497, n_2501;
  wire n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509;
  wire n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517;
  wire n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525;
  wire n_2528, n_2530, n_2531, n_2533, n_2534, n_2535, n_2536, n_2537;
  wire n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545;
  wire n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553;
  wire n_2554, n_2555, n_2558, n_2562, n_2563, n_2564, n_2565, n_2566;
  wire n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574;
  wire n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2586;
  wire n_2589, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598;
  wire n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606;
  wire n_2607, n_2608, n_2609, n_2610, n_2614, n_2617, n_2618, n_2620;
  wire n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628;
  wire n_2629, n_2630, n_2631, n_2632, n_2633, n_2642, n_2644, n_2645;
  wire n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653;
  wire n_2654, n_2655, n_2656, n_2657, n_2664, n_2665, n_2666, n_2667;
  wire n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675;
  wire n_2676, n_2677, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691;
  wire n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2704, n_2705;
  wire n_2706, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713, n_2720;
  wire n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728;
  wire n_2729, n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2746;
  wire n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2756;
  wire n_2757, n_2758, n_2759, n_2760, n_2761, n_2766, n_2767, n_2768;
  wire n_2769, n_2771, n_2772, n_2773, n_2776, n_2777, n_2788, n_2789;
  wire n_2791, n_2793, n_2794, n_2795, n_2796, n_2797, n_2799, n_2800;
  wire n_2801, n_2802, n_2803, n_2805, n_2806, n_2807, n_2808, n_2809;
  wire n_2811, n_2812, n_2813, n_2814, n_2815, n_2817, n_2818, n_2819;
  wire n_2820, n_2821, n_2823, n_2824, n_2825, n_2826, n_2827, n_2829;
  wire n_2830, n_2831, n_2832, n_2833, n_2835, n_2836, n_2837, n_2838;
  wire n_2839, n_2841, n_2842, n_2843, n_2844, n_2845, n_2847, n_2848;
  wire n_2849, n_2850, n_2851, n_2853, n_2854, n_2855, n_2856, n_2857;
  wire n_2859, n_2860, n_2861, n_2862, n_2863, n_2865, n_2866, n_2867;
  wire n_2868, n_2869, n_2871, n_2872, n_2873, n_2874, n_2875, n_2877;
  wire n_2878, n_2879, n_2880, n_2881, n_2883, n_2884, n_2885, n_2886;
  wire n_2887, n_2889, n_2890, n_2891, n_2892, n_2893, n_2895, n_2896;
  wire n_2897, n_2898, n_2899, n_2901, n_2902, n_2903, n_2904, n_2905;
  wire n_2907, n_2908, n_2909, n_2910, n_2911, n_2913, n_2914, n_2915;
  wire n_2916, n_2917, n_2919, n_2920, n_2921, n_2922, n_2923, n_2925;
  wire n_2926, n_2927, n_2928, n_2929, n_2931, n_2932, n_2933, n_2934;
  wire n_2935, n_2937, n_2938, n_2939, n_2940, n_2941, n_2943, n_2944;
  wire n_2945, n_2946, n_2947, n_2949, n_2950, n_2951, n_2952, n_2953;
  wire n_2955, n_2956, n_2957, n_2958, n_2959, n_2961, n_2962, n_2963;
  wire n_2964, n_2965, n_2967, n_2968, n_2969, n_2970, n_2971, n_2973;
  wire n_2974, n_2975, n_2976, n_2977, n_2979, n_2980, n_2981, n_2982;
  wire n_2983, n_2985, n_2986, n_2987, n_2988, n_2989, n_2991, n_2992;
  wire n_2993, n_2994, n_2995, n_2997, n_2998, n_2999, n_3000, n_3001;
  wire n_3003, n_3004, n_3007, n_3010, n_3012, n_3013, n_3015, n_3016;
  wire n_3018, n_3019, n_3020, n_3022, n_3023, n_3025, n_3026, n_3027;
  wire n_3029, n_3030, n_3032, n_3033, n_3034, n_3036, n_3037, n_3039;
  wire n_3040, n_3041, n_3043, n_3044, n_3046, n_3047, n_3048, n_3050;
  wire n_3051, n_3053, n_3054, n_3055, n_3057, n_3058, n_3060, n_3061;
  wire n_3062, n_3064, n_3065, n_3067, n_3068, n_3069, n_3071, n_3072;
  wire n_3074, n_3075, n_3076, n_3078, n_3079, n_3081, n_3082, n_3083;
  wire n_3085, n_3086, n_3088, n_3089, n_3090, n_3092, n_3093, n_3095;
  wire n_3096, n_3097, n_3099, n_3100, n_3102, n_3103, n_3104, n_3106;
  wire n_3107, n_3109, n_3110, n_3111, n_3113, n_3114, n_3116, n_3117;
  wire n_3118, n_3120, n_3121, n_3123, n_3124, n_3125, n_3127, n_3128;
  wire n_3130, n_3131, n_3132, n_3133, n_3136, n_3137, n_3138, n_3139;
  wire n_3140, n_3141, n_3143, n_3144, n_3145, n_3146, n_3147, n_3149;
  wire n_3150, n_3151, n_3152, n_3153, n_3155, n_3156, n_3157, n_3158;
  wire n_3159, n_3161, n_3162, n_3163, n_3164, n_3165, n_3167, n_3168;
  wire n_3169, n_3170, n_3171, n_3173, n_3174, n_3175, n_3176, n_3177;
  wire n_3179, n_3180, n_3181, n_3182, n_3183, n_3185, n_3186, n_3187;
  wire n_3188, n_3189, n_3190, n_3191, n_3193, n_3194, n_3196, n_3197;
  wire n_3198, n_3200, n_3201, n_3203, n_3204, n_3205, n_3207, n_3208;
  wire n_3210, n_3211, n_3212, n_3214, n_3215, n_3216, n_3217, n_3218;
  wire n_3219, n_3221, n_3222, n_3223, n_3224, n_3225, n_3227, n_3228;
  wire n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, n_3237;
  wire n_3239, n_3240, n_3242, n_3244, n_3245, n_3247, n_3249, n_3250;
  wire n_3252, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260;
  wire n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268;
  wire n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, n_3276;
  wire n_3277, n_3278, n_3279, n_3280, n_3281, n_3285, n_3286, n_3288;
  wire n_3290, n_3291, n_3293, n_3295, n_3296, n_3298, n_3300, n_3301;
  wire n_3303, n_3305, n_3306, n_3308, n_3310, n_3311, n_3313, n_3315;
  wire n_3316, n_3318, n_3320, n_3321, n_3323, n_3325, n_3326, n_3328;
  wire n_3330, n_3331, n_3333, n_3335, n_3336, n_3338, n_3340, n_3341;
  wire n_3343, n_3345, n_3346, n_3348, n_3350, n_3351, n_3353, n_3355;
  wire n_3356, n_3358, n_3360, n_3361, n_3363, n_3365, n_3366, n_3368;
  wire n_3370, n_3371, n_3373, n_3375, n_3378, n_3379, n_3381, n_3382;
  wire n_3383, n_3385, n_3386, n_3387, n_3389, n_3390, n_3391, n_3393;
  wire n_3394, n_3395, n_3397, n_3398, n_3399, n_3401, n_3402, n_3403;
  wire n_3405, n_3406, n_3407, n_3409, n_3410, n_3411, n_3413, n_3414;
  wire n_3415, n_3417, n_3418, n_3419, n_3421, n_3422, n_3423, n_3425;
  wire n_3426, n_3427, n_3429, n_3430, n_3431, n_3433, n_3434, n_3435;
  wire n_3437, n_3438, n_3439, n_3441, n_3442, n_3443, n_3445, n_3446;
  wire n_3447, n_3449, n_3450, n_3451, n_3453, n_3454, n_3455, n_3457;
  wire n_3458, n_3459, n_3461, n_3462, n_3463, n_3465, n_3466, n_3467;
  wire n_3469, n_3470, n_3471, n_3473, n_3474, n_3475, n_3477, n_3478;
  wire n_3479, n_3481, n_3482, n_3483, n_3485, n_3486, n_3487, n_3489;
  wire n_3490, n_3491, n_3493, n_3494, n_3495, n_3497, n_3498, n_3499;
  wire n_3501, n_3502, n_3503, n_3505, n_3506, n_3507, n_3509, n_3510;
  wire n_3511, n_3513, n_3514, n_3515, n_3517, n_3518, n_3519, n_3521;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g452 (n_205, A[0], A[4]);
  and g2 (n_128, A[0], A[4]);
  xor g453 (n_1050, A[1], A[3]);
  xor g454 (n_204, n_1050, A[5]);
  nand g3 (n_1051, A[1], A[3]);
  nand g455 (n_1052, A[5], A[3]);
  nand g456 (n_1053, A[1], A[5]);
  nand g457 (n_127, n_1051, n_1052, n_1053);
  xor g458 (n_287, A[0], A[6]);
  and g459 (n_288, A[0], A[6]);
  xor g460 (n_1054, A[4], A[2]);
  xor g461 (n_203, n_1054, n_287);
  nand g462 (n_1055, A[4], A[2]);
  nand g4 (n_1056, n_287, A[2]);
  nand g5 (n_1057, A[4], n_287);
  nand g463 (n_126, n_1055, n_1056, n_1057);
  xor g464 (n_1058, A[1], A[7]);
  xor g465 (n_289, n_1058, A[5]);
  nand g466 (n_1059, A[1], A[7]);
  nand g467 (n_1060, A[5], A[7]);
  nand g6 (n_291, n_1059, n_1060, n_1053);
  xor g469 (n_1062, A[3], n_288);
  xor g470 (n_202, n_1062, n_289);
  nand g471 (n_1063, A[3], n_288);
  nand g472 (n_1064, n_289, n_288);
  nand g473 (n_1065, A[3], n_289);
  nand g474 (n_125, n_1063, n_1064, n_1065);
  xor g475 (n_290, A[0], A[8]);
  and g476 (n_293, A[0], A[8]);
  xor g477 (n_1066, A[2], A[6]);
  xor g478 (n_292, n_1066, A[4]);
  nand g479 (n_1067, A[2], A[6]);
  nand g480 (n_1068, A[4], A[6]);
  nand g482 (n_294, n_1067, n_1068, n_1055);
  xor g483 (n_1070, n_290, n_291);
  xor g484 (n_201, n_1070, n_292);
  nand g485 (n_1071, n_290, n_291);
  nand g486 (n_1072, n_292, n_291);
  nand g487 (n_1073, n_290, n_292);
  nand g488 (n_124, n_1071, n_1072, n_1073);
  xor g489 (n_1074, A[1], A[9]);
  xor g490 (n_295, n_1074, A[3]);
  nand g491 (n_1075, A[1], A[9]);
  nand g492 (n_1076, A[3], A[9]);
  nand g494 (n_298, n_1075, n_1076, n_1051);
  xor g495 (n_1078, A[7], A[5]);
  xor g496 (n_296, n_1078, n_293);
  nand g498 (n_1080, n_293, A[5]);
  nand g499 (n_1081, A[7], n_293);
  nand g500 (n_300, n_1060, n_1080, n_1081);
  xor g501 (n_1082, n_294, n_295);
  xor g502 (n_200, n_1082, n_296);
  nand g503 (n_1083, n_294, n_295);
  nand g504 (n_1084, n_296, n_295);
  nand g505 (n_1085, n_294, n_296);
  nand g506 (n_123, n_1083, n_1084, n_1085);
  xor g510 (n_299, n_1054, A[10]);
  nand g512 (n_1088, A[10], A[2]);
  nand g513 (n_1089, A[4], A[10]);
  nand g514 (n_303, n_1055, n_1088, n_1089);
  xor g515 (n_1090, A[6], n_290);
  xor g516 (n_301, n_1090, n_298);
  nand g517 (n_1091, A[6], n_290);
  nand g518 (n_1092, n_298, n_290);
  nand g519 (n_1093, A[6], n_298);
  nand g520 (n_306, n_1091, n_1092, n_1093);
  xor g521 (n_1094, n_299, n_300);
  xor g522 (n_199, n_1094, n_301);
  nand g523 (n_1095, n_299, n_300);
  nand g524 (n_1096, n_301, n_300);
  nand g525 (n_1097, n_299, n_301);
  nand g526 (n_122, n_1095, n_1096, n_1097);
  xor g528 (n_304, n_1074, A[5]);
  nand g530 (n_1100, A[5], A[9]);
  nand g532 (n_309, n_1075, n_1100, n_1053);
  xor g533 (n_1102, A[3], A[11]);
  xor g534 (n_305, n_1102, A[7]);
  nand g535 (n_1103, A[3], A[11]);
  nand g536 (n_1104, A[7], A[11]);
  nand g537 (n_1105, A[3], A[7]);
  nand g538 (n_310, n_1103, n_1104, n_1105);
  xor g539 (n_1106, n_293, n_303);
  xor g540 (n_307, n_1106, n_304);
  nand g541 (n_1107, n_293, n_303);
  nand g542 (n_1108, n_304, n_303);
  nand g543 (n_1109, n_293, n_304);
  nand g544 (n_314, n_1107, n_1108, n_1109);
  xor g545 (n_1110, n_305, n_306);
  xor g546 (n_198, n_1110, n_307);
  nand g547 (n_1111, n_305, n_306);
  nand g548 (n_1112, n_307, n_306);
  nand g549 (n_1113, n_305, n_307);
  nand g550 (n_121, n_1111, n_1112, n_1113);
  xor g551 (n_308, A[0], A[10]);
  and g552 (n_315, A[0], A[10]);
  xor g553 (n_1114, A[6], A[4]);
  xor g554 (n_133, n_1114, A[12]);
  nand g556 (n_1116, A[12], A[4]);
  nand g557 (n_1117, A[6], A[12]);
  nand g558 (n_316, n_1068, n_1116, n_1117);
  xor g559 (n_1118, A[2], A[8]);
  xor g560 (n_312, n_1118, n_308);
  nand g561 (n_1119, A[2], A[8]);
  nand g562 (n_1120, n_308, A[8]);
  nand g563 (n_1121, A[2], n_308);
  nand g564 (n_319, n_1119, n_1120, n_1121);
  xor g565 (n_1122, n_309, n_310);
  xor g566 (n_313, n_1122, n_133);
  nand g567 (n_1123, n_309, n_310);
  nand g568 (n_1124, n_133, n_310);
  nand g569 (n_1125, n_309, n_133);
  nand g570 (n_321, n_1123, n_1124, n_1125);
  xor g571 (n_1126, n_312, n_313);
  xor g572 (n_197, n_1126, n_314);
  nand g573 (n_1127, n_312, n_313);
  nand g574 (n_1128, n_314, n_313);
  nand g575 (n_1129, n_312, n_314);
  nand g576 (n_120, n_1127, n_1128, n_1129);
  xor g577 (n_1130, A[1], A[11]);
  xor g578 (n_318, n_1130, A[7]);
  nand g579 (n_1131, A[1], A[11]);
  nand g582 (n_324, n_1131, n_1104, n_1059);
  xor g583 (n_1134, A[5], A[13]);
  xor g584 (n_317, n_1134, A[3]);
  nand g585 (n_1135, A[5], A[13]);
  nand g586 (n_1136, A[3], A[13]);
  nand g588 (n_325, n_1135, n_1136, n_1052);
  xor g589 (n_1138, A[9], n_315);
  xor g590 (n_320, n_1138, n_316);
  nand g591 (n_1139, A[9], n_315);
  nand g592 (n_1140, n_316, n_315);
  nand g593 (n_1141, A[9], n_316);
  nand g594 (n_328, n_1139, n_1140, n_1141);
  xor g595 (n_1142, n_317, n_318);
  xor g596 (n_322, n_1142, n_319);
  nand g597 (n_1143, n_317, n_318);
  nand g598 (n_1144, n_319, n_318);
  nand g599 (n_1145, n_317, n_319);
  nand g600 (n_330, n_1143, n_1144, n_1145);
  xor g601 (n_1146, n_320, n_321);
  xor g602 (n_196, n_1146, n_322);
  nand g603 (n_1147, n_320, n_321);
  nand g604 (n_1148, n_322, n_321);
  nand g605 (n_1149, n_320, n_322);
  nand g606 (n_119, n_1147, n_1148, n_1149);
  xor g607 (n_323, A[0], A[14]);
  and g608 (n_332, A[0], A[14]);
  xor g609 (n_1150, A[12], A[8]);
  xor g610 (n_327, n_1150, A[6]);
  nand g611 (n_1151, A[12], A[8]);
  nand g612 (n_1152, A[6], A[8]);
  nand g614 (n_333, n_1151, n_1152, n_1117);
  xor g615 (n_1154, A[10], A[4]);
  xor g616 (n_326, n_1154, A[2]);
  xor g621 (n_1158, n_323, n_324);
  xor g622 (n_329, n_1158, n_325);
  nand g623 (n_1159, n_323, n_324);
  nand g624 (n_1160, n_325, n_324);
  nand g625 (n_1161, n_323, n_325);
  nand g626 (n_338, n_1159, n_1160, n_1161);
  xor g627 (n_1162, n_326, n_327);
  xor g628 (n_331, n_1162, n_328);
  nand g629 (n_1163, n_326, n_327);
  nand g630 (n_1164, n_328, n_327);
  nand g631 (n_1165, n_326, n_328);
  nand g632 (n_341, n_1163, n_1164, n_1165);
  xor g633 (n_1166, n_329, n_330);
  xor g634 (n_195, n_1166, n_331);
  nand g635 (n_1167, n_329, n_330);
  nand g636 (n_1168, n_331, n_330);
  nand g637 (n_1169, n_329, n_331);
  nand g638 (n_118, n_1167, n_1168, n_1169);
  xor g639 (n_1170, A[1], A[15]);
  xor g640 (n_335, n_1170, A[13]);
  nand g641 (n_1171, A[1], A[15]);
  nand g642 (n_1172, A[13], A[15]);
  nand g643 (n_1173, A[1], A[13]);
  nand g644 (n_343, n_1171, n_1172, n_1173);
  xor g645 (n_1174, A[9], A[7]);
  xor g646 (n_336, n_1174, A[11]);
  nand g647 (n_1175, A[9], A[7]);
  nand g649 (n_1177, A[9], A[11]);
  nand g650 (n_344, n_1175, n_1104, n_1177);
  xor g651 (n_1178, A[5], A[3]);
  xor g652 (n_337, n_1178, n_332);
  nand g654 (n_1180, n_332, A[3]);
  nand g655 (n_1181, A[5], n_332);
  nand g656 (n_347, n_1052, n_1180, n_1181);
  xor g657 (n_1182, n_333, n_303);
  xor g658 (n_339, n_1182, n_335);
  nand g659 (n_1183, n_333, n_303);
  nand g660 (n_1184, n_335, n_303);
  nand g661 (n_1185, n_333, n_335);
  nand g662 (n_349, n_1183, n_1184, n_1185);
  xor g663 (n_1186, n_336, n_337);
  xor g664 (n_340, n_1186, n_338);
  nand g665 (n_1187, n_336, n_337);
  nand g666 (n_1188, n_338, n_337);
  nand g667 (n_1189, n_336, n_338);
  nand g668 (n_351, n_1187, n_1188, n_1189);
  xor g669 (n_1190, n_339, n_340);
  xor g670 (n_194, n_1190, n_341);
  nand g671 (n_1191, n_339, n_340);
  nand g672 (n_1192, n_341, n_340);
  nand g673 (n_1193, n_339, n_341);
  nand g674 (n_117, n_1191, n_1192, n_1193);
  xor g675 (n_342, A[0], A[16]);
  and g676 (n_353, A[0], A[16]);
  xor g677 (n_1194, A[14], A[2]);
  xor g678 (n_346, n_1194, A[10]);
  nand g679 (n_1195, A[14], A[2]);
  nand g681 (n_1197, A[14], A[10]);
  nand g682 (n_354, n_1195, n_1088, n_1197);
  xor g689 (n_1202, A[4], n_342);
  xor g690 (n_348, n_1202, n_343);
  nand g691 (n_1203, A[4], n_342);
  nand g692 (n_1204, n_343, n_342);
  nand g693 (n_1205, A[4], n_343);
  nand g694 (n_359, n_1203, n_1204, n_1205);
  xor g695 (n_1206, n_344, n_327);
  xor g696 (n_350, n_1206, n_346);
  nand g697 (n_1207, n_344, n_327);
  nand g698 (n_1208, n_346, n_327);
  nand g699 (n_1209, n_344, n_346);
  nand g700 (n_361, n_1207, n_1208, n_1209);
  xor g701 (n_1210, n_347, n_348);
  xor g702 (n_352, n_1210, n_349);
  nand g703 (n_1211, n_347, n_348);
  nand g704 (n_1212, n_349, n_348);
  nand g705 (n_1213, n_347, n_349);
  nand g706 (n_363, n_1211, n_1212, n_1213);
  xor g707 (n_1214, n_350, n_351);
  xor g708 (n_193, n_1214, n_352);
  nand g709 (n_1215, n_350, n_351);
  nand g710 (n_1216, n_352, n_351);
  nand g711 (n_1217, n_350, n_352);
  nand g712 (n_116, n_1215, n_1216, n_1217);
  xor g713 (n_1218, A[1], A[17]);
  xor g714 (n_357, n_1218, A[15]);
  nand g715 (n_1219, A[1], A[17]);
  nand g716 (n_1220, A[15], A[17]);
  nand g718 (n_366, n_1219, n_1220, n_1171);
  xor g720 (n_358, n_1102, A[9]);
  nand g724 (n_368, n_1103, n_1177, n_1076);
  xor g725 (n_1226, A[13], A[7]);
  xor g726 (n_356, n_1226, A[5]);
  nand g727 (n_1227, A[13], A[7]);
  nand g730 (n_367, n_1227, n_1060, n_1135);
  xor g731 (n_1230, n_353, n_354);
  xor g732 (n_360, n_1230, n_333);
  nand g733 (n_1231, n_353, n_354);
  nand g734 (n_1232, n_333, n_354);
  nand g735 (n_1233, n_353, n_333);
  nand g736 (n_372, n_1231, n_1232, n_1233);
  xor g737 (n_1234, n_356, n_357);
  xor g738 (n_362, n_1234, n_358);
  nand g739 (n_1235, n_356, n_357);
  nand g740 (n_1236, n_358, n_357);
  nand g741 (n_1237, n_356, n_358);
  nand g742 (n_374, n_1235, n_1236, n_1237);
  xor g743 (n_1238, n_359, n_360);
  xor g744 (n_364, n_1238, n_361);
  nand g745 (n_1239, n_359, n_360);
  nand g746 (n_1240, n_361, n_360);
  nand g747 (n_1241, n_359, n_361);
  nand g748 (n_376, n_1239, n_1240, n_1241);
  xor g749 (n_1242, n_362, n_363);
  xor g750 (n_192, n_1242, n_364);
  nand g751 (n_1243, n_362, n_363);
  nand g752 (n_1244, n_364, n_363);
  nand g753 (n_1245, n_362, n_364);
  nand g754 (n_115, n_1243, n_1244, n_1245);
  xor g755 (n_365, A[0], A[18]);
  and g756 (n_378, A[0], A[18]);
  xor g757 (n_1246, A[12], A[4]);
  xor g758 (n_369, n_1246, A[2]);
  nand g761 (n_1249, A[12], A[2]);
  nand g762 (n_379, n_1116, n_1055, n_1249);
  xor g763 (n_1250, A[16], A[10]);
  xor g764 (n_370, n_1250, A[14]);
  nand g765 (n_1251, A[16], A[10]);
  nand g767 (n_1253, A[16], A[14]);
  nand g768 (n_380, n_1251, n_1197, n_1253);
  xor g769 (n_1254, A[8], A[6]);
  xor g770 (n_371, n_1254, n_365);
  nand g772 (n_1256, n_365, A[6]);
  nand g773 (n_1257, A[8], n_365);
  nand g774 (n_384, n_1152, n_1256, n_1257);
  xor g775 (n_1258, n_366, n_367);
  xor g776 (n_373, n_1258, n_368);
  nand g777 (n_1259, n_366, n_367);
  nand g778 (n_1260, n_368, n_367);
  nand g779 (n_1261, n_366, n_368);
  nand g780 (n_386, n_1259, n_1260, n_1261);
  xor g781 (n_1262, n_369, n_370);
  xor g782 (n_375, n_1262, n_371);
  nand g783 (n_1263, n_369, n_370);
  nand g784 (n_1264, n_371, n_370);
  nand g785 (n_1265, n_369, n_371);
  nand g786 (n_387, n_1263, n_1264, n_1265);
  xor g787 (n_1266, n_372, n_373);
  xor g788 (n_377, n_1266, n_374);
  nand g789 (n_1267, n_372, n_373);
  nand g790 (n_1268, n_374, n_373);
  nand g791 (n_1269, n_372, n_374);
  nand g792 (n_390, n_1267, n_1268, n_1269);
  xor g793 (n_1270, n_375, n_376);
  xor g794 (n_191, n_1270, n_377);
  nand g795 (n_1271, n_375, n_376);
  nand g796 (n_1272, n_377, n_376);
  nand g797 (n_1273, n_375, n_377);
  nand g798 (n_114, n_1271, n_1272, n_1273);
  xor g799 (n_1274, A[1], A[19]);
  xor g800 (n_382, n_1274, A[13]);
  nand g801 (n_1275, A[1], A[19]);
  nand g802 (n_1276, A[13], A[19]);
  nand g804 (n_392, n_1275, n_1276, n_1173);
  xor g806 (n_383, n_1178, A[17]);
  nand g808 (n_1280, A[17], A[3]);
  nand g809 (n_1281, A[5], A[17]);
  nand g810 (n_129, n_1052, n_1280, n_1281);
  xor g811 (n_1282, A[11], A[15]);
  xor g812 (n_381, n_1282, A[9]);
  nand g813 (n_1283, A[11], A[15]);
  nand g814 (n_1284, A[9], A[15]);
  nand g816 (n_130, n_1283, n_1284, n_1177);
  xor g817 (n_1286, A[7], n_378);
  xor g818 (n_385, n_1286, n_379);
  nand g819 (n_1287, A[7], n_378);
  nand g820 (n_1288, n_379, n_378);
  nand g821 (n_1289, A[7], n_379);
  nand g822 (n_393, n_1287, n_1288, n_1289);
  xor g823 (n_1290, n_380, n_381);
  xor g824 (n_388, n_1290, n_382);
  nand g825 (n_1291, n_380, n_381);
  nand g826 (n_1292, n_382, n_381);
  nand g827 (n_1293, n_380, n_382);
  nand g828 (n_395, n_1291, n_1292, n_1293);
  xor g829 (n_1294, n_383, n_384);
  xor g830 (n_389, n_1294, n_385);
  nand g831 (n_1295, n_383, n_384);
  nand g832 (n_1296, n_385, n_384);
  nand g833 (n_1297, n_383, n_385);
  nand g834 (n_397, n_1295, n_1296, n_1297);
  xor g835 (n_1298, n_386, n_387);
  xor g836 (n_391, n_1298, n_388);
  nand g837 (n_1299, n_386, n_387);
  nand g838 (n_1300, n_388, n_387);
  nand g839 (n_1301, n_386, n_388);
  nand g840 (n_399, n_1299, n_1300, n_1301);
  xor g841 (n_1302, n_389, n_390);
  xor g842 (n_190, n_1302, n_391);
  nand g843 (n_1303, n_389, n_390);
  nand g844 (n_1304, n_391, n_390);
  nand g845 (n_1305, n_389, n_391);
  nand g846 (n_113, n_1303, n_1304, n_1305);
  xor g847 (n_1306, A[20], A[18]);
  xor g848 (n_132, n_1306, A[14]);
  nand g849 (n_1307, A[20], A[18]);
  nand g850 (n_1308, A[14], A[18]);
  nand g851 (n_1309, A[20], A[14]);
  nand g852 (n_401, n_1307, n_1308, n_1309);
  xor g859 (n_1314, A[2], A[16]);
  xor g860 (n_131, n_1314, A[10]);
  nand g861 (n_1315, A[2], A[16]);
  nand g864 (n_403, n_1315, n_1251, n_1088);
  xor g865 (n_1318, A[8], n_392);
  xor g866 (n_394, n_1318, n_129);
  nand g867 (n_1319, A[8], n_392);
  nand g868 (n_1320, n_129, n_392);
  nand g869 (n_1321, A[8], n_129);
  nand g870 (n_407, n_1319, n_1320, n_1321);
  xor g871 (n_1322, n_130, n_131);
  xor g872 (n_396, n_1322, n_132);
  nand g873 (n_1323, n_130, n_131);
  nand g874 (n_1324, n_132, n_131);
  nand g875 (n_1325, n_130, n_132);
  nand g876 (n_409, n_1323, n_1324, n_1325);
  xor g877 (n_1326, n_133, n_393);
  xor g878 (n_398, n_1326, n_394);
  nand g879 (n_1327, n_133, n_393);
  nand g880 (n_1328, n_394, n_393);
  nand g881 (n_1329, n_133, n_394);
  nand g882 (n_411, n_1327, n_1328, n_1329);
  xor g883 (n_1330, n_395, n_396);
  xor g884 (n_400, n_1330, n_397);
  nand g885 (n_1331, n_395, n_396);
  nand g886 (n_1332, n_397, n_396);
  nand g887 (n_1333, n_395, n_397);
  nand g888 (n_413, n_1331, n_1332, n_1333);
  xor g889 (n_1334, n_398, n_399);
  xor g890 (n_189, n_1334, n_400);
  nand g891 (n_1335, n_398, n_399);
  nand g892 (n_1336, n_400, n_399);
  nand g893 (n_1337, n_398, n_400);
  nand g894 (n_112, n_1335, n_1336, n_1337);
  xor g895 (n_1338, A[21], A[19]);
  xor g896 (n_405, n_1338, A[15]);
  nand g897 (n_1339, A[21], A[19]);
  nand g898 (n_1340, A[15], A[19]);
  nand g899 (n_1341, A[21], A[15]);
  nand g900 (n_415, n_1339, n_1340, n_1341);
  xor g902 (n_406, n_1078, A[13]);
  xor g907 (n_1346, A[3], A[17]);
  xor g908 (n_404, n_1346, A[11]);
  nand g910 (n_1348, A[11], A[17]);
  nand g912 (n_417, n_1280, n_1348, n_1103);
  xor g913 (n_1350, A[9], n_401);
  xor g914 (n_408, n_1350, n_316);
  nand g915 (n_1351, A[9], n_401);
  nand g916 (n_1352, n_316, n_401);
  nand g918 (n_421, n_1351, n_1352, n_1141);
  xor g919 (n_1354, n_403, n_404);
  xor g920 (n_410, n_1354, n_405);
  nand g921 (n_1355, n_403, n_404);
  nand g922 (n_1356, n_405, n_404);
  nand g923 (n_1357, n_403, n_405);
  nand g924 (n_423, n_1355, n_1356, n_1357);
  xor g925 (n_1358, n_406, n_407);
  xor g926 (n_412, n_1358, n_408);
  nand g927 (n_1359, n_406, n_407);
  nand g928 (n_1360, n_408, n_407);
  nand g929 (n_1361, n_406, n_408);
  nand g930 (n_425, n_1359, n_1360, n_1361);
  xor g931 (n_1362, n_409, n_410);
  xor g932 (n_414, n_1362, n_411);
  nand g933 (n_1363, n_409, n_410);
  nand g934 (n_1364, n_411, n_410);
  nand g935 (n_1365, n_409, n_411);
  nand g936 (n_428, n_1363, n_1364, n_1365);
  xor g937 (n_1366, n_412, n_413);
  xor g938 (n_188, n_1366, n_414);
  nand g939 (n_1367, n_412, n_413);
  nand g940 (n_1368, n_414, n_413);
  nand g941 (n_1369, n_412, n_414);
  nand g942 (n_111, n_1367, n_1368, n_1369);
  xor g943 (n_1370, A[22], A[20]);
  xor g944 (n_419, n_1370, A[16]);
  nand g945 (n_1371, A[22], A[20]);
  nand g946 (n_1372, A[16], A[20]);
  nand g947 (n_1373, A[22], A[16]);
  nand g948 (n_429, n_1371, n_1372, n_1373);
  xor g950 (n_420, n_1254, A[14]);
  nand g952 (n_1376, A[14], A[6]);
  nand g953 (n_1377, A[8], A[14]);
  nand g954 (n_430, n_1152, n_1376, n_1377);
  xor g955 (n_1378, A[4], A[18]);
  xor g956 (n_418, n_1378, A[12]);
  nand g957 (n_1379, A[4], A[18]);
  nand g958 (n_1380, A[12], A[18]);
  nand g960 (n_431, n_1379, n_1380, n_1116);
  xor g961 (n_1382, A[10], n_415);
  xor g962 (n_422, n_1382, n_367);
  nand g963 (n_1383, A[10], n_415);
  nand g964 (n_1384, n_367, n_415);
  nand g965 (n_1385, A[10], n_367);
  nand g966 (n_435, n_1383, n_1384, n_1385);
  xor g967 (n_1386, n_417, n_418);
  xor g968 (n_424, n_1386, n_419);
  nand g969 (n_1387, n_417, n_418);
  nand g970 (n_1388, n_419, n_418);
  nand g971 (n_1389, n_417, n_419);
  nand g972 (n_437, n_1387, n_1388, n_1389);
  xor g973 (n_1390, n_420, n_421);
  xor g974 (n_426, n_1390, n_422);
  nand g975 (n_1391, n_420, n_421);
  nand g976 (n_1392, n_422, n_421);
  nand g977 (n_1393, n_420, n_422);
  nand g978 (n_439, n_1391, n_1392, n_1393);
  xor g979 (n_1394, n_423, n_424);
  xor g980 (n_427, n_1394, n_425);
  nand g981 (n_1395, n_423, n_424);
  nand g982 (n_1396, n_425, n_424);
  nand g983 (n_1397, n_423, n_425);
  nand g984 (n_442, n_1395, n_1396, n_1397);
  xor g985 (n_1398, n_426, n_427);
  xor g986 (n_187, n_1398, n_428);
  nand g987 (n_1399, n_426, n_427);
  nand g988 (n_1400, n_428, n_427);
  nand g989 (n_1401, n_426, n_428);
  nand g990 (n_110, n_1399, n_1400, n_1401);
  xor g991 (n_1402, A[23], A[21]);
  xor g992 (n_433, n_1402, A[17]);
  nand g993 (n_1403, A[23], A[21]);
  nand g994 (n_1404, A[17], A[21]);
  nand g995 (n_1405, A[23], A[17]);
  nand g996 (n_443, n_1403, n_1404, n_1405);
  xor g998 (n_434, n_1174, A[15]);
  nand g1000 (n_1408, A[15], A[7]);
  nand g1002 (n_444, n_1175, n_1408, n_1284);
  xor g1003 (n_1410, A[5], A[19]);
  xor g1004 (n_432, n_1410, A[13]);
  nand g1005 (n_1411, A[5], A[19]);
  nand g1008 (n_445, n_1411, n_1276, n_1135);
  xor g1009 (n_1414, A[11], n_429);
  xor g1010 (n_436, n_1414, n_430);
  nand g1011 (n_1415, A[11], n_429);
  nand g1012 (n_1416, n_430, n_429);
  nand g1013 (n_1417, A[11], n_430);
  nand g1014 (n_449, n_1415, n_1416, n_1417);
  xor g1015 (n_1418, n_431, n_432);
  xor g1016 (n_438, n_1418, n_433);
  nand g1017 (n_1419, n_431, n_432);
  nand g1018 (n_1420, n_433, n_432);
  nand g1019 (n_1421, n_431, n_433);
  nand g1020 (n_451, n_1419, n_1420, n_1421);
  xor g1021 (n_1422, n_434, n_435);
  xor g1022 (n_440, n_1422, n_436);
  nand g1023 (n_1423, n_434, n_435);
  nand g1024 (n_1424, n_436, n_435);
  nand g1025 (n_1425, n_434, n_436);
  nand g1026 (n_453, n_1423, n_1424, n_1425);
  xor g1027 (n_1426, n_437, n_438);
  xor g1028 (n_441, n_1426, n_439);
  nand g1029 (n_1427, n_437, n_438);
  nand g1030 (n_1428, n_439, n_438);
  nand g1031 (n_1429, n_437, n_439);
  nand g1032 (n_456, n_1427, n_1428, n_1429);
  xor g1033 (n_1430, n_440, n_441);
  xor g1034 (n_186, n_1430, n_442);
  nand g1035 (n_1431, n_440, n_441);
  nand g1036 (n_1432, n_442, n_441);
  nand g1037 (n_1433, n_440, n_442);
  nand g1038 (n_109, n_1431, n_1432, n_1433);
  xor g1039 (n_1434, A[24], A[22]);
  xor g1040 (n_447, n_1434, A[18]);
  nand g1041 (n_1435, A[24], A[22]);
  nand g1042 (n_1436, A[18], A[22]);
  nand g1043 (n_1437, A[24], A[18]);
  nand g1044 (n_457, n_1435, n_1436, n_1437);
  xor g1045 (n_1438, A[10], A[8]);
  xor g1046 (n_448, n_1438, A[16]);
  nand g1047 (n_1439, A[10], A[8]);
  nand g1048 (n_1440, A[16], A[8]);
  nand g1050 (n_458, n_1439, n_1440, n_1251);
  xor g1051 (n_1442, A[6], A[20]);
  xor g1052 (n_446, n_1442, A[14]);
  nand g1053 (n_1443, A[6], A[20]);
  nand g1056 (n_459, n_1443, n_1309, n_1376);
  xor g1057 (n_1446, A[12], n_443);
  xor g1058 (n_450, n_1446, n_444);
  nand g1059 (n_1447, A[12], n_443);
  nand g1060 (n_1448, n_444, n_443);
  nand g1061 (n_1449, A[12], n_444);
  nand g1062 (n_461, n_1447, n_1448, n_1449);
  xor g1063 (n_1450, n_445, n_446);
  xor g1064 (n_452, n_1450, n_447);
  nand g1065 (n_1451, n_445, n_446);
  nand g1066 (n_1452, n_447, n_446);
  nand g1067 (n_1453, n_445, n_447);
  nand g1068 (n_463, n_1451, n_1452, n_1453);
  xor g1069 (n_1454, n_448, n_449);
  xor g1070 (n_454, n_1454, n_450);
  nand g1071 (n_1455, n_448, n_449);
  nand g1072 (n_1456, n_450, n_449);
  nand g1073 (n_1457, n_448, n_450);
  nand g1074 (n_465, n_1455, n_1456, n_1457);
  xor g1075 (n_1458, n_451, n_452);
  xor g1076 (n_455, n_1458, n_453);
  nand g1077 (n_1459, n_451, n_452);
  nand g1078 (n_1460, n_453, n_452);
  nand g1079 (n_1461, n_451, n_453);
  nand g1080 (n_468, n_1459, n_1460, n_1461);
  xor g1081 (n_1462, n_454, n_455);
  xor g1082 (n_185, n_1462, n_456);
  nand g1083 (n_1463, n_454, n_455);
  nand g1084 (n_1464, n_456, n_455);
  nand g1085 (n_1465, n_454, n_456);
  nand g1086 (n_108, n_1463, n_1464, n_1465);
  xor g1087 (n_1466, A[25], A[23]);
  xor g1088 (n_207, n_1466, A[19]);
  nand g1089 (n_1467, A[25], A[23]);
  nand g1090 (n_1468, A[19], A[23]);
  nand g1091 (n_1469, A[25], A[19]);
  nand g1092 (n_469, n_1467, n_1468, n_1469);
  xor g1093 (n_1470, A[11], A[9]);
  xor g1094 (n_460, n_1470, A[17]);
  nand g1096 (n_1472, A[17], A[9]);
  nand g1098 (n_470, n_1177, n_1472, n_1348);
  xor g1099 (n_1474, A[7], A[21]);
  xor g1100 (n_206, n_1474, A[15]);
  nand g1101 (n_1475, A[7], A[21]);
  nand g1104 (n_471, n_1475, n_1341, n_1408);
  xor g1105 (n_1478, A[13], n_457);
  xor g1106 (n_462, n_1478, n_458);
  nand g1107 (n_1479, A[13], n_457);
  nand g1108 (n_1480, n_458, n_457);
  nand g1109 (n_1481, A[13], n_458);
  nand g1110 (n_475, n_1479, n_1480, n_1481);
  xor g1111 (n_1482, n_459, n_206);
  xor g1112 (n_464, n_1482, n_207);
  nand g1113 (n_1483, n_459, n_206);
  nand g1114 (n_1484, n_207, n_206);
  nand g1115 (n_1485, n_459, n_207);
  nand g1116 (n_477, n_1483, n_1484, n_1485);
  xor g1117 (n_1486, n_460, n_461);
  xor g1118 (n_466, n_1486, n_462);
  nand g1119 (n_1487, n_460, n_461);
  nand g1120 (n_1488, n_462, n_461);
  nand g1121 (n_1489, n_460, n_462);
  nand g1122 (n_479, n_1487, n_1488, n_1489);
  xor g1123 (n_1490, n_463, n_464);
  xor g1124 (n_467, n_1490, n_465);
  nand g1125 (n_1491, n_463, n_464);
  nand g1126 (n_1492, n_465, n_464);
  nand g1127 (n_1493, n_463, n_465);
  nand g1128 (n_482, n_1491, n_1492, n_1493);
  xor g1129 (n_1494, n_466, n_467);
  xor g1130 (n_184, n_1494, n_468);
  nand g1131 (n_1495, n_466, n_467);
  nand g1132 (n_1496, n_468, n_467);
  nand g1133 (n_1497, n_466, n_468);
  nand g1134 (n_107, n_1495, n_1496, n_1497);
  xor g1135 (n_1498, A[26], A[24]);
  xor g1136 (n_473, n_1498, A[20]);
  nand g1137 (n_1499, A[26], A[24]);
  nand g1138 (n_1500, A[20], A[24]);
  nand g1139 (n_1501, A[26], A[20]);
  nand g1140 (n_483, n_1499, n_1500, n_1501);
  xor g1141 (n_1502, A[12], A[10]);
  xor g1142 (n_474, n_1502, A[18]);
  nand g1143 (n_1503, A[12], A[10]);
  nand g1144 (n_1504, A[18], A[10]);
  nand g1146 (n_484, n_1503, n_1504, n_1380);
  xor g1147 (n_1506, A[8], A[22]);
  xor g1148 (n_472, n_1506, A[16]);
  nand g1149 (n_1507, A[8], A[22]);
  nand g1152 (n_485, n_1507, n_1373, n_1440);
  xor g1153 (n_1510, A[14], n_469);
  xor g1154 (n_476, n_1510, n_470);
  nand g1155 (n_1511, A[14], n_469);
  nand g1156 (n_1512, n_470, n_469);
  nand g1157 (n_1513, A[14], n_470);
  nand g1158 (n_489, n_1511, n_1512, n_1513);
  xor g1159 (n_1514, n_471, n_472);
  xor g1160 (n_478, n_1514, n_473);
  nand g1161 (n_1515, n_471, n_472);
  nand g1162 (n_1516, n_473, n_472);
  nand g1163 (n_1517, n_471, n_473);
  nand g1164 (n_491, n_1515, n_1516, n_1517);
  xor g1165 (n_1518, n_474, n_475);
  xor g1166 (n_480, n_1518, n_476);
  nand g1167 (n_1519, n_474, n_475);
  nand g1168 (n_1520, n_476, n_475);
  nand g1169 (n_1521, n_474, n_476);
  nand g1170 (n_493, n_1519, n_1520, n_1521);
  xor g1171 (n_1522, n_477, n_478);
  xor g1172 (n_481, n_1522, n_479);
  nand g1173 (n_1523, n_477, n_478);
  nand g1174 (n_1524, n_479, n_478);
  nand g1175 (n_1525, n_477, n_479);
  nand g1176 (n_496, n_1523, n_1524, n_1525);
  xor g1177 (n_1526, n_480, n_481);
  xor g1178 (n_183, n_1526, n_482);
  nand g1179 (n_1527, n_480, n_481);
  nand g1180 (n_1528, n_482, n_481);
  nand g1181 (n_1529, n_480, n_482);
  nand g1182 (n_106, n_1527, n_1528, n_1529);
  xor g1183 (n_1530, A[27], A[25]);
  xor g1184 (n_487, n_1530, A[21]);
  nand g1185 (n_1531, A[27], A[25]);
  nand g1186 (n_1532, A[21], A[25]);
  nand g1187 (n_1533, A[27], A[21]);
  nand g1188 (n_497, n_1531, n_1532, n_1533);
  xor g1189 (n_1534, A[13], A[11]);
  xor g1190 (n_488, n_1534, A[19]);
  nand g1191 (n_1535, A[13], A[11]);
  nand g1192 (n_1536, A[19], A[11]);
  nand g1194 (n_498, n_1535, n_1536, n_1276);
  xor g1195 (n_1538, A[9], A[23]);
  xor g1196 (n_486, n_1538, A[17]);
  nand g1197 (n_1539, A[9], A[23]);
  nand g1200 (n_499, n_1539, n_1405, n_1472);
  xor g1201 (n_1542, A[15], n_483);
  xor g1202 (n_490, n_1542, n_484);
  nand g1203 (n_1543, A[15], n_483);
  nand g1204 (n_1544, n_484, n_483);
  nand g1205 (n_1545, A[15], n_484);
  nand g1206 (n_503, n_1543, n_1544, n_1545);
  xor g1207 (n_1546, n_485, n_486);
  xor g1208 (n_492, n_1546, n_487);
  nand g1209 (n_1547, n_485, n_486);
  nand g1210 (n_1548, n_487, n_486);
  nand g1211 (n_1549, n_485, n_487);
  nand g1212 (n_505, n_1547, n_1548, n_1549);
  xor g1213 (n_1550, n_488, n_489);
  xor g1214 (n_494, n_1550, n_490);
  nand g1215 (n_1551, n_488, n_489);
  nand g1216 (n_1552, n_490, n_489);
  nand g1217 (n_1553, n_488, n_490);
  nand g1218 (n_507, n_1551, n_1552, n_1553);
  xor g1219 (n_1554, n_491, n_492);
  xor g1220 (n_495, n_1554, n_493);
  nand g1221 (n_1555, n_491, n_492);
  nand g1222 (n_1556, n_493, n_492);
  nand g1223 (n_1557, n_491, n_493);
  nand g1224 (n_510, n_1555, n_1556, n_1557);
  xor g1225 (n_1558, n_494, n_495);
  xor g1226 (n_182, n_1558, n_496);
  nand g1227 (n_1559, n_494, n_495);
  nand g1228 (n_1560, n_496, n_495);
  nand g1229 (n_1561, n_494, n_496);
  nand g1230 (n_105, n_1559, n_1560, n_1561);
  xor g1231 (n_1562, A[28], A[26]);
  xor g1232 (n_501, n_1562, A[22]);
  nand g1233 (n_1563, A[28], A[26]);
  nand g1234 (n_1564, A[22], A[26]);
  nand g1235 (n_1565, A[28], A[22]);
  nand g1236 (n_511, n_1563, n_1564, n_1565);
  xor g1237 (n_1566, A[14], A[12]);
  xor g1238 (n_502, n_1566, A[20]);
  nand g1239 (n_1567, A[14], A[12]);
  nand g1240 (n_1568, A[20], A[12]);
  nand g1242 (n_512, n_1567, n_1568, n_1309);
  xor g1243 (n_1570, A[10], A[24]);
  xor g1244 (n_500, n_1570, A[18]);
  nand g1245 (n_1571, A[10], A[24]);
  nand g1248 (n_513, n_1571, n_1437, n_1504);
  xor g1249 (n_1574, A[16], n_497);
  xor g1250 (n_504, n_1574, n_498);
  nand g1251 (n_1575, A[16], n_497);
  nand g1252 (n_1576, n_498, n_497);
  nand g1253 (n_1577, A[16], n_498);
  nand g1254 (n_517, n_1575, n_1576, n_1577);
  xor g1255 (n_1578, n_499, n_500);
  xor g1256 (n_506, n_1578, n_501);
  nand g1257 (n_1579, n_499, n_500);
  nand g1258 (n_1580, n_501, n_500);
  nand g1259 (n_1581, n_499, n_501);
  nand g1260 (n_519, n_1579, n_1580, n_1581);
  xor g1261 (n_1582, n_502, n_503);
  xor g1262 (n_508, n_1582, n_504);
  nand g1263 (n_1583, n_502, n_503);
  nand g1264 (n_1584, n_504, n_503);
  nand g1265 (n_1585, n_502, n_504);
  nand g1266 (n_521, n_1583, n_1584, n_1585);
  xor g1267 (n_1586, n_505, n_506);
  xor g1268 (n_509, n_1586, n_507);
  nand g1269 (n_1587, n_505, n_506);
  nand g1270 (n_1588, n_507, n_506);
  nand g1271 (n_1589, n_505, n_507);
  nand g1272 (n_524, n_1587, n_1588, n_1589);
  xor g1273 (n_1590, n_508, n_509);
  xor g1274 (n_181, n_1590, n_510);
  nand g1275 (n_1591, n_508, n_509);
  nand g1276 (n_1592, n_510, n_509);
  nand g1277 (n_1593, n_508, n_510);
  nand g1278 (n_104, n_1591, n_1592, n_1593);
  xor g1279 (n_1594, A[29], A[27]);
  xor g1280 (n_515, n_1594, A[23]);
  nand g1281 (n_1595, A[29], A[27]);
  nand g1282 (n_1596, A[23], A[27]);
  nand g1283 (n_1597, A[29], A[23]);
  nand g1284 (n_525, n_1595, n_1596, n_1597);
  xor g1285 (n_1598, A[15], A[13]);
  xor g1286 (n_516, n_1598, A[21]);
  nand g1288 (n_1600, A[21], A[13]);
  nand g1290 (n_526, n_1172, n_1600, n_1341);
  xor g1291 (n_1602, A[11], A[25]);
  xor g1292 (n_514, n_1602, A[19]);
  nand g1293 (n_1603, A[11], A[25]);
  nand g1296 (n_527, n_1603, n_1469, n_1536);
  xor g1297 (n_1606, A[17], n_511);
  xor g1298 (n_518, n_1606, n_512);
  nand g1299 (n_1607, A[17], n_511);
  nand g1300 (n_1608, n_512, n_511);
  nand g1301 (n_1609, A[17], n_512);
  nand g1302 (n_531, n_1607, n_1608, n_1609);
  xor g1303 (n_1610, n_513, n_514);
  xor g1304 (n_520, n_1610, n_515);
  nand g1305 (n_1611, n_513, n_514);
  nand g1306 (n_1612, n_515, n_514);
  nand g1307 (n_1613, n_513, n_515);
  nand g1308 (n_533, n_1611, n_1612, n_1613);
  xor g1309 (n_1614, n_516, n_517);
  xor g1310 (n_522, n_1614, n_518);
  nand g1311 (n_1615, n_516, n_517);
  nand g1312 (n_1616, n_518, n_517);
  nand g1313 (n_1617, n_516, n_518);
  nand g1314 (n_535, n_1615, n_1616, n_1617);
  xor g1315 (n_1618, n_519, n_520);
  xor g1316 (n_523, n_1618, n_521);
  nand g1317 (n_1619, n_519, n_520);
  nand g1318 (n_1620, n_521, n_520);
  nand g1319 (n_1621, n_519, n_521);
  nand g1320 (n_538, n_1619, n_1620, n_1621);
  xor g1321 (n_1622, n_522, n_523);
  xor g1322 (n_180, n_1622, n_524);
  nand g1323 (n_1623, n_522, n_523);
  nand g1324 (n_1624, n_524, n_523);
  nand g1325 (n_1625, n_522, n_524);
  nand g1326 (n_103, n_1623, n_1624, n_1625);
  xor g1327 (n_1626, A[30], A[28]);
  xor g1328 (n_529, n_1626, A[24]);
  nand g1329 (n_1627, A[30], A[28]);
  nand g1330 (n_1628, A[24], A[28]);
  nand g1331 (n_1629, A[30], A[24]);
  nand g1332 (n_539, n_1627, n_1628, n_1629);
  xor g1333 (n_1630, A[16], A[14]);
  xor g1334 (n_530, n_1630, A[22]);
  nand g1336 (n_1632, A[22], A[14]);
  nand g1338 (n_540, n_1253, n_1632, n_1373);
  xor g1339 (n_1634, A[12], A[26]);
  xor g1340 (n_528, n_1634, A[20]);
  nand g1341 (n_1635, A[12], A[26]);
  nand g1344 (n_541, n_1635, n_1501, n_1568);
  xor g1345 (n_1638, A[18], n_525);
  xor g1346 (n_532, n_1638, n_526);
  nand g1347 (n_1639, A[18], n_525);
  nand g1348 (n_1640, n_526, n_525);
  nand g1349 (n_1641, A[18], n_526);
  nand g1350 (n_545, n_1639, n_1640, n_1641);
  xor g1351 (n_1642, n_527, n_528);
  xor g1352 (n_534, n_1642, n_529);
  nand g1353 (n_1643, n_527, n_528);
  nand g1354 (n_1644, n_529, n_528);
  nand g1355 (n_1645, n_527, n_529);
  nand g1356 (n_547, n_1643, n_1644, n_1645);
  xor g1357 (n_1646, n_530, n_531);
  xor g1358 (n_536, n_1646, n_532);
  nand g1359 (n_1647, n_530, n_531);
  nand g1360 (n_1648, n_532, n_531);
  nand g1361 (n_1649, n_530, n_532);
  nand g1362 (n_549, n_1647, n_1648, n_1649);
  xor g1363 (n_1650, n_533, n_534);
  xor g1364 (n_537, n_1650, n_535);
  nand g1365 (n_1651, n_533, n_534);
  nand g1366 (n_1652, n_535, n_534);
  nand g1367 (n_1653, n_533, n_535);
  nand g1368 (n_552, n_1651, n_1652, n_1653);
  xor g1369 (n_1654, n_536, n_537);
  xor g1370 (n_179, n_1654, n_538);
  nand g1371 (n_1655, n_536, n_537);
  nand g1372 (n_1656, n_538, n_537);
  nand g1373 (n_1657, n_536, n_538);
  nand g1374 (n_102, n_1655, n_1656, n_1657);
  xor g1375 (n_1658, A[31], A[29]);
  xor g1376 (n_543, n_1658, A[25]);
  nand g1377 (n_1659, A[31], A[29]);
  nand g1378 (n_1660, A[25], A[29]);
  nand g1379 (n_1661, A[31], A[25]);
  nand g1380 (n_553, n_1659, n_1660, n_1661);
  xor g1381 (n_1662, A[17], A[15]);
  xor g1382 (n_544, n_1662, A[23]);
  nand g1384 (n_1664, A[23], A[15]);
  nand g1386 (n_554, n_1220, n_1664, n_1405);
  xor g1387 (n_1666, A[13], A[27]);
  xor g1388 (n_542, n_1666, A[21]);
  nand g1389 (n_1667, A[13], A[27]);
  nand g1392 (n_555, n_1667, n_1533, n_1600);
  xor g1393 (n_1670, A[19], n_539);
  xor g1394 (n_546, n_1670, n_540);
  nand g1395 (n_1671, A[19], n_539);
  nand g1396 (n_1672, n_540, n_539);
  nand g1397 (n_1673, A[19], n_540);
  nand g1398 (n_559, n_1671, n_1672, n_1673);
  xor g1399 (n_1674, n_541, n_542);
  xor g1400 (n_548, n_1674, n_543);
  nand g1401 (n_1675, n_541, n_542);
  nand g1402 (n_1676, n_543, n_542);
  nand g1403 (n_1677, n_541, n_543);
  nand g1404 (n_561, n_1675, n_1676, n_1677);
  xor g1405 (n_1678, n_544, n_545);
  xor g1406 (n_550, n_1678, n_546);
  nand g1407 (n_1679, n_544, n_545);
  nand g1408 (n_1680, n_546, n_545);
  nand g1409 (n_1681, n_544, n_546);
  nand g1410 (n_563, n_1679, n_1680, n_1681);
  xor g1411 (n_1682, n_547, n_548);
  xor g1412 (n_551, n_1682, n_549);
  nand g1413 (n_1683, n_547, n_548);
  nand g1414 (n_1684, n_549, n_548);
  nand g1415 (n_1685, n_547, n_549);
  nand g1416 (n_566, n_1683, n_1684, n_1685);
  xor g1417 (n_1686, n_550, n_551);
  xor g1418 (n_178, n_1686, n_552);
  nand g1419 (n_1687, n_550, n_551);
  nand g1420 (n_1688, n_552, n_551);
  nand g1421 (n_1689, n_550, n_552);
  nand g1422 (n_101, n_1687, n_1688, n_1689);
  xor g1423 (n_1690, A[32], A[30]);
  xor g1424 (n_557, n_1690, A[26]);
  nand g1425 (n_1691, A[32], A[30]);
  nand g1426 (n_1692, A[26], A[30]);
  nand g1427 (n_1693, A[32], A[26]);
  nand g1428 (n_567, n_1691, n_1692, n_1693);
  xor g1429 (n_1694, A[18], A[16]);
  xor g1430 (n_558, n_1694, A[24]);
  nand g1431 (n_1695, A[18], A[16]);
  nand g1432 (n_1696, A[24], A[16]);
  nand g1434 (n_568, n_1695, n_1696, n_1437);
  xor g1435 (n_1698, A[14], A[28]);
  xor g1436 (n_556, n_1698, A[22]);
  nand g1437 (n_1699, A[14], A[28]);
  nand g1440 (n_569, n_1699, n_1565, n_1632);
  xor g1441 (n_1702, A[20], n_553);
  xor g1442 (n_560, n_1702, n_554);
  nand g1443 (n_1703, A[20], n_553);
  nand g1444 (n_1704, n_554, n_553);
  nand g1445 (n_1705, A[20], n_554);
  nand g1446 (n_573, n_1703, n_1704, n_1705);
  xor g1447 (n_1706, n_555, n_556);
  xor g1448 (n_562, n_1706, n_557);
  nand g1449 (n_1707, n_555, n_556);
  nand g1450 (n_1708, n_557, n_556);
  nand g1451 (n_1709, n_555, n_557);
  nand g1452 (n_575, n_1707, n_1708, n_1709);
  xor g1453 (n_1710, n_558, n_559);
  xor g1454 (n_564, n_1710, n_560);
  nand g1455 (n_1711, n_558, n_559);
  nand g1456 (n_1712, n_560, n_559);
  nand g1457 (n_1713, n_558, n_560);
  nand g1458 (n_577, n_1711, n_1712, n_1713);
  xor g1459 (n_1714, n_561, n_562);
  xor g1460 (n_565, n_1714, n_563);
  nand g1461 (n_1715, n_561, n_562);
  nand g1462 (n_1716, n_563, n_562);
  nand g1463 (n_1717, n_561, n_563);
  nand g1464 (n_580, n_1715, n_1716, n_1717);
  xor g1465 (n_1718, n_564, n_565);
  xor g1466 (n_177, n_1718, n_566);
  nand g1467 (n_1719, n_564, n_565);
  nand g1468 (n_1720, n_566, n_565);
  nand g1469 (n_1721, n_564, n_566);
  nand g1470 (n_100, n_1719, n_1720, n_1721);
  xor g1471 (n_1722, A[33], A[31]);
  xor g1472 (n_571, n_1722, A[27]);
  nand g1473 (n_1723, A[33], A[31]);
  nand g1474 (n_1724, A[27], A[31]);
  nand g1475 (n_1725, A[33], A[27]);
  nand g1476 (n_581, n_1723, n_1724, n_1725);
  xor g1477 (n_1726, A[19], A[17]);
  xor g1478 (n_572, n_1726, A[25]);
  nand g1479 (n_1727, A[19], A[17]);
  nand g1480 (n_1728, A[25], A[17]);
  nand g1482 (n_582, n_1727, n_1728, n_1469);
  xor g1483 (n_1730, A[15], A[29]);
  xor g1484 (n_570, n_1730, A[23]);
  nand g1485 (n_1731, A[15], A[29]);
  nand g1488 (n_583, n_1731, n_1597, n_1664);
  xor g1489 (n_1734, A[21], n_567);
  xor g1490 (n_574, n_1734, n_568);
  nand g1491 (n_1735, A[21], n_567);
  nand g1492 (n_1736, n_568, n_567);
  nand g1493 (n_1737, A[21], n_568);
  nand g1494 (n_587, n_1735, n_1736, n_1737);
  xor g1495 (n_1738, n_569, n_570);
  xor g1496 (n_576, n_1738, n_571);
  nand g1497 (n_1739, n_569, n_570);
  nand g1498 (n_1740, n_571, n_570);
  nand g1499 (n_1741, n_569, n_571);
  nand g1500 (n_589, n_1739, n_1740, n_1741);
  xor g1501 (n_1742, n_572, n_573);
  xor g1502 (n_578, n_1742, n_574);
  nand g1503 (n_1743, n_572, n_573);
  nand g1504 (n_1744, n_574, n_573);
  nand g1505 (n_1745, n_572, n_574);
  nand g1506 (n_591, n_1743, n_1744, n_1745);
  xor g1507 (n_1746, n_575, n_576);
  xor g1508 (n_579, n_1746, n_577);
  nand g1509 (n_1747, n_575, n_576);
  nand g1510 (n_1748, n_577, n_576);
  nand g1511 (n_1749, n_575, n_577);
  nand g1512 (n_594, n_1747, n_1748, n_1749);
  xor g1513 (n_1750, n_578, n_579);
  xor g1514 (n_176, n_1750, n_580);
  nand g1515 (n_1751, n_578, n_579);
  nand g1516 (n_1752, n_580, n_579);
  nand g1517 (n_1753, n_578, n_580);
  nand g1518 (n_99, n_1751, n_1752, n_1753);
  xor g1519 (n_1754, A[34], A[32]);
  xor g1520 (n_585, n_1754, A[28]);
  nand g1521 (n_1755, A[34], A[32]);
  nand g1522 (n_1756, A[28], A[32]);
  nand g1523 (n_1757, A[34], A[28]);
  nand g1524 (n_595, n_1755, n_1756, n_1757);
  xor g1526 (n_586, n_1306, A[26]);
  nand g1528 (n_1760, A[26], A[18]);
  nand g1530 (n_596, n_1307, n_1760, n_1501);
  xor g1531 (n_1762, A[16], A[30]);
  xor g1532 (n_584, n_1762, A[24]);
  nand g1533 (n_1763, A[16], A[30]);
  nand g1536 (n_597, n_1763, n_1629, n_1696);
  xor g1537 (n_1766, A[22], n_581);
  xor g1538 (n_588, n_1766, n_582);
  nand g1539 (n_1767, A[22], n_581);
  nand g1540 (n_1768, n_582, n_581);
  nand g1541 (n_1769, A[22], n_582);
  nand g1542 (n_601, n_1767, n_1768, n_1769);
  xor g1543 (n_1770, n_583, n_584);
  xor g1544 (n_590, n_1770, n_585);
  nand g1545 (n_1771, n_583, n_584);
  nand g1546 (n_1772, n_585, n_584);
  nand g1547 (n_1773, n_583, n_585);
  nand g1548 (n_603, n_1771, n_1772, n_1773);
  xor g1549 (n_1774, n_586, n_587);
  xor g1550 (n_592, n_1774, n_588);
  nand g1551 (n_1775, n_586, n_587);
  nand g1552 (n_1776, n_588, n_587);
  nand g1553 (n_1777, n_586, n_588);
  nand g1554 (n_605, n_1775, n_1776, n_1777);
  xor g1555 (n_1778, n_589, n_590);
  xor g1556 (n_593, n_1778, n_591);
  nand g1557 (n_1779, n_589, n_590);
  nand g1558 (n_1780, n_591, n_590);
  nand g1559 (n_1781, n_589, n_591);
  nand g1560 (n_608, n_1779, n_1780, n_1781);
  xor g1561 (n_1782, n_592, n_593);
  xor g1562 (n_175, n_1782, n_594);
  nand g1563 (n_1783, n_592, n_593);
  nand g1564 (n_1784, n_594, n_593);
  nand g1565 (n_1785, n_592, n_594);
  nand g1566 (n_98, n_1783, n_1784, n_1785);
  xor g1567 (n_1786, A[35], A[33]);
  xor g1568 (n_599, n_1786, A[29]);
  nand g1569 (n_1787, A[35], A[33]);
  nand g1570 (n_1788, A[29], A[33]);
  nand g1571 (n_1789, A[35], A[29]);
  nand g1572 (n_609, n_1787, n_1788, n_1789);
  xor g1574 (n_600, n_1338, A[27]);
  nand g1576 (n_1792, A[27], A[19]);
  nand g1578 (n_610, n_1339, n_1792, n_1533);
  xor g1579 (n_1794, A[17], A[31]);
  xor g1580 (n_598, n_1794, A[25]);
  nand g1581 (n_1795, A[17], A[31]);
  nand g1584 (n_611, n_1795, n_1661, n_1728);
  xor g1585 (n_1798, A[23], n_595);
  xor g1586 (n_602, n_1798, n_596);
  nand g1587 (n_1799, A[23], n_595);
  nand g1588 (n_1800, n_596, n_595);
  nand g1589 (n_1801, A[23], n_596);
  nand g1590 (n_615, n_1799, n_1800, n_1801);
  xor g1591 (n_1802, n_597, n_598);
  xor g1592 (n_604, n_1802, n_599);
  nand g1593 (n_1803, n_597, n_598);
  nand g1594 (n_1804, n_599, n_598);
  nand g1595 (n_1805, n_597, n_599);
  nand g1596 (n_617, n_1803, n_1804, n_1805);
  xor g1597 (n_1806, n_600, n_601);
  xor g1598 (n_606, n_1806, n_602);
  nand g1599 (n_1807, n_600, n_601);
  nand g1600 (n_1808, n_602, n_601);
  nand g1601 (n_1809, n_600, n_602);
  nand g1602 (n_619, n_1807, n_1808, n_1809);
  xor g1603 (n_1810, n_603, n_604);
  xor g1604 (n_607, n_1810, n_605);
  nand g1605 (n_1811, n_603, n_604);
  nand g1606 (n_1812, n_605, n_604);
  nand g1607 (n_1813, n_603, n_605);
  nand g1608 (n_622, n_1811, n_1812, n_1813);
  xor g1609 (n_1814, n_606, n_607);
  xor g1610 (n_174, n_1814, n_608);
  nand g1611 (n_1815, n_606, n_607);
  nand g1612 (n_1816, n_608, n_607);
  nand g1613 (n_1817, n_606, n_608);
  nand g1614 (n_97, n_1815, n_1816, n_1817);
  xor g1615 (n_1818, A[36], A[34]);
  xor g1616 (n_613, n_1818, A[30]);
  nand g1617 (n_1819, A[36], A[34]);
  nand g1618 (n_1820, A[30], A[34]);
  nand g1619 (n_1821, A[36], A[30]);
  nand g1620 (n_623, n_1819, n_1820, n_1821);
  xor g1622 (n_614, n_1370, A[28]);
  nand g1624 (n_1824, A[28], A[20]);
  nand g1626 (n_624, n_1371, n_1824, n_1565);
  xor g1627 (n_1826, A[18], A[32]);
  xor g1628 (n_612, n_1826, A[26]);
  nand g1629 (n_1827, A[18], A[32]);
  nand g1632 (n_625, n_1827, n_1693, n_1760);
  xor g1633 (n_1830, A[24], n_609);
  xor g1634 (n_616, n_1830, n_610);
  nand g1635 (n_1831, A[24], n_609);
  nand g1636 (n_1832, n_610, n_609);
  nand g1637 (n_1833, A[24], n_610);
  nand g1638 (n_629, n_1831, n_1832, n_1833);
  xor g1639 (n_1834, n_611, n_612);
  xor g1640 (n_618, n_1834, n_613);
  nand g1641 (n_1835, n_611, n_612);
  nand g1642 (n_1836, n_613, n_612);
  nand g1643 (n_1837, n_611, n_613);
  nand g1644 (n_631, n_1835, n_1836, n_1837);
  xor g1645 (n_1838, n_614, n_615);
  xor g1646 (n_620, n_1838, n_616);
  nand g1647 (n_1839, n_614, n_615);
  nand g1648 (n_1840, n_616, n_615);
  nand g1649 (n_1841, n_614, n_616);
  nand g1650 (n_633, n_1839, n_1840, n_1841);
  xor g1651 (n_1842, n_617, n_618);
  xor g1652 (n_621, n_1842, n_619);
  nand g1653 (n_1843, n_617, n_618);
  nand g1654 (n_1844, n_619, n_618);
  nand g1655 (n_1845, n_617, n_619);
  nand g1656 (n_636, n_1843, n_1844, n_1845);
  xor g1657 (n_1846, n_620, n_621);
  xor g1658 (n_173, n_1846, n_622);
  nand g1659 (n_1847, n_620, n_621);
  nand g1660 (n_1848, n_622, n_621);
  nand g1661 (n_1849, n_620, n_622);
  nand g1662 (n_96, n_1847, n_1848, n_1849);
  xor g1663 (n_1850, A[37], A[35]);
  xor g1664 (n_627, n_1850, A[31]);
  nand g1665 (n_1851, A[37], A[35]);
  nand g1666 (n_1852, A[31], A[35]);
  nand g1667 (n_1853, A[37], A[31]);
  nand g1668 (n_637, n_1851, n_1852, n_1853);
  xor g1670 (n_628, n_1402, A[29]);
  nand g1672 (n_1856, A[29], A[21]);
  nand g1674 (n_638, n_1403, n_1856, n_1597);
  xor g1675 (n_1858, A[19], A[33]);
  xor g1676 (n_626, n_1858, A[27]);
  nand g1677 (n_1859, A[19], A[33]);
  nand g1680 (n_639, n_1859, n_1725, n_1792);
  xor g1681 (n_1862, A[25], n_623);
  xor g1682 (n_630, n_1862, n_624);
  nand g1683 (n_1863, A[25], n_623);
  nand g1684 (n_1864, n_624, n_623);
  nand g1685 (n_1865, A[25], n_624);
  nand g1686 (n_643, n_1863, n_1864, n_1865);
  xor g1687 (n_1866, n_625, n_626);
  xor g1688 (n_632, n_1866, n_627);
  nand g1689 (n_1867, n_625, n_626);
  nand g1690 (n_1868, n_627, n_626);
  nand g1691 (n_1869, n_625, n_627);
  nand g1692 (n_645, n_1867, n_1868, n_1869);
  xor g1693 (n_1870, n_628, n_629);
  xor g1694 (n_634, n_1870, n_630);
  nand g1695 (n_1871, n_628, n_629);
  nand g1696 (n_1872, n_630, n_629);
  nand g1697 (n_1873, n_628, n_630);
  nand g1698 (n_647, n_1871, n_1872, n_1873);
  xor g1699 (n_1874, n_631, n_632);
  xor g1700 (n_635, n_1874, n_633);
  nand g1701 (n_1875, n_631, n_632);
  nand g1702 (n_1876, n_633, n_632);
  nand g1703 (n_1877, n_631, n_633);
  nand g1704 (n_650, n_1875, n_1876, n_1877);
  xor g1705 (n_1878, n_634, n_635);
  xor g1706 (n_172, n_1878, n_636);
  nand g1707 (n_1879, n_634, n_635);
  nand g1708 (n_1880, n_636, n_635);
  nand g1709 (n_1881, n_634, n_636);
  nand g1710 (n_95, n_1879, n_1880, n_1881);
  xor g1711 (n_1882, A[38], A[36]);
  xor g1712 (n_641, n_1882, A[32]);
  nand g1713 (n_1883, A[38], A[36]);
  nand g1714 (n_1884, A[32], A[36]);
  nand g1715 (n_1885, A[38], A[32]);
  nand g1716 (n_651, n_1883, n_1884, n_1885);
  xor g1718 (n_642, n_1434, A[30]);
  nand g1720 (n_1888, A[30], A[22]);
  nand g1722 (n_652, n_1435, n_1888, n_1629);
  xor g1723 (n_1890, A[20], A[34]);
  xor g1724 (n_640, n_1890, A[28]);
  nand g1725 (n_1891, A[20], A[34]);
  nand g1728 (n_653, n_1891, n_1757, n_1824);
  xor g1729 (n_1894, A[26], n_637);
  xor g1730 (n_644, n_1894, n_638);
  nand g1731 (n_1895, A[26], n_637);
  nand g1732 (n_1896, n_638, n_637);
  nand g1733 (n_1897, A[26], n_638);
  nand g1734 (n_657, n_1895, n_1896, n_1897);
  xor g1735 (n_1898, n_639, n_640);
  xor g1736 (n_646, n_1898, n_641);
  nand g1737 (n_1899, n_639, n_640);
  nand g1738 (n_1900, n_641, n_640);
  nand g1739 (n_1901, n_639, n_641);
  nand g1740 (n_659, n_1899, n_1900, n_1901);
  xor g1741 (n_1902, n_642, n_643);
  xor g1742 (n_648, n_1902, n_644);
  nand g1743 (n_1903, n_642, n_643);
  nand g1744 (n_1904, n_644, n_643);
  nand g1745 (n_1905, n_642, n_644);
  nand g1746 (n_661, n_1903, n_1904, n_1905);
  xor g1747 (n_1906, n_645, n_646);
  xor g1748 (n_649, n_1906, n_647);
  nand g1749 (n_1907, n_645, n_646);
  nand g1750 (n_1908, n_647, n_646);
  nand g1751 (n_1909, n_645, n_647);
  nand g1752 (n_664, n_1907, n_1908, n_1909);
  xor g1753 (n_1910, n_648, n_649);
  xor g1754 (n_171, n_1910, n_650);
  nand g1755 (n_1911, n_648, n_649);
  nand g1756 (n_1912, n_650, n_649);
  nand g1757 (n_1913, n_648, n_650);
  nand g1758 (n_94, n_1911, n_1912, n_1913);
  xor g1759 (n_1914, A[39], A[37]);
  xor g1760 (n_655, n_1914, A[33]);
  nand g1761 (n_1915, A[39], A[37]);
  nand g1762 (n_1916, A[33], A[37]);
  nand g1763 (n_1917, A[39], A[33]);
  nand g1764 (n_665, n_1915, n_1916, n_1917);
  xor g1766 (n_656, n_1466, A[31]);
  nand g1768 (n_1920, A[31], A[23]);
  nand g1770 (n_666, n_1467, n_1920, n_1661);
  xor g1771 (n_1922, A[21], A[35]);
  xor g1772 (n_654, n_1922, A[29]);
  nand g1773 (n_1923, A[21], A[35]);
  nand g1776 (n_667, n_1923, n_1789, n_1856);
  xor g1777 (n_1926, A[27], n_651);
  xor g1778 (n_658, n_1926, n_652);
  nand g1779 (n_1927, A[27], n_651);
  nand g1780 (n_1928, n_652, n_651);
  nand g1781 (n_1929, A[27], n_652);
  nand g1782 (n_671, n_1927, n_1928, n_1929);
  xor g1783 (n_1930, n_653, n_654);
  xor g1784 (n_660, n_1930, n_655);
  nand g1785 (n_1931, n_653, n_654);
  nand g1786 (n_1932, n_655, n_654);
  nand g1787 (n_1933, n_653, n_655);
  nand g1788 (n_673, n_1931, n_1932, n_1933);
  xor g1789 (n_1934, n_656, n_657);
  xor g1790 (n_662, n_1934, n_658);
  nand g1791 (n_1935, n_656, n_657);
  nand g1792 (n_1936, n_658, n_657);
  nand g1793 (n_1937, n_656, n_658);
  nand g1794 (n_675, n_1935, n_1936, n_1937);
  xor g1795 (n_1938, n_659, n_660);
  xor g1796 (n_663, n_1938, n_661);
  nand g1797 (n_1939, n_659, n_660);
  nand g1798 (n_1940, n_661, n_660);
  nand g1799 (n_1941, n_659, n_661);
  nand g1800 (n_678, n_1939, n_1940, n_1941);
  xor g1801 (n_1942, n_662, n_663);
  xor g1802 (n_170, n_1942, n_664);
  nand g1803 (n_1943, n_662, n_663);
  nand g1804 (n_1944, n_664, n_663);
  nand g1805 (n_1945, n_662, n_664);
  nand g1806 (n_93, n_1943, n_1944, n_1945);
  xor g1807 (n_1946, A[40], A[38]);
  xor g1808 (n_669, n_1946, A[34]);
  nand g1809 (n_1947, A[40], A[38]);
  nand g1810 (n_1948, A[34], A[38]);
  nand g1811 (n_1949, A[40], A[34]);
  nand g1812 (n_679, n_1947, n_1948, n_1949);
  xor g1814 (n_670, n_1498, A[32]);
  nand g1816 (n_1952, A[32], A[24]);
  nand g1818 (n_680, n_1499, n_1952, n_1693);
  xor g1819 (n_1954, A[22], A[36]);
  xor g1820 (n_668, n_1954, A[30]);
  nand g1821 (n_1955, A[22], A[36]);
  nand g1824 (n_681, n_1955, n_1821, n_1888);
  xor g1825 (n_1958, A[28], n_665);
  xor g1826 (n_672, n_1958, n_666);
  nand g1827 (n_1959, A[28], n_665);
  nand g1828 (n_1960, n_666, n_665);
  nand g1829 (n_1961, A[28], n_666);
  nand g1830 (n_685, n_1959, n_1960, n_1961);
  xor g1831 (n_1962, n_667, n_668);
  xor g1832 (n_674, n_1962, n_669);
  nand g1833 (n_1963, n_667, n_668);
  nand g1834 (n_1964, n_669, n_668);
  nand g1835 (n_1965, n_667, n_669);
  nand g1836 (n_687, n_1963, n_1964, n_1965);
  xor g1837 (n_1966, n_670, n_671);
  xor g1838 (n_676, n_1966, n_672);
  nand g1839 (n_1967, n_670, n_671);
  nand g1840 (n_1968, n_672, n_671);
  nand g1841 (n_1969, n_670, n_672);
  nand g1842 (n_689, n_1967, n_1968, n_1969);
  xor g1843 (n_1970, n_673, n_674);
  xor g1844 (n_677, n_1970, n_675);
  nand g1845 (n_1971, n_673, n_674);
  nand g1846 (n_1972, n_675, n_674);
  nand g1847 (n_1973, n_673, n_675);
  nand g1848 (n_692, n_1971, n_1972, n_1973);
  xor g1849 (n_1974, n_676, n_677);
  xor g1850 (n_169, n_1974, n_678);
  nand g1851 (n_1975, n_676, n_677);
  nand g1852 (n_1976, n_678, n_677);
  nand g1853 (n_1977, n_676, n_678);
  nand g1854 (n_92, n_1975, n_1976, n_1977);
  xor g1855 (n_1978, A[41], A[39]);
  xor g1856 (n_683, n_1978, A[35]);
  nand g1857 (n_1979, A[41], A[39]);
  nand g1858 (n_1980, A[35], A[39]);
  nand g1859 (n_1981, A[41], A[35]);
  nand g1860 (n_693, n_1979, n_1980, n_1981);
  xor g1862 (n_684, n_1530, A[33]);
  nand g1864 (n_1984, A[33], A[25]);
  nand g1866 (n_694, n_1531, n_1984, n_1725);
  xor g1867 (n_1986, A[23], A[37]);
  xor g1868 (n_682, n_1986, A[31]);
  nand g1869 (n_1987, A[23], A[37]);
  nand g1872 (n_695, n_1987, n_1853, n_1920);
  xor g1873 (n_1990, A[29], n_679);
  xor g1874 (n_686, n_1990, n_680);
  nand g1875 (n_1991, A[29], n_679);
  nand g1876 (n_1992, n_680, n_679);
  nand g1877 (n_1993, A[29], n_680);
  nand g1878 (n_699, n_1991, n_1992, n_1993);
  xor g1879 (n_1994, n_681, n_682);
  xor g1880 (n_688, n_1994, n_683);
  nand g1881 (n_1995, n_681, n_682);
  nand g1882 (n_1996, n_683, n_682);
  nand g1883 (n_1997, n_681, n_683);
  nand g1884 (n_701, n_1995, n_1996, n_1997);
  xor g1885 (n_1998, n_684, n_685);
  xor g1886 (n_690, n_1998, n_686);
  nand g1887 (n_1999, n_684, n_685);
  nand g1888 (n_2000, n_686, n_685);
  nand g1889 (n_2001, n_684, n_686);
  nand g1890 (n_703, n_1999, n_2000, n_2001);
  xor g1891 (n_2002, n_687, n_688);
  xor g1892 (n_691, n_2002, n_689);
  nand g1893 (n_2003, n_687, n_688);
  nand g1894 (n_2004, n_689, n_688);
  nand g1895 (n_2005, n_687, n_689);
  nand g1896 (n_706, n_2003, n_2004, n_2005);
  xor g1897 (n_2006, n_690, n_691);
  xor g1898 (n_168, n_2006, n_692);
  nand g1899 (n_2007, n_690, n_691);
  nand g1900 (n_2008, n_692, n_691);
  nand g1901 (n_2009, n_690, n_692);
  nand g1902 (n_91, n_2007, n_2008, n_2009);
  xor g1903 (n_2010, A[42], A[40]);
  xor g1904 (n_697, n_2010, A[36]);
  nand g1905 (n_2011, A[42], A[40]);
  nand g1906 (n_2012, A[36], A[40]);
  nand g1907 (n_2013, A[42], A[36]);
  nand g1908 (n_707, n_2011, n_2012, n_2013);
  xor g1910 (n_698, n_1562, A[34]);
  nand g1912 (n_2016, A[34], A[26]);
  nand g1914 (n_708, n_1563, n_2016, n_1757);
  xor g1915 (n_2018, A[24], A[38]);
  xor g1916 (n_696, n_2018, A[32]);
  nand g1917 (n_2019, A[24], A[38]);
  nand g1920 (n_709, n_2019, n_1885, n_1952);
  xor g1921 (n_2022, A[30], n_693);
  xor g1922 (n_700, n_2022, n_694);
  nand g1923 (n_2023, A[30], n_693);
  nand g1924 (n_2024, n_694, n_693);
  nand g1925 (n_2025, A[30], n_694);
  nand g1926 (n_713, n_2023, n_2024, n_2025);
  xor g1927 (n_2026, n_695, n_696);
  xor g1928 (n_702, n_2026, n_697);
  nand g1929 (n_2027, n_695, n_696);
  nand g1930 (n_2028, n_697, n_696);
  nand g1931 (n_2029, n_695, n_697);
  nand g1932 (n_715, n_2027, n_2028, n_2029);
  xor g1933 (n_2030, n_698, n_699);
  xor g1934 (n_704, n_2030, n_700);
  nand g1935 (n_2031, n_698, n_699);
  nand g1936 (n_2032, n_700, n_699);
  nand g1937 (n_2033, n_698, n_700);
  nand g1938 (n_717, n_2031, n_2032, n_2033);
  xor g1939 (n_2034, n_701, n_702);
  xor g1940 (n_705, n_2034, n_703);
  nand g1941 (n_2035, n_701, n_702);
  nand g1942 (n_2036, n_703, n_702);
  nand g1943 (n_2037, n_701, n_703);
  nand g1944 (n_720, n_2035, n_2036, n_2037);
  xor g1945 (n_2038, n_704, n_705);
  xor g1946 (n_167, n_2038, n_706);
  nand g1947 (n_2039, n_704, n_705);
  nand g1948 (n_2040, n_706, n_705);
  nand g1949 (n_2041, n_704, n_706);
  nand g1950 (n_90, n_2039, n_2040, n_2041);
  xor g1951 (n_2042, A[43], A[41]);
  xor g1952 (n_711, n_2042, A[37]);
  nand g1953 (n_2043, A[43], A[41]);
  nand g1954 (n_2044, A[37], A[41]);
  nand g1955 (n_2045, A[43], A[37]);
  nand g1956 (n_721, n_2043, n_2044, n_2045);
  xor g1958 (n_712, n_1594, A[35]);
  nand g1960 (n_2048, A[35], A[27]);
  nand g1962 (n_722, n_1595, n_2048, n_1789);
  xor g1963 (n_2050, A[25], A[39]);
  xor g1964 (n_710, n_2050, A[33]);
  nand g1965 (n_2051, A[25], A[39]);
  nand g1968 (n_723, n_2051, n_1917, n_1984);
  xor g1969 (n_2054, A[31], n_707);
  xor g1970 (n_714, n_2054, n_708);
  nand g1971 (n_2055, A[31], n_707);
  nand g1972 (n_2056, n_708, n_707);
  nand g1973 (n_2057, A[31], n_708);
  nand g1974 (n_727, n_2055, n_2056, n_2057);
  xor g1975 (n_2058, n_709, n_710);
  xor g1976 (n_716, n_2058, n_711);
  nand g1977 (n_2059, n_709, n_710);
  nand g1978 (n_2060, n_711, n_710);
  nand g1979 (n_2061, n_709, n_711);
  nand g1980 (n_729, n_2059, n_2060, n_2061);
  xor g1981 (n_2062, n_712, n_713);
  xor g1982 (n_718, n_2062, n_714);
  nand g1983 (n_2063, n_712, n_713);
  nand g1984 (n_2064, n_714, n_713);
  nand g1985 (n_2065, n_712, n_714);
  nand g1986 (n_731, n_2063, n_2064, n_2065);
  xor g1987 (n_2066, n_715, n_716);
  xor g1988 (n_719, n_2066, n_717);
  nand g1989 (n_2067, n_715, n_716);
  nand g1990 (n_2068, n_717, n_716);
  nand g1991 (n_2069, n_715, n_717);
  nand g1992 (n_734, n_2067, n_2068, n_2069);
  xor g1993 (n_2070, n_718, n_719);
  xor g1994 (n_166, n_2070, n_720);
  nand g1995 (n_2071, n_718, n_719);
  nand g1996 (n_2072, n_720, n_719);
  nand g1997 (n_2073, n_718, n_720);
  nand g1998 (n_89, n_2071, n_2072, n_2073);
  xor g1999 (n_2074, A[44], A[42]);
  xor g2000 (n_725, n_2074, A[38]);
  nand g2001 (n_2075, A[44], A[42]);
  nand g2002 (n_2076, A[38], A[42]);
  nand g2003 (n_2077, A[44], A[38]);
  nand g2004 (n_735, n_2075, n_2076, n_2077);
  xor g2006 (n_726, n_1626, A[36]);
  nand g2008 (n_2080, A[36], A[28]);
  nand g2010 (n_736, n_1627, n_2080, n_1821);
  xor g2011 (n_2082, A[26], A[40]);
  xor g2012 (n_724, n_2082, A[34]);
  nand g2013 (n_2083, A[26], A[40]);
  nand g2016 (n_737, n_2083, n_1949, n_2016);
  xor g2017 (n_2086, A[32], n_721);
  xor g2018 (n_728, n_2086, n_722);
  nand g2019 (n_2087, A[32], n_721);
  nand g2020 (n_2088, n_722, n_721);
  nand g2021 (n_2089, A[32], n_722);
  nand g2022 (n_741, n_2087, n_2088, n_2089);
  xor g2023 (n_2090, n_723, n_724);
  xor g2024 (n_730, n_2090, n_725);
  nand g2025 (n_2091, n_723, n_724);
  nand g2026 (n_2092, n_725, n_724);
  nand g2027 (n_2093, n_723, n_725);
  nand g2028 (n_743, n_2091, n_2092, n_2093);
  xor g2029 (n_2094, n_726, n_727);
  xor g2030 (n_732, n_2094, n_728);
  nand g2031 (n_2095, n_726, n_727);
  nand g2032 (n_2096, n_728, n_727);
  nand g2033 (n_2097, n_726, n_728);
  nand g2034 (n_745, n_2095, n_2096, n_2097);
  xor g2035 (n_2098, n_729, n_730);
  xor g2036 (n_733, n_2098, n_731);
  nand g2037 (n_2099, n_729, n_730);
  nand g2038 (n_2100, n_731, n_730);
  nand g2039 (n_2101, n_729, n_731);
  nand g2040 (n_748, n_2099, n_2100, n_2101);
  xor g2041 (n_2102, n_732, n_733);
  xor g2042 (n_165, n_2102, n_734);
  nand g2043 (n_2103, n_732, n_733);
  nand g2044 (n_2104, n_734, n_733);
  nand g2045 (n_2105, n_732, n_734);
  nand g2046 (n_88, n_2103, n_2104, n_2105);
  xor g2047 (n_2106, A[45], A[43]);
  xor g2048 (n_739, n_2106, A[39]);
  nand g2049 (n_2107, A[45], A[43]);
  nand g2050 (n_2108, A[39], A[43]);
  nand g2051 (n_2109, A[45], A[39]);
  nand g2052 (n_749, n_2107, n_2108, n_2109);
  xor g2054 (n_740, n_1658, A[37]);
  nand g2056 (n_2112, A[37], A[29]);
  nand g2058 (n_750, n_1659, n_2112, n_1853);
  xor g2059 (n_2114, A[27], A[41]);
  xor g2060 (n_738, n_2114, A[35]);
  nand g2061 (n_2115, A[27], A[41]);
  nand g2064 (n_751, n_2115, n_1981, n_2048);
  xor g2065 (n_2118, A[33], n_735);
  xor g2066 (n_742, n_2118, n_736);
  nand g2067 (n_2119, A[33], n_735);
  nand g2068 (n_2120, n_736, n_735);
  nand g2069 (n_2121, A[33], n_736);
  nand g2070 (n_755, n_2119, n_2120, n_2121);
  xor g2071 (n_2122, n_737, n_738);
  xor g2072 (n_744, n_2122, n_739);
  nand g2073 (n_2123, n_737, n_738);
  nand g2074 (n_2124, n_739, n_738);
  nand g2075 (n_2125, n_737, n_739);
  nand g2076 (n_757, n_2123, n_2124, n_2125);
  xor g2077 (n_2126, n_740, n_741);
  xor g2078 (n_746, n_2126, n_742);
  nand g2079 (n_2127, n_740, n_741);
  nand g2080 (n_2128, n_742, n_741);
  nand g2081 (n_2129, n_740, n_742);
  nand g2082 (n_759, n_2127, n_2128, n_2129);
  xor g2083 (n_2130, n_743, n_744);
  xor g2084 (n_747, n_2130, n_745);
  nand g2085 (n_2131, n_743, n_744);
  nand g2086 (n_2132, n_745, n_744);
  nand g2087 (n_2133, n_743, n_745);
  nand g2088 (n_762, n_2131, n_2132, n_2133);
  xor g2089 (n_2134, n_746, n_747);
  xor g2090 (n_164, n_2134, n_748);
  nand g2091 (n_2135, n_746, n_747);
  nand g2092 (n_2136, n_748, n_747);
  nand g2093 (n_2137, n_746, n_748);
  nand g2094 (n_87, n_2135, n_2136, n_2137);
  xor g2095 (n_2138, A[46], A[44]);
  xor g2096 (n_753, n_2138, A[40]);
  nand g2097 (n_2139, A[46], A[44]);
  nand g2098 (n_2140, A[40], A[44]);
  nand g2099 (n_2141, A[46], A[40]);
  nand g2100 (n_763, n_2139, n_2140, n_2141);
  xor g2102 (n_754, n_1690, A[38]);
  nand g2104 (n_2144, A[38], A[30]);
  nand g2106 (n_764, n_1691, n_2144, n_1885);
  xor g2107 (n_2146, A[28], A[42]);
  xor g2108 (n_752, n_2146, A[36]);
  nand g2109 (n_2147, A[28], A[42]);
  nand g2112 (n_765, n_2147, n_2013, n_2080);
  xor g2113 (n_2150, A[34], n_749);
  xor g2114 (n_756, n_2150, n_750);
  nand g2115 (n_2151, A[34], n_749);
  nand g2116 (n_2152, n_750, n_749);
  nand g2117 (n_2153, A[34], n_750);
  nand g2118 (n_769, n_2151, n_2152, n_2153);
  xor g2119 (n_2154, n_751, n_752);
  xor g2120 (n_758, n_2154, n_753);
  nand g2121 (n_2155, n_751, n_752);
  nand g2122 (n_2156, n_753, n_752);
  nand g2123 (n_2157, n_751, n_753);
  nand g2124 (n_771, n_2155, n_2156, n_2157);
  xor g2125 (n_2158, n_754, n_755);
  xor g2126 (n_760, n_2158, n_756);
  nand g2127 (n_2159, n_754, n_755);
  nand g2128 (n_2160, n_756, n_755);
  nand g2129 (n_2161, n_754, n_756);
  nand g2130 (n_773, n_2159, n_2160, n_2161);
  xor g2131 (n_2162, n_757, n_758);
  xor g2132 (n_761, n_2162, n_759);
  nand g2133 (n_2163, n_757, n_758);
  nand g2134 (n_2164, n_759, n_758);
  nand g2135 (n_2165, n_757, n_759);
  nand g2136 (n_776, n_2163, n_2164, n_2165);
  xor g2137 (n_2166, n_760, n_761);
  xor g2138 (n_163, n_2166, n_762);
  nand g2139 (n_2167, n_760, n_761);
  nand g2140 (n_2168, n_762, n_761);
  nand g2141 (n_2169, n_760, n_762);
  nand g2142 (n_86, n_2167, n_2168, n_2169);
  xor g2143 (n_2170, A[47], A[45]);
  xor g2144 (n_767, n_2170, A[41]);
  nand g2145 (n_2171, A[47], A[45]);
  nand g2146 (n_2172, A[41], A[45]);
  nand g2147 (n_2173, A[47], A[41]);
  nand g2148 (n_777, n_2171, n_2172, n_2173);
  xor g2150 (n_768, n_1722, A[39]);
  nand g2152 (n_2176, A[39], A[31]);
  nand g2154 (n_778, n_1723, n_2176, n_1917);
  xor g2155 (n_2178, A[29], A[43]);
  xor g2156 (n_766, n_2178, A[37]);
  nand g2157 (n_2179, A[29], A[43]);
  nand g2160 (n_779, n_2179, n_2045, n_2112);
  xor g2161 (n_2182, A[35], n_763);
  xor g2162 (n_770, n_2182, n_764);
  nand g2163 (n_2183, A[35], n_763);
  nand g2164 (n_2184, n_764, n_763);
  nand g2165 (n_2185, A[35], n_764);
  nand g2166 (n_783, n_2183, n_2184, n_2185);
  xor g2167 (n_2186, n_765, n_766);
  xor g2168 (n_772, n_2186, n_767);
  nand g2169 (n_2187, n_765, n_766);
  nand g2170 (n_2188, n_767, n_766);
  nand g2171 (n_2189, n_765, n_767);
  nand g2172 (n_785, n_2187, n_2188, n_2189);
  xor g2173 (n_2190, n_768, n_769);
  xor g2174 (n_774, n_2190, n_770);
  nand g2175 (n_2191, n_768, n_769);
  nand g2176 (n_2192, n_770, n_769);
  nand g2177 (n_2193, n_768, n_770);
  nand g2178 (n_787, n_2191, n_2192, n_2193);
  xor g2179 (n_2194, n_771, n_772);
  xor g2180 (n_775, n_2194, n_773);
  nand g2181 (n_2195, n_771, n_772);
  nand g2182 (n_2196, n_773, n_772);
  nand g2183 (n_2197, n_771, n_773);
  nand g2184 (n_790, n_2195, n_2196, n_2197);
  xor g2185 (n_2198, n_774, n_775);
  xor g2186 (n_162, n_2198, n_776);
  nand g2187 (n_2199, n_774, n_775);
  nand g2188 (n_2200, n_776, n_775);
  nand g2189 (n_2201, n_774, n_776);
  nand g2190 (n_85, n_2199, n_2200, n_2201);
  xor g2191 (n_2202, A[48], A[46]);
  xor g2192 (n_781, n_2202, A[42]);
  nand g2193 (n_2203, A[48], A[46]);
  nand g2194 (n_2204, A[42], A[46]);
  nand g2195 (n_2205, A[48], A[42]);
  nand g2196 (n_791, n_2203, n_2204, n_2205);
  xor g2198 (n_782, n_1754, A[40]);
  nand g2200 (n_2208, A[40], A[32]);
  nand g2202 (n_792, n_1755, n_2208, n_1949);
  xor g2203 (n_2210, A[30], A[44]);
  xor g2204 (n_780, n_2210, A[38]);
  nand g2205 (n_2211, A[30], A[44]);
  nand g2208 (n_793, n_2211, n_2077, n_2144);
  xor g2209 (n_2214, A[36], n_777);
  xor g2210 (n_784, n_2214, n_778);
  nand g2211 (n_2215, A[36], n_777);
  nand g2212 (n_2216, n_778, n_777);
  nand g2213 (n_2217, A[36], n_778);
  nand g2214 (n_797, n_2215, n_2216, n_2217);
  xor g2215 (n_2218, n_779, n_780);
  xor g2216 (n_786, n_2218, n_781);
  nand g2217 (n_2219, n_779, n_780);
  nand g2218 (n_2220, n_781, n_780);
  nand g2219 (n_2221, n_779, n_781);
  nand g2220 (n_799, n_2219, n_2220, n_2221);
  xor g2221 (n_2222, n_782, n_783);
  xor g2222 (n_788, n_2222, n_784);
  nand g2223 (n_2223, n_782, n_783);
  nand g2224 (n_2224, n_784, n_783);
  nand g2225 (n_2225, n_782, n_784);
  nand g2226 (n_801, n_2223, n_2224, n_2225);
  xor g2227 (n_2226, n_785, n_786);
  xor g2228 (n_789, n_2226, n_787);
  nand g2229 (n_2227, n_785, n_786);
  nand g2230 (n_2228, n_787, n_786);
  nand g2231 (n_2229, n_785, n_787);
  nand g2232 (n_804, n_2227, n_2228, n_2229);
  xor g2233 (n_2230, n_788, n_789);
  xor g2234 (n_161, n_2230, n_790);
  nand g2235 (n_2231, n_788, n_789);
  nand g2236 (n_2232, n_790, n_789);
  nand g2237 (n_2233, n_788, n_790);
  nand g2238 (n_84, n_2231, n_2232, n_2233);
  xor g2239 (n_2234, A[49], A[47]);
  xor g2240 (n_795, n_2234, A[43]);
  nand g2241 (n_2235, A[49], A[47]);
  nand g2242 (n_2236, A[43], A[47]);
  nand g2243 (n_2237, A[49], A[43]);
  nand g2244 (n_805, n_2235, n_2236, n_2237);
  xor g2246 (n_796, n_1786, A[41]);
  nand g2248 (n_2240, A[41], A[33]);
  nand g2250 (n_806, n_1787, n_2240, n_1981);
  xor g2251 (n_2242, A[31], A[45]);
  xor g2252 (n_794, n_2242, A[39]);
  nand g2253 (n_2243, A[31], A[45]);
  nand g2256 (n_807, n_2243, n_2109, n_2176);
  xor g2257 (n_2246, A[37], n_791);
  xor g2258 (n_798, n_2246, n_792);
  nand g2259 (n_2247, A[37], n_791);
  nand g2260 (n_2248, n_792, n_791);
  nand g2261 (n_2249, A[37], n_792);
  nand g2262 (n_811, n_2247, n_2248, n_2249);
  xor g2263 (n_2250, n_793, n_794);
  xor g2264 (n_800, n_2250, n_795);
  nand g2265 (n_2251, n_793, n_794);
  nand g2266 (n_2252, n_795, n_794);
  nand g2267 (n_2253, n_793, n_795);
  nand g2268 (n_813, n_2251, n_2252, n_2253);
  xor g2269 (n_2254, n_796, n_797);
  xor g2270 (n_802, n_2254, n_798);
  nand g2271 (n_2255, n_796, n_797);
  nand g2272 (n_2256, n_798, n_797);
  nand g2273 (n_2257, n_796, n_798);
  nand g2274 (n_815, n_2255, n_2256, n_2257);
  xor g2275 (n_2258, n_799, n_800);
  xor g2276 (n_803, n_2258, n_801);
  nand g2277 (n_2259, n_799, n_800);
  nand g2278 (n_2260, n_801, n_800);
  nand g2279 (n_2261, n_799, n_801);
  nand g2280 (n_818, n_2259, n_2260, n_2261);
  xor g2281 (n_2262, n_802, n_803);
  xor g2282 (n_160, n_2262, n_804);
  nand g2283 (n_2263, n_802, n_803);
  nand g2284 (n_2264, n_804, n_803);
  nand g2285 (n_2265, n_802, n_804);
  nand g2286 (n_83, n_2263, n_2264, n_2265);
  xor g2287 (n_2266, A[50], A[48]);
  xor g2288 (n_809, n_2266, A[44]);
  nand g2289 (n_2267, A[50], A[48]);
  nand g2290 (n_2268, A[44], A[48]);
  nand g2291 (n_2269, A[50], A[44]);
  nand g2292 (n_819, n_2267, n_2268, n_2269);
  xor g2294 (n_810, n_1818, A[42]);
  nand g2296 (n_2272, A[42], A[34]);
  nand g2298 (n_820, n_1819, n_2272, n_2013);
  xor g2299 (n_2274, A[32], A[46]);
  xor g2300 (n_808, n_2274, A[40]);
  nand g2301 (n_2275, A[32], A[46]);
  nand g2304 (n_821, n_2275, n_2141, n_2208);
  xor g2305 (n_2278, A[38], n_805);
  xor g2306 (n_812, n_2278, n_806);
  nand g2307 (n_2279, A[38], n_805);
  nand g2308 (n_2280, n_806, n_805);
  nand g2309 (n_2281, A[38], n_806);
  nand g2310 (n_825, n_2279, n_2280, n_2281);
  xor g2311 (n_2282, n_807, n_808);
  xor g2312 (n_814, n_2282, n_809);
  nand g2313 (n_2283, n_807, n_808);
  nand g2314 (n_2284, n_809, n_808);
  nand g2315 (n_2285, n_807, n_809);
  nand g2316 (n_827, n_2283, n_2284, n_2285);
  xor g2317 (n_2286, n_810, n_811);
  xor g2318 (n_816, n_2286, n_812);
  nand g2319 (n_2287, n_810, n_811);
  nand g2320 (n_2288, n_812, n_811);
  nand g2321 (n_2289, n_810, n_812);
  nand g2322 (n_829, n_2287, n_2288, n_2289);
  xor g2323 (n_2290, n_813, n_814);
  xor g2324 (n_817, n_2290, n_815);
  nand g2325 (n_2291, n_813, n_814);
  nand g2326 (n_2292, n_815, n_814);
  nand g2327 (n_2293, n_813, n_815);
  nand g2328 (n_832, n_2291, n_2292, n_2293);
  xor g2329 (n_2294, n_816, n_817);
  xor g2330 (n_159, n_2294, n_818);
  nand g2331 (n_2295, n_816, n_817);
  nand g2332 (n_2296, n_818, n_817);
  nand g2333 (n_2297, n_816, n_818);
  nand g2334 (n_82, n_2295, n_2296, n_2297);
  xor g2335 (n_2298, A[51], A[49]);
  xor g2336 (n_823, n_2298, A[45]);
  nand g2337 (n_2299, A[51], A[49]);
  nand g2338 (n_2300, A[45], A[49]);
  nand g2339 (n_2301, A[51], A[45]);
  nand g2340 (n_833, n_2299, n_2300, n_2301);
  xor g2342 (n_824, n_1850, A[43]);
  nand g2344 (n_2304, A[43], A[35]);
  nand g2346 (n_834, n_1851, n_2304, n_2045);
  xor g2347 (n_2306, A[33], A[47]);
  xor g2348 (n_822, n_2306, A[41]);
  nand g2349 (n_2307, A[33], A[47]);
  nand g2352 (n_835, n_2307, n_2173, n_2240);
  xor g2353 (n_2310, A[39], n_819);
  xor g2354 (n_826, n_2310, n_820);
  nand g2355 (n_2311, A[39], n_819);
  nand g2356 (n_2312, n_820, n_819);
  nand g2357 (n_2313, A[39], n_820);
  nand g2358 (n_839, n_2311, n_2312, n_2313);
  xor g2359 (n_2314, n_821, n_822);
  xor g2360 (n_828, n_2314, n_823);
  nand g2361 (n_2315, n_821, n_822);
  nand g2362 (n_2316, n_823, n_822);
  nand g2363 (n_2317, n_821, n_823);
  nand g2364 (n_841, n_2315, n_2316, n_2317);
  xor g2365 (n_2318, n_824, n_825);
  xor g2366 (n_830, n_2318, n_826);
  nand g2367 (n_2319, n_824, n_825);
  nand g2368 (n_2320, n_826, n_825);
  nand g2369 (n_2321, n_824, n_826);
  nand g2370 (n_843, n_2319, n_2320, n_2321);
  xor g2371 (n_2322, n_827, n_828);
  xor g2372 (n_831, n_2322, n_829);
  nand g2373 (n_2323, n_827, n_828);
  nand g2374 (n_2324, n_829, n_828);
  nand g2375 (n_2325, n_827, n_829);
  nand g2376 (n_846, n_2323, n_2324, n_2325);
  xor g2377 (n_2326, n_830, n_831);
  xor g2378 (n_158, n_2326, n_832);
  nand g2379 (n_2327, n_830, n_831);
  nand g2380 (n_2328, n_832, n_831);
  nand g2381 (n_2329, n_830, n_832);
  nand g2382 (n_81, n_2327, n_2328, n_2329);
  xor g2383 (n_2330, A[52], A[50]);
  xor g2384 (n_837, n_2330, A[46]);
  nand g2385 (n_2331, A[52], A[50]);
  nand g2386 (n_2332, A[46], A[50]);
  nand g2387 (n_2333, A[52], A[46]);
  nand g2388 (n_847, n_2331, n_2332, n_2333);
  xor g2390 (n_838, n_1882, A[44]);
  nand g2392 (n_2336, A[44], A[36]);
  nand g2394 (n_848, n_1883, n_2336, n_2077);
  xor g2395 (n_2338, A[34], A[48]);
  xor g2396 (n_836, n_2338, A[42]);
  nand g2397 (n_2339, A[34], A[48]);
  nand g2400 (n_849, n_2339, n_2205, n_2272);
  xor g2401 (n_2342, A[40], n_833);
  xor g2402 (n_840, n_2342, n_834);
  nand g2403 (n_2343, A[40], n_833);
  nand g2404 (n_2344, n_834, n_833);
  nand g2405 (n_2345, A[40], n_834);
  nand g2406 (n_853, n_2343, n_2344, n_2345);
  xor g2407 (n_2346, n_835, n_836);
  xor g2408 (n_842, n_2346, n_837);
  nand g2409 (n_2347, n_835, n_836);
  nand g2410 (n_2348, n_837, n_836);
  nand g2411 (n_2349, n_835, n_837);
  nand g2412 (n_855, n_2347, n_2348, n_2349);
  xor g2413 (n_2350, n_838, n_839);
  xor g2414 (n_844, n_2350, n_840);
  nand g2415 (n_2351, n_838, n_839);
  nand g2416 (n_2352, n_840, n_839);
  nand g2417 (n_2353, n_838, n_840);
  nand g2418 (n_857, n_2351, n_2352, n_2353);
  xor g2419 (n_2354, n_841, n_842);
  xor g2420 (n_845, n_2354, n_843);
  nand g2421 (n_2355, n_841, n_842);
  nand g2422 (n_2356, n_843, n_842);
  nand g2423 (n_2357, n_841, n_843);
  nand g2424 (n_860, n_2355, n_2356, n_2357);
  xor g2425 (n_2358, n_844, n_845);
  xor g2426 (n_157, n_2358, n_846);
  nand g2427 (n_2359, n_844, n_845);
  nand g2428 (n_2360, n_846, n_845);
  nand g2429 (n_2361, n_844, n_846);
  nand g2430 (n_80, n_2359, n_2360, n_2361);
  xor g2431 (n_2362, A[53], A[51]);
  xor g2432 (n_851, n_2362, A[47]);
  nand g2433 (n_2363, A[53], A[51]);
  nand g2434 (n_2364, A[47], A[51]);
  nand g2435 (n_2365, A[53], A[47]);
  nand g2436 (n_861, n_2363, n_2364, n_2365);
  xor g2438 (n_852, n_1914, A[45]);
  nand g2440 (n_2368, A[45], A[37]);
  nand g2442 (n_862, n_1915, n_2368, n_2109);
  xor g2443 (n_2370, A[35], A[49]);
  xor g2444 (n_850, n_2370, A[43]);
  nand g2445 (n_2371, A[35], A[49]);
  nand g2448 (n_863, n_2371, n_2237, n_2304);
  xor g2449 (n_2374, A[41], n_847);
  xor g2450 (n_854, n_2374, n_848);
  nand g2451 (n_2375, A[41], n_847);
  nand g2452 (n_2376, n_848, n_847);
  nand g2453 (n_2377, A[41], n_848);
  nand g2454 (n_867, n_2375, n_2376, n_2377);
  xor g2455 (n_2378, n_849, n_850);
  xor g2456 (n_856, n_2378, n_851);
  nand g2457 (n_2379, n_849, n_850);
  nand g2458 (n_2380, n_851, n_850);
  nand g2459 (n_2381, n_849, n_851);
  nand g2460 (n_869, n_2379, n_2380, n_2381);
  xor g2461 (n_2382, n_852, n_853);
  xor g2462 (n_858, n_2382, n_854);
  nand g2463 (n_2383, n_852, n_853);
  nand g2464 (n_2384, n_854, n_853);
  nand g2465 (n_2385, n_852, n_854);
  nand g2466 (n_871, n_2383, n_2384, n_2385);
  xor g2467 (n_2386, n_855, n_856);
  xor g2468 (n_859, n_2386, n_857);
  nand g2469 (n_2387, n_855, n_856);
  nand g2470 (n_2388, n_857, n_856);
  nand g2471 (n_2389, n_855, n_857);
  nand g2472 (n_874, n_2387, n_2388, n_2389);
  xor g2473 (n_2390, n_858, n_859);
  xor g2474 (n_156, n_2390, n_860);
  nand g2475 (n_2391, n_858, n_859);
  nand g2476 (n_2392, n_860, n_859);
  nand g2477 (n_2393, n_858, n_860);
  nand g2478 (n_79, n_2391, n_2392, n_2393);
  xor g2479 (n_2394, A[54], A[52]);
  xor g2480 (n_865, n_2394, A[48]);
  nand g2481 (n_2395, A[54], A[52]);
  nand g2482 (n_2396, A[48], A[52]);
  nand g2483 (n_2397, A[54], A[48]);
  nand g2484 (n_875, n_2395, n_2396, n_2397);
  xor g2486 (n_866, n_1946, A[46]);
  nand g2488 (n_2400, A[46], A[38]);
  nand g2490 (n_876, n_1947, n_2400, n_2141);
  xor g2491 (n_2402, A[36], A[50]);
  xor g2492 (n_864, n_2402, A[44]);
  nand g2493 (n_2403, A[36], A[50]);
  nand g2496 (n_877, n_2403, n_2269, n_2336);
  xor g2497 (n_2406, A[42], n_861);
  xor g2498 (n_868, n_2406, n_862);
  nand g2499 (n_2407, A[42], n_861);
  nand g2500 (n_2408, n_862, n_861);
  nand g2501 (n_2409, A[42], n_862);
  nand g2502 (n_881, n_2407, n_2408, n_2409);
  xor g2503 (n_2410, n_863, n_864);
  xor g2504 (n_870, n_2410, n_865);
  nand g2505 (n_2411, n_863, n_864);
  nand g2506 (n_2412, n_865, n_864);
  nand g2507 (n_2413, n_863, n_865);
  nand g2508 (n_883, n_2411, n_2412, n_2413);
  xor g2509 (n_2414, n_866, n_867);
  xor g2510 (n_872, n_2414, n_868);
  nand g2511 (n_2415, n_866, n_867);
  nand g2512 (n_2416, n_868, n_867);
  nand g2513 (n_2417, n_866, n_868);
  nand g2514 (n_885, n_2415, n_2416, n_2417);
  xor g2515 (n_2418, n_869, n_870);
  xor g2516 (n_873, n_2418, n_871);
  nand g2517 (n_2419, n_869, n_870);
  nand g2518 (n_2420, n_871, n_870);
  nand g2519 (n_2421, n_869, n_871);
  nand g2520 (n_888, n_2419, n_2420, n_2421);
  xor g2521 (n_2422, n_872, n_873);
  xor g2522 (n_155, n_2422, n_874);
  nand g2523 (n_2423, n_872, n_873);
  nand g2524 (n_2424, n_874, n_873);
  nand g2525 (n_2425, n_872, n_874);
  nand g2526 (n_78, n_2423, n_2424, n_2425);
  xor g2527 (n_2426, A[55], A[53]);
  xor g2528 (n_879, n_2426, A[49]);
  nand g2529 (n_2427, A[55], A[53]);
  nand g2530 (n_2428, A[49], A[53]);
  nand g2531 (n_2429, A[55], A[49]);
  nand g2532 (n_892, n_2427, n_2428, n_2429);
  xor g2534 (n_880, n_1978, A[47]);
  nand g2536 (n_2432, A[47], A[39]);
  nand g2538 (n_893, n_1979, n_2432, n_2173);
  xor g2539 (n_2434, A[37], A[51]);
  xor g2540 (n_878, n_2434, A[45]);
  nand g2541 (n_2435, A[37], A[51]);
  nand g2544 (n_891, n_2435, n_2301, n_2368);
  xor g2545 (n_2438, A[43], n_875);
  xor g2546 (n_882, n_2438, n_876);
  nand g2547 (n_2439, A[43], n_875);
  nand g2548 (n_2440, n_876, n_875);
  nand g2549 (n_2441, A[43], n_876);
  nand g2550 (n_897, n_2439, n_2440, n_2441);
  xor g2551 (n_2442, n_877, n_878);
  xor g2552 (n_884, n_2442, n_879);
  nand g2553 (n_2443, n_877, n_878);
  nand g2554 (n_2444, n_879, n_878);
  nand g2555 (n_2445, n_877, n_879);
  nand g2556 (n_899, n_2443, n_2444, n_2445);
  xor g2557 (n_2446, n_880, n_881);
  xor g2558 (n_886, n_2446, n_882);
  nand g2559 (n_2447, n_880, n_881);
  nand g2560 (n_2448, n_882, n_881);
  nand g2561 (n_2449, n_880, n_882);
  nand g2562 (n_901, n_2447, n_2448, n_2449);
  xor g2563 (n_2450, n_883, n_884);
  xor g2564 (n_887, n_2450, n_885);
  nand g2565 (n_2451, n_883, n_884);
  nand g2566 (n_2452, n_885, n_884);
  nand g2567 (n_2453, n_883, n_885);
  nand g2568 (n_904, n_2451, n_2452, n_2453);
  xor g2569 (n_2454, n_886, n_887);
  xor g2570 (n_154, n_2454, n_888);
  nand g2571 (n_2455, n_886, n_887);
  nand g2572 (n_2456, n_888, n_887);
  nand g2573 (n_2457, n_886, n_888);
  nand g2574 (n_77, n_2455, n_2456, n_2457);
  xor g2577 (n_2458, A[56], A[50]);
  xor g2578 (n_895, n_2458, A[42]);
  nand g2579 (n_2459, A[56], A[50]);
  nand g2580 (n_2460, A[42], A[50]);
  nand g2581 (n_2461, A[56], A[42]);
  nand g2582 (n_909, n_2459, n_2460, n_2461);
  xor g2583 (n_2462, A[40], A[54]);
  xor g2584 (n_896, n_2462, A[38]);
  nand g2585 (n_2463, A[40], A[54]);
  nand g2586 (n_2464, A[38], A[54]);
  nand g2588 (n_910, n_2463, n_2464, n_1947);
  xor g2589 (n_2466, A[48], A[52]);
  xor g2590 (n_894, n_2466, A[46]);
  nand g2594 (n_908, n_2396, n_2333, n_2203);
  xor g2595 (n_2470, A[44], n_891);
  xor g2596 (n_898, n_2470, n_892);
  nand g2597 (n_2471, A[44], n_891);
  nand g2598 (n_2472, n_892, n_891);
  nand g2599 (n_2473, A[44], n_892);
  nand g2600 (n_914, n_2471, n_2472, n_2473);
  xor g2601 (n_2474, n_893, n_894);
  xor g2602 (n_900, n_2474, n_895);
  nand g2603 (n_2475, n_893, n_894);
  nand g2604 (n_2476, n_895, n_894);
  nand g2605 (n_2477, n_893, n_895);
  nand g2606 (n_916, n_2475, n_2476, n_2477);
  xor g2607 (n_2478, n_896, n_897);
  xor g2608 (n_902, n_2478, n_898);
  nand g2609 (n_2479, n_896, n_897);
  nand g2610 (n_2480, n_898, n_897);
  nand g2611 (n_2481, n_896, n_898);
  nand g2612 (n_918, n_2479, n_2480, n_2481);
  xor g2613 (n_2482, n_899, n_900);
  xor g2614 (n_903, n_2482, n_901);
  nand g2615 (n_2483, n_899, n_900);
  nand g2616 (n_2484, n_901, n_900);
  nand g2617 (n_2485, n_899, n_901);
  nand g2618 (n_921, n_2483, n_2484, n_2485);
  xor g2619 (n_2486, n_902, n_903);
  xor g2620 (n_153, n_2486, n_904);
  nand g2621 (n_2487, n_902, n_903);
  nand g2622 (n_2488, n_904, n_903);
  nand g2623 (n_2489, n_902, n_904);
  nand g2624 (n_76, n_2487, n_2488, n_2489);
  xor g2627 (n_2490, A[49], A[41]);
  xor g2628 (n_912, n_2490, A[39]);
  nand g2629 (n_2491, A[49], A[41]);
  nand g2631 (n_2493, A[49], A[39]);
  nand g2632 (n_923, n_2491, n_1979, n_2493);
  xor g2633 (n_2494, A[56], A[55]);
  xor g2634 (n_913, n_2494, A[47]);
  nand g2635 (n_2495, A[56], A[55]);
  nand g2636 (n_2496, A[47], A[55]);
  nand g2637 (n_2497, A[56], A[47]);
  nand g2638 (n_924, n_2495, n_2496, n_2497);
  xor g2640 (n_911, n_2362, A[45]);
  nand g2643 (n_2501, A[53], A[45]);
  nand g2644 (n_925, n_2363, n_2301, n_2501);
  xor g2645 (n_2502, A[43], n_908);
  xor g2646 (n_915, n_2502, n_909);
  nand g2647 (n_2503, A[43], n_908);
  nand g2648 (n_2504, n_909, n_908);
  nand g2649 (n_2505, A[43], n_909);
  nand g2650 (n_929, n_2503, n_2504, n_2505);
  xor g2651 (n_2506, n_910, n_911);
  xor g2652 (n_917, n_2506, n_912);
  nand g2653 (n_2507, n_910, n_911);
  nand g2654 (n_2508, n_912, n_911);
  nand g2655 (n_2509, n_910, n_912);
  nand g2656 (n_931, n_2507, n_2508, n_2509);
  xor g2657 (n_2510, n_913, n_914);
  xor g2658 (n_919, n_2510, n_915);
  nand g2659 (n_2511, n_913, n_914);
  nand g2660 (n_2512, n_915, n_914);
  nand g2661 (n_2513, n_913, n_915);
  nand g2662 (n_933, n_2511, n_2512, n_2513);
  xor g2663 (n_2514, n_916, n_917);
  xor g2664 (n_920, n_2514, n_918);
  nand g2665 (n_2515, n_916, n_917);
  nand g2666 (n_2516, n_918, n_917);
  nand g2667 (n_2517, n_916, n_918);
  nand g2668 (n_936, n_2515, n_2516, n_2517);
  xor g2669 (n_2518, n_919, n_920);
  xor g2670 (n_152, n_2518, n_921);
  nand g2671 (n_2519, n_919, n_920);
  nand g2672 (n_2520, n_921, n_920);
  nand g2673 (n_2521, n_919, n_921);
  nand g2674 (n_75, n_2519, n_2520, n_2521);
  xor g2676 (n_927, n_2522, A[50]);
  nand g2678 (n_2524, A[50], A[54]);
  nand g2680 (n_939, n_2523, n_2524, n_2525);
  xor g2682 (n_928, n_2010, A[48]);
  nand g2684 (n_2528, A[48], A[40]);
  nand g2686 (n_940, n_2011, n_2528, n_2205);
  xor g2688 (n_926, n_2530, A[46]);
  nand g2692 (n_941, n_2531, n_2333, n_2533);
  xor g2693 (n_2534, A[44], n_923);
  xor g2694 (n_930, n_2534, n_924);
  nand g2695 (n_2535, A[44], n_923);
  nand g2696 (n_2536, n_924, n_923);
  nand g2697 (n_2537, A[44], n_924);
  nand g2698 (n_945, n_2535, n_2536, n_2537);
  xor g2699 (n_2538, n_925, n_926);
  xor g2700 (n_932, n_2538, n_927);
  nand g2701 (n_2539, n_925, n_926);
  nand g2702 (n_2540, n_927, n_926);
  nand g2703 (n_2541, n_925, n_927);
  nand g2704 (n_947, n_2539, n_2540, n_2541);
  xor g2705 (n_2542, n_928, n_929);
  xor g2706 (n_934, n_2542, n_930);
  nand g2707 (n_2543, n_928, n_929);
  nand g2708 (n_2544, n_930, n_929);
  nand g2709 (n_2545, n_928, n_930);
  nand g2710 (n_949, n_2543, n_2544, n_2545);
  xor g2711 (n_2546, n_931, n_932);
  xor g2712 (n_935, n_2546, n_933);
  nand g2713 (n_2547, n_931, n_932);
  nand g2714 (n_2548, n_933, n_932);
  nand g2715 (n_2549, n_931, n_933);
  nand g2716 (n_951, n_2547, n_2548, n_2549);
  xor g2717 (n_2550, n_934, n_935);
  xor g2718 (n_151, n_2550, n_936);
  nand g2719 (n_2551, n_934, n_935);
  nand g2720 (n_2552, n_936, n_935);
  nand g2721 (n_2553, n_934, n_936);
  nand g2722 (n_74, n_2551, n_2552, n_2553);
  xor g2725 (n_2554, A[53], A[41]);
  xor g2726 (n_943, n_2554, A[49]);
  nand g2727 (n_2555, A[53], A[41]);
  nand g2730 (n_954, n_2555, n_2491, n_2428);
  xor g2731 (n_2558, A[47], A[51]);
  xor g2732 (n_942, n_2558, A[45]);
  nand g2736 (n_953, n_2364, n_2301, n_2171);
  xor g2738 (n_944, n_2562, n_939);
  nand g2741 (n_2565, A[43], n_939);
  nand g2742 (n_958, n_2563, n_2564, n_2565);
  xor g2743 (n_2566, n_940, n_941);
  xor g2744 (n_946, n_2566, n_942);
  nand g2745 (n_2567, n_940, n_941);
  nand g2746 (n_2568, n_942, n_941);
  nand g2747 (n_2569, n_940, n_942);
  nand g2748 (n_960, n_2567, n_2568, n_2569);
  xor g2749 (n_2570, n_943, n_944);
  xor g2750 (n_948, n_2570, n_945);
  nand g2751 (n_2571, n_943, n_944);
  nand g2752 (n_2572, n_945, n_944);
  nand g2753 (n_2573, n_943, n_945);
  nand g2754 (n_961, n_2571, n_2572, n_2573);
  xor g2755 (n_2574, n_946, n_947);
  xor g2756 (n_950, n_2574, n_948);
  nand g2757 (n_2575, n_946, n_947);
  nand g2758 (n_2576, n_948, n_947);
  nand g2759 (n_2577, n_946, n_948);
  nand g2760 (n_964, n_2575, n_2576, n_2577);
  xor g2761 (n_2578, n_949, n_950);
  xor g2762 (n_150, n_2578, n_951);
  nand g2763 (n_2579, n_949, n_950);
  nand g2764 (n_2580, n_951, n_950);
  nand g2765 (n_2581, n_949, n_951);
  nand g2766 (n_73, n_2579, n_2580, n_2581);
  xor g2773 (n_2586, A[42], A[48]);
  xor g2774 (n_956, n_2586, A[52]);
  nand g2777 (n_2589, A[42], A[52]);
  nand g2778 (n_968, n_2205, n_2396, n_2589);
  xor g2780 (n_957, n_2138, A[55]);
  nand g2782 (n_2592, A[55], A[44]);
  nand g2783 (n_2593, A[46], A[55]);
  nand g2784 (n_971, n_2139, n_2592, n_2593);
  xor g2785 (n_2594, n_953, n_954);
  xor g2786 (n_959, n_2594, n_927);
  nand g2787 (n_2595, n_953, n_954);
  nand g2788 (n_2596, n_927, n_954);
  nand g2789 (n_2597, n_953, n_927);
  nand g2790 (n_973, n_2595, n_2596, n_2597);
  xor g2791 (n_2598, n_956, n_957);
  xor g2792 (n_962, n_2598, n_958);
  nand g2793 (n_2599, n_956, n_957);
  nand g2794 (n_2600, n_958, n_957);
  nand g2795 (n_2601, n_956, n_958);
  nand g2796 (n_975, n_2599, n_2600, n_2601);
  xor g2797 (n_2602, n_959, n_960);
  xor g2798 (n_963, n_2602, n_961);
  nand g2799 (n_2603, n_959, n_960);
  nand g2800 (n_2604, n_961, n_960);
  nand g2801 (n_2605, n_959, n_961);
  nand g2802 (n_977, n_2603, n_2604, n_2605);
  xor g2803 (n_2606, n_962, n_963);
  xor g2804 (n_149, n_2606, n_964);
  nand g2805 (n_2607, n_962, n_963);
  nand g2806 (n_2608, n_964, n_963);
  nand g2807 (n_2609, n_962, n_964);
  nand g2808 (n_148, n_2607, n_2608, n_2609);
  xor g2811 (n_2610, A[53], A[49]);
  xor g2812 (n_970, n_2610, A[47]);
  nand g2816 (n_979, n_2428, n_2235, n_2365);
  xor g2817 (n_2614, A[51], A[45]);
  xor g2818 (n_969, n_2614, A[43]);
  nand g2821 (n_2617, A[51], A[43]);
  nand g2822 (n_980, n_2301, n_2107, n_2617);
  xor g2824 (n_972, n_2618, n_968);
  nand g2826 (n_2620, n_968, n_939);
  nand g2828 (n_984, n_2564, n_2620, n_2621);
  xor g2829 (n_2622, n_969, n_970);
  xor g2830 (n_974, n_2622, n_971);
  nand g2831 (n_2623, n_969, n_970);
  nand g2832 (n_2624, n_971, n_970);
  nand g2833 (n_2625, n_969, n_971);
  nand g2834 (n_985, n_2623, n_2624, n_2625);
  xor g2835 (n_2626, n_972, n_973);
  xor g2836 (n_976, n_2626, n_974);
  nand g2837 (n_2627, n_972, n_973);
  nand g2838 (n_2628, n_974, n_973);
  nand g2839 (n_2629, n_972, n_974);
  nand g2840 (n_988, n_2627, n_2628, n_2629);
  xor g2841 (n_2630, n_975, n_976);
  xor g2842 (n_72, n_2630, n_977);
  nand g2843 (n_2631, n_975, n_976);
  nand g2844 (n_2632, n_977, n_976);
  nand g2845 (n_2633, n_975, n_977);
  nand g2846 (n_71, n_2631, n_2632, n_2633);
  xor g2859 (n_2642, A[44], A[55]);
  xor g2860 (n_983, n_2642, n_979);
  nand g2862 (n_2644, n_979, A[55]);
  nand g2863 (n_2645, A[44], n_979);
  nand g2864 (n_995, n_2592, n_2644, n_2645);
  xor g2865 (n_2646, n_980, n_894);
  xor g2866 (n_986, n_2646, n_927);
  nand g2867 (n_2647, n_980, n_894);
  nand g2868 (n_2648, n_927, n_894);
  nand g2869 (n_2649, n_980, n_927);
  nand g2870 (n_996, n_2647, n_2648, n_2649);
  xor g2871 (n_2650, n_983, n_984);
  xor g2872 (n_987, n_2650, n_985);
  nand g2873 (n_2651, n_983, n_984);
  nand g2874 (n_2652, n_985, n_984);
  nand g2875 (n_2653, n_983, n_985);
  nand g2876 (n_999, n_2651, n_2652, n_2653);
  xor g2877 (n_2654, n_986, n_987);
  xor g2878 (n_147, n_2654, n_988);
  nand g2879 (n_2655, n_986, n_987);
  nand g2880 (n_2656, n_988, n_987);
  nand g2881 (n_2657, n_986, n_988);
  nand g2882 (n_70, n_2655, n_2656, n_2657);
  xor g2886 (n_993, n_2234, A[55]);
  nand g2890 (n_1001, n_2235, n_2496, n_2429);
  nand g2896 (n_1004, n_2301, n_2664, n_2665);
  xor g2897 (n_2666, n_908, n_939);
  xor g2898 (n_997, n_2666, n_993);
  nand g2899 (n_2667, n_908, n_939);
  nand g2900 (n_2668, n_993, n_939);
  nand g2901 (n_2669, n_908, n_993);
  nand g2902 (n_1006, n_2667, n_2668, n_2669);
  xor g2903 (n_2670, n_994, n_995);
  xor g2904 (n_998, n_2670, n_996);
  nand g2905 (n_2671, n_994, n_995);
  nand g2906 (n_2672, n_996, n_995);
  nand g2907 (n_2673, n_994, n_996);
  nand g2908 (n_1008, n_2671, n_2672, n_2673);
  xor g2909 (n_2674, n_997, n_998);
  xor g2910 (n_146, n_2674, n_999);
  nand g2911 (n_2675, n_997, n_998);
  nand g2912 (n_2676, n_999, n_998);
  nand g2913 (n_2677, n_997, n_999);
  nand g2914 (n_69, n_2675, n_2676, n_2677);
  xor g2927 (n_2686, A[53], n_1001);
  xor g2928 (n_1005, n_2686, n_894);
  nand g2929 (n_2687, A[53], n_1001);
  nand g2930 (n_2688, n_894, n_1001);
  nand g2931 (n_2689, A[53], n_894);
  nand g2932 (n_1015, n_2687, n_2688, n_2689);
  xor g2933 (n_2690, n_927, n_1004);
  xor g2934 (n_1007, n_2690, n_1005);
  nand g2935 (n_2691, n_927, n_1004);
  nand g2936 (n_2692, n_1005, n_1004);
  nand g2937 (n_2693, n_927, n_1005);
  nand g2938 (n_1017, n_2691, n_2692, n_2693);
  xor g2939 (n_2694, n_1006, n_1007);
  xor g2940 (n_145, n_2694, n_1008);
  nand g2941 (n_2695, n_1006, n_1007);
  nand g2942 (n_2696, n_1008, n_1007);
  nand g2943 (n_2697, n_1006, n_1008);
  nand g2944 (n_68, n_2695, n_2696, n_2697);
  nand g2957 (n_2705, A[51], n_908);
  nand g2958 (n_1022, n_2664, n_2704, n_2705);
  xor g2959 (n_2706, n_939, n_993);
  xor g2960 (n_1016, n_2706, n_1014);
  nand g2962 (n_2708, n_1014, n_993);
  nand g2963 (n_2709, n_939, n_1014);
  nand g2964 (n_1024, n_2668, n_2708, n_2709);
  xor g2965 (n_2710, n_1015, n_1016);
  xor g2966 (n_144, n_2710, n_1017);
  nand g2967 (n_2711, n_1015, n_1016);
  nand g2968 (n_2712, n_1017, n_1016);
  nand g2969 (n_2713, n_1015, n_1017);
  nand g2970 (n_143, n_2711, n_2712, n_2713);
  xor g2978 (n_1021, n_2466, A[53]);
  nand g2980 (n_2720, A[53], A[52]);
  nand g2981 (n_2721, A[48], A[53]);
  nand g2982 (n_1029, n_2396, n_2720, n_2721);
  xor g2983 (n_2722, n_1001, n_927);
  xor g2984 (n_1023, n_2722, n_1021);
  nand g2985 (n_2723, n_1001, n_927);
  nand g2986 (n_2724, n_1021, n_927);
  nand g2987 (n_2725, n_1001, n_1021);
  nand g2988 (n_1031, n_2723, n_2724, n_2725);
  xor g2989 (n_2726, n_1022, n_1023);
  xor g2990 (n_67, n_2726, n_1024);
  nand g2991 (n_2727, n_1022, n_1023);
  nand g2992 (n_2728, n_1024, n_1023);
  nand g2993 (n_2729, n_1022, n_1024);
  nand g2994 (n_142, n_2727, n_2728, n_2729);
  xor g2998 (n_1028, n_2610, A[51]);
  nand g3002 (n_1033, n_2428, n_2363, n_2299);
  xor g3004 (n_1030, n_2618, n_1028);
  nand g3006 (n_2736, n_1028, n_939);
  nand g3008 (n_1036, n_2564, n_2736, n_2737);
  xor g3009 (n_2738, n_1029, n_1030);
  xor g3010 (n_66, n_2738, n_1031);
  nand g3011 (n_2739, n_1029, n_1030);
  nand g3012 (n_2740, n_1031, n_1030);
  nand g3013 (n_2741, n_1029, n_1031);
  nand g3014 (n_141, n_2739, n_2740, n_2741);
  xor g3021 (n_2746, A[52], A[55]);
  xor g3022 (n_1035, n_2746, n_1033);
  nand g3023 (n_2747, A[52], A[55]);
  nand g3024 (n_2748, n_1033, A[55]);
  nand g3025 (n_2749, A[52], n_1033);
  nand g3026 (n_1041, n_2747, n_2748, n_2749);
  xor g3027 (n_2750, n_927, n_1035);
  xor g3028 (n_65, n_2750, n_1036);
  nand g3029 (n_2751, n_927, n_1035);
  nand g3030 (n_2752, n_1036, n_1035);
  nand g3031 (n_2753, n_927, n_1036);
  nand g3032 (n_140, n_2751, n_2752, n_2753);
  nand g3040 (n_1044, n_2363, n_2756, n_2757);
  xor g3041 (n_2758, n_939, n_1040);
  xor g3042 (n_64, n_2758, n_1041);
  nand g3043 (n_2759, n_939, n_1040);
  nand g3044 (n_2760, n_1041, n_1040);
  nand g3045 (n_2761, n_939, n_1041);
  nand g3046 (n_139, n_2759, n_2760, n_2761);
  xor g3048 (n_1043, n_2522, A[52]);
  nand g3052 (n_1047, n_2523, n_2395, n_2531);
  xor g3053 (n_2766, A[55], n_1043);
  xor g3054 (n_63, n_2766, n_1044);
  nand g3055 (n_2767, A[55], n_1043);
  nand g3056 (n_2768, n_1044, n_1043);
  nand g3057 (n_2769, A[55], n_1044);
  nand g3058 (n_138, n_2767, n_2768, n_2769);
  nand g3065 (n_2773, A[55], n_1047);
  nand g3066 (n_137, n_2771, n_2772, n_2773);
  xor g3068 (n_61, n_2522, A[53]);
  nand g3070 (n_2776, A[53], A[54]);
  nand g3072 (n_136, n_2523, n_2776, n_2777);
  nor g11 (n_2793, A[0], A[2]);
  nand g12 (n_2788, A[0], A[2]);
  nor g13 (n_2789, A[1], A[3]);
  nor g15 (n_2799, A[2], n_205);
  nand g16 (n_2794, A[2], n_205);
  nor g17 (n_2795, n_128, n_204);
  nand g18 (n_2796, n_128, n_204);
  nor g19 (n_2805, n_127, n_203);
  nand g20 (n_2800, n_127, n_203);
  nor g21 (n_2801, n_126, n_202);
  nand g22 (n_2802, n_126, n_202);
  nor g23 (n_2811, n_125, n_201);
  nand g24 (n_2806, n_125, n_201);
  nor g25 (n_2807, n_124, n_200);
  nand g26 (n_2808, n_124, n_200);
  nor g27 (n_2817, n_123, n_199);
  nand g28 (n_2812, n_123, n_199);
  nor g29 (n_2813, n_122, n_198);
  nand g30 (n_2814, n_122, n_198);
  nor g31 (n_2823, n_121, n_197);
  nand g32 (n_2818, n_121, n_197);
  nor g33 (n_2819, n_120, n_196);
  nand g34 (n_2820, n_120, n_196);
  nor g35 (n_2829, n_119, n_195);
  nand g36 (n_2824, n_119, n_195);
  nor g37 (n_2825, n_118, n_194);
  nand g38 (n_2826, n_118, n_194);
  nor g39 (n_2835, n_117, n_193);
  nand g40 (n_2830, n_117, n_193);
  nor g41 (n_2831, n_116, n_192);
  nand g42 (n_2832, n_116, n_192);
  nor g43 (n_2841, n_115, n_191);
  nand g44 (n_2836, n_115, n_191);
  nor g45 (n_2837, n_114, n_190);
  nand g46 (n_2838, n_114, n_190);
  nor g47 (n_2847, n_113, n_189);
  nand g48 (n_2842, n_113, n_189);
  nor g49 (n_2843, n_112, n_188);
  nand g50 (n_2844, n_112, n_188);
  nor g51 (n_2853, n_111, n_187);
  nand g52 (n_2848, n_111, n_187);
  nor g53 (n_2849, n_110, n_186);
  nand g54 (n_2850, n_110, n_186);
  nor g55 (n_2859, n_109, n_185);
  nand g56 (n_2854, n_109, n_185);
  nor g57 (n_2855, n_108, n_184);
  nand g58 (n_2856, n_108, n_184);
  nor g59 (n_2865, n_107, n_183);
  nand g60 (n_2860, n_107, n_183);
  nor g61 (n_2861, n_106, n_182);
  nand g62 (n_2862, n_106, n_182);
  nor g63 (n_2871, n_105, n_181);
  nand g64 (n_2866, n_105, n_181);
  nor g65 (n_2867, n_104, n_180);
  nand g66 (n_2868, n_104, n_180);
  nor g67 (n_2877, n_103, n_179);
  nand g68 (n_2872, n_103, n_179);
  nor g69 (n_2873, n_102, n_178);
  nand g70 (n_2874, n_102, n_178);
  nor g71 (n_2883, n_101, n_177);
  nand g72 (n_2878, n_101, n_177);
  nor g73 (n_2879, n_100, n_176);
  nand g74 (n_2880, n_100, n_176);
  nor g75 (n_2889, n_99, n_175);
  nand g76 (n_2884, n_99, n_175);
  nor g77 (n_2885, n_98, n_174);
  nand g78 (n_2886, n_98, n_174);
  nor g79 (n_2895, n_97, n_173);
  nand g80 (n_2890, n_97, n_173);
  nor g81 (n_2891, n_96, n_172);
  nand g82 (n_2892, n_96, n_172);
  nor g83 (n_2901, n_95, n_171);
  nand g84 (n_2896, n_95, n_171);
  nor g85 (n_2897, n_94, n_170);
  nand g86 (n_2898, n_94, n_170);
  nor g87 (n_2907, n_93, n_169);
  nand g88 (n_2902, n_93, n_169);
  nor g89 (n_2903, n_92, n_168);
  nand g90 (n_2904, n_92, n_168);
  nor g91 (n_2913, n_91, n_167);
  nand g92 (n_2908, n_91, n_167);
  nor g93 (n_2909, n_90, n_166);
  nand g94 (n_2910, n_90, n_166);
  nor g95 (n_2919, n_89, n_165);
  nand g96 (n_2914, n_89, n_165);
  nor g97 (n_2915, n_88, n_164);
  nand g98 (n_2916, n_88, n_164);
  nor g99 (n_2925, n_87, n_163);
  nand g100 (n_2920, n_87, n_163);
  nor g101 (n_2921, n_86, n_162);
  nand g102 (n_2922, n_86, n_162);
  nor g103 (n_2931, n_85, n_161);
  nand g104 (n_2926, n_85, n_161);
  nor g105 (n_2927, n_84, n_160);
  nand g106 (n_2928, n_84, n_160);
  nor g107 (n_2937, n_83, n_159);
  nand g108 (n_2932, n_83, n_159);
  nor g109 (n_2933, n_82, n_158);
  nand g110 (n_2934, n_82, n_158);
  nor g111 (n_2943, n_81, n_157);
  nand g112 (n_2938, n_81, n_157);
  nor g113 (n_2939, n_80, n_156);
  nand g114 (n_2940, n_80, n_156);
  nor g115 (n_2949, n_79, n_155);
  nand g116 (n_2944, n_79, n_155);
  nor g117 (n_2945, n_78, n_154);
  nand g118 (n_2946, n_78, n_154);
  nor g119 (n_2955, n_77, n_153);
  nand g120 (n_2950, n_77, n_153);
  nor g121 (n_2951, n_76, n_152);
  nand g122 (n_2952, n_76, n_152);
  nor g123 (n_2961, n_75, n_151);
  nand g124 (n_2956, n_75, n_151);
  nor g125 (n_2957, n_74, n_150);
  nand g126 (n_2958, n_74, n_150);
  nor g127 (n_2967, n_73, n_149);
  nand g128 (n_2962, n_73, n_149);
  nor g129 (n_2963, n_72, n_148);
  nand g130 (n_2964, n_72, n_148);
  nor g131 (n_2973, n_71, n_147);
  nand g132 (n_2968, n_71, n_147);
  nor g133 (n_2969, n_70, n_146);
  nand g134 (n_2970, n_70, n_146);
  nor g135 (n_2979, n_69, n_145);
  nand g136 (n_2974, n_69, n_145);
  nor g137 (n_2975, n_68, n_144);
  nand g138 (n_2976, n_68, n_144);
  nor g139 (n_2985, n_67, n_143);
  nand g140 (n_2980, n_67, n_143);
  nor g141 (n_2981, n_66, n_142);
  nand g142 (n_2982, n_66, n_142);
  nor g143 (n_2991, n_65, n_141);
  nand g144 (n_2986, n_65, n_141);
  nor g145 (n_2987, n_64, n_140);
  nand g146 (n_2988, n_64, n_140);
  nor g147 (n_2997, n_63, n_139);
  nand g148 (n_2992, n_63, n_139);
  nor g149 (n_2993, n_62, n_138);
  nand g150 (n_2994, n_62, n_138);
  nor g151 (n_3003, n_61, n_137);
  nand g152 (n_2998, n_61, n_137);
  nor g162 (n_2791, n_2788, n_2789);
  nor g166 (n_2797, n_2794, n_2795);
  nor g169 (n_3018, n_2799, n_2795);
  nor g170 (n_2803, n_2800, n_2801);
  nor g173 (n_3012, n_2805, n_2801);
  nor g174 (n_2809, n_2806, n_2807);
  nor g177 (n_3025, n_2811, n_2807);
  nor g178 (n_2815, n_2812, n_2813);
  nor g181 (n_3019, n_2817, n_2813);
  nor g182 (n_2821, n_2818, n_2819);
  nor g185 (n_3032, n_2823, n_2819);
  nor g186 (n_2827, n_2824, n_2825);
  nor g189 (n_3026, n_2829, n_2825);
  nor g190 (n_2833, n_2830, n_2831);
  nor g193 (n_3039, n_2835, n_2831);
  nor g194 (n_2839, n_2836, n_2837);
  nor g197 (n_3033, n_2841, n_2837);
  nor g198 (n_2845, n_2842, n_2843);
  nor g201 (n_3046, n_2847, n_2843);
  nor g202 (n_2851, n_2848, n_2849);
  nor g205 (n_3040, n_2853, n_2849);
  nor g206 (n_2857, n_2854, n_2855);
  nor g209 (n_3053, n_2859, n_2855);
  nor g210 (n_2863, n_2860, n_2861);
  nor g213 (n_3047, n_2865, n_2861);
  nor g214 (n_2869, n_2866, n_2867);
  nor g217 (n_3060, n_2871, n_2867);
  nor g218 (n_2875, n_2872, n_2873);
  nor g221 (n_3054, n_2877, n_2873);
  nor g222 (n_2881, n_2878, n_2879);
  nor g225 (n_3067, n_2883, n_2879);
  nor g226 (n_2887, n_2884, n_2885);
  nor g229 (n_3061, n_2889, n_2885);
  nor g230 (n_2893, n_2890, n_2891);
  nor g233 (n_3074, n_2895, n_2891);
  nor g234 (n_2899, n_2896, n_2897);
  nor g237 (n_3068, n_2901, n_2897);
  nor g238 (n_2905, n_2902, n_2903);
  nor g241 (n_3081, n_2907, n_2903);
  nor g242 (n_2911, n_2908, n_2909);
  nor g245 (n_3075, n_2913, n_2909);
  nor g246 (n_2917, n_2914, n_2915);
  nor g249 (n_3088, n_2919, n_2915);
  nor g250 (n_2923, n_2920, n_2921);
  nor g253 (n_3082, n_2925, n_2921);
  nor g254 (n_2929, n_2926, n_2927);
  nor g257 (n_3095, n_2931, n_2927);
  nor g258 (n_2935, n_2932, n_2933);
  nor g261 (n_3089, n_2937, n_2933);
  nor g262 (n_2941, n_2938, n_2939);
  nor g265 (n_3102, n_2943, n_2939);
  nor g266 (n_2947, n_2944, n_2945);
  nor g269 (n_3096, n_2949, n_2945);
  nor g270 (n_2953, n_2950, n_2951);
  nor g273 (n_3109, n_2955, n_2951);
  nor g274 (n_2959, n_2956, n_2957);
  nor g277 (n_3103, n_2961, n_2957);
  nor g278 (n_2965, n_2962, n_2963);
  nor g281 (n_3116, n_2967, n_2963);
  nor g282 (n_2971, n_2968, n_2969);
  nor g285 (n_3110, n_2973, n_2969);
  nor g286 (n_2977, n_2974, n_2975);
  nor g289 (n_3123, n_2979, n_2975);
  nor g290 (n_2983, n_2980, n_2981);
  nor g293 (n_3117, n_2985, n_2981);
  nor g294 (n_2989, n_2986, n_2987);
  nor g297 (n_3130, n_2991, n_2987);
  nor g298 (n_2995, n_2992, n_2993);
  nor g301 (n_3124, n_2997, n_2993);
  nor g302 (n_3001, n_2998, n_2999);
  nor g305 (n_3132, n_3003, n_2999);
  nand g316 (n_3133, n_3018, n_3012);
  nand g321 (n_3143, n_3025, n_3019);
  nand g326 (n_3138, n_3032, n_3026);
  nand g331 (n_3149, n_3039, n_3033);
  nand g336 (n_3144, n_3046, n_3040);
  nand g341 (n_3155, n_3053, n_3047);
  nand g346 (n_3150, n_3060, n_3054);
  nand g351 (n_3161, n_3067, n_3061);
  nand g356 (n_3156, n_3074, n_3068);
  nand g361 (n_3167, n_3081, n_3075);
  nand g366 (n_3162, n_3088, n_3082);
  nand g371 (n_3173, n_3095, n_3089);
  nand g376 (n_3168, n_3102, n_3096);
  nand g381 (n_3179, n_3109, n_3103);
  nand g386 (n_3174, n_3116, n_3110);
  nand g391 (n_3185, n_3123, n_3117);
  nand g396 (n_3180, n_3130, n_3124);
  nand g404 (n_3187, n_3136, n_3137);
  nor g405 (n_3141, n_3138, n_3139);
  nor g408 (n_3186, n_3143, n_3138);
  nor g409 (n_3147, n_3144, n_3145);
  nor g412 (n_3196, n_3149, n_3144);
  nor g413 (n_3153, n_3150, n_3151);
  nor g416 (n_3190, n_3155, n_3150);
  nor g417 (n_3159, n_3156, n_3157);
  nor g420 (n_3203, n_3161, n_3156);
  nor g421 (n_3165, n_3162, n_3163);
  nor g424 (n_3197, n_3167, n_3162);
  nor g425 (n_3171, n_3168, n_3169);
  nor g428 (n_3210, n_3173, n_3168);
  nor g429 (n_3177, n_3174, n_3175);
  nor g432 (n_3204, n_3179, n_3174);
  nor g433 (n_3183, n_3180, n_3181);
  nor g436 (n_3232, n_3185, n_3180);
  nand g437 (n_3189, n_3186, n_3187);
  nand g438 (n_3212, n_3188, n_3189);
  nand g443 (n_3211, n_3196, n_3190);
  nand g448 (n_3221, n_3203, n_3197);
  nand g3081 (n_3216, n_3210, n_3204);
  nand g3084 (n_3223, n_3214, n_3215);
  nor g3085 (n_3219, n_3216, n_3217);
  nor g3088 (n_3222, n_3221, n_3216);
  nand g3089 (n_3225, n_3222, n_3223);
  nand g3090 (n_3233, n_3224, n_3225);
  nand g3093 (n_3230, n_3217, n_3227);
  nand g3094 (n_3228, n_3196, n_3212);
  nand g3095 (n_3240, n_3191, n_3228);
  nand g3096 (n_3229, n_3203, n_3223);
  nand g3097 (n_3245, n_3198, n_3229);
  nand g3098 (n_3231, n_3210, n_3230);
  nand g3099 (n_3250, n_3205, n_3231);
  nand g3100 (n_3235, n_3232, n_3233);
  nand g3101 (n_3255, n_3234, n_3235);
  nand g3104 (n_3258, n_3139, n_3237);
  nand g3107 (n_3261, n_3145, n_3239);
  nand g3110 (n_3264, n_3151, n_3242);
  nand g3113 (n_3267, n_3157, n_3244);
  nand g3116 (n_3270, n_3163, n_3247);
  nand g3119 (n_3273, n_3169, n_3249);
  nand g3122 (n_3276, n_3175, n_3252);
  nand g3125 (n_3279, n_3181, n_3254);
  nand g3127 (n_3286, n_3013, n_3256);
  nand g3128 (n_3257, n_3025, n_3187);
  nand g3129 (n_3291, n_3020, n_3257);
  nand g3130 (n_3259, n_3032, n_3258);
  nand g3131 (n_3296, n_3027, n_3259);
  nand g3132 (n_3260, n_3039, n_3212);
  nand g3133 (n_3301, n_3034, n_3260);
  nand g3134 (n_3262, n_3046, n_3261);
  nand g3135 (n_3306, n_3041, n_3262);
  nand g3136 (n_3263, n_3053, n_3240);
  nand g3137 (n_3311, n_3048, n_3263);
  nand g3138 (n_3265, n_3060, n_3264);
  nand g3139 (n_3316, n_3055, n_3265);
  nand g3140 (n_3266, n_3067, n_3223);
  nand g3141 (n_3321, n_3062, n_3266);
  nand g3142 (n_3268, n_3074, n_3267);
  nand g3143 (n_3326, n_3069, n_3268);
  nand g3144 (n_3269, n_3081, n_3245);
  nand g3145 (n_3331, n_3076, n_3269);
  nand g3146 (n_3271, n_3088, n_3270);
  nand g3147 (n_3336, n_3083, n_3271);
  nand g3148 (n_3272, n_3095, n_3230);
  nand g3149 (n_3341, n_3090, n_3272);
  nand g3150 (n_3274, n_3102, n_3273);
  nand g3151 (n_3346, n_3097, n_3274);
  nand g3152 (n_3275, n_3109, n_3250);
  nand g3153 (n_3351, n_3104, n_3275);
  nand g3154 (n_3277, n_3116, n_3276);
  nand g3155 (n_3356, n_3111, n_3277);
  nand g3156 (n_3278, n_3123, n_3233);
  nand g3157 (n_3361, n_3118, n_3278);
  nand g3158 (n_3280, n_3130, n_3279);
  nand g3159 (n_3366, n_3125, n_3280);
  nand g3160 (n_3281, n_3132, n_3255);
  nand g3161 (n_3371, n_3131, n_3281);
  nand g3167 (n_3381, n_2794, n_3285);
  nand g3170 (n_3385, n_2800, n_3288);
  nand g3173 (n_3389, n_2806, n_3290);
  nand g3176 (n_3393, n_2812, n_3293);
  nand g3179 (n_3397, n_2818, n_3295);
  nand g3182 (n_3401, n_2824, n_3298);
  nand g3185 (n_3405, n_2830, n_3300);
  nand g3188 (n_3409, n_2836, n_3303);
  nand g3191 (n_3413, n_2842, n_3305);
  nand g3194 (n_3417, n_2848, n_3308);
  nand g3197 (n_3421, n_2854, n_3310);
  nand g3200 (n_3425, n_2860, n_3313);
  nand g3203 (n_3429, n_2866, n_3315);
  nand g3206 (n_3433, n_2872, n_3318);
  nand g3209 (n_3437, n_2878, n_3320);
  nand g3212 (n_3441, n_2884, n_3323);
  nand g3215 (n_3445, n_2890, n_3325);
  nand g3218 (n_3449, n_2896, n_3328);
  nand g3221 (n_3453, n_2902, n_3330);
  nand g3224 (n_3457, n_2908, n_3333);
  nand g3227 (n_3461, n_2914, n_3335);
  nand g3230 (n_3465, n_2920, n_3338);
  nand g3233 (n_3469, n_2926, n_3340);
  nand g3236 (n_3473, n_2932, n_3343);
  nand g3239 (n_3477, n_2938, n_3345);
  nand g3242 (n_3481, n_2944, n_3348);
  nand g3245 (n_3485, n_2950, n_3350);
  nand g3248 (n_3489, n_2956, n_3353);
  nand g3251 (n_3493, n_2962, n_3355);
  nand g3254 (n_3497, n_2968, n_3358);
  nand g3257 (n_3501, n_2974, n_3360);
  nand g3260 (n_3505, n_2980, n_3363);
  nand g3263 (n_3509, n_2986, n_3365);
  nand g3266 (n_3513, n_2992, n_3368);
  nand g3269 (n_3517, n_2998, n_3370);
  nand g3272 (n_3521, n_3004, n_3373);
  xnor g3284 (Z[5], n_3381, n_3382);
  xnor g3286 (Z[6], n_3286, n_3383);
  xnor g3289 (Z[7], n_3385, n_3386);
  xnor g3291 (Z[8], n_3187, n_3387);
  xnor g3294 (Z[9], n_3389, n_3390);
  xnor g3296 (Z[10], n_3291, n_3391);
  xnor g3299 (Z[11], n_3393, n_3394);
  xnor g3301 (Z[12], n_3258, n_3395);
  xnor g3304 (Z[13], n_3397, n_3398);
  xnor g3306 (Z[14], n_3296, n_3399);
  xnor g3309 (Z[15], n_3401, n_3402);
  xnor g3311 (Z[16], n_3212, n_3403);
  xnor g3314 (Z[17], n_3405, n_3406);
  xnor g3316 (Z[18], n_3301, n_3407);
  xnor g3319 (Z[19], n_3409, n_3410);
  xnor g3321 (Z[20], n_3261, n_3411);
  xnor g3324 (Z[21], n_3413, n_3414);
  xnor g3326 (Z[22], n_3306, n_3415);
  xnor g3329 (Z[23], n_3417, n_3418);
  xnor g3331 (Z[24], n_3240, n_3419);
  xnor g3334 (Z[25], n_3421, n_3422);
  xnor g3336 (Z[26], n_3311, n_3423);
  xnor g3339 (Z[27], n_3425, n_3426);
  xnor g3341 (Z[28], n_3264, n_3427);
  xnor g3344 (Z[29], n_3429, n_3430);
  xnor g3346 (Z[30], n_3316, n_3431);
  xnor g3349 (Z[31], n_3433, n_3434);
  xnor g3351 (Z[32], n_3223, n_3435);
  xnor g3354 (Z[33], n_3437, n_3438);
  xnor g3356 (Z[34], n_3321, n_3439);
  xnor g3359 (Z[35], n_3441, n_3442);
  xnor g3361 (Z[36], n_3267, n_3443);
  xnor g3364 (Z[37], n_3445, n_3446);
  xnor g3366 (Z[38], n_3326, n_3447);
  xnor g3369 (Z[39], n_3449, n_3450);
  xnor g3371 (Z[40], n_3245, n_3451);
  xnor g3374 (Z[41], n_3453, n_3454);
  xnor g3376 (Z[42], n_3331, n_3455);
  xnor g3379 (Z[43], n_3457, n_3458);
  xnor g3381 (Z[44], n_3270, n_3459);
  xnor g3384 (Z[45], n_3461, n_3462);
  xnor g3386 (Z[46], n_3336, n_3463);
  xnor g3389 (Z[47], n_3465, n_3466);
  xnor g3391 (Z[48], n_3230, n_3467);
  xnor g3394 (Z[49], n_3469, n_3470);
  xnor g3396 (Z[50], n_3341, n_3471);
  xnor g3399 (Z[51], n_3473, n_3474);
  xnor g3401 (Z[52], n_3273, n_3475);
  xnor g3404 (Z[53], n_3477, n_3478);
  xnor g3406 (Z[54], n_3346, n_3479);
  xnor g3409 (Z[55], n_3481, n_3482);
  xnor g3411 (Z[56], n_3250, n_3483);
  xnor g3414 (Z[57], n_3485, n_3486);
  xnor g3416 (Z[58], n_3351, n_3487);
  xnor g3419 (Z[59], n_3489, n_3490);
  xnor g3421 (Z[60], n_3276, n_3491);
  xnor g3424 (Z[61], n_3493, n_3494);
  xnor g3426 (Z[62], n_3356, n_3495);
  xnor g3429 (Z[63], n_3497, n_3498);
  xnor g3431 (Z[64], n_3233, n_3499);
  xnor g3434 (Z[65], n_3501, n_3502);
  xnor g3436 (Z[66], n_3361, n_3503);
  xnor g3439 (Z[67], n_3505, n_3506);
  xnor g3441 (Z[68], n_3279, n_3507);
  xnor g3444 (Z[69], n_3509, n_3510);
  xnor g3446 (Z[70], n_3366, n_3511);
  xnor g3449 (Z[71], n_3513, n_3514);
  xnor g3451 (Z[72], n_3255, n_3515);
  xnor g3454 (Z[73], n_3517, n_3518);
  xnor g3456 (Z[74], n_3371, n_3519);
  xnor g3464 (n_2522, A[56], A[54]);
  or g3465 (n_2523, wc, A[56]);
  not gc (wc, A[54]);
  or g3466 (n_2525, wc0, A[56]);
  not gc0 (wc0, A[50]);
  xnor g3467 (n_2562, A[55], A[43]);
  or g3468 (n_2563, wc1, A[55]);
  not gc1 (wc1, A[43]);
  xnor g3469 (n_994, n_2614, A[53]);
  or g3470 (n_2664, wc2, A[53]);
  not gc2 (wc2, A[51]);
  or g3471 (n_2665, wc3, A[53]);
  not gc3 (wc3, A[45]);
  xnor g3473 (n_1040, n_2362, A[55]);
  or g3474 (n_2756, wc4, A[55]);
  not gc4 (wc4, A[51]);
  or g3475 (n_2757, wc5, A[55]);
  not gc5 (wc5, A[53]);
  or g3476 (n_2531, wc6, A[56]);
  not gc6 (wc6, A[52]);
  or g3478 (n_2771, A[53], wc7);
  not gc7 (wc7, A[55]);
  or g3479 (n_2777, wc8, A[56]);
  not gc8 (wc8, A[53]);
  and g3480 (n_3007, wc9, A[56]);
  not gc9 (wc9, A[55]);
  or g3481 (n_3004, wc10, A[56]);
  not gc10 (wc10, A[55]);
  or g3482 (n_2621, A[55], wc11);
  not gc11 (wc11, n_968);
  xnor g3483 (n_1014, n_2362, n_908);
  or g3484 (n_2704, A[53], wc12);
  not gc12 (wc12, n_908);
  or g3485 (n_2737, A[55], wc13);
  not gc13 (wc13, n_1028);
  and g3486 (n_3010, wc14, n_1051);
  not gc14 (wc14, n_2791);
  or g3488 (n_3375, wc15, n_2793);
  not gc15 (wc15, n_2788);
  or g3489 (n_3378, n_2789, wc16);
  not gc16 (wc16, n_1051);
  xnor g3490 (n_2530, A[56], A[52]);
  or g3491 (n_2533, wc17, A[56]);
  not gc17 (wc17, A[46]);
  or g3492 (n_2564, A[55], wc18);
  not gc18 (wc18, n_939);
  xnor g3493 (n_2618, n_939, A[55]);
  xnor g3494 (n_62, n_2426, n_1047);
  or g3495 (n_2772, A[53], wc19);
  not gc19 (wc19, n_1047);
  and g3496 (n_2999, A[55], wc20);
  not gc20 (wc20, n_136);
  or g3497 (n_3000, A[55], wc21);
  not gc21 (wc21, n_136);
  or g3498 (n_3379, wc22, n_2799);
  not gc22 (wc22, n_2794);
  or g3499 (n_3519, wc23, n_3007);
  not gc23 (wc23, n_3004);
  and g3500 (n_3013, wc24, n_2796);
  not gc24 (wc24, n_2797);
  not g3501 (Z[2], n_3375);
  or g3502 (n_3382, wc25, n_2795);
  not gc25 (wc25, n_2796);
  or g3503 (n_3383, wc26, n_2805);
  not gc26 (wc26, n_2800);
  and g3504 (n_3015, wc27, n_2802);
  not gc27 (wc27, n_2803);
  or g3507 (n_3386, wc28, n_2801);
  not gc28 (wc28, n_2802);
  or g3508 (n_3518, wc29, n_2999);
  not gc29 (wc29, n_3000);
  and g3509 (n_3020, wc30, n_2808);
  not gc30 (wc30, n_2809);
  and g3510 (n_3016, wc31, n_3012);
  not gc31 (wc31, n_3013);
  or g3511 (n_3256, n_3010, wc32);
  not gc32 (wc32, n_3018);
  or g3512 (n_3285, n_2799, n_3010);
  xor g3513 (Z[3], n_2788, n_3378);
  xor g3514 (Z[4], n_3010, n_3379);
  or g3515 (n_3387, wc33, n_2811);
  not gc33 (wc33, n_2806);
  or g3516 (n_3390, wc34, n_2807);
  not gc34 (wc34, n_2808);
  and g3517 (n_3131, n_3000, wc35);
  not gc35 (wc35, n_3001);
  and g3518 (n_3136, wc36, n_3015);
  not gc36 (wc36, n_3016);
  or g3519 (n_3137, n_3133, n_3010);
  or g3520 (n_3391, wc37, n_2817);
  not gc37 (wc37, n_2812);
  or g3521 (n_3514, wc38, n_2993);
  not gc38 (wc38, n_2994);
  or g3522 (n_3515, wc39, n_3003);
  not gc39 (wc39, n_2998);
  and g3523 (n_3022, wc40, n_2814);
  not gc40 (wc40, n_2815);
  and g3524 (n_3027, wc41, n_2820);
  not gc41 (wc41, n_2821);
  and g3525 (n_3127, wc42, n_2994);
  not gc42 (wc42, n_2995);
  or g3526 (n_3288, wc43, n_2805);
  not gc43 (wc43, n_3286);
  or g3527 (n_3394, wc44, n_2813);
  not gc44 (wc44, n_2814);
  or g3528 (n_3395, wc45, n_2823);
  not gc45 (wc45, n_2818);
  or g3529 (n_3398, wc46, n_2819);
  not gc46 (wc46, n_2820);
  or g3530 (n_3511, wc47, n_2997);
  not gc47 (wc47, n_2992);
  and g3531 (n_3029, wc48, n_2826);
  not gc48 (wc48, n_2827);
  and g3532 (n_3125, wc49, n_2988);
  not gc49 (wc49, n_2989);
  and g3533 (n_3023, wc50, n_3019);
  not gc50 (wc50, n_3020);
  or g3534 (n_3290, wc51, n_2811);
  not gc51 (wc51, n_3187);
  or g3535 (n_3399, wc52, n_2829);
  not gc52 (wc52, n_2824);
  or g3536 (n_3402, wc53, n_2825);
  not gc53 (wc53, n_2826);
  or g3537 (n_3506, wc54, n_2981);
  not gc54 (wc54, n_2982);
  or g3538 (n_3507, wc55, n_2991);
  not gc55 (wc55, n_2986);
  or g3539 (n_3510, wc56, n_2987);
  not gc56 (wc56, n_2988);
  and g3540 (n_3034, wc57, n_2832);
  not gc57 (wc57, n_2833);
  and g3541 (n_3036, wc58, n_2838);
  not gc58 (wc58, n_2839);
  and g3542 (n_3120, wc59, n_2982);
  not gc59 (wc59, n_2983);
  and g3543 (n_3139, wc60, n_3022);
  not gc60 (wc60, n_3023);
  and g3544 (n_3030, wc61, n_3026);
  not gc61 (wc61, n_3027);
  and g3545 (n_3128, wc62, n_3124);
  not gc62 (wc62, n_3125);
  or g3546 (n_3237, wc63, n_3143);
  not gc63 (wc63, n_3187);
  or g3547 (n_3403, wc64, n_2835);
  not gc64 (wc64, n_2830);
  or g3548 (n_3406, wc65, n_2831);
  not gc65 (wc65, n_2832);
  or g3549 (n_3407, wc66, n_2841);
  not gc66 (wc66, n_2836);
  or g3550 (n_3410, wc67, n_2837);
  not gc67 (wc67, n_2838);
  or g3551 (n_3411, wc68, n_2847);
  not gc68 (wc68, n_2842);
  or g3552 (n_3503, wc69, n_2985);
  not gc69 (wc69, n_2980);
  and g3553 (n_3041, wc70, n_2844);
  not gc70 (wc70, n_2845);
  and g3554 (n_3118, wc71, n_2976);
  not gc71 (wc71, n_2977);
  and g3555 (n_3140, wc72, n_3029);
  not gc72 (wc72, n_3030);
  and g3556 (n_3037, wc73, n_3033);
  not gc73 (wc73, n_3034);
  and g3557 (n_3182, wc74, n_3127);
  not gc74 (wc74, n_3128);
  or g3558 (n_3293, wc75, n_2817);
  not gc75 (wc75, n_3291);
  or g3559 (n_3414, wc76, n_2843);
  not gc76 (wc76, n_2844);
  or g3560 (n_3415, wc77, n_2853);
  not gc77 (wc77, n_2848);
  or g3561 (n_3498, wc78, n_2969);
  not gc78 (wc78, n_2970);
  or g3562 (n_3499, wc79, n_2979);
  not gc79 (wc79, n_2974);
  or g3563 (n_3502, wc80, n_2975);
  not gc80 (wc80, n_2976);
  and g3564 (n_3043, wc81, n_2850);
  not gc81 (wc81, n_2851);
  and g3565 (n_3048, wc82, n_2856);
  not gc82 (wc82, n_2857);
  and g3566 (n_3050, wc83, n_2862);
  not gc83 (wc83, n_2863);
  and g3567 (n_3055, wc84, n_2868);
  not gc84 (wc84, n_2869);
  and g3568 (n_3057, wc85, n_2874);
  not gc85 (wc85, n_2875);
  and g3569 (n_3062, wc86, n_2880);
  not gc86 (wc86, n_2881);
  and g3570 (n_3064, wc87, n_2886);
  not gc87 (wc87, n_2887);
  and g3571 (n_3069, wc88, n_2892);
  not gc88 (wc88, n_2893);
  and g3572 (n_3071, wc89, n_2898);
  not gc89 (wc89, n_2899);
  and g3573 (n_3076, wc90, n_2904);
  not gc90 (wc90, n_2905);
  and g3574 (n_3078, wc91, n_2910);
  not gc91 (wc91, n_2911);
  and g3575 (n_3083, wc92, n_2916);
  not gc92 (wc92, n_2917);
  and g3576 (n_3085, wc93, n_2922);
  not gc93 (wc93, n_2923);
  and g3577 (n_3090, wc94, n_2928);
  not gc94 (wc94, n_2929);
  and g3578 (n_3092, wc95, n_2934);
  not gc95 (wc95, n_2935);
  and g3579 (n_3097, wc96, n_2940);
  not gc96 (wc96, n_2941);
  and g3580 (n_3099, wc97, n_2946);
  not gc97 (wc97, n_2947);
  and g3581 (n_3104, wc98, n_2952);
  not gc98 (wc98, n_2953);
  and g3582 (n_3145, wc99, n_3036);
  not gc99 (wc99, n_3037);
  and g3583 (n_3121, wc100, n_3117);
  not gc100 (wc100, n_3118);
  or g3584 (n_3295, wc101, n_2823);
  not gc101 (wc101, n_3258);
  or g3585 (n_3418, wc102, n_2849);
  not gc102 (wc102, n_2850);
  or g3586 (n_3419, wc103, n_2859);
  not gc103 (wc103, n_2854);
  or g3587 (n_3422, wc104, n_2855);
  not gc104 (wc104, n_2856);
  or g3588 (n_3423, wc105, n_2865);
  not gc105 (wc105, n_2860);
  or g3589 (n_3426, wc106, n_2861);
  not gc106 (wc106, n_2862);
  or g3590 (n_3427, wc107, n_2871);
  not gc107 (wc107, n_2866);
  or g3591 (n_3430, wc108, n_2867);
  not gc108 (wc108, n_2868);
  or g3592 (n_3431, wc109, n_2877);
  not gc109 (wc109, n_2872);
  or g3593 (n_3434, wc110, n_2873);
  not gc110 (wc110, n_2874);
  or g3594 (n_3435, wc111, n_2883);
  not gc111 (wc111, n_2878);
  or g3595 (n_3438, wc112, n_2879);
  not gc112 (wc112, n_2880);
  or g3596 (n_3439, wc113, n_2889);
  not gc113 (wc113, n_2884);
  or g3597 (n_3442, wc114, n_2885);
  not gc114 (wc114, n_2886);
  or g3598 (n_3443, wc115, n_2895);
  not gc115 (wc115, n_2890);
  or g3599 (n_3446, wc116, n_2891);
  not gc116 (wc116, n_2892);
  or g3600 (n_3447, wc117, n_2901);
  not gc117 (wc117, n_2896);
  or g3601 (n_3450, wc118, n_2897);
  not gc118 (wc118, n_2898);
  or g3602 (n_3451, wc119, n_2907);
  not gc119 (wc119, n_2902);
  or g3603 (n_3454, wc120, n_2903);
  not gc120 (wc120, n_2904);
  or g3604 (n_3455, wc121, n_2913);
  not gc121 (wc121, n_2908);
  or g3605 (n_3458, wc122, n_2909);
  not gc122 (wc122, n_2910);
  or g3606 (n_3459, wc123, n_2919);
  not gc123 (wc123, n_2914);
  or g3607 (n_3462, wc124, n_2915);
  not gc124 (wc124, n_2916);
  or g3608 (n_3463, wc125, n_2925);
  not gc125 (wc125, n_2920);
  or g3609 (n_3466, wc126, n_2921);
  not gc126 (wc126, n_2922);
  or g3610 (n_3467, wc127, n_2931);
  not gc127 (wc127, n_2926);
  or g3611 (n_3470, wc128, n_2927);
  not gc128 (wc128, n_2928);
  or g3612 (n_3471, wc129, n_2937);
  not gc129 (wc129, n_2932);
  or g3613 (n_3474, wc130, n_2933);
  not gc130 (wc130, n_2934);
  or g3614 (n_3475, wc131, n_2943);
  not gc131 (wc131, n_2938);
  or g3615 (n_3478, wc132, n_2939);
  not gc132 (wc132, n_2940);
  or g3616 (n_3479, wc133, n_2949);
  not gc133 (wc133, n_2944);
  or g3617 (n_3482, wc134, n_2945);
  not gc134 (wc134, n_2946);
  or g3618 (n_3483, wc135, n_2955);
  not gc135 (wc135, n_2950);
  or g3619 (n_3486, wc136, n_2951);
  not gc136 (wc136, n_2952);
  and g3620 (n_3106, wc137, n_2958);
  not gc137 (wc137, n_2959);
  and g3621 (n_3044, wc138, n_3040);
  not gc138 (wc138, n_3041);
  and g3622 (n_3051, wc139, n_3047);
  not gc139 (wc139, n_3048);
  and g3623 (n_3058, wc140, n_3054);
  not gc140 (wc140, n_3055);
  and g3624 (n_3065, wc141, n_3061);
  not gc141 (wc141, n_3062);
  and g3625 (n_3072, wc142, n_3068);
  not gc142 (wc142, n_3069);
  and g3626 (n_3079, wc143, n_3075);
  not gc143 (wc143, n_3076);
  and g3627 (n_3086, wc144, n_3082);
  not gc144 (wc144, n_3083);
  and g3628 (n_3093, wc145, n_3089);
  not gc145 (wc145, n_3090);
  and g3629 (n_3100, wc146, n_3096);
  not gc146 (wc146, n_3097);
  and g3630 (n_3181, wc147, n_3120);
  not gc147 (wc147, n_3121);
  and g3631 (n_3188, n_3140, wc148);
  not gc148 (wc148, n_3141);
  or g3632 (n_3487, wc149, n_2961);
  not gc149 (wc149, n_2956);
  or g3633 (n_3490, wc150, n_2957);
  not gc150 (wc150, n_2958);
  and g3634 (n_3111, wc151, n_2964);
  not gc151 (wc151, n_2965);
  and g3635 (n_3146, wc152, n_3043);
  not gc152 (wc152, n_3044);
  and g3636 (n_3151, wc153, n_3050);
  not gc153 (wc153, n_3051);
  and g3637 (n_3152, wc154, n_3057);
  not gc154 (wc154, n_3058);
  and g3638 (n_3157, wc155, n_3064);
  not gc155 (wc155, n_3065);
  and g3639 (n_3158, wc156, n_3071);
  not gc156 (wc156, n_3072);
  and g3640 (n_3163, wc157, n_3078);
  not gc157 (wc157, n_3079);
  and g3641 (n_3164, wc158, n_3085);
  not gc158 (wc158, n_3086);
  and g3642 (n_3169, wc159, n_3092);
  not gc159 (wc159, n_3093);
  and g3643 (n_3170, wc160, n_3099);
  not gc160 (wc160, n_3100);
  and g3644 (n_3107, wc161, n_3103);
  not gc161 (wc161, n_3104);
  or g3645 (n_3298, wc162, n_2829);
  not gc162 (wc162, n_3296);
  or g3646 (n_3491, wc163, n_2967);
  not gc163 (wc163, n_2962);
  or g3647 (n_3494, wc164, n_2963);
  not gc164 (wc164, n_2964);
  and g3648 (n_3113, wc165, n_2970);
  not gc165 (wc165, n_2971);
  and g3649 (n_3175, wc166, n_3106);
  not gc166 (wc166, n_3107);
  and g3650 (n_3234, n_3182, wc167);
  not gc167 (wc167, n_3183);
  or g3651 (n_3239, wc168, n_3149);
  not gc168 (wc168, n_3212);
  or g3652 (n_3300, wc169, n_2835);
  not gc169 (wc169, n_3212);
  or g3653 (n_3495, wc170, n_2973);
  not gc170 (wc170, n_2968);
  and g3654 (n_3114, wc171, n_3110);
  not gc171 (wc171, n_3111);
  and g3655 (n_3191, n_3146, wc172);
  not gc172 (wc172, n_3147);
  and g3656 (n_3193, n_3152, wc173);
  not gc173 (wc173, n_3153);
  and g3657 (n_3198, n_3158, wc174);
  not gc174 (wc174, n_3159);
  and g3658 (n_3200, n_3164, wc175);
  not gc175 (wc175, n_3165);
  and g3659 (n_3205, n_3170, wc176);
  not gc176 (wc176, n_3171);
  or g3660 (n_3215, n_3211, wc177);
  not gc177 (wc177, n_3212);
  and g3661 (n_3176, wc178, n_3113);
  not gc178 (wc178, n_3114);
  and g3662 (n_3194, wc179, n_3190);
  not gc179 (wc179, n_3191);
  and g3663 (n_3201, wc180, n_3197);
  not gc180 (wc180, n_3198);
  or g3664 (n_3303, wc181, n_2841);
  not gc181 (wc181, n_3301);
  or g3665 (n_3305, wc182, n_2847);
  not gc182 (wc182, n_3261);
  and g3666 (n_3214, wc183, n_3193);
  not gc183 (wc183, n_3194);
  and g3667 (n_3217, wc184, n_3200);
  not gc184 (wc184, n_3201);
  and g3668 (n_3208, wc185, n_3204);
  not gc185 (wc185, n_3205);
  or g3669 (n_3242, wc186, n_3155);
  not gc186 (wc186, n_3240);
  or g3670 (n_3310, wc187, n_2859);
  not gc187 (wc187, n_3240);
  and g3671 (n_3207, n_3176, wc188);
  not gc188 (wc188, n_3177);
  or g3672 (n_3308, wc189, n_2853);
  not gc189 (wc189, n_3306);
  or g3673 (n_3227, wc190, n_3221);
  not gc190 (wc190, n_3223);
  or g3674 (n_3244, wc191, n_3161);
  not gc191 (wc191, n_3223);
  or g3675 (n_3313, wc192, n_2865);
  not gc192 (wc192, n_3311);
  or g3676 (n_3315, wc193, n_2871);
  not gc193 (wc193, n_3264);
  or g3677 (n_3320, wc194, n_2883);
  not gc194 (wc194, n_3223);
  and g3678 (n_3218, n_3207, wc195);
  not gc195 (wc195, n_3208);
  or g3679 (n_3247, wc196, n_3167);
  not gc196 (wc196, n_3245);
  or g3680 (n_3249, wc197, n_3173);
  not gc197 (wc197, n_3230);
  or g3681 (n_3318, wc198, n_2877);
  not gc198 (wc198, n_3316);
  or g3682 (n_3323, wc199, n_2889);
  not gc199 (wc199, n_3321);
  or g3683 (n_3325, wc200, n_2895);
  not gc200 (wc200, n_3267);
  or g3684 (n_3330, wc201, n_2907);
  not gc201 (wc201, n_3245);
  or g3685 (n_3340, wc202, n_2931);
  not gc202 (wc202, n_3230);
  and g3686 (n_3224, n_3218, wc203);
  not gc203 (wc203, n_3219);
  or g3687 (n_3252, wc204, n_3179);
  not gc204 (wc204, n_3250);
  or g3688 (n_3328, wc205, n_2901);
  not gc205 (wc205, n_3326);
  or g3689 (n_3333, wc206, n_2913);
  not gc206 (wc206, n_3331);
  or g3690 (n_3335, wc207, n_2919);
  not gc207 (wc207, n_3270);
  or g3691 (n_3343, wc208, n_2937);
  not gc208 (wc208, n_3341);
  or g3692 (n_3345, wc209, n_2943);
  not gc209 (wc209, n_3273);
  or g3693 (n_3350, wc210, n_2955);
  not gc210 (wc210, n_3250);
  or g3694 (n_3254, wc211, n_3185);
  not gc211 (wc211, n_3233);
  or g3695 (n_3360, wc212, n_2979);
  not gc212 (wc212, n_3233);
  or g3696 (n_3338, wc213, n_2925);
  not gc213 (wc213, n_3336);
  or g3697 (n_3348, wc214, n_2949);
  not gc214 (wc214, n_3346);
  or g3698 (n_3353, wc215, n_2961);
  not gc215 (wc215, n_3351);
  or g3699 (n_3355, wc216, n_2967);
  not gc216 (wc216, n_3276);
  or g3700 (n_3363, wc217, n_2985);
  not gc217 (wc217, n_3361);
  or g3701 (n_3365, wc218, n_2991);
  not gc218 (wc218, n_3279);
  or g3702 (n_3370, wc219, n_3003);
  not gc219 (wc219, n_3255);
  or g3703 (n_3358, wc220, n_2973);
  not gc220 (wc220, n_3356);
  or g3704 (n_3368, wc221, n_2997);
  not gc221 (wc221, n_3366);
  or g3705 (n_3373, n_3007, wc222);
  not gc222 (wc222, n_3371);
  not g3706 (Z[75], n_3521);
endmodule

module mult_signed_const_12824_GENERIC(A, Z);
  input [56:0] A;
  output [75:0] Z;
  wire [56:0] A;
  wire [75:0] Z;
  mult_signed_const_12824_GENERIC_REAL g1(.A ({A[56:2], A[0], A[0]}),
       .Z (Z));
endmodule

module mult_signed_const_13291_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [58:0] A;
  output [77:0] Z;
  wire [58:0] A;
  wire [77:0] Z;
  wire n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78;
  wire n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_374, n_375, n_376, n_377, n_378;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_388, n_390;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_401, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_441, n_442, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451;
  wire n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459;
  wire n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467;
  wire n_468, n_470, n_471, n_472, n_473, n_474, n_475, n_476;
  wire n_478, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_591, n_592, n_593, n_594;
  wire n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602;
  wire n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612;
  wire n_613, n_614, n_615, n_616, n_618, n_619, n_620, n_621;
  wire n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629;
  wire n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637;
  wire n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645;
  wire n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
  wire n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669;
  wire n_670, n_671, n_672, n_674, n_675, n_676, n_678, n_679;
  wire n_680, n_681, n_682, n_683, n_684, n_685, n_686, n_690;
  wire n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699;
  wire n_700, n_701, n_704, n_705, n_706, n_707, n_708, n_709;
  wire n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717;
  wire n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725;
  wire n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733;
  wire n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741;
  wire n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749;
  wire n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_758;
  wire n_759, n_760, n_762, n_763, n_764, n_765, n_766, n_767;
  wire n_768, n_769, n_770, n_773, n_776, n_777, n_778, n_779;
  wire n_780, n_781, n_782, n_783, n_784, n_786, n_788, n_789;
  wire n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797;
  wire n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805;
  wire n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813;
  wire n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821;
  wire n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_830;
  wire n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838;
  wire n_839, n_840, n_841, n_842, n_844, n_845, n_846, n_847;
  wire n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855;
  wire n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863;
  wire n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871;
  wire n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879;
  wire n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887;
  wire n_888, n_889, n_890, n_891, n_892, n_893, n_894, n_895;
  wire n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903;
  wire n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911;
  wire n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919;
  wire n_920, n_921, n_922, n_923, n_924, n_927, n_928, n_929;
  wire n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937;
  wire n_938, n_939, n_940, n_944, n_945, n_946, n_947, n_948;
  wire n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956;
  wire n_957, n_959, n_960, n_961, n_962, n_963, n_964, n_965;
  wire n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_975;
  wire n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983;
  wire n_984, n_985, n_986, n_987, n_989, n_990, n_992, n_993;
  wire n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1004;
  wire n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012;
  wire n_1013, n_1015, n_1016, n_1019, n_1020, n_1021, n_1022, n_1023;
  wire n_1024, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035;
  wire n_1037, n_1040, n_1041, n_1042, n_1043, n_1044, n_1050, n_1051;
  wire n_1052, n_1053, n_1057, n_1058, n_1059, n_1060, n_1064, n_1065;
  wire n_1066, n_1067, n_1069, n_1071, n_1072, n_1076, n_1077, n_1079;
  wire n_1080, n_1083, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091;
  wire n_1092, n_1093, n_1094, n_1095, n_1096, n_1098, n_1099, n_1100;
  wire n_1101, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111;
  wire n_1112, n_1114, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121;
  wire n_1122, n_1124, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131;
  wire n_1132, n_1133, n_1136, n_1138, n_1139, n_1140, n_1141, n_1142;
  wire n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1152;
  wire n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163;
  wire n_1164, n_1165, n_1166, n_1167, n_1170, n_1171, n_1172, n_1174;
  wire n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182;
  wire n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1190, n_1191;
  wire n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200;
  wire n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208;
  wire n_1209, n_1210, n_1211, n_1213, n_1214, n_1216, n_1217, n_1218;
  wire n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226;
  wire n_1227, n_1228, n_1229, n_1230, n_1233, n_1234, n_1235, n_1236;
  wire n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
  wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253;
  wire n_1254, n_1255, n_1256, n_1262, n_1263, n_1266, n_1267, n_1268;
  wire n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276;
  wire n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284;
  wire n_1285, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298;
  wire n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306;
  wire n_1307, n_1308, n_1309, n_1318, n_1319, n_1321, n_1322, n_1323;
  wire n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332;
  wire n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340;
  wire n_1341, n_1344, n_1345, n_1350, n_1351, n_1352, n_1354, n_1355;
  wire n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363;
  wire n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371;
  wire n_1372, n_1373, n_1374, n_1376, n_1377, n_1382, n_1383, n_1384;
  wire n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393;
  wire n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401;
  wire n_1402, n_1403, n_1404, n_1405, n_1408, n_1409, n_1412, n_1413;
  wire n_1414, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424;
  wire n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432;
  wire n_1433, n_1434, n_1435, n_1436, n_1437, n_1440, n_1441, n_1444;
  wire n_1445, n_1446, n_1447, n_1448, n_1450, n_1451, n_1452, n_1453;
  wire n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461;
  wire n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469;
  wire n_1472, n_1473, n_1474, n_1475, n_1477, n_1478, n_1480, n_1481;
  wire n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489;
  wire n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
  wire n_1498, n_1499, n_1500, n_1501, n_1504, n_1505, n_1510, n_1512;
  wire n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520;
  wire n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528;
  wire n_1529, n_1530, n_1531, n_1532, n_1533, n_1538, n_1539, n_1542;
  wire n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552;
  wire n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560;
  wire n_1561, n_1562, n_1563, n_1564, n_1565, n_1570, n_1571, n_1572;
  wire n_1574, n_1577, n_1578, n_1579, n_1581, n_1582, n_1583, n_1584;
  wire n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592;
  wire n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1601;
  wire n_1602, n_1603, n_1604, n_1605, n_1606, n_1609, n_1610, n_1611;
  wire n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619;
  wire n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627;
  wire n_1628, n_1629, n_1630, n_1631, n_1633, n_1634, n_1635, n_1636;
  wire n_1637, n_1638, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646;
  wire n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654;
  wire n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662;
  wire n_1663, n_1665, n_1666, n_1668, n_1669, n_1670, n_1672, n_1674;
  wire n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682;
  wire n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690;
  wire n_1691, n_1692, n_1693, n_1694, n_1695, n_1697, n_1698, n_1700;
  wire n_1701, n_1702, n_1704, n_1706, n_1707, n_1708, n_1709, n_1710;
  wire n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718;
  wire n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726;
  wire n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1738;
  wire n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746;
  wire n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754;
  wire n_1755, n_1756, n_1757, n_1758, n_1761, n_1762, n_1763, n_1764;
  wire n_1765, n_1766, n_1767, n_1770, n_1771, n_1772, n_1773, n_1774;
  wire n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782;
  wire n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1794;
  wire n_1795, n_1798, n_1799, n_1800, n_1802, n_1803, n_1804, n_1805;
  wire n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813;
  wire n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821;
  wire n_1826, n_1827, n_1830, n_1831, n_1832, n_1834, n_1835, n_1837;
  wire n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845;
  wire n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853;
  wire n_1856, n_1857, n_1858, n_1860, n_1861, n_1862, n_1864, n_1865;
  wire n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873;
  wire n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881;
  wire n_1882, n_1883, n_1884, n_1885, n_1888, n_1889, n_1890, n_1892;
  wire n_1893, n_1894, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901;
  wire n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909;
  wire n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917;
  wire n_1920, n_1921, n_1922, n_1923, n_1925, n_1926, n_1928, n_1929;
  wire n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937;
  wire n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945;
  wire n_1946, n_1947, n_1948, n_1949, n_1952, n_1953, n_1954, n_1955;
  wire n_1957, n_1958, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965;
  wire n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973;
  wire n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981;
  wire n_1990, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999;
  wire n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007;
  wire n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2022, n_2025;
  wire n_2026, n_2027, n_2029, n_2030, n_2031, n_2032, n_2034, n_2035;
  wire n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043;
  wire n_2044, n_2045, n_2048, n_2049, n_2050, n_2051, n_2054, n_2055;
  wire n_2056, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064;
  wire n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072;
  wire n_2073, n_2074, n_2075, n_2076, n_2077, n_2080, n_2081, n_2082;
  wire n_2083, n_2086, n_2087, n_2088, n_2090, n_2091, n_2092, n_2093;
  wire n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101;
  wire n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109;
  wire n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119;
  wire n_2120, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128;
  wire n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136;
  wire n_2137, n_2138, n_2139, n_2140, n_2141, n_2144, n_2145, n_2146;
  wire n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2154, n_2155;
  wire n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163;
  wire n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171;
  wire n_2172, n_2173, n_2178, n_2179, n_2180, n_2181, n_2186, n_2187;
  wire n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195;
  wire n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203;
  wire n_2204, n_2205, n_2210, n_2211, n_2212, n_2213, n_2218, n_2219;
  wire n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228;
  wire n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236;
  wire n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2245;
  wire n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253;
  wire n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261;
  wire n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269;
  wire n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2277, n_2278;
  wire n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286;
  wire n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294;
  wire n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302;
  wire n_2303, n_2304, n_2305, n_2306, n_2308, n_2310, n_2314, n_2315;
  wire n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323;
  wire n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331;
  wire n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2340;
  wire n_2342, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352;
  wire n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360;
  wire n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368;
  wire n_2369, n_2370, n_2372, n_2374, n_2375, n_2378, n_2379, n_2380;
  wire n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388;
  wire n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396;
  wire n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2404, n_2406;
  wire n_2407, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416;
  wire n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424;
  wire n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432;
  wire n_2433, n_2434, n_2436, n_2438, n_2439, n_2442, n_2443, n_2444;
  wire n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452;
  wire n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460;
  wire n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2468, n_2470;
  wire n_2471, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480;
  wire n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488;
  wire n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496;
  wire n_2497, n_2498, n_2499, n_2500, n_2502, n_2503, n_2506, n_2507;
  wire n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515;
  wire n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523;
  wire n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531;
  wire n_2532, n_2534, n_2535, n_2538, n_2539, n_2540, n_2541, n_2542;
  wire n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550;
  wire n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558;
  wire n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2566, n_2570;
  wire n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578;
  wire n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586;
  wire n_2587, n_2588, n_2589, n_2590, n_2591, n_2593, n_2594, n_2595;
  wire n_2596, n_2597, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606;
  wire n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614;
  wire n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622;
  wire n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2630, n_2631;
  wire n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640;
  wire n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648;
  wire n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2658;
  wire n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668;
  wire n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676;
  wire n_2677, n_2678, n_2679, n_2680, n_2681, n_2686, n_2689, n_2690;
  wire n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698;
  wire n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706;
  wire n_2707, n_2708, n_2709, n_2710, n_2714, n_2716, n_2717, n_2718;
  wire n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727;
  wire n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2742, n_2744;
  wire n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752;
  wire n_2753, n_2754, n_2755, n_2756, n_2757, n_2764, n_2765, n_2766;
  wire n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774;
  wire n_2775, n_2776, n_2777, n_2786, n_2787, n_2788, n_2789, n_2790;
  wire n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2804;
  wire n_2805, n_2806, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813;
  wire n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827;
  wire n_2828, n_2829, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841;
  wire n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853;
  wire n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2866, n_2867;
  wire n_2868, n_2869, n_2871, n_2872, n_2873, n_2876, n_2877, n_2889;
  wire n_2891, n_2893, n_2894, n_2895, n_2896, n_2897, n_2899, n_2900;
  wire n_2901, n_2902, n_2903, n_2905, n_2906, n_2907, n_2908, n_2909;
  wire n_2911, n_2912, n_2913, n_2914, n_2915, n_2917, n_2918, n_2919;
  wire n_2920, n_2921, n_2923, n_2924, n_2925, n_2926, n_2927, n_2929;
  wire n_2930, n_2931, n_2932, n_2933, n_2935, n_2936, n_2937, n_2938;
  wire n_2939, n_2941, n_2942, n_2943, n_2944, n_2945, n_2947, n_2948;
  wire n_2949, n_2950, n_2951, n_2953, n_2954, n_2955, n_2956, n_2957;
  wire n_2959, n_2960, n_2961, n_2962, n_2963, n_2965, n_2966, n_2967;
  wire n_2968, n_2969, n_2971, n_2972, n_2973, n_2974, n_2975, n_2977;
  wire n_2978, n_2979, n_2980, n_2981, n_2983, n_2984, n_2985, n_2986;
  wire n_2987, n_2989, n_2990, n_2991, n_2992, n_2993, n_2995, n_2996;
  wire n_2997, n_2998, n_2999, n_3001, n_3002, n_3003, n_3004, n_3005;
  wire n_3007, n_3008, n_3009, n_3010, n_3011, n_3013, n_3014, n_3015;
  wire n_3016, n_3017, n_3019, n_3020, n_3021, n_3022, n_3023, n_3025;
  wire n_3026, n_3027, n_3028, n_3029, n_3031, n_3032, n_3033, n_3034;
  wire n_3035, n_3037, n_3038, n_3039, n_3040, n_3041, n_3043, n_3044;
  wire n_3045, n_3046, n_3047, n_3049, n_3050, n_3051, n_3052, n_3053;
  wire n_3055, n_3056, n_3057, n_3058, n_3059, n_3061, n_3062, n_3063;
  wire n_3064, n_3065, n_3067, n_3068, n_3069, n_3070, n_3071, n_3073;
  wire n_3074, n_3075, n_3076, n_3077, n_3079, n_3080, n_3081, n_3082;
  wire n_3083, n_3085, n_3086, n_3087, n_3088, n_3089, n_3091, n_3092;
  wire n_3093, n_3094, n_3095, n_3097, n_3098, n_3099, n_3100, n_3101;
  wire n_3103, n_3104, n_3105, n_3106, n_3107, n_3109, n_3110, n_3113;
  wire n_3118, n_3120, n_3121, n_3123, n_3125, n_3127, n_3128, n_3130;
  wire n_3131, n_3133, n_3135, n_3137, n_3138, n_3140, n_3141, n_3143;
  wire n_3145, n_3147, n_3148, n_3150, n_3151, n_3153, n_3155, n_3157;
  wire n_3158, n_3160, n_3161, n_3163, n_3165, n_3167, n_3168, n_3170;
  wire n_3171, n_3173, n_3175, n_3177, n_3178, n_3180, n_3181, n_3183;
  wire n_3185, n_3187, n_3188, n_3190, n_3191, n_3193, n_3195, n_3197;
  wire n_3198, n_3200, n_3201, n_3203, n_3205, n_3207, n_3208, n_3210;
  wire n_3211, n_3213, n_3215, n_3217, n_3218, n_3220, n_3221, n_3223;
  wire n_3225, n_3227, n_3228, n_3230, n_3231, n_3233, n_3235, n_3237;
  wire n_3238, n_3240, n_3241, n_3243, n_3245, n_3247, n_3248, n_3250;
  wire n_3251, n_3253, n_3255, n_3257, n_3258, n_3260, n_3261, n_3263;
  wire n_3265, n_3267, n_3268, n_3270, n_3271, n_3273, n_3275, n_3277;
  wire n_3278, n_3280, n_3281, n_3283, n_3285, n_3287, n_3288, n_3290;
  wire n_3291, n_3293, n_3295, n_3297, n_3298, n_3302, n_3303, n_3304;
  wire n_3306, n_3307, n_3308, n_3310, n_3311, n_3312, n_3313, n_3315;
  wire n_3317, n_3319, n_3320, n_3321, n_3323, n_3324, n_3325, n_3327;
  wire n_3328, n_3330, n_3332, n_3334, n_3335, n_3336, n_3338, n_3339;
  wire n_3340, n_3342, n_3343, n_3345, n_3347, n_3349, n_3350, n_3351;
  wire n_3353, n_3354, n_3355, n_3357, n_3358, n_3360, n_3362, n_3364;
  wire n_3365, n_3366, n_3368, n_3369, n_3370, n_3372, n_3373, n_3375;
  wire n_3377, n_3379, n_3380, n_3381, n_3383, n_3384, n_3385, n_3387;
  wire n_3388, n_3390, n_3392, n_3394, n_3395, n_3396, n_3398, n_3399;
  wire n_3400, n_3402, n_3403, n_3405, n_3407, n_3409, n_3410, n_3411;
  wire n_3413, n_3414, n_3415, n_3417, n_3418, n_3420, n_3422, n_3424;
  wire n_3425, n_3426, n_3428, n_3429, n_3430, n_3432, n_3433, n_3435;
  wire n_3436, n_3438, n_3439, n_3440, n_3442, n_3443, n_3445, n_3446;
  wire n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454;
  wire n_3455, n_3456, n_3457, n_3458, n_3459, n_3461, n_3464, n_3466;
  wire n_3467, n_3468, n_3471, n_3474, n_3476, n_3477, n_3479, n_3481;
  wire n_3482, n_3484, n_3486, n_3487, n_3489, n_3491, n_3492, n_3494;
  wire n_3495, n_3497, n_3500, n_3502, n_3503, n_3504, n_3507, n_3510;
  wire n_3512, n_3513, n_3515, n_3517, n_3518, n_3520, n_3522, n_3523;
  wire n_3525, n_3527, n_3528, n_3530, n_3531, n_3533, n_3536, n_3538;
  wire n_3539, n_3540, n_3543, n_3546, n_3548, n_3549, n_3551, n_3553;
  wire n_3554, n_3556, n_3558, n_3559, n_3561, n_3563, n_3564, n_3566;
  wire n_3567, n_3569, n_3572, n_3574, n_3575, n_3576, n_3579, n_3582;
  wire n_3584, n_3585, n_3587, n_3589, n_3590, n_3591, n_3593, n_3594;
  wire n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603;
  wire n_3604, n_3605, n_3606, n_3607, n_3609, n_3610, n_3611, n_3613;
  wire n_3614, n_3615, n_3617, n_3618, n_3619, n_3621, n_3622, n_3623;
  wire n_3625, n_3626, n_3627, n_3629, n_3630, n_3631, n_3633, n_3634;
  wire n_3635, n_3637, n_3638, n_3639, n_3640, n_3642, n_3644, n_3646;
  wire n_3647, n_3648, n_3650, n_3652, n_3654, n_3655, n_3657, n_3659;
  wire n_3660, n_3662, n_3664, n_3665, n_3668, n_3670, n_3671, n_3672;
  wire n_3674, n_3675, n_3676, n_3678, n_3679, n_3680, n_3682, n_3683;
  wire n_3684, n_3686, n_3687, n_3688, n_3690, n_3691, n_3692, n_3694;
  wire n_3695, n_3696, n_3698, n_3699, n_3700, n_3702, n_3704, n_3705;
  wire n_3706, n_3708, n_3709, n_3711, n_3712, n_3713, n_3714, n_3715;
  wire n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3724;
  wire n_3725, n_3726, n_3728, n_3729, n_3730, n_3732, n_3733, n_3734;
  wire n_3736, n_3737, n_3738, n_3740, n_3741, n_3742, n_3744, n_3745;
  wire n_3746, n_3748, n_3749, n_3751, n_3752, n_3753, n_3754, n_3755;
  wire n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, n_3762, n_3763;
  wire n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771;
  wire n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779;
  wire n_3780, n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787;
  wire n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795;
  wire n_3796, n_3797, n_3798, n_3799, n_3800, n_3802, n_3803, n_3804;
  wire n_3806, n_3807, n_3809, n_3810, n_3811, n_3812, n_3813, n_3814;
  wire n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, n_3822, n_3823;
  wire n_3824, n_3826, n_3827, n_3828, n_3830, n_3831, n_3832, n_3834;
  wire n_3835, n_3836, n_3838, n_3839, n_3841, n_3844, n_3845, n_3847;
  wire n_3848, n_3849, n_3850, n_3852, n_3853, n_3854, n_3856, n_3857;
  wire n_3858, n_3859, n_3861, n_3862, n_3864, n_3865, n_3867, n_3868;
  wire n_3869, n_3870, n_3872, n_3873, n_3874, n_3876, n_3877, n_3878;
  wire n_3879, n_3881, n_3882, n_3884, n_3885, n_3887, n_3888, n_3889;
  wire n_3890, n_3892, n_3893, n_3894, n_3895, n_3897, n_3898, n_3899;
  wire n_3900, n_3902, n_3903, n_3905, n_3906, n_3908, n_3909, n_3910;
  wire n_3911, n_3913, n_3914, n_3915, n_3917, n_3918, n_3919, n_3920;
  wire n_3922, n_3923, n_3925, n_3926, n_3928, n_3929, n_3930, n_3931;
  wire n_3933, n_3934, n_3935, n_3936, n_3938, n_3939, n_3940, n_3941;
  wire n_3943, n_3944, n_3946, n_3947, n_3949, n_3950, n_3951, n_3952;
  wire n_3954, n_3955, n_3957, n_3958, n_3960, n_3961, n_3962, n_3963;
  wire n_3965, n_3966, n_3968, n_3969, n_3971, n_3972, n_3973, n_3974;
  wire n_3976, n_3977, n_3978, n_3979, n_3981, n_3982, n_3983, n_3984;
  wire n_3986, n_3987, n_3989, n_3990, n_3992, n_3993, n_3994, n_3995;
  wire n_3997, n_3998, n_3999, n_4001, n_4002, n_4003, n_4004, n_4006;
  wire n_4007, n_4009, n_4010, n_4012, n_4013, n_4014, n_4015, n_4017;
  wire n_4018, n_4019, n_4020, n_4022, n_4023, n_4024, n_4025, n_4027;
  wire n_4028, n_4030, n_4031, n_4033;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g468 (n_211, A[4], A[0]);
  and g2 (n_132, A[4], A[0]);
  xor g469 (n_1086, A[1], A[3]);
  xor g470 (n_210, n_1086, A[5]);
  nand g3 (n_1087, A[1], A[3]);
  nand g471 (n_1088, A[5], A[3]);
  nand g472 (n_1089, A[1], A[5]);
  nand g473 (n_131, n_1087, n_1088, n_1089);
  xor g474 (n_295, A[6], A[4]);
  and g475 (n_296, A[6], A[4]);
  xor g476 (n_1090, A[0], A[2]);
  xor g477 (n_209, n_1090, n_295);
  nand g478 (n_1091, A[0], A[2]);
  nand g4 (n_1092, n_295, A[2]);
  nand g5 (n_1093, A[0], n_295);
  nand g479 (n_130, n_1091, n_1092, n_1093);
  xor g480 (n_1094, A[1], A[7]);
  xor g481 (n_297, n_1094, A[5]);
  nand g482 (n_1095, A[1], A[7]);
  nand g483 (n_1096, A[5], A[7]);
  nand g6 (n_299, n_1095, n_1096, n_1089);
  xor g485 (n_1098, A[3], n_296);
  xor g486 (n_208, n_1098, n_297);
  nand g487 (n_1099, A[3], n_296);
  nand g488 (n_1100, n_297, n_296);
  nand g489 (n_1101, A[3], n_297);
  nand g490 (n_129, n_1099, n_1100, n_1101);
  xor g491 (n_298, A[8], A[6]);
  and g492 (n_301, A[8], A[6]);
  xor g494 (n_300, n_1090, A[4]);
  nand g497 (n_1105, A[2], A[4]);
  xor g499 (n_1106, n_298, n_299);
  xor g500 (n_207, n_1106, n_300);
  nand g501 (n_1107, n_298, n_299);
  nand g502 (n_1108, n_300, n_299);
  nand g503 (n_1109, n_298, n_300);
  nand g504 (n_128, n_1107, n_1108, n_1109);
  xor g505 (n_1110, A[1], A[9]);
  xor g506 (n_303, n_1110, A[3]);
  nand g507 (n_1111, A[1], A[9]);
  nand g508 (n_1112, A[3], A[9]);
  nand g510 (n_306, n_1111, n_1112, n_1087);
  xor g511 (n_1114, A[7], A[5]);
  xor g512 (n_304, n_1114, n_301);
  nand g514 (n_1116, n_301, A[5]);
  nand g515 (n_1117, A[7], n_301);
  nand g516 (n_308, n_1096, n_1116, n_1117);
  xor g517 (n_1118, n_302, n_303);
  xor g518 (n_206, n_1118, n_304);
  nand g519 (n_1119, n_302, n_303);
  nand g520 (n_1120, n_304, n_303);
  nand g521 (n_1121, n_302, n_304);
  nand g522 (n_127, n_1119, n_1120, n_1121);
  xor g523 (n_305, A[10], A[8]);
  and g524 (n_310, A[10], A[8]);
  xor g525 (n_1122, A[4], A[2]);
  xor g526 (n_307, n_1122, A[6]);
  nand g528 (n_1124, A[6], A[2]);
  xor g531 (n_1126, A[0], n_305);
  xor g532 (n_309, n_1126, n_306);
  nand g533 (n_1127, A[0], n_305);
  nand g534 (n_1128, n_306, n_305);
  nand g535 (n_1129, A[0], n_306);
  nand g536 (n_314, n_1127, n_1128, n_1129);
  xor g537 (n_1130, n_307, n_308);
  xor g538 (n_205, n_1130, n_309);
  nand g539 (n_1131, n_307, n_308);
  nand g540 (n_1132, n_309, n_308);
  nand g541 (n_1133, n_307, n_309);
  nand g542 (n_126, n_1131, n_1132, n_1133);
  xor g544 (n_312, n_1110, A[5]);
  nand g546 (n_1136, A[5], A[9]);
  nand g548 (n_317, n_1111, n_1136, n_1089);
  xor g549 (n_1138, A[3], A[11]);
  xor g550 (n_313, n_1138, A[7]);
  nand g551 (n_1139, A[3], A[11]);
  nand g552 (n_1140, A[7], A[11]);
  nand g553 (n_1141, A[3], A[7]);
  nand g554 (n_318, n_1139, n_1140, n_1141);
  xor g555 (n_1142, n_310, n_311);
  xor g556 (n_315, n_1142, n_312);
  nand g557 (n_1143, n_310, n_311);
  nand g558 (n_1144, n_312, n_311);
  nand g559 (n_1145, n_310, n_312);
  nand g560 (n_322, n_1143, n_1144, n_1145);
  xor g561 (n_1146, n_313, n_314);
  xor g562 (n_204, n_1146, n_315);
  nand g563 (n_1147, n_313, n_314);
  nand g564 (n_1148, n_315, n_314);
  nand g565 (n_1149, n_313, n_315);
  nand g566 (n_125, n_1147, n_1148, n_1149);
  xor g567 (n_316, A[12], A[10]);
  and g568 (n_323, A[12], A[10]);
  xor g570 (n_319, n_295, A[8]);
  nand g572 (n_1152, A[8], A[4]);
  xor g576 (n_320, n_1090, n_316);
  nand g578 (n_1156, n_316, A[0]);
  nand g579 (n_1157, A[2], n_316);
  nand g580 (n_327, n_1091, n_1156, n_1157);
  xor g581 (n_1158, n_317, n_318);
  xor g582 (n_321, n_1158, n_319);
  nand g583 (n_1159, n_317, n_318);
  nand g584 (n_1160, n_319, n_318);
  nand g585 (n_1161, n_317, n_319);
  nand g586 (n_329, n_1159, n_1160, n_1161);
  xor g587 (n_1162, n_320, n_321);
  xor g588 (n_203, n_1162, n_322);
  nand g589 (n_1163, n_320, n_321);
  nand g590 (n_1164, n_322, n_321);
  nand g591 (n_1165, n_320, n_322);
  nand g592 (n_124, n_1163, n_1164, n_1165);
  xor g593 (n_1166, A[1], A[11]);
  xor g594 (n_326, n_1166, A[7]);
  nand g595 (n_1167, A[1], A[11]);
  nand g598 (n_332, n_1167, n_1140, n_1095);
  xor g599 (n_1170, A[5], A[13]);
  xor g600 (n_325, n_1170, A[3]);
  nand g601 (n_1171, A[5], A[13]);
  nand g602 (n_1172, A[3], A[13]);
  nand g604 (n_333, n_1171, n_1172, n_1088);
  xor g605 (n_1174, A[9], n_323);
  xor g606 (n_328, n_1174, n_324);
  nand g607 (n_1175, A[9], n_323);
  nand g608 (n_1176, n_324, n_323);
  nand g609 (n_1177, A[9], n_324);
  nand g610 (n_336, n_1175, n_1176, n_1177);
  xor g611 (n_1178, n_325, n_326);
  xor g612 (n_330, n_1178, n_327);
  nand g613 (n_1179, n_325, n_326);
  nand g614 (n_1180, n_327, n_326);
  nand g615 (n_1181, n_325, n_327);
  nand g616 (n_338, n_1179, n_1180, n_1181);
  xor g617 (n_1182, n_328, n_329);
  xor g618 (n_202, n_1182, n_330);
  nand g619 (n_1183, n_328, n_329);
  nand g620 (n_1184, n_330, n_329);
  nand g621 (n_1185, n_328, n_330);
  nand g622 (n_123, n_1183, n_1184, n_1185);
  xor g623 (n_331, A[14], A[12]);
  and g624 (n_340, A[14], A[12]);
  xor g625 (n_1186, A[8], A[0]);
  xor g626 (n_335, n_1186, A[6]);
  nand g627 (n_1187, A[8], A[0]);
  nand g628 (n_1188, A[6], A[0]);
  xor g631 (n_1190, A[10], A[4]);
  xor g632 (n_334, n_1190, A[2]);
  nand g633 (n_1191, A[10], A[4]);
  nand g635 (n_1193, A[10], A[2]);
  nand g636 (n_343, n_1191, n_1105, n_1193);
  xor g637 (n_1194, n_331, n_332);
  xor g638 (n_337, n_1194, n_333);
  nand g639 (n_1195, n_331, n_332);
  nand g640 (n_1196, n_333, n_332);
  nand g641 (n_1197, n_331, n_333);
  nand g642 (n_346, n_1195, n_1196, n_1197);
  xor g643 (n_1198, n_334, n_335);
  xor g644 (n_339, n_1198, n_336);
  nand g645 (n_1199, n_334, n_335);
  nand g646 (n_1200, n_336, n_335);
  nand g647 (n_1201, n_334, n_336);
  nand g648 (n_349, n_1199, n_1200, n_1201);
  xor g649 (n_1202, n_337, n_338);
  xor g650 (n_201, n_1202, n_339);
  nand g651 (n_1203, n_337, n_338);
  nand g652 (n_1204, n_339, n_338);
  nand g653 (n_1205, n_337, n_339);
  nand g654 (n_122, n_1203, n_1204, n_1205);
  xor g655 (n_1206, A[1], A[15]);
  xor g656 (n_341, n_1206, A[13]);
  nand g657 (n_1207, A[1], A[15]);
  nand g658 (n_1208, A[13], A[15]);
  nand g659 (n_1209, A[1], A[13]);
  nand g660 (n_351, n_1207, n_1208, n_1209);
  xor g661 (n_1210, A[9], A[7]);
  xor g662 (n_344, n_1210, A[11]);
  nand g663 (n_1211, A[9], A[7]);
  nand g665 (n_1213, A[9], A[11]);
  nand g666 (n_352, n_1211, n_1140, n_1213);
  xor g667 (n_1214, A[5], A[3]);
  xor g668 (n_345, n_1214, n_340);
  nand g670 (n_1216, n_340, A[3]);
  nand g671 (n_1217, A[5], n_340);
  nand g672 (n_355, n_1088, n_1216, n_1217);
  xor g673 (n_1218, n_341, n_342);
  xor g674 (n_347, n_1218, n_343);
  nand g675 (n_1219, n_341, n_342);
  nand g676 (n_1220, n_343, n_342);
  nand g677 (n_1221, n_341, n_343);
  nand g678 (n_357, n_1219, n_1220, n_1221);
  xor g679 (n_1222, n_344, n_345);
  xor g680 (n_348, n_1222, n_346);
  nand g681 (n_1223, n_344, n_345);
  nand g682 (n_1224, n_346, n_345);
  nand g683 (n_1225, n_344, n_346);
  nand g684 (n_359, n_1223, n_1224, n_1225);
  xor g685 (n_1226, n_347, n_348);
  xor g686 (n_200, n_1226, n_349);
  nand g687 (n_1227, n_347, n_348);
  nand g688 (n_1228, n_349, n_348);
  nand g689 (n_1229, n_347, n_349);
  nand g690 (n_121, n_1227, n_1228, n_1229);
  xor g691 (n_350, A[16], A[14]);
  and g692 (n_361, A[16], A[14]);
  xor g693 (n_1230, A[10], A[2]);
  xor g694 (n_354, n_1230, A[0]);
  nand g697 (n_1233, A[10], A[0]);
  nand g698 (n_363, n_1193, n_1091, n_1233);
  xor g699 (n_1234, A[8], A[12]);
  xor g700 (n_353, n_1234, A[6]);
  nand g701 (n_1235, A[8], A[12]);
  nand g702 (n_1236, A[6], A[12]);
  xor g705 (n_1238, A[4], n_350);
  xor g706 (n_356, n_1238, n_351);
  nand g707 (n_1239, A[4], n_350);
  nand g708 (n_1240, n_351, n_350);
  nand g709 (n_1241, A[4], n_351);
  nand g710 (n_367, n_1239, n_1240, n_1241);
  xor g711 (n_1242, n_352, n_353);
  xor g712 (n_358, n_1242, n_354);
  nand g713 (n_1243, n_352, n_353);
  nand g714 (n_1244, n_354, n_353);
  nand g715 (n_1245, n_352, n_354);
  nand g716 (n_368, n_1243, n_1244, n_1245);
  xor g717 (n_1246, n_355, n_356);
  xor g718 (n_360, n_1246, n_357);
  nand g719 (n_1247, n_355, n_356);
  nand g720 (n_1248, n_357, n_356);
  nand g721 (n_1249, n_355, n_357);
  nand g722 (n_371, n_1247, n_1248, n_1249);
  xor g723 (n_1250, n_358, n_359);
  xor g724 (n_199, n_1250, n_360);
  nand g725 (n_1251, n_358, n_359);
  nand g726 (n_1252, n_360, n_359);
  nand g727 (n_1253, n_358, n_360);
  nand g728 (n_120, n_1251, n_1252, n_1253);
  xor g729 (n_1254, A[1], A[17]);
  xor g730 (n_362, n_1254, A[15]);
  nand g731 (n_1255, A[1], A[17]);
  nand g732 (n_1256, A[15], A[17]);
  nand g734 (n_374, n_1255, n_1256, n_1207);
  xor g736 (n_366, n_1138, A[9]);
  nand g740 (n_376, n_1139, n_1213, n_1112);
  xor g741 (n_1262, A[13], A[7]);
  xor g742 (n_365, n_1262, A[5]);
  nand g743 (n_1263, A[13], A[7]);
  nand g746 (n_375, n_1263, n_1096, n_1171);
  xor g747 (n_1266, n_361, n_362);
  xor g748 (n_369, n_1266, n_363);
  nand g749 (n_1267, n_361, n_362);
  nand g750 (n_1268, n_363, n_362);
  nand g751 (n_1269, n_361, n_363);
  nand g752 (n_380, n_1267, n_1268, n_1269);
  xor g753 (n_1270, n_364, n_365);
  xor g754 (n_370, n_1270, n_366);
  nand g755 (n_1271, n_364, n_365);
  nand g756 (n_1272, n_366, n_365);
  nand g757 (n_1273, n_364, n_366);
  nand g758 (n_382, n_1271, n_1272, n_1273);
  xor g759 (n_1274, n_367, n_368);
  xor g760 (n_372, n_1274, n_369);
  nand g761 (n_1275, n_367, n_368);
  nand g762 (n_1276, n_369, n_368);
  nand g763 (n_1277, n_367, n_369);
  nand g764 (n_384, n_1275, n_1276, n_1277);
  xor g765 (n_1278, n_370, n_371);
  xor g766 (n_198, n_1278, n_372);
  nand g767 (n_1279, n_370, n_371);
  nand g768 (n_1280, n_372, n_371);
  nand g769 (n_1281, n_370, n_372);
  nand g770 (n_119, n_1279, n_1280, n_1281);
  xor g773 (n_1282, A[18], A[12]);
  xor g774 (n_378, n_1282, A[4]);
  nand g775 (n_1283, A[18], A[12]);
  nand g776 (n_1284, A[4], A[12]);
  nand g777 (n_1285, A[18], A[4]);
  nand g778 (n_388, n_1283, n_1284, n_1285);
  xor g786 (n_377, n_298, n_350);
  nand g788 (n_1292, n_350, A[6]);
  nand g789 (n_1293, A[8], n_350);
  xor g791 (n_1294, n_374, n_375);
  xor g792 (n_381, n_1294, n_376);
  nand g793 (n_1295, n_374, n_375);
  nand g794 (n_1296, n_376, n_375);
  nand g795 (n_1297, n_374, n_376);
  nand g796 (n_393, n_1295, n_1296, n_1297);
  xor g797 (n_1298, n_377, n_378);
  xor g798 (n_383, n_1298, n_354);
  nand g799 (n_1299, n_377, n_378);
  nand g800 (n_1300, n_354, n_378);
  nand g801 (n_1301, n_377, n_354);
  nand g802 (n_395, n_1299, n_1300, n_1301);
  xor g803 (n_1302, n_380, n_381);
  xor g804 (n_385, n_1302, n_382);
  nand g805 (n_1303, n_380, n_381);
  nand g806 (n_1304, n_382, n_381);
  nand g807 (n_1305, n_380, n_382);
  nand g808 (n_398, n_1303, n_1304, n_1305);
  xor g809 (n_1306, n_383, n_384);
  xor g810 (n_197, n_1306, n_385);
  nand g811 (n_1307, n_383, n_384);
  nand g812 (n_1308, n_385, n_384);
  nand g813 (n_1309, n_383, n_385);
  nand g814 (n_118, n_1307, n_1308, n_1309);
  xor g827 (n_1318, A[19], A[11]);
  xor g828 (n_392, n_1318, A[9]);
  nand g829 (n_1319, A[19], A[11]);
  nand g831 (n_1321, A[19], A[9]);
  nand g832 (n_403, n_1319, n_1213, n_1321);
  xor g833 (n_1322, A[7], n_361);
  xor g834 (n_394, n_1322, n_362);
  nand g835 (n_1323, A[7], n_361);
  nand g837 (n_1325, A[7], n_362);
  nand g838 (n_134, n_1323, n_1267, n_1325);
  xor g839 (n_1326, n_388, n_363);
  xor g840 (n_396, n_1326, n_390);
  nand g841 (n_1327, n_388, n_363);
  nand g842 (n_1328, n_390, n_363);
  nand g843 (n_1329, n_388, n_390);
  nand g844 (n_137, n_1327, n_1328, n_1329);
  xor g845 (n_1330, n_325, n_392);
  xor g846 (n_397, n_1330, n_393);
  nand g847 (n_1331, n_325, n_392);
  nand g848 (n_1332, n_393, n_392);
  nand g849 (n_1333, n_325, n_393);
  nand g850 (n_405, n_1331, n_1332, n_1333);
  xor g851 (n_1334, n_394, n_395);
  xor g852 (n_399, n_1334, n_396);
  nand g853 (n_1335, n_394, n_395);
  nand g854 (n_1336, n_396, n_395);
  nand g855 (n_1337, n_394, n_396);
  nand g856 (n_407, n_1335, n_1336, n_1337);
  xor g857 (n_1338, n_397, n_398);
  xor g858 (n_196, n_1338, n_399);
  nand g859 (n_1339, n_397, n_398);
  nand g860 (n_1340, n_399, n_398);
  nand g861 (n_1341, n_397, n_399);
  nand g862 (n_117, n_1339, n_1340, n_1341);
  xor g864 (n_401, n_350, A[18]);
  nand g866 (n_1344, A[18], A[14]);
  nand g867 (n_1345, A[16], A[18]);
  xor g870 (n_133, n_295, A[12]);
  xor g875 (n_1350, A[2], A[20]);
  xor g876 (n_404, n_1350, A[10]);
  nand g877 (n_1351, A[2], A[20]);
  nand g878 (n_1352, A[10], A[20]);
  nand g880 (n_412, n_1351, n_1352, n_1193);
  xor g881 (n_1354, A[8], n_374);
  xor g882 (n_135, n_1354, n_401);
  nand g883 (n_1355, A[8], n_374);
  nand g884 (n_1356, n_401, n_374);
  nand g885 (n_1357, A[8], n_401);
  nand g886 (n_415, n_1355, n_1356, n_1357);
  xor g887 (n_1358, n_333, n_403);
  xor g888 (n_136, n_1358, n_404);
  nand g889 (n_1359, n_333, n_403);
  nand g890 (n_1360, n_404, n_403);
  nand g891 (n_1361, n_333, n_404);
  nand g892 (n_417, n_1359, n_1360, n_1361);
  xor g893 (n_1362, n_133, n_134);
  xor g894 (n_406, n_1362, n_135);
  nand g895 (n_1363, n_133, n_134);
  nand g896 (n_1364, n_135, n_134);
  nand g897 (n_1365, n_133, n_135);
  nand g898 (n_419, n_1363, n_1364, n_1365);
  xor g899 (n_1366, n_136, n_137);
  xor g900 (n_408, n_1366, n_405);
  nand g901 (n_1367, n_136, n_137);
  nand g902 (n_1368, n_405, n_137);
  nand g903 (n_1369, n_136, n_405);
  nand g904 (n_422, n_1367, n_1368, n_1369);
  xor g905 (n_1370, n_406, n_407);
  xor g906 (n_195, n_1370, n_408);
  nand g907 (n_1371, n_406, n_407);
  nand g908 (n_1372, n_408, n_407);
  nand g909 (n_1373, n_406, n_408);
  nand g910 (n_116, n_1371, n_1372, n_1373);
  xor g911 (n_1374, A[17], A[15]);
  xor g912 (n_409, n_1374, A[19]);
  nand g914 (n_1376, A[19], A[15]);
  nand g915 (n_1377, A[17], A[19]);
  nand g916 (n_424, n_1256, n_1376, n_1377);
  xor g918 (n_414, n_1114, A[13]);
  xor g923 (n_1382, A[3], A[21]);
  xor g924 (n_413, n_1382, A[11]);
  nand g925 (n_1383, A[3], A[21]);
  nand g926 (n_1384, A[11], A[21]);
  nand g928 (n_426, n_1383, n_1384, n_1139);
  xor g929 (n_1386, A[9], n_409);
  xor g930 (n_418, n_1386, n_410);
  nand g931 (n_1387, A[9], n_409);
  nand g932 (n_1388, n_410, n_409);
  nand g933 (n_1389, A[9], n_410);
  nand g934 (n_429, n_1387, n_1388, n_1389);
  xor g935 (n_1390, n_411, n_412);
  xor g936 (n_416, n_1390, n_413);
  nand g937 (n_1391, n_411, n_412);
  nand g938 (n_1392, n_413, n_412);
  nand g939 (n_1393, n_411, n_413);
  nand g940 (n_431, n_1391, n_1392, n_1393);
  xor g941 (n_1394, n_414, n_415);
  xor g942 (n_420, n_1394, n_416);
  nand g943 (n_1395, n_414, n_415);
  nand g944 (n_1396, n_416, n_415);
  nand g945 (n_1397, n_414, n_416);
  nand g946 (n_433, n_1395, n_1396, n_1397);
  xor g947 (n_1398, n_417, n_418);
  xor g948 (n_421, n_1398, n_419);
  nand g949 (n_1399, n_417, n_418);
  nand g950 (n_1400, n_419, n_418);
  nand g951 (n_1401, n_417, n_419);
  nand g952 (n_435, n_1399, n_1400, n_1401);
  xor g953 (n_1402, n_420, n_421);
  xor g954 (n_194, n_1402, n_422);
  nand g955 (n_1403, n_420, n_421);
  nand g956 (n_1404, n_422, n_421);
  nand g957 (n_1405, n_420, n_422);
  nand g958 (n_115, n_1403, n_1404, n_1405);
  xor g960 (n_423, n_350, A[20]);
  nand g962 (n_1408, A[20], A[14]);
  nand g963 (n_1409, A[16], A[20]);
  xor g966 (n_428, n_298, A[22]);
  nand g968 (n_1412, A[22], A[6]);
  nand g969 (n_1413, A[8], A[22]);
  xor g971 (n_1414, A[4], A[18]);
  xor g972 (n_427, n_1414, A[12]);
  xor g977 (n_1418, A[10], n_423);
  xor g978 (n_432, n_1418, n_424);
  nand g979 (n_1419, A[10], n_423);
  nand g980 (n_1420, n_424, n_423);
  nand g981 (n_1421, A[10], n_424);
  nand g982 (n_443, n_1419, n_1420, n_1421);
  xor g983 (n_1422, n_375, n_426);
  xor g984 (n_430, n_1422, n_427);
  nand g985 (n_1423, n_375, n_426);
  nand g986 (n_1424, n_427, n_426);
  nand g987 (n_1425, n_375, n_427);
  nand g988 (n_445, n_1423, n_1424, n_1425);
  xor g989 (n_1426, n_428, n_429);
  xor g990 (n_434, n_1426, n_430);
  nand g991 (n_1427, n_428, n_429);
  nand g992 (n_1428, n_430, n_429);
  nand g993 (n_1429, n_428, n_430);
  nand g994 (n_447, n_1427, n_1428, n_1429);
  xor g995 (n_1430, n_431, n_432);
  xor g996 (n_436, n_1430, n_433);
  nand g997 (n_1431, n_431, n_432);
  nand g998 (n_1432, n_433, n_432);
  nand g999 (n_1433, n_431, n_433);
  nand g1000 (n_450, n_1431, n_1432, n_1433);
  xor g1001 (n_1434, n_434, n_435);
  xor g1002 (n_193, n_1434, n_436);
  nand g1003 (n_1435, n_434, n_435);
  nand g1004 (n_1436, n_436, n_435);
  nand g1005 (n_1437, n_434, n_436);
  nand g1006 (n_114, n_1435, n_1436, n_1437);
  xor g1008 (n_437, n_1374, A[21]);
  nand g1010 (n_1440, A[21], A[15]);
  nand g1011 (n_1441, A[17], A[21]);
  nand g1012 (n_452, n_1256, n_1440, n_1441);
  xor g1014 (n_442, n_1210, A[23]);
  nand g1016 (n_1444, A[23], A[7]);
  nand g1017 (n_1445, A[9], A[23]);
  nand g1018 (n_453, n_1211, n_1444, n_1445);
  xor g1019 (n_1446, A[5], A[19]);
  xor g1020 (n_441, n_1446, A[13]);
  nand g1021 (n_1447, A[5], A[19]);
  nand g1022 (n_1448, A[13], A[19]);
  nand g1024 (n_454, n_1447, n_1448, n_1171);
  xor g1025 (n_1450, A[11], n_437);
  xor g1026 (n_446, n_1450, n_438);
  nand g1027 (n_1451, A[11], n_437);
  nand g1028 (n_1452, n_438, n_437);
  nand g1029 (n_1453, A[11], n_438);
  nand g1030 (n_457, n_1451, n_1452, n_1453);
  xor g1031 (n_1454, n_439, n_388);
  xor g1032 (n_444, n_1454, n_441);
  nand g1033 (n_1455, n_439, n_388);
  nand g1034 (n_1456, n_441, n_388);
  nand g1035 (n_1457, n_439, n_441);
  nand g1036 (n_458, n_1455, n_1456, n_1457);
  xor g1037 (n_1458, n_442, n_443);
  xor g1038 (n_448, n_1458, n_444);
  nand g1039 (n_1459, n_442, n_443);
  nand g1040 (n_1460, n_444, n_443);
  nand g1041 (n_1461, n_442, n_444);
  nand g1042 (n_461, n_1459, n_1460, n_1461);
  xor g1043 (n_1462, n_445, n_446);
  xor g1044 (n_449, n_1462, n_447);
  nand g1045 (n_1463, n_445, n_446);
  nand g1046 (n_1464, n_447, n_446);
  nand g1047 (n_1465, n_445, n_447);
  nand g1048 (n_464, n_1463, n_1464, n_1465);
  xor g1049 (n_1466, n_448, n_449);
  xor g1050 (n_192, n_1466, n_450);
  nand g1051 (n_1467, n_448, n_449);
  nand g1052 (n_1468, n_450, n_449);
  nand g1053 (n_1469, n_448, n_450);
  nand g1054 (n_113, n_1467, n_1468, n_1469);
  xor g1056 (n_451, n_350, A[24]);
  nand g1058 (n_1472, A[24], A[14]);
  nand g1059 (n_1473, A[16], A[24]);
  xor g1061 (n_1474, A[18], A[10]);
  xor g1062 (n_455, n_1474, A[8]);
  nand g1063 (n_1475, A[18], A[10]);
  nand g1065 (n_1477, A[18], A[8]);
  xor g1067 (n_1478, A[22], A[6]);
  xor g1068 (n_456, n_1478, A[20]);
  nand g1070 (n_1480, A[20], A[6]);
  nand g1071 (n_1481, A[22], A[20]);
  nand g1072 (n_468, n_1412, n_1480, n_1481);
  xor g1073 (n_1482, A[12], n_451);
  xor g1074 (n_460, n_1482, n_452);
  nand g1075 (n_1483, A[12], n_451);
  nand g1076 (n_1484, n_452, n_451);
  nand g1077 (n_1485, A[12], n_452);
  nand g1078 (n_471, n_1483, n_1484, n_1485);
  xor g1079 (n_1486, n_453, n_454);
  xor g1080 (n_459, n_1486, n_455);
  nand g1081 (n_1487, n_453, n_454);
  nand g1082 (n_1488, n_455, n_454);
  nand g1083 (n_1489, n_453, n_455);
  nand g1084 (n_472, n_1487, n_1488, n_1489);
  xor g1085 (n_1490, n_456, n_457);
  xor g1086 (n_462, n_1490, n_458);
  nand g1087 (n_1491, n_456, n_457);
  nand g1088 (n_1492, n_458, n_457);
  nand g1089 (n_1493, n_456, n_458);
  nand g1090 (n_213, n_1491, n_1492, n_1493);
  xor g1091 (n_1494, n_459, n_460);
  xor g1092 (n_463, n_1494, n_461);
  nand g1093 (n_1495, n_459, n_460);
  nand g1094 (n_1496, n_461, n_460);
  nand g1095 (n_1497, n_459, n_461);
  nand g1096 (n_476, n_1495, n_1496, n_1497);
  xor g1097 (n_1498, n_462, n_463);
  xor g1098 (n_191, n_1498, n_464);
  nand g1099 (n_1499, n_462, n_463);
  nand g1100 (n_1500, n_464, n_463);
  nand g1101 (n_1501, n_462, n_464);
  nand g1102 (n_112, n_1499, n_1500, n_1501);
  xor g1104 (n_465, n_1374, A[25]);
  nand g1106 (n_1504, A[25], A[15]);
  nand g1107 (n_1505, A[17], A[25]);
  nand g1108 (n_478, n_1256, n_1504, n_1505);
  xor g1115 (n_1510, A[23], A[7]);
  xor g1116 (n_470, n_1510, A[21]);
  nand g1118 (n_1512, A[21], A[7]);
  nand g1119 (n_1513, A[23], A[21]);
  nand g1120 (n_480, n_1444, n_1512, n_1513);
  xor g1121 (n_1514, A[13], n_465);
  xor g1122 (n_212, n_1514, n_466);
  nand g1123 (n_1515, A[13], n_465);
  nand g1124 (n_1516, n_466, n_465);
  nand g1125 (n_1517, A[13], n_466);
  nand g1126 (n_483, n_1515, n_1516, n_1517);
  xor g1127 (n_1518, n_467, n_468);
  xor g1128 (n_473, n_1518, n_392);
  nand g1129 (n_1519, n_467, n_468);
  nand g1130 (n_1520, n_392, n_468);
  nand g1131 (n_1521, n_467, n_392);
  nand g1132 (n_484, n_1519, n_1520, n_1521);
  xor g1133 (n_1522, n_470, n_471);
  xor g1134 (n_474, n_1522, n_472);
  nand g1135 (n_1523, n_470, n_471);
  nand g1136 (n_1524, n_472, n_471);
  nand g1137 (n_1525, n_470, n_472);
  nand g1138 (n_487, n_1523, n_1524, n_1525);
  xor g1139 (n_1526, n_473, n_212);
  xor g1140 (n_475, n_1526, n_213);
  nand g1141 (n_1527, n_473, n_212);
  nand g1142 (n_1528, n_213, n_212);
  nand g1143 (n_1529, n_473, n_213);
  nand g1144 (n_490, n_1527, n_1528, n_1529);
  xor g1145 (n_1530, n_474, n_475);
  xor g1146 (n_190, n_1530, n_476);
  nand g1147 (n_1531, n_474, n_475);
  nand g1148 (n_1532, n_476, n_475);
  nand g1149 (n_1533, n_474, n_476);
  nand g1150 (n_111, n_1531, n_1532, n_1533);
  xor g1157 (n_1538, A[20], A[12]);
  xor g1158 (n_481, n_1538, A[10]);
  nand g1159 (n_1539, A[20], A[12]);
  xor g1163 (n_1542, A[18], A[8]);
  xor g1164 (n_482, n_1542, A[22]);
  nand g1167 (n_1545, A[18], A[22]);
  nand g1168 (n_494, n_1477, n_1413, n_1545);
  xor g1169 (n_1546, A[26], n_451);
  xor g1170 (n_486, n_1546, n_478);
  nand g1171 (n_1547, A[26], n_451);
  nand g1172 (n_1548, n_478, n_451);
  nand g1173 (n_1549, A[26], n_478);
  nand g1174 (n_497, n_1547, n_1548, n_1549);
  xor g1175 (n_1550, n_403, n_480);
  xor g1176 (n_485, n_1550, n_481);
  nand g1177 (n_1551, n_403, n_480);
  nand g1178 (n_1552, n_481, n_480);
  nand g1179 (n_1553, n_403, n_481);
  nand g1180 (n_498, n_1551, n_1552, n_1553);
  xor g1181 (n_1554, n_482, n_483);
  xor g1182 (n_488, n_1554, n_484);
  nand g1183 (n_1555, n_482, n_483);
  nand g1184 (n_1556, n_484, n_483);
  nand g1185 (n_1557, n_482, n_484);
  nand g1186 (n_501, n_1555, n_1556, n_1557);
  xor g1187 (n_1558, n_485, n_486);
  xor g1188 (n_489, n_1558, n_487);
  nand g1189 (n_1559, n_485, n_486);
  nand g1190 (n_1560, n_487, n_486);
  nand g1191 (n_1561, n_485, n_487);
  nand g1192 (n_504, n_1559, n_1560, n_1561);
  xor g1193 (n_1562, n_488, n_489);
  xor g1194 (n_189, n_1562, n_490);
  nand g1195 (n_1563, n_488, n_489);
  nand g1196 (n_1564, n_490, n_489);
  nand g1197 (n_1565, n_488, n_490);
  nand g1198 (n_110, n_1563, n_1564, n_1565);
  xor g1205 (n_1570, A[21], A[13]);
  xor g1206 (n_495, n_1570, A[11]);
  nand g1207 (n_1571, A[21], A[13]);
  nand g1208 (n_1572, A[11], A[13]);
  nand g1210 (n_507, n_1571, n_1572, n_1384);
  xor g1211 (n_1574, A[19], A[9]);
  xor g1212 (n_496, n_1574, A[23]);
  nand g1215 (n_1577, A[19], A[23]);
  nand g1216 (n_508, n_1321, n_1445, n_1577);
  xor g1217 (n_1578, A[27], n_465);
  xor g1218 (n_500, n_1578, n_466);
  nand g1219 (n_1579, A[27], n_465);
  nand g1221 (n_1581, A[27], n_466);
  nand g1222 (n_511, n_1579, n_1516, n_1581);
  xor g1223 (n_1582, n_493, n_494);
  xor g1224 (n_499, n_1582, n_495);
  nand g1225 (n_1583, n_493, n_494);
  nand g1226 (n_1584, n_495, n_494);
  nand g1227 (n_1585, n_493, n_495);
  nand g1228 (n_512, n_1583, n_1584, n_1585);
  xor g1229 (n_1586, n_496, n_497);
  xor g1230 (n_502, n_1586, n_498);
  nand g1231 (n_1587, n_496, n_497);
  nand g1232 (n_1588, n_498, n_497);
  nand g1233 (n_1589, n_496, n_498);
  nand g1234 (n_515, n_1587, n_1588, n_1589);
  xor g1235 (n_1590, n_499, n_500);
  xor g1236 (n_503, n_1590, n_501);
  nand g1237 (n_1591, n_499, n_500);
  nand g1238 (n_1592, n_501, n_500);
  nand g1239 (n_1593, n_499, n_501);
  nand g1240 (n_518, n_1591, n_1592, n_1593);
  xor g1241 (n_1594, n_502, n_503);
  xor g1242 (n_188, n_1594, n_504);
  nand g1243 (n_1595, n_502, n_503);
  nand g1244 (n_1596, n_504, n_503);
  nand g1245 (n_1597, n_502, n_504);
  nand g1246 (n_109, n_1595, n_1596, n_1597);
  xor g1247 (n_1598, A[28], A[14]);
  xor g1248 (n_505, n_1598, A[16]);
  nand g1249 (n_1599, A[28], A[14]);
  nand g1251 (n_1601, A[28], A[16]);
  xor g1253 (n_1602, A[26], A[22]);
  xor g1254 (n_509, n_1602, A[12]);
  nand g1255 (n_1603, A[26], A[22]);
  nand g1256 (n_1604, A[12], A[22]);
  nand g1257 (n_1605, A[26], A[12]);
  nand g1258 (n_521, n_1603, n_1604, n_1605);
  xor g1259 (n_1606, A[20], A[10]);
  xor g1260 (n_510, n_1606, A[18]);
  nand g1263 (n_1609, A[20], A[18]);
  nand g1264 (n_522, n_1352, n_1475, n_1609);
  xor g1265 (n_1610, A[24], n_505);
  xor g1266 (n_514, n_1610, n_478);
  nand g1267 (n_1611, A[24], n_505);
  nand g1268 (n_1612, n_478, n_505);
  nand g1269 (n_1613, A[24], n_478);
  nand g1270 (n_525, n_1611, n_1612, n_1613);
  xor g1271 (n_1614, n_507, n_508);
  xor g1272 (n_513, n_1614, n_509);
  nand g1273 (n_1615, n_507, n_508);
  nand g1274 (n_1616, n_509, n_508);
  nand g1275 (n_1617, n_507, n_509);
  nand g1276 (n_528, n_1615, n_1616, n_1617);
  xor g1277 (n_1618, n_510, n_511);
  xor g1278 (n_516, n_1618, n_512);
  nand g1279 (n_1619, n_510, n_511);
  nand g1280 (n_1620, n_512, n_511);
  nand g1281 (n_1621, n_510, n_512);
  nand g1282 (n_529, n_1619, n_1620, n_1621);
  xor g1283 (n_1622, n_513, n_514);
  xor g1284 (n_517, n_1622, n_515);
  nand g1285 (n_1623, n_513, n_514);
  nand g1286 (n_1624, n_515, n_514);
  nand g1287 (n_1625, n_513, n_515);
  nand g1288 (n_532, n_1623, n_1624, n_1625);
  xor g1289 (n_1626, n_516, n_517);
  xor g1290 (n_187, n_1626, n_518);
  nand g1291 (n_1627, n_516, n_517);
  nand g1292 (n_1628, n_518, n_517);
  nand g1293 (n_1629, n_516, n_518);
  nand g1294 (n_108, n_1627, n_1628, n_1629);
  xor g1295 (n_1630, A[29], A[15]);
  xor g1296 (n_520, n_1630, A[17]);
  nand g1297 (n_1631, A[29], A[15]);
  nand g1299 (n_1633, A[29], A[17]);
  nand g1300 (n_533, n_1631, n_1256, n_1633);
  xor g1301 (n_1634, A[27], A[23]);
  xor g1302 (n_523, n_1634, A[13]);
  nand g1303 (n_1635, A[27], A[23]);
  nand g1304 (n_1636, A[13], A[23]);
  nand g1305 (n_1637, A[27], A[13]);
  nand g1306 (n_535, n_1635, n_1636, n_1637);
  xor g1307 (n_1638, A[21], A[11]);
  xor g1308 (n_524, n_1638, A[19]);
  nand g1311 (n_1641, A[21], A[19]);
  nand g1312 (n_536, n_1384, n_1319, n_1641);
  xor g1313 (n_1642, A[25], n_519);
  xor g1314 (n_526, n_1642, n_520);
  nand g1315 (n_1643, A[25], n_519);
  nand g1316 (n_1644, n_520, n_519);
  nand g1317 (n_1645, A[25], n_520);
  nand g1318 (n_539, n_1643, n_1644, n_1645);
  xor g1319 (n_1646, n_521, n_522);
  xor g1320 (n_527, n_1646, n_523);
  nand g1321 (n_1647, n_521, n_522);
  nand g1322 (n_1648, n_523, n_522);
  nand g1323 (n_1649, n_521, n_523);
  nand g1324 (n_542, n_1647, n_1648, n_1649);
  xor g1325 (n_1650, n_524, n_525);
  xor g1326 (n_530, n_1650, n_526);
  nand g1327 (n_1651, n_524, n_525);
  nand g1328 (n_1652, n_526, n_525);
  nand g1329 (n_1653, n_524, n_526);
  nand g1330 (n_543, n_1651, n_1652, n_1653);
  xor g1331 (n_1654, n_527, n_528);
  xor g1332 (n_531, n_1654, n_529);
  nand g1333 (n_1655, n_527, n_528);
  nand g1334 (n_1656, n_529, n_528);
  nand g1335 (n_1657, n_527, n_529);
  nand g1336 (n_546, n_1655, n_1656, n_1657);
  xor g1337 (n_1658, n_530, n_531);
  xor g1338 (n_186, n_1658, n_532);
  nand g1339 (n_1659, n_530, n_531);
  nand g1340 (n_1660, n_532, n_531);
  nand g1341 (n_1661, n_530, n_532);
  nand g1342 (n_107, n_1659, n_1660, n_1661);
  xor g1343 (n_1662, A[30], A[28]);
  xor g1344 (n_534, n_1662, A[16]);
  nand g1345 (n_1663, A[30], A[28]);
  nand g1347 (n_1665, A[30], A[16]);
  nand g1348 (n_547, n_1663, n_1601, n_1665);
  xor g1349 (n_1666, A[14], A[24]);
  xor g1350 (n_538, n_1666, A[22]);
  nand g1352 (n_1668, A[22], A[24]);
  nand g1353 (n_1669, A[14], A[22]);
  nand g1354 (n_549, n_1472, n_1668, n_1669);
  xor g1355 (n_1670, A[12], A[26]);
  xor g1356 (n_537, n_1670, A[20]);
  nand g1358 (n_1672, A[20], A[26]);
  nand g1360 (n_550, n_1605, n_1672, n_1539);
  xor g1361 (n_1674, A[18], n_533);
  xor g1362 (n_540, n_1674, n_534);
  nand g1363 (n_1675, A[18], n_533);
  nand g1364 (n_1676, n_534, n_533);
  nand g1365 (n_1677, A[18], n_534);
  nand g1366 (n_553, n_1675, n_1676, n_1677);
  xor g1367 (n_1678, n_535, n_536);
  xor g1368 (n_541, n_1678, n_537);
  nand g1369 (n_1679, n_535, n_536);
  nand g1370 (n_1680, n_537, n_536);
  nand g1371 (n_1681, n_535, n_537);
  nand g1372 (n_556, n_1679, n_1680, n_1681);
  xor g1373 (n_1682, n_538, n_539);
  xor g1374 (n_544, n_1682, n_540);
  nand g1375 (n_1683, n_538, n_539);
  nand g1376 (n_1684, n_540, n_539);
  nand g1377 (n_1685, n_538, n_540);
  nand g1378 (n_557, n_1683, n_1684, n_1685);
  xor g1379 (n_1686, n_541, n_542);
  xor g1380 (n_545, n_1686, n_543);
  nand g1381 (n_1687, n_541, n_542);
  nand g1382 (n_1688, n_543, n_542);
  nand g1383 (n_1689, n_541, n_543);
  nand g1384 (n_560, n_1687, n_1688, n_1689);
  xor g1385 (n_1690, n_544, n_545);
  xor g1386 (n_185, n_1690, n_546);
  nand g1387 (n_1691, n_544, n_545);
  nand g1388 (n_1692, n_546, n_545);
  nand g1389 (n_1693, n_544, n_546);
  nand g1390 (n_106, n_1691, n_1692, n_1693);
  xor g1391 (n_1694, A[31], A[29]);
  xor g1392 (n_548, n_1694, A[17]);
  nand g1393 (n_1695, A[31], A[29]);
  nand g1395 (n_1697, A[31], A[17]);
  nand g1396 (n_561, n_1695, n_1633, n_1697);
  xor g1397 (n_1698, A[15], A[25]);
  xor g1398 (n_552, n_1698, A[23]);
  nand g1400 (n_1700, A[23], A[25]);
  nand g1401 (n_1701, A[15], A[23]);
  nand g1402 (n_563, n_1504, n_1700, n_1701);
  xor g1403 (n_1702, A[13], A[27]);
  xor g1404 (n_551, n_1702, A[21]);
  nand g1406 (n_1704, A[21], A[27]);
  nand g1408 (n_564, n_1637, n_1704, n_1571);
  xor g1409 (n_1706, A[19], n_547);
  xor g1410 (n_554, n_1706, n_548);
  nand g1411 (n_1707, A[19], n_547);
  nand g1412 (n_1708, n_548, n_547);
  nand g1413 (n_1709, A[19], n_548);
  nand g1414 (n_567, n_1707, n_1708, n_1709);
  xor g1415 (n_1710, n_549, n_550);
  xor g1416 (n_555, n_1710, n_551);
  nand g1417 (n_1711, n_549, n_550);
  nand g1418 (n_1712, n_551, n_550);
  nand g1419 (n_1713, n_549, n_551);
  nand g1420 (n_570, n_1711, n_1712, n_1713);
  xor g1421 (n_1714, n_552, n_553);
  xor g1422 (n_558, n_1714, n_554);
  nand g1423 (n_1715, n_552, n_553);
  nand g1424 (n_1716, n_554, n_553);
  nand g1425 (n_1717, n_552, n_554);
  nand g1426 (n_571, n_1715, n_1716, n_1717);
  xor g1427 (n_1718, n_555, n_556);
  xor g1428 (n_559, n_1718, n_557);
  nand g1429 (n_1719, n_555, n_556);
  nand g1430 (n_1720, n_557, n_556);
  nand g1431 (n_1721, n_555, n_557);
  nand g1432 (n_574, n_1719, n_1720, n_1721);
  xor g1433 (n_1722, n_558, n_559);
  xor g1434 (n_184, n_1722, n_560);
  nand g1435 (n_1723, n_558, n_559);
  nand g1436 (n_1724, n_560, n_559);
  nand g1437 (n_1725, n_558, n_560);
  nand g1438 (n_105, n_1723, n_1724, n_1725);
  xor g1439 (n_1726, A[30], A[16]);
  xor g1440 (n_562, n_1726, A[14]);
  nand g1443 (n_1729, A[30], A[14]);
  xor g1445 (n_1730, A[28], A[32]);
  xor g1446 (n_565, n_1730, A[18]);
  nand g1447 (n_1731, A[28], A[32]);
  nand g1448 (n_1732, A[18], A[32]);
  nand g1449 (n_1733, A[28], A[18]);
  nand g1450 (n_577, n_1731, n_1732, n_1733);
  xor g1451 (n_1734, A[26], A[24]);
  xor g1452 (n_566, n_1734, A[22]);
  nand g1453 (n_1735, A[26], A[24]);
  nand g1456 (n_578, n_1735, n_1668, n_1603);
  xor g1457 (n_1738, A[20], n_561);
  xor g1458 (n_568, n_1738, n_562);
  nand g1459 (n_1739, A[20], n_561);
  nand g1460 (n_1740, n_562, n_561);
  nand g1461 (n_1741, A[20], n_562);
  nand g1462 (n_581, n_1739, n_1740, n_1741);
  xor g1463 (n_1742, n_563, n_564);
  xor g1464 (n_569, n_1742, n_565);
  nand g1465 (n_1743, n_563, n_564);
  nand g1466 (n_1744, n_565, n_564);
  nand g1467 (n_1745, n_563, n_565);
  nand g1468 (n_584, n_1743, n_1744, n_1745);
  xor g1469 (n_1746, n_566, n_567);
  xor g1470 (n_572, n_1746, n_568);
  nand g1471 (n_1747, n_566, n_567);
  nand g1472 (n_1748, n_568, n_567);
  nand g1473 (n_1749, n_566, n_568);
  nand g1474 (n_585, n_1747, n_1748, n_1749);
  xor g1475 (n_1750, n_569, n_570);
  xor g1476 (n_573, n_1750, n_571);
  nand g1477 (n_1751, n_569, n_570);
  nand g1478 (n_1752, n_571, n_570);
  nand g1479 (n_1753, n_569, n_571);
  nand g1480 (n_588, n_1751, n_1752, n_1753);
  xor g1481 (n_1754, n_572, n_573);
  xor g1482 (n_183, n_1754, n_574);
  nand g1483 (n_1755, n_572, n_573);
  nand g1484 (n_1756, n_574, n_573);
  nand g1485 (n_1757, n_572, n_574);
  nand g1486 (n_104, n_1755, n_1756, n_1757);
  xor g1487 (n_1758, A[31], A[17]);
  xor g1488 (n_576, n_1758, A[15]);
  nand g1491 (n_1761, A[31], A[15]);
  nand g1492 (n_589, n_1697, n_1256, n_1761);
  xor g1493 (n_1762, A[29], A[33]);
  xor g1494 (n_579, n_1762, A[19]);
  nand g1495 (n_1763, A[29], A[33]);
  nand g1496 (n_1764, A[19], A[33]);
  nand g1497 (n_1765, A[29], A[19]);
  nand g1498 (n_591, n_1763, n_1764, n_1765);
  xor g1499 (n_1766, A[27], A[25]);
  xor g1500 (n_580, n_1766, A[23]);
  nand g1501 (n_1767, A[27], A[25]);
  nand g1504 (n_592, n_1767, n_1700, n_1635);
  xor g1505 (n_1770, A[21], n_575);
  xor g1506 (n_582, n_1770, n_576);
  nand g1507 (n_1771, A[21], n_575);
  nand g1508 (n_1772, n_576, n_575);
  nand g1509 (n_1773, A[21], n_576);
  nand g1510 (n_595, n_1771, n_1772, n_1773);
  xor g1511 (n_1774, n_577, n_578);
  xor g1512 (n_583, n_1774, n_579);
  nand g1513 (n_1775, n_577, n_578);
  nand g1514 (n_1776, n_579, n_578);
  nand g1515 (n_1777, n_577, n_579);
  nand g1516 (n_598, n_1775, n_1776, n_1777);
  xor g1517 (n_1778, n_580, n_581);
  xor g1518 (n_586, n_1778, n_582);
  nand g1519 (n_1779, n_580, n_581);
  nand g1520 (n_1780, n_582, n_581);
  nand g1521 (n_1781, n_580, n_582);
  nand g1522 (n_599, n_1779, n_1780, n_1781);
  xor g1523 (n_1782, n_583, n_584);
  xor g1524 (n_587, n_1782, n_585);
  nand g1525 (n_1783, n_583, n_584);
  nand g1526 (n_1784, n_585, n_584);
  nand g1527 (n_1785, n_583, n_585);
  nand g1528 (n_602, n_1783, n_1784, n_1785);
  xor g1529 (n_1786, n_586, n_587);
  xor g1530 (n_182, n_1786, n_588);
  nand g1531 (n_1787, n_586, n_587);
  nand g1532 (n_1788, n_588, n_587);
  nand g1533 (n_1789, n_586, n_588);
  nand g1534 (n_103, n_1787, n_1788, n_1789);
  xor g1541 (n_1794, A[32], A[20]);
  xor g1542 (n_594, n_1794, A[18]);
  nand g1543 (n_1795, A[32], A[20]);
  nand g1546 (n_605, n_1795, n_1609, n_1732);
  xor g1547 (n_1798, A[26], A[34]);
  xor g1548 (n_593, n_1798, A[24]);
  nand g1549 (n_1799, A[26], A[34]);
  nand g1550 (n_1800, A[24], A[34]);
  nand g1552 (n_606, n_1799, n_1800, n_1735);
  xor g1553 (n_1802, A[22], n_589);
  xor g1554 (n_596, n_1802, n_534);
  nand g1555 (n_1803, A[22], n_589);
  nand g1556 (n_1804, n_534, n_589);
  nand g1557 (n_1805, A[22], n_534);
  nand g1558 (n_609, n_1803, n_1804, n_1805);
  xor g1559 (n_1806, n_591, n_592);
  xor g1560 (n_597, n_1806, n_593);
  nand g1561 (n_1807, n_591, n_592);
  nand g1562 (n_1808, n_593, n_592);
  nand g1563 (n_1809, n_591, n_593);
  nand g1564 (n_612, n_1807, n_1808, n_1809);
  xor g1565 (n_1810, n_594, n_595);
  xor g1566 (n_600, n_1810, n_596);
  nand g1567 (n_1811, n_594, n_595);
  nand g1568 (n_1812, n_596, n_595);
  nand g1569 (n_1813, n_594, n_596);
  nand g1570 (n_613, n_1811, n_1812, n_1813);
  xor g1571 (n_1814, n_597, n_598);
  xor g1572 (n_601, n_1814, n_599);
  nand g1573 (n_1815, n_597, n_598);
  nand g1574 (n_1816, n_599, n_598);
  nand g1575 (n_1817, n_597, n_599);
  nand g1576 (n_616, n_1815, n_1816, n_1817);
  xor g1577 (n_1818, n_600, n_601);
  xor g1578 (n_181, n_1818, n_602);
  nand g1579 (n_1819, n_600, n_601);
  nand g1580 (n_1820, n_602, n_601);
  nand g1581 (n_1821, n_600, n_602);
  nand g1582 (n_102, n_1819, n_1820, n_1821);
  xor g1589 (n_1826, A[33], A[21]);
  xor g1590 (n_608, n_1826, A[19]);
  nand g1591 (n_1827, A[33], A[21]);
  nand g1594 (n_619, n_1827, n_1641, n_1764);
  xor g1595 (n_1830, A[27], A[35]);
  xor g1596 (n_607, n_1830, A[25]);
  nand g1597 (n_1831, A[27], A[35]);
  nand g1598 (n_1832, A[25], A[35]);
  nand g1600 (n_620, n_1831, n_1832, n_1767);
  xor g1601 (n_1834, A[23], n_547);
  xor g1602 (n_610, n_1834, n_548);
  nand g1603 (n_1835, A[23], n_547);
  nand g1605 (n_1837, A[23], n_548);
  nand g1606 (n_623, n_1835, n_1708, n_1837);
  xor g1607 (n_1838, n_605, n_606);
  xor g1608 (n_611, n_1838, n_607);
  nand g1609 (n_1839, n_605, n_606);
  nand g1610 (n_1840, n_607, n_606);
  nand g1611 (n_1841, n_605, n_607);
  nand g1612 (n_626, n_1839, n_1840, n_1841);
  xor g1613 (n_1842, n_608, n_609);
  xor g1614 (n_614, n_1842, n_610);
  nand g1615 (n_1843, n_608, n_609);
  nand g1616 (n_1844, n_610, n_609);
  nand g1617 (n_1845, n_608, n_610);
  nand g1618 (n_627, n_1843, n_1844, n_1845);
  xor g1619 (n_1846, n_611, n_612);
  xor g1620 (n_615, n_1846, n_613);
  nand g1621 (n_1847, n_611, n_612);
  nand g1622 (n_1848, n_613, n_612);
  nand g1623 (n_1849, n_611, n_613);
  nand g1624 (n_630, n_1847, n_1848, n_1849);
  xor g1625 (n_1850, n_614, n_615);
  xor g1626 (n_180, n_1850, n_616);
  nand g1627 (n_1851, n_614, n_615);
  nand g1628 (n_1852, n_616, n_615);
  nand g1629 (n_1853, n_614, n_616);
  nand g1630 (n_101, n_1851, n_1852, n_1853);
  xor g1632 (n_618, n_1662, A[34]);
  nand g1634 (n_1856, A[34], A[28]);
  nand g1635 (n_1857, A[30], A[34]);
  nand g1636 (n_632, n_1663, n_1856, n_1857);
  xor g1637 (n_1858, A[22], A[20]);
  xor g1638 (n_622, n_1858, A[36]);
  nand g1640 (n_1860, A[36], A[20]);
  nand g1641 (n_1861, A[22], A[36]);
  nand g1642 (n_633, n_1481, n_1860, n_1861);
  xor g1643 (n_1862, A[18], A[32]);
  xor g1644 (n_621, n_1862, A[26]);
  nand g1646 (n_1864, A[26], A[32]);
  nand g1647 (n_1865, A[18], A[26]);
  nand g1648 (n_634, n_1732, n_1864, n_1865);
  xor g1649 (n_1866, A[24], n_561);
  xor g1650 (n_624, n_1866, n_618);
  nand g1651 (n_1867, A[24], n_561);
  nand g1652 (n_1868, n_618, n_561);
  nand g1653 (n_1869, A[24], n_618);
  nand g1654 (n_637, n_1867, n_1868, n_1869);
  xor g1655 (n_1870, n_619, n_620);
  xor g1656 (n_625, n_1870, n_621);
  nand g1657 (n_1871, n_619, n_620);
  nand g1658 (n_1872, n_621, n_620);
  nand g1659 (n_1873, n_619, n_621);
  nand g1660 (n_639, n_1871, n_1872, n_1873);
  xor g1661 (n_1874, n_622, n_623);
  xor g1662 (n_628, n_1874, n_624);
  nand g1663 (n_1875, n_622, n_623);
  nand g1664 (n_1876, n_624, n_623);
  nand g1665 (n_1877, n_622, n_624);
  nand g1666 (n_641, n_1875, n_1876, n_1877);
  xor g1667 (n_1878, n_625, n_626);
  xor g1668 (n_629, n_1878, n_627);
  nand g1669 (n_1879, n_625, n_626);
  nand g1670 (n_1880, n_627, n_626);
  nand g1671 (n_1881, n_625, n_627);
  nand g1672 (n_644, n_1879, n_1880, n_1881);
  xor g1673 (n_1882, n_628, n_629);
  xor g1674 (n_179, n_1882, n_630);
  nand g1675 (n_1883, n_628, n_629);
  nand g1676 (n_1884, n_630, n_629);
  nand g1677 (n_1885, n_628, n_630);
  nand g1678 (n_100, n_1883, n_1884, n_1885);
  xor g1680 (n_631, n_1694, A[35]);
  nand g1682 (n_1888, A[35], A[29]);
  nand g1683 (n_1889, A[31], A[35]);
  nand g1684 (n_646, n_1695, n_1888, n_1889);
  xor g1685 (n_1890, A[23], A[21]);
  xor g1686 (n_636, n_1890, A[37]);
  nand g1688 (n_1892, A[37], A[21]);
  nand g1689 (n_1893, A[23], A[37]);
  nand g1690 (n_647, n_1513, n_1892, n_1893);
  xor g1691 (n_1894, A[19], A[33]);
  xor g1692 (n_635, n_1894, A[27]);
  nand g1694 (n_1896, A[27], A[33]);
  nand g1695 (n_1897, A[19], A[27]);
  nand g1696 (n_648, n_1764, n_1896, n_1897);
  xor g1697 (n_1898, A[25], n_631);
  xor g1698 (n_640, n_1898, n_632);
  nand g1699 (n_1899, A[25], n_631);
  nand g1700 (n_1900, n_632, n_631);
  nand g1701 (n_1901, A[25], n_632);
  nand g1702 (n_651, n_1899, n_1900, n_1901);
  xor g1703 (n_1902, n_633, n_634);
  xor g1704 (n_638, n_1902, n_635);
  nand g1705 (n_1903, n_633, n_634);
  nand g1706 (n_1904, n_635, n_634);
  nand g1707 (n_1905, n_633, n_635);
  nand g1708 (n_652, n_1903, n_1904, n_1905);
  xor g1709 (n_1906, n_636, n_637);
  xor g1710 (n_642, n_1906, n_638);
  nand g1711 (n_1907, n_636, n_637);
  nand g1712 (n_1908, n_638, n_637);
  nand g1713 (n_1909, n_636, n_638);
  nand g1714 (n_655, n_1907, n_1908, n_1909);
  xor g1715 (n_1910, n_639, n_640);
  xor g1716 (n_643, n_1910, n_641);
  nand g1717 (n_1911, n_639, n_640);
  nand g1718 (n_1912, n_641, n_640);
  nand g1719 (n_1913, n_639, n_641);
  nand g1720 (n_657, n_1911, n_1912, n_1913);
  xor g1721 (n_1914, n_642, n_643);
  xor g1722 (n_178, n_1914, n_644);
  nand g1723 (n_1915, n_642, n_643);
  nand g1724 (n_1916, n_644, n_643);
  nand g1725 (n_1917, n_642, n_644);
  nand g1726 (n_99, n_1915, n_1916, n_1917);
  xor g1728 (n_645, n_1662, A[38]);
  nand g1730 (n_1920, A[38], A[28]);
  nand g1731 (n_1921, A[30], A[38]);
  nand g1732 (n_660, n_1663, n_1920, n_1921);
  xor g1733 (n_1922, A[32], A[24]);
  xor g1734 (n_649, n_1922, A[22]);
  nand g1735 (n_1923, A[32], A[24]);
  nand g1737 (n_1925, A[32], A[22]);
  nand g1738 (n_661, n_1923, n_1668, n_1925);
  xor g1739 (n_1926, A[36], A[20]);
  xor g1740 (n_650, n_1926, A[34]);
  nand g1742 (n_1928, A[34], A[20]);
  nand g1743 (n_1929, A[36], A[34]);
  nand g1744 (n_662, n_1860, n_1928, n_1929);
  xor g1745 (n_1930, A[26], n_645);
  xor g1746 (n_654, n_1930, n_646);
  nand g1747 (n_1931, A[26], n_645);
  nand g1748 (n_1932, n_646, n_645);
  nand g1749 (n_1933, A[26], n_646);
  nand g1750 (n_665, n_1931, n_1932, n_1933);
  xor g1751 (n_1934, n_647, n_648);
  xor g1752 (n_653, n_1934, n_649);
  nand g1753 (n_1935, n_647, n_648);
  nand g1754 (n_1936, n_649, n_648);
  nand g1755 (n_1937, n_647, n_649);
  nand g1756 (n_666, n_1935, n_1936, n_1937);
  xor g1757 (n_1938, n_650, n_651);
  xor g1758 (n_656, n_1938, n_652);
  nand g1759 (n_1939, n_650, n_651);
  nand g1760 (n_1940, n_652, n_651);
  nand g1761 (n_1941, n_650, n_652);
  nand g1762 (n_669, n_1939, n_1940, n_1941);
  xor g1763 (n_1942, n_653, n_654);
  xor g1764 (n_658, n_1942, n_655);
  nand g1765 (n_1943, n_653, n_654);
  nand g1766 (n_1944, n_655, n_654);
  nand g1767 (n_1945, n_653, n_655);
  nand g1768 (n_672, n_1943, n_1944, n_1945);
  xor g1769 (n_1946, n_656, n_657);
  xor g1770 (n_177, n_1946, n_658);
  nand g1771 (n_1947, n_656, n_657);
  nand g1772 (n_1948, n_658, n_657);
  nand g1773 (n_1949, n_656, n_658);
  nand g1774 (n_98, n_1947, n_1948, n_1949);
  xor g1776 (n_659, n_1694, A[39]);
  nand g1778 (n_1952, A[39], A[29]);
  nand g1779 (n_1953, A[31], A[39]);
  nand g1780 (n_674, n_1695, n_1952, n_1953);
  xor g1781 (n_1954, A[33], A[25]);
  xor g1782 (n_663, n_1954, A[23]);
  nand g1783 (n_1955, A[33], A[25]);
  nand g1785 (n_1957, A[33], A[23]);
  nand g1786 (n_675, n_1955, n_1700, n_1957);
  xor g1787 (n_1958, A[37], A[21]);
  xor g1788 (n_664, n_1958, A[35]);
  nand g1790 (n_1960, A[35], A[21]);
  nand g1791 (n_1961, A[37], A[35]);
  nand g1792 (n_676, n_1892, n_1960, n_1961);
  xor g1793 (n_1962, A[27], n_659);
  xor g1794 (n_668, n_1962, n_660);
  nand g1795 (n_1963, A[27], n_659);
  nand g1796 (n_1964, n_660, n_659);
  nand g1797 (n_1965, A[27], n_660);
  nand g1798 (n_679, n_1963, n_1964, n_1965);
  xor g1799 (n_1966, n_661, n_662);
  xor g1800 (n_667, n_1966, n_663);
  nand g1801 (n_1967, n_661, n_662);
  nand g1802 (n_1968, n_663, n_662);
  nand g1803 (n_1969, n_661, n_663);
  nand g1804 (n_680, n_1967, n_1968, n_1969);
  xor g1805 (n_1970, n_664, n_665);
  xor g1806 (n_670, n_1970, n_666);
  nand g1807 (n_1971, n_664, n_665);
  nand g1808 (n_1972, n_666, n_665);
  nand g1809 (n_1973, n_664, n_666);
  nand g1810 (n_683, n_1971, n_1972, n_1973);
  xor g1811 (n_1974, n_667, n_668);
  xor g1812 (n_671, n_1974, n_669);
  nand g1813 (n_1975, n_667, n_668);
  nand g1814 (n_1976, n_669, n_668);
  nand g1815 (n_1977, n_667, n_669);
  nand g1816 (n_686, n_1975, n_1976, n_1977);
  xor g1817 (n_1978, n_670, n_671);
  xor g1818 (n_176, n_1978, n_672);
  nand g1819 (n_1979, n_670, n_671);
  nand g1820 (n_1980, n_672, n_671);
  nand g1821 (n_1981, n_670, n_672);
  nand g1822 (n_97, n_1979, n_1980, n_1981);
  xor g1835 (n_1990, A[32], A[22]);
  xor g1836 (n_678, n_1990, A[36]);
  nand g1839 (n_1993, A[32], A[36]);
  nand g1840 (n_690, n_1925, n_1861, n_1993);
  xor g1841 (n_1994, A[40], n_645);
  xor g1842 (n_682, n_1994, n_674);
  nand g1843 (n_1995, A[40], n_645);
  nand g1844 (n_1996, n_674, n_645);
  nand g1845 (n_1997, A[40], n_674);
  nand g1846 (n_693, n_1995, n_1996, n_1997);
  xor g1847 (n_1998, n_675, n_676);
  xor g1848 (n_681, n_1998, n_593);
  nand g1849 (n_1999, n_675, n_676);
  nand g1850 (n_2000, n_593, n_676);
  nand g1851 (n_2001, n_675, n_593);
  nand g1852 (n_694, n_1999, n_2000, n_2001);
  xor g1853 (n_2002, n_678, n_679);
  xor g1854 (n_684, n_2002, n_680);
  nand g1855 (n_2003, n_678, n_679);
  nand g1856 (n_2004, n_680, n_679);
  nand g1857 (n_2005, n_678, n_680);
  nand g1858 (n_697, n_2003, n_2004, n_2005);
  xor g1859 (n_2006, n_681, n_682);
  xor g1860 (n_685, n_2006, n_683);
  nand g1861 (n_2007, n_681, n_682);
  nand g1862 (n_2008, n_683, n_682);
  nand g1863 (n_2009, n_681, n_683);
  nand g1864 (n_700, n_2007, n_2008, n_2009);
  xor g1865 (n_2010, n_684, n_685);
  xor g1866 (n_175, n_2010, n_686);
  nand g1867 (n_2011, n_684, n_685);
  nand g1868 (n_2012, n_686, n_685);
  nand g1869 (n_2013, n_684, n_686);
  nand g1870 (n_96, n_2011, n_2012, n_2013);
  xor g1883 (n_2022, A[33], A[23]);
  xor g1884 (n_692, n_2022, A[37]);
  nand g1887 (n_2025, A[33], A[37]);
  nand g1888 (n_704, n_1957, n_1893, n_2025);
  xor g1889 (n_2026, A[41], n_659);
  xor g1890 (n_696, n_2026, n_660);
  nand g1891 (n_2027, A[41], n_659);
  nand g1893 (n_2029, A[41], n_660);
  nand g1894 (n_707, n_2027, n_1964, n_2029);
  xor g1895 (n_2030, n_606, n_690);
  xor g1896 (n_695, n_2030, n_607);
  nand g1897 (n_2031, n_606, n_690);
  nand g1898 (n_2032, n_607, n_690);
  nand g1900 (n_709, n_2031, n_2032, n_1840);
  xor g1901 (n_2034, n_692, n_693);
  xor g1902 (n_698, n_2034, n_694);
  nand g1903 (n_2035, n_692, n_693);
  nand g1904 (n_2036, n_694, n_693);
  nand g1905 (n_2037, n_692, n_694);
  nand g1906 (n_711, n_2035, n_2036, n_2037);
  xor g1907 (n_2038, n_695, n_696);
  xor g1908 (n_699, n_2038, n_697);
  nand g1909 (n_2039, n_695, n_696);
  nand g1910 (n_2040, n_697, n_696);
  nand g1911 (n_2041, n_695, n_697);
  nand g1912 (n_714, n_2039, n_2040, n_2041);
  xor g1913 (n_2042, n_698, n_699);
  xor g1914 (n_174, n_2042, n_700);
  nand g1915 (n_2043, n_698, n_699);
  nand g1916 (n_2044, n_700, n_699);
  nand g1917 (n_2045, n_698, n_700);
  nand g1918 (n_95, n_2043, n_2044, n_2045);
  xor g1920 (n_701, n_1662, A[40]);
  nand g1922 (n_2048, A[40], A[28]);
  nand g1923 (n_2049, A[30], A[40]);
  nand g1924 (n_716, n_1663, n_2048, n_2049);
  xor g1925 (n_2050, A[36], A[26]);
  xor g1926 (n_706, n_2050, A[34]);
  nand g1927 (n_2051, A[36], A[26]);
  nand g1930 (n_717, n_2051, n_1799, n_1929);
  xor g1931 (n_2054, A[24], A[42]);
  xor g1932 (n_705, n_2054, A[32]);
  nand g1933 (n_2055, A[24], A[42]);
  nand g1934 (n_2056, A[32], A[42]);
  nand g1936 (n_718, n_2055, n_2056, n_1923);
  xor g1937 (n_2058, A[38], n_701);
  xor g1938 (n_710, n_2058, n_674);
  nand g1939 (n_2059, A[38], n_701);
  nand g1940 (n_2060, n_674, n_701);
  nand g1941 (n_2061, A[38], n_674);
  nand g1942 (n_721, n_2059, n_2060, n_2061);
  xor g1943 (n_2062, n_620, n_704);
  xor g1944 (n_708, n_2062, n_705);
  nand g1945 (n_2063, n_620, n_704);
  nand g1946 (n_2064, n_705, n_704);
  nand g1947 (n_2065, n_620, n_705);
  nand g1948 (n_723, n_2063, n_2064, n_2065);
  xor g1949 (n_2066, n_706, n_707);
  xor g1950 (n_712, n_2066, n_708);
  nand g1951 (n_2067, n_706, n_707);
  nand g1952 (n_2068, n_708, n_707);
  nand g1953 (n_2069, n_706, n_708);
  nand g1954 (n_725, n_2067, n_2068, n_2069);
  xor g1955 (n_2070, n_709, n_710);
  xor g1956 (n_713, n_2070, n_711);
  nand g1957 (n_2071, n_709, n_710);
  nand g1958 (n_2072, n_711, n_710);
  nand g1959 (n_2073, n_709, n_711);
  nand g1960 (n_728, n_2071, n_2072, n_2073);
  xor g1961 (n_2074, n_712, n_713);
  xor g1962 (n_173, n_2074, n_714);
  nand g1963 (n_2075, n_712, n_713);
  nand g1964 (n_2076, n_714, n_713);
  nand g1965 (n_2077, n_712, n_714);
  nand g1966 (n_94, n_2075, n_2076, n_2077);
  xor g1968 (n_715, n_1694, A[41]);
  nand g1970 (n_2080, A[41], A[29]);
  nand g1971 (n_2081, A[31], A[41]);
  nand g1972 (n_730, n_1695, n_2080, n_2081);
  xor g1973 (n_2082, A[37], A[27]);
  xor g1974 (n_720, n_2082, A[35]);
  nand g1975 (n_2083, A[37], A[27]);
  nand g1978 (n_731, n_2083, n_1831, n_1961);
  xor g1979 (n_2086, A[25], A[43]);
  xor g1980 (n_719, n_2086, A[33]);
  nand g1981 (n_2087, A[25], A[43]);
  nand g1982 (n_2088, A[33], A[43]);
  nand g1984 (n_732, n_2087, n_2088, n_1955);
  xor g1985 (n_2090, A[39], n_715);
  xor g1986 (n_724, n_2090, n_716);
  nand g1987 (n_2091, A[39], n_715);
  nand g1988 (n_2092, n_716, n_715);
  nand g1989 (n_2093, A[39], n_716);
  nand g1990 (n_735, n_2091, n_2092, n_2093);
  xor g1991 (n_2094, n_717, n_718);
  xor g1992 (n_722, n_2094, n_719);
  nand g1993 (n_2095, n_717, n_718);
  nand g1994 (n_2096, n_719, n_718);
  nand g1995 (n_2097, n_717, n_719);
  nand g1996 (n_737, n_2095, n_2096, n_2097);
  xor g1997 (n_2098, n_720, n_721);
  xor g1998 (n_726, n_2098, n_722);
  nand g1999 (n_2099, n_720, n_721);
  nand g2000 (n_2100, n_722, n_721);
  nand g2001 (n_2101, n_720, n_722);
  nand g2002 (n_739, n_2099, n_2100, n_2101);
  xor g2003 (n_2102, n_723, n_724);
  xor g2004 (n_727, n_2102, n_725);
  nand g2005 (n_2103, n_723, n_724);
  nand g2006 (n_2104, n_725, n_724);
  nand g2007 (n_2105, n_723, n_725);
  nand g2008 (n_742, n_2103, n_2104, n_2105);
  xor g2009 (n_2106, n_726, n_727);
  xor g2010 (n_172, n_2106, n_728);
  nand g2011 (n_2107, n_726, n_727);
  nand g2012 (n_2108, n_728, n_727);
  nand g2013 (n_2109, n_726, n_728);
  nand g2014 (n_93, n_2107, n_2108, n_2109);
  xor g2016 (n_729, n_1662, A[44]);
  nand g2018 (n_2112, A[44], A[28]);
  nand g2019 (n_2113, A[30], A[44]);
  nand g2020 (n_744, n_1663, n_2112, n_2113);
  xor g2021 (n_2114, A[38], A[42]);
  xor g2022 (n_734, n_2114, A[36]);
  nand g2023 (n_2115, A[38], A[42]);
  nand g2024 (n_2116, A[36], A[42]);
  nand g2025 (n_2117, A[38], A[36]);
  nand g2026 (n_745, n_2115, n_2116, n_2117);
  xor g2027 (n_2118, A[26], A[40]);
  xor g2028 (n_733, n_2118, A[34]);
  nand g2029 (n_2119, A[26], A[40]);
  nand g2030 (n_2120, A[34], A[40]);
  nand g2032 (n_746, n_2119, n_2120, n_1799);
  xor g2033 (n_2122, A[32], n_729);
  xor g2034 (n_738, n_2122, n_730);
  nand g2035 (n_2123, A[32], n_729);
  nand g2036 (n_2124, n_730, n_729);
  nand g2037 (n_2125, A[32], n_730);
  nand g2038 (n_749, n_2123, n_2124, n_2125);
  xor g2039 (n_2126, n_731, n_732);
  xor g2040 (n_736, n_2126, n_733);
  nand g2041 (n_2127, n_731, n_732);
  nand g2042 (n_2128, n_733, n_732);
  nand g2043 (n_2129, n_731, n_733);
  nand g2044 (n_751, n_2127, n_2128, n_2129);
  xor g2045 (n_2130, n_734, n_735);
  xor g2046 (n_740, n_2130, n_736);
  nand g2047 (n_2131, n_734, n_735);
  nand g2048 (n_2132, n_736, n_735);
  nand g2049 (n_2133, n_734, n_736);
  nand g2050 (n_753, n_2131, n_2132, n_2133);
  xor g2051 (n_2134, n_737, n_738);
  xor g2052 (n_741, n_2134, n_739);
  nand g2053 (n_2135, n_737, n_738);
  nand g2054 (n_2136, n_739, n_738);
  nand g2055 (n_2137, n_737, n_739);
  nand g2056 (n_756, n_2135, n_2136, n_2137);
  xor g2057 (n_2138, n_740, n_741);
  xor g2058 (n_171, n_2138, n_742);
  nand g2059 (n_2139, n_740, n_741);
  nand g2060 (n_2140, n_742, n_741);
  nand g2061 (n_2141, n_740, n_742);
  nand g2062 (n_92, n_2139, n_2140, n_2141);
  xor g2064 (n_743, n_1694, A[45]);
  nand g2066 (n_2144, A[45], A[29]);
  nand g2067 (n_2145, A[31], A[45]);
  nand g2068 (n_758, n_1695, n_2144, n_2145);
  xor g2069 (n_2146, A[39], A[43]);
  xor g2070 (n_748, n_2146, A[37]);
  nand g2071 (n_2147, A[39], A[43]);
  nand g2072 (n_2148, A[37], A[43]);
  nand g2073 (n_2149, A[39], A[37]);
  nand g2074 (n_759, n_2147, n_2148, n_2149);
  xor g2075 (n_2150, A[27], A[41]);
  xor g2076 (n_747, n_2150, A[35]);
  nand g2077 (n_2151, A[27], A[41]);
  nand g2078 (n_2152, A[35], A[41]);
  nand g2080 (n_760, n_2151, n_2152, n_1831);
  xor g2081 (n_2154, A[33], n_743);
  xor g2082 (n_752, n_2154, n_744);
  nand g2083 (n_2155, A[33], n_743);
  nand g2084 (n_2156, n_744, n_743);
  nand g2085 (n_2157, A[33], n_744);
  nand g2086 (n_763, n_2155, n_2156, n_2157);
  xor g2087 (n_2158, n_745, n_746);
  xor g2088 (n_750, n_2158, n_747);
  nand g2089 (n_2159, n_745, n_746);
  nand g2090 (n_2160, n_747, n_746);
  nand g2091 (n_2161, n_745, n_747);
  nand g2092 (n_765, n_2159, n_2160, n_2161);
  xor g2093 (n_2162, n_748, n_749);
  xor g2094 (n_754, n_2162, n_750);
  nand g2095 (n_2163, n_748, n_749);
  nand g2096 (n_2164, n_750, n_749);
  nand g2097 (n_2165, n_748, n_750);
  nand g2098 (n_767, n_2163, n_2164, n_2165);
  xor g2099 (n_2166, n_751, n_752);
  xor g2100 (n_755, n_2166, n_753);
  nand g2101 (n_2167, n_751, n_752);
  nand g2102 (n_2168, n_753, n_752);
  nand g2103 (n_2169, n_751, n_753);
  nand g2104 (n_770, n_2167, n_2168, n_2169);
  xor g2105 (n_2170, n_754, n_755);
  xor g2106 (n_170, n_2170, n_756);
  nand g2107 (n_2171, n_754, n_755);
  nand g2108 (n_2172, n_756, n_755);
  nand g2109 (n_2173, n_754, n_756);
  nand g2110 (n_91, n_2171, n_2172, n_2173);
  xor g2117 (n_2178, A[32], A[40]);
  xor g2118 (n_762, n_2178, A[46]);
  nand g2119 (n_2179, A[32], A[40]);
  nand g2120 (n_2180, A[46], A[40]);
  nand g2121 (n_2181, A[32], A[46]);
  nand g2122 (n_773, n_2179, n_2180, n_2181);
  xor g2129 (n_2186, A[34], n_729);
  xor g2130 (n_766, n_2186, n_758);
  nand g2131 (n_2187, A[34], n_729);
  nand g2132 (n_2188, n_758, n_729);
  nand g2133 (n_2189, A[34], n_758);
  nand g2134 (n_777, n_2187, n_2188, n_2189);
  xor g2135 (n_2190, n_759, n_760);
  xor g2136 (n_764, n_2190, n_734);
  nand g2137 (n_2191, n_759, n_760);
  nand g2138 (n_2192, n_734, n_760);
  nand g2139 (n_2193, n_759, n_734);
  nand g2140 (n_779, n_2191, n_2192, n_2193);
  xor g2141 (n_2194, n_762, n_763);
  xor g2142 (n_768, n_2194, n_764);
  nand g2143 (n_2195, n_762, n_763);
  nand g2144 (n_2196, n_764, n_763);
  nand g2145 (n_2197, n_762, n_764);
  nand g2146 (n_781, n_2195, n_2196, n_2197);
  xor g2147 (n_2198, n_765, n_766);
  xor g2148 (n_769, n_2198, n_767);
  nand g2149 (n_2199, n_765, n_766);
  nand g2150 (n_2200, n_767, n_766);
  nand g2151 (n_2201, n_765, n_767);
  nand g2152 (n_784, n_2199, n_2200, n_2201);
  xor g2153 (n_2202, n_768, n_769);
  xor g2154 (n_169, n_2202, n_770);
  nand g2155 (n_2203, n_768, n_769);
  nand g2156 (n_2204, n_770, n_769);
  nand g2157 (n_2205, n_768, n_770);
  nand g2158 (n_90, n_2203, n_2204, n_2205);
  xor g2165 (n_2210, A[33], A[41]);
  xor g2166 (n_776, n_2210, A[47]);
  nand g2167 (n_2211, A[33], A[41]);
  nand g2168 (n_2212, A[47], A[41]);
  nand g2169 (n_2213, A[33], A[47]);
  nand g2170 (n_786, n_2211, n_2212, n_2213);
  xor g2177 (n_2218, A[35], n_743);
  xor g2178 (n_780, n_2218, n_744);
  nand g2179 (n_2219, A[35], n_743);
  nand g2181 (n_2221, A[35], n_744);
  nand g2182 (n_791, n_2219, n_2156, n_2221);
  xor g2183 (n_2222, n_773, n_745);
  xor g2184 (n_778, n_2222, n_748);
  nand g2185 (n_2223, n_773, n_745);
  nand g2186 (n_2224, n_748, n_745);
  nand g2187 (n_2225, n_773, n_748);
  nand g2188 (n_793, n_2223, n_2224, n_2225);
  xor g2189 (n_2226, n_776, n_777);
  xor g2190 (n_782, n_2226, n_778);
  nand g2191 (n_2227, n_776, n_777);
  nand g2192 (n_2228, n_778, n_777);
  nand g2193 (n_2229, n_776, n_778);
  nand g2194 (n_795, n_2227, n_2228, n_2229);
  xor g2195 (n_2230, n_779, n_780);
  xor g2196 (n_783, n_2230, n_781);
  nand g2197 (n_2231, n_779, n_780);
  nand g2198 (n_2232, n_781, n_780);
  nand g2199 (n_2233, n_779, n_781);
  nand g2200 (n_798, n_2231, n_2232, n_2233);
  xor g2201 (n_2234, n_782, n_783);
  xor g2202 (n_168, n_2234, n_784);
  nand g2203 (n_2235, n_782, n_783);
  nand g2204 (n_2236, n_784, n_783);
  nand g2205 (n_2237, n_782, n_784);
  nand g2206 (n_89, n_2235, n_2236, n_2237);
  xor g2207 (n_2238, A[30], A[48]);
  xor g2208 (n_789, n_2238, A[42]);
  nand g2209 (n_2239, A[30], A[48]);
  nand g2210 (n_2240, A[42], A[48]);
  nand g2211 (n_2241, A[30], A[42]);
  nand g2212 (n_799, n_2239, n_2240, n_2241);
  xor g2213 (n_2242, A[34], A[32]);
  xor g2214 (n_790, n_2242, A[46]);
  nand g2215 (n_2243, A[34], A[32]);
  nand g2217 (n_2245, A[34], A[46]);
  nand g2218 (n_800, n_2243, n_2181, n_2245);
  xor g2219 (n_2246, A[40], A[44]);
  xor g2220 (n_788, n_2246, A[38]);
  nand g2221 (n_2247, A[40], A[44]);
  nand g2222 (n_2248, A[38], A[44]);
  nand g2223 (n_2249, A[40], A[38]);
  nand g2224 (n_801, n_2247, n_2248, n_2249);
  xor g2225 (n_2250, A[36], n_758);
  xor g2226 (n_792, n_2250, n_786);
  nand g2227 (n_2251, A[36], n_758);
  nand g2228 (n_2252, n_786, n_758);
  nand g2229 (n_2253, A[36], n_786);
  nand g2230 (n_805, n_2251, n_2252, n_2253);
  xor g2231 (n_2254, n_759, n_788);
  xor g2232 (n_794, n_2254, n_789);
  nand g2233 (n_2255, n_759, n_788);
  nand g2234 (n_2256, n_789, n_788);
  nand g2235 (n_2257, n_759, n_789);
  nand g2236 (n_807, n_2255, n_2256, n_2257);
  xor g2237 (n_2258, n_790, n_791);
  xor g2238 (n_796, n_2258, n_792);
  nand g2239 (n_2259, n_790, n_791);
  nand g2240 (n_2260, n_792, n_791);
  nand g2241 (n_2261, n_790, n_792);
  nand g2242 (n_809, n_2259, n_2260, n_2261);
  xor g2243 (n_2262, n_793, n_794);
  xor g2244 (n_797, n_2262, n_795);
  nand g2245 (n_2263, n_793, n_794);
  nand g2246 (n_2264, n_795, n_794);
  nand g2247 (n_2265, n_793, n_795);
  nand g2248 (n_812, n_2263, n_2264, n_2265);
  xor g2249 (n_2266, n_796, n_797);
  xor g2250 (n_167, n_2266, n_798);
  nand g2251 (n_2267, n_796, n_797);
  nand g2252 (n_2268, n_798, n_797);
  nand g2253 (n_2269, n_796, n_798);
  nand g2254 (n_88, n_2267, n_2268, n_2269);
  xor g2255 (n_2270, A[31], A[49]);
  xor g2256 (n_803, n_2270, A[43]);
  nand g2257 (n_2271, A[31], A[49]);
  nand g2258 (n_2272, A[43], A[49]);
  nand g2259 (n_2273, A[31], A[43]);
  nand g2260 (n_813, n_2271, n_2272, n_2273);
  xor g2261 (n_2274, A[35], A[33]);
  xor g2262 (n_804, n_2274, A[47]);
  nand g2263 (n_2275, A[35], A[33]);
  nand g2265 (n_2277, A[35], A[47]);
  nand g2266 (n_814, n_2275, n_2213, n_2277);
  xor g2267 (n_2278, A[41], A[45]);
  xor g2268 (n_802, n_2278, A[39]);
  nand g2269 (n_2279, A[41], A[45]);
  nand g2270 (n_2280, A[39], A[45]);
  nand g2271 (n_2281, A[41], A[39]);
  nand g2272 (n_815, n_2279, n_2280, n_2281);
  xor g2273 (n_2282, A[37], n_799);
  xor g2274 (n_806, n_2282, n_800);
  nand g2275 (n_2283, A[37], n_799);
  nand g2276 (n_2284, n_800, n_799);
  nand g2277 (n_2285, A[37], n_800);
  nand g2278 (n_819, n_2283, n_2284, n_2285);
  xor g2279 (n_2286, n_801, n_802);
  xor g2280 (n_808, n_2286, n_803);
  nand g2281 (n_2287, n_801, n_802);
  nand g2282 (n_2288, n_803, n_802);
  nand g2283 (n_2289, n_801, n_803);
  nand g2284 (n_821, n_2287, n_2288, n_2289);
  xor g2285 (n_2290, n_804, n_805);
  xor g2286 (n_810, n_2290, n_806);
  nand g2287 (n_2291, n_804, n_805);
  nand g2288 (n_2292, n_806, n_805);
  nand g2289 (n_2293, n_804, n_806);
  nand g2290 (n_823, n_2291, n_2292, n_2293);
  xor g2291 (n_2294, n_807, n_808);
  xor g2292 (n_811, n_2294, n_809);
  nand g2293 (n_2295, n_807, n_808);
  nand g2294 (n_2296, n_809, n_808);
  nand g2295 (n_2297, n_807, n_809);
  nand g2296 (n_826, n_2295, n_2296, n_2297);
  xor g2297 (n_2298, n_810, n_811);
  xor g2298 (n_166, n_2298, n_812);
  nand g2299 (n_2299, n_810, n_811);
  nand g2300 (n_2300, n_812, n_811);
  nand g2301 (n_2301, n_810, n_812);
  nand g2302 (n_87, n_2299, n_2300, n_2301);
  xor g2303 (n_2302, A[50], A[48]);
  xor g2304 (n_817, n_2302, A[44]);
  nand g2305 (n_2303, A[50], A[48]);
  nand g2306 (n_2304, A[44], A[48]);
  nand g2307 (n_2305, A[50], A[44]);
  nand g2308 (n_827, n_2303, n_2304, n_2305);
  xor g2309 (n_2306, A[36], A[34]);
  xor g2310 (n_818, n_2306, A[42]);
  nand g2312 (n_2308, A[42], A[34]);
  nand g2314 (n_828, n_1929, n_2308, n_2116);
  xor g2315 (n_2310, A[32], A[46]);
  xor g2316 (n_816, n_2310, A[40]);
  xor g2321 (n_2314, A[38], n_813);
  xor g2322 (n_820, n_2314, n_814);
  nand g2323 (n_2315, A[38], n_813);
  nand g2324 (n_2316, n_814, n_813);
  nand g2325 (n_2317, A[38], n_814);
  nand g2326 (n_833, n_2315, n_2316, n_2317);
  xor g2327 (n_2318, n_815, n_816);
  xor g2328 (n_822, n_2318, n_817);
  nand g2329 (n_2319, n_815, n_816);
  nand g2330 (n_2320, n_817, n_816);
  nand g2331 (n_2321, n_815, n_817);
  nand g2332 (n_835, n_2319, n_2320, n_2321);
  xor g2333 (n_2322, n_818, n_819);
  xor g2334 (n_824, n_2322, n_820);
  nand g2335 (n_2323, n_818, n_819);
  nand g2336 (n_2324, n_820, n_819);
  nand g2337 (n_2325, n_818, n_820);
  nand g2338 (n_837, n_2323, n_2324, n_2325);
  xor g2339 (n_2326, n_821, n_822);
  xor g2340 (n_825, n_2326, n_823);
  nand g2341 (n_2327, n_821, n_822);
  nand g2342 (n_2328, n_823, n_822);
  nand g2343 (n_2329, n_821, n_823);
  nand g2344 (n_840, n_2327, n_2328, n_2329);
  xor g2345 (n_2330, n_824, n_825);
  xor g2346 (n_165, n_2330, n_826);
  nand g2347 (n_2331, n_824, n_825);
  nand g2348 (n_2332, n_826, n_825);
  nand g2349 (n_2333, n_824, n_826);
  nand g2350 (n_86, n_2331, n_2332, n_2333);
  xor g2351 (n_2334, A[51], A[49]);
  xor g2352 (n_831, n_2334, A[45]);
  nand g2353 (n_2335, A[51], A[49]);
  nand g2354 (n_2336, A[45], A[49]);
  nand g2355 (n_2337, A[51], A[45]);
  nand g2356 (n_841, n_2335, n_2336, n_2337);
  xor g2357 (n_2338, A[37], A[35]);
  xor g2358 (n_832, n_2338, A[43]);
  nand g2360 (n_2340, A[43], A[35]);
  nand g2362 (n_842, n_1961, n_2340, n_2148);
  xor g2363 (n_2342, A[33], A[47]);
  xor g2364 (n_830, n_2342, A[41]);
  xor g2369 (n_2346, A[39], n_827);
  xor g2370 (n_834, n_2346, n_828);
  nand g2371 (n_2347, A[39], n_827);
  nand g2372 (n_2348, n_828, n_827);
  nand g2373 (n_2349, A[39], n_828);
  nand g2374 (n_847, n_2347, n_2348, n_2349);
  xor g2375 (n_2350, n_773, n_830);
  xor g2376 (n_836, n_2350, n_831);
  nand g2377 (n_2351, n_773, n_830);
  nand g2378 (n_2352, n_831, n_830);
  nand g2379 (n_2353, n_773, n_831);
  nand g2380 (n_849, n_2351, n_2352, n_2353);
  xor g2381 (n_2354, n_832, n_833);
  xor g2382 (n_838, n_2354, n_834);
  nand g2383 (n_2355, n_832, n_833);
  nand g2384 (n_2356, n_834, n_833);
  nand g2385 (n_2357, n_832, n_834);
  nand g2386 (n_851, n_2355, n_2356, n_2357);
  xor g2387 (n_2358, n_835, n_836);
  xor g2388 (n_839, n_2358, n_837);
  nand g2389 (n_2359, n_835, n_836);
  nand g2390 (n_2360, n_837, n_836);
  nand g2391 (n_2361, n_835, n_837);
  nand g2392 (n_854, n_2359, n_2360, n_2361);
  xor g2393 (n_2362, n_838, n_839);
  xor g2394 (n_164, n_2362, n_840);
  nand g2395 (n_2363, n_838, n_839);
  nand g2396 (n_2364, n_840, n_839);
  nand g2397 (n_2365, n_838, n_840);
  nand g2398 (n_85, n_2363, n_2364, n_2365);
  xor g2399 (n_2366, A[52], A[50]);
  xor g2400 (n_845, n_2366, A[46]);
  nand g2401 (n_2367, A[52], A[50]);
  nand g2402 (n_2368, A[46], A[50]);
  nand g2403 (n_2369, A[52], A[46]);
  nand g2404 (n_855, n_2367, n_2368, n_2369);
  xor g2405 (n_2370, A[38], A[36]);
  xor g2406 (n_846, n_2370, A[44]);
  nand g2408 (n_2372, A[44], A[36]);
  nand g2410 (n_856, n_2117, n_2372, n_2248);
  xor g2411 (n_2374, A[34], A[48]);
  xor g2412 (n_844, n_2374, A[42]);
  nand g2413 (n_2375, A[34], A[48]);
  nand g2416 (n_857, n_2375, n_2240, n_2308);
  xor g2417 (n_2378, A[40], n_841);
  xor g2418 (n_848, n_2378, n_842);
  nand g2419 (n_2379, A[40], n_841);
  nand g2420 (n_2380, n_842, n_841);
  nand g2421 (n_2381, A[40], n_842);
  nand g2422 (n_861, n_2379, n_2380, n_2381);
  xor g2423 (n_2382, n_786, n_844);
  xor g2424 (n_850, n_2382, n_845);
  nand g2425 (n_2383, n_786, n_844);
  nand g2426 (n_2384, n_845, n_844);
  nand g2427 (n_2385, n_786, n_845);
  nand g2428 (n_863, n_2383, n_2384, n_2385);
  xor g2429 (n_2386, n_846, n_847);
  xor g2430 (n_852, n_2386, n_848);
  nand g2431 (n_2387, n_846, n_847);
  nand g2432 (n_2388, n_848, n_847);
  nand g2433 (n_2389, n_846, n_848);
  nand g2434 (n_865, n_2387, n_2388, n_2389);
  xor g2435 (n_2390, n_849, n_850);
  xor g2436 (n_853, n_2390, n_851);
  nand g2437 (n_2391, n_849, n_850);
  nand g2438 (n_2392, n_851, n_850);
  nand g2439 (n_2393, n_849, n_851);
  nand g2440 (n_868, n_2391, n_2392, n_2393);
  xor g2441 (n_2394, n_852, n_853);
  xor g2442 (n_163, n_2394, n_854);
  nand g2443 (n_2395, n_852, n_853);
  nand g2444 (n_2396, n_854, n_853);
  nand g2445 (n_2397, n_852, n_854);
  nand g2446 (n_84, n_2395, n_2396, n_2397);
  xor g2447 (n_2398, A[53], A[51]);
  xor g2448 (n_859, n_2398, A[47]);
  nand g2449 (n_2399, A[53], A[51]);
  nand g2450 (n_2400, A[47], A[51]);
  nand g2451 (n_2401, A[53], A[47]);
  nand g2452 (n_869, n_2399, n_2400, n_2401);
  xor g2453 (n_2402, A[39], A[37]);
  xor g2454 (n_860, n_2402, A[45]);
  nand g2456 (n_2404, A[45], A[37]);
  nand g2458 (n_870, n_2149, n_2404, n_2280);
  xor g2459 (n_2406, A[35], A[49]);
  xor g2460 (n_858, n_2406, A[43]);
  nand g2461 (n_2407, A[35], A[49]);
  nand g2464 (n_871, n_2407, n_2272, n_2340);
  xor g2465 (n_2410, A[41], n_855);
  xor g2466 (n_862, n_2410, n_856);
  nand g2467 (n_2411, A[41], n_855);
  nand g2468 (n_2412, n_856, n_855);
  nand g2469 (n_2413, A[41], n_856);
  nand g2470 (n_875, n_2411, n_2412, n_2413);
  xor g2471 (n_2414, n_857, n_858);
  xor g2472 (n_864, n_2414, n_859);
  nand g2473 (n_2415, n_857, n_858);
  nand g2474 (n_2416, n_859, n_858);
  nand g2475 (n_2417, n_857, n_859);
  nand g2476 (n_877, n_2415, n_2416, n_2417);
  xor g2477 (n_2418, n_860, n_861);
  xor g2478 (n_866, n_2418, n_862);
  nand g2479 (n_2419, n_860, n_861);
  nand g2480 (n_2420, n_862, n_861);
  nand g2481 (n_2421, n_860, n_862);
  nand g2482 (n_879, n_2419, n_2420, n_2421);
  xor g2483 (n_2422, n_863, n_864);
  xor g2484 (n_867, n_2422, n_865);
  nand g2485 (n_2423, n_863, n_864);
  nand g2486 (n_2424, n_865, n_864);
  nand g2487 (n_2425, n_863, n_865);
  nand g2488 (n_882, n_2423, n_2424, n_2425);
  xor g2489 (n_2426, n_866, n_867);
  xor g2490 (n_162, n_2426, n_868);
  nand g2491 (n_2427, n_866, n_867);
  nand g2492 (n_2428, n_868, n_867);
  nand g2493 (n_2429, n_866, n_868);
  nand g2494 (n_83, n_2427, n_2428, n_2429);
  xor g2495 (n_2430, A[54], A[52]);
  xor g2496 (n_873, n_2430, A[48]);
  nand g2497 (n_2431, A[54], A[52]);
  nand g2498 (n_2432, A[48], A[52]);
  nand g2499 (n_2433, A[54], A[48]);
  nand g2500 (n_883, n_2431, n_2432, n_2433);
  xor g2501 (n_2434, A[40], A[38]);
  xor g2502 (n_874, n_2434, A[46]);
  nand g2504 (n_2436, A[46], A[38]);
  nand g2506 (n_884, n_2249, n_2436, n_2180);
  xor g2507 (n_2438, A[36], A[50]);
  xor g2508 (n_872, n_2438, A[44]);
  nand g2509 (n_2439, A[36], A[50]);
  nand g2512 (n_885, n_2439, n_2305, n_2372);
  xor g2513 (n_2442, A[42], n_869);
  xor g2514 (n_876, n_2442, n_870);
  nand g2515 (n_2443, A[42], n_869);
  nand g2516 (n_2444, n_870, n_869);
  nand g2517 (n_2445, A[42], n_870);
  nand g2518 (n_889, n_2443, n_2444, n_2445);
  xor g2519 (n_2446, n_871, n_872);
  xor g2520 (n_878, n_2446, n_873);
  nand g2521 (n_2447, n_871, n_872);
  nand g2522 (n_2448, n_873, n_872);
  nand g2523 (n_2449, n_871, n_873);
  nand g2524 (n_891, n_2447, n_2448, n_2449);
  xor g2525 (n_2450, n_874, n_875);
  xor g2526 (n_880, n_2450, n_876);
  nand g2527 (n_2451, n_874, n_875);
  nand g2528 (n_2452, n_876, n_875);
  nand g2529 (n_2453, n_874, n_876);
  nand g2530 (n_893, n_2451, n_2452, n_2453);
  xor g2531 (n_2454, n_877, n_878);
  xor g2532 (n_881, n_2454, n_879);
  nand g2533 (n_2455, n_877, n_878);
  nand g2534 (n_2456, n_879, n_878);
  nand g2535 (n_2457, n_877, n_879);
  nand g2536 (n_896, n_2455, n_2456, n_2457);
  xor g2537 (n_2458, n_880, n_881);
  xor g2538 (n_161, n_2458, n_882);
  nand g2539 (n_2459, n_880, n_881);
  nand g2540 (n_2460, n_882, n_881);
  nand g2541 (n_2461, n_880, n_882);
  nand g2542 (n_82, n_2459, n_2460, n_2461);
  xor g2543 (n_2462, A[55], A[53]);
  xor g2544 (n_887, n_2462, A[49]);
  nand g2545 (n_2463, A[55], A[53]);
  nand g2546 (n_2464, A[49], A[53]);
  nand g2547 (n_2465, A[55], A[49]);
  nand g2548 (n_897, n_2463, n_2464, n_2465);
  xor g2549 (n_2466, A[41], A[39]);
  xor g2550 (n_888, n_2466, A[47]);
  nand g2552 (n_2468, A[47], A[39]);
  nand g2554 (n_898, n_2281, n_2468, n_2212);
  xor g2555 (n_2470, A[37], A[51]);
  xor g2556 (n_886, n_2470, A[45]);
  nand g2557 (n_2471, A[37], A[51]);
  nand g2560 (n_899, n_2471, n_2337, n_2404);
  xor g2561 (n_2474, A[43], n_883);
  xor g2562 (n_890, n_2474, n_884);
  nand g2563 (n_2475, A[43], n_883);
  nand g2564 (n_2476, n_884, n_883);
  nand g2565 (n_2477, A[43], n_884);
  nand g2566 (n_903, n_2475, n_2476, n_2477);
  xor g2567 (n_2478, n_885, n_886);
  xor g2568 (n_892, n_2478, n_887);
  nand g2569 (n_2479, n_885, n_886);
  nand g2570 (n_2480, n_887, n_886);
  nand g2571 (n_2481, n_885, n_887);
  nand g2572 (n_905, n_2479, n_2480, n_2481);
  xor g2573 (n_2482, n_888, n_889);
  xor g2574 (n_894, n_2482, n_890);
  nand g2575 (n_2483, n_888, n_889);
  nand g2576 (n_2484, n_890, n_889);
  nand g2577 (n_2485, n_888, n_890);
  nand g2578 (n_907, n_2483, n_2484, n_2485);
  xor g2579 (n_2486, n_891, n_892);
  xor g2580 (n_895, n_2486, n_893);
  nand g2581 (n_2487, n_891, n_892);
  nand g2582 (n_2488, n_893, n_892);
  nand g2583 (n_2489, n_891, n_893);
  nand g2584 (n_910, n_2487, n_2488, n_2489);
  xor g2585 (n_2490, n_894, n_895);
  xor g2586 (n_160, n_2490, n_896);
  nand g2587 (n_2491, n_894, n_895);
  nand g2588 (n_2492, n_896, n_895);
  nand g2589 (n_2493, n_894, n_896);
  nand g2590 (n_81, n_2491, n_2492, n_2493);
  xor g2591 (n_2494, A[56], A[54]);
  xor g2592 (n_901, n_2494, A[50]);
  nand g2593 (n_2495, A[56], A[54]);
  nand g2594 (n_2496, A[50], A[54]);
  nand g2595 (n_2497, A[56], A[50]);
  nand g2596 (n_911, n_2495, n_2496, n_2497);
  xor g2597 (n_2498, A[42], A[40]);
  xor g2598 (n_902, n_2498, A[48]);
  nand g2599 (n_2499, A[42], A[40]);
  nand g2600 (n_2500, A[48], A[40]);
  nand g2602 (n_912, n_2499, n_2500, n_2240);
  xor g2603 (n_2502, A[38], A[52]);
  xor g2604 (n_900, n_2502, A[46]);
  nand g2605 (n_2503, A[38], A[52]);
  nand g2608 (n_913, n_2503, n_2369, n_2436);
  xor g2609 (n_2506, A[44], n_897);
  xor g2610 (n_904, n_2506, n_898);
  nand g2611 (n_2507, A[44], n_897);
  nand g2612 (n_2508, n_898, n_897);
  nand g2613 (n_2509, A[44], n_898);
  nand g2614 (n_917, n_2507, n_2508, n_2509);
  xor g2615 (n_2510, n_899, n_900);
  xor g2616 (n_906, n_2510, n_901);
  nand g2617 (n_2511, n_899, n_900);
  nand g2618 (n_2512, n_901, n_900);
  nand g2619 (n_2513, n_899, n_901);
  nand g2620 (n_919, n_2511, n_2512, n_2513);
  xor g2621 (n_2514, n_902, n_903);
  xor g2622 (n_908, n_2514, n_904);
  nand g2623 (n_2515, n_902, n_903);
  nand g2624 (n_2516, n_904, n_903);
  nand g2625 (n_2517, n_902, n_904);
  nand g2626 (n_921, n_2515, n_2516, n_2517);
  xor g2627 (n_2518, n_905, n_906);
  xor g2628 (n_909, n_2518, n_907);
  nand g2629 (n_2519, n_905, n_906);
  nand g2630 (n_2520, n_907, n_906);
  nand g2631 (n_2521, n_905, n_907);
  nand g2632 (n_924, n_2519, n_2520, n_2521);
  xor g2633 (n_2522, n_908, n_909);
  xor g2634 (n_159, n_2522, n_910);
  nand g2635 (n_2523, n_908, n_909);
  nand g2636 (n_2524, n_910, n_909);
  nand g2637 (n_2525, n_908, n_910);
  nand g2638 (n_80, n_2523, n_2524, n_2525);
  xor g2639 (n_2526, A[57], A[55]);
  xor g2640 (n_915, n_2526, A[51]);
  nand g2641 (n_2527, A[57], A[55]);
  nand g2642 (n_2528, A[51], A[55]);
  nand g2643 (n_2529, A[57], A[51]);
  nand g2644 (n_928, n_2527, n_2528, n_2529);
  xor g2645 (n_2530, A[43], A[41]);
  xor g2646 (n_916, n_2530, A[49]);
  nand g2647 (n_2531, A[43], A[41]);
  nand g2648 (n_2532, A[49], A[41]);
  nand g2650 (n_929, n_2531, n_2532, n_2272);
  xor g2651 (n_2534, A[39], A[53]);
  xor g2652 (n_914, n_2534, A[47]);
  nand g2653 (n_2535, A[39], A[53]);
  nand g2656 (n_927, n_2535, n_2401, n_2468);
  xor g2657 (n_2538, A[45], n_911);
  xor g2658 (n_918, n_2538, n_912);
  nand g2659 (n_2539, A[45], n_911);
  nand g2660 (n_2540, n_912, n_911);
  nand g2661 (n_2541, A[45], n_912);
  nand g2662 (n_933, n_2539, n_2540, n_2541);
  xor g2663 (n_2542, n_913, n_914);
  xor g2664 (n_920, n_2542, n_915);
  nand g2665 (n_2543, n_913, n_914);
  nand g2666 (n_2544, n_915, n_914);
  nand g2667 (n_2545, n_913, n_915);
  nand g2668 (n_935, n_2543, n_2544, n_2545);
  xor g2669 (n_2546, n_916, n_917);
  xor g2670 (n_922, n_2546, n_918);
  nand g2671 (n_2547, n_916, n_917);
  nand g2672 (n_2548, n_918, n_917);
  nand g2673 (n_2549, n_916, n_918);
  nand g2674 (n_937, n_2547, n_2548, n_2549);
  xor g2675 (n_2550, n_919, n_920);
  xor g2676 (n_923, n_2550, n_921);
  nand g2677 (n_2551, n_919, n_920);
  nand g2678 (n_2552, n_921, n_920);
  nand g2679 (n_2553, n_919, n_921);
  nand g2680 (n_940, n_2551, n_2552, n_2553);
  xor g2681 (n_2554, n_922, n_923);
  xor g2682 (n_158, n_2554, n_924);
  nand g2683 (n_2555, n_922, n_923);
  nand g2684 (n_2556, n_924, n_923);
  nand g2685 (n_2557, n_922, n_924);
  nand g2686 (n_79, n_2555, n_2556, n_2557);
  xor g2689 (n_2558, A[58], A[52]);
  xor g2690 (n_931, n_2558, A[44]);
  nand g2691 (n_2559, A[58], A[52]);
  nand g2692 (n_2560, A[44], A[52]);
  nand g2693 (n_2561, A[58], A[44]);
  nand g2694 (n_945, n_2559, n_2560, n_2561);
  xor g2695 (n_2562, A[42], A[56]);
  xor g2696 (n_932, n_2562, A[40]);
  nand g2697 (n_2563, A[42], A[56]);
  nand g2698 (n_2564, A[40], A[56]);
  nand g2700 (n_946, n_2563, n_2564, n_2499);
  xor g2701 (n_2566, A[50], A[54]);
  xor g2702 (n_930, n_2566, A[48]);
  nand g2706 (n_944, n_2496, n_2433, n_2303);
  xor g2707 (n_2570, A[46], n_927);
  xor g2708 (n_934, n_2570, n_928);
  nand g2709 (n_2571, A[46], n_927);
  nand g2710 (n_2572, n_928, n_927);
  nand g2711 (n_2573, A[46], n_928);
  nand g2712 (n_950, n_2571, n_2572, n_2573);
  xor g2713 (n_2574, n_929, n_930);
  xor g2714 (n_936, n_2574, n_931);
  nand g2715 (n_2575, n_929, n_930);
  nand g2716 (n_2576, n_931, n_930);
  nand g2717 (n_2577, n_929, n_931);
  nand g2718 (n_952, n_2575, n_2576, n_2577);
  xor g2719 (n_2578, n_932, n_933);
  xor g2720 (n_938, n_2578, n_934);
  nand g2721 (n_2579, n_932, n_933);
  nand g2722 (n_2580, n_934, n_933);
  nand g2723 (n_2581, n_932, n_934);
  nand g2724 (n_954, n_2579, n_2580, n_2581);
  xor g2725 (n_2582, n_935, n_936);
  xor g2726 (n_939, n_2582, n_937);
  nand g2727 (n_2583, n_935, n_936);
  nand g2728 (n_2584, n_937, n_936);
  nand g2729 (n_2585, n_935, n_937);
  nand g2730 (n_957, n_2583, n_2584, n_2585);
  xor g2731 (n_2586, n_938, n_939);
  xor g2732 (n_157, n_2586, n_940);
  nand g2733 (n_2587, n_938, n_939);
  nand g2734 (n_2588, n_940, n_939);
  nand g2735 (n_2589, n_938, n_940);
  nand g2736 (n_78, n_2587, n_2588, n_2589);
  xor g2739 (n_2590, A[51], A[43]);
  xor g2740 (n_948, n_2590, A[41]);
  nand g2741 (n_2591, A[51], A[43]);
  nand g2743 (n_2593, A[51], A[41]);
  nand g2744 (n_959, n_2591, n_2531, n_2593);
  xor g2745 (n_2594, A[58], A[57]);
  xor g2746 (n_949, n_2594, A[49]);
  nand g2747 (n_2595, A[58], A[57]);
  nand g2748 (n_2596, A[49], A[57]);
  nand g2749 (n_2597, A[58], A[49]);
  nand g2750 (n_960, n_2595, n_2596, n_2597);
  xor g2752 (n_947, n_2462, A[47]);
  nand g2755 (n_2601, A[55], A[47]);
  nand g2756 (n_961, n_2463, n_2401, n_2601);
  xor g2757 (n_2602, A[45], n_944);
  xor g2758 (n_951, n_2602, n_945);
  nand g2759 (n_2603, A[45], n_944);
  nand g2760 (n_2604, n_945, n_944);
  nand g2761 (n_2605, A[45], n_945);
  nand g2762 (n_965, n_2603, n_2604, n_2605);
  xor g2763 (n_2606, n_946, n_947);
  xor g2764 (n_953, n_2606, n_948);
  nand g2765 (n_2607, n_946, n_947);
  nand g2766 (n_2608, n_948, n_947);
  nand g2767 (n_2609, n_946, n_948);
  nand g2768 (n_967, n_2607, n_2608, n_2609);
  xor g2769 (n_2610, n_949, n_950);
  xor g2770 (n_955, n_2610, n_951);
  nand g2771 (n_2611, n_949, n_950);
  nand g2772 (n_2612, n_951, n_950);
  nand g2773 (n_2613, n_949, n_951);
  nand g2774 (n_969, n_2611, n_2612, n_2613);
  xor g2775 (n_2614, n_952, n_953);
  xor g2776 (n_956, n_2614, n_954);
  nand g2777 (n_2615, n_952, n_953);
  nand g2778 (n_2616, n_954, n_953);
  nand g2779 (n_2617, n_952, n_954);
  nand g2780 (n_972, n_2615, n_2616, n_2617);
  xor g2781 (n_2618, n_955, n_956);
  xor g2782 (n_156, n_2618, n_957);
  nand g2783 (n_2619, n_955, n_956);
  nand g2784 (n_2620, n_957, n_956);
  nand g2785 (n_2621, n_955, n_957);
  nand g2786 (n_77, n_2619, n_2620, n_2621);
  xor g2788 (n_963, n_2622, A[52]);
  nand g2790 (n_2624, A[52], A[56]);
  nand g2792 (n_975, n_2623, n_2624, n_2625);
  xor g2793 (n_2626, A[44], A[42]);
  xor g2794 (n_964, n_2626, A[50]);
  nand g2795 (n_2627, A[44], A[42]);
  nand g2796 (n_2628, A[50], A[42]);
  nand g2798 (n_976, n_2627, n_2628, n_2305);
  xor g2800 (n_962, n_2630, A[48]);
  nand g2804 (n_977, n_2631, n_2433, n_2633);
  xor g2805 (n_2634, A[46], n_959);
  xor g2806 (n_966, n_2634, n_960);
  nand g2807 (n_2635, A[46], n_959);
  nand g2808 (n_2636, n_960, n_959);
  nand g2809 (n_2637, A[46], n_960);
  nand g2810 (n_981, n_2635, n_2636, n_2637);
  xor g2811 (n_2638, n_961, n_962);
  xor g2812 (n_968, n_2638, n_963);
  nand g2813 (n_2639, n_961, n_962);
  nand g2814 (n_2640, n_963, n_962);
  nand g2815 (n_2641, n_961, n_963);
  nand g2816 (n_983, n_2639, n_2640, n_2641);
  xor g2817 (n_2642, n_964, n_965);
  xor g2818 (n_970, n_2642, n_966);
  nand g2819 (n_2643, n_964, n_965);
  nand g2820 (n_2644, n_966, n_965);
  nand g2821 (n_2645, n_964, n_966);
  nand g2822 (n_985, n_2643, n_2644, n_2645);
  xor g2823 (n_2646, n_967, n_968);
  xor g2824 (n_971, n_2646, n_969);
  nand g2825 (n_2647, n_967, n_968);
  nand g2826 (n_2648, n_969, n_968);
  nand g2827 (n_2649, n_967, n_969);
  nand g2828 (n_987, n_2647, n_2648, n_2649);
  xor g2829 (n_2650, n_970, n_971);
  xor g2830 (n_155, n_2650, n_972);
  nand g2831 (n_2651, n_970, n_971);
  nand g2832 (n_2652, n_972, n_971);
  nand g2833 (n_2653, n_970, n_972);
  nand g2834 (n_76, n_2651, n_2652, n_2653);
  xor g2837 (n_2654, A[55], A[43]);
  xor g2838 (n_979, n_2654, A[51]);
  nand g2839 (n_2655, A[55], A[43]);
  nand g2842 (n_990, n_2655, n_2591, n_2528);
  xor g2843 (n_2658, A[49], A[53]);
  xor g2844 (n_978, n_2658, A[47]);
  nand g2847 (n_2661, A[49], A[47]);
  nand g2848 (n_989, n_2464, n_2401, n_2661);
  xor g2850 (n_980, n_2662, n_975);
  nand g2853 (n_2665, A[45], n_975);
  nand g2854 (n_994, n_2663, n_2664, n_2665);
  xor g2855 (n_2666, n_976, n_977);
  xor g2856 (n_982, n_2666, n_978);
  nand g2857 (n_2667, n_976, n_977);
  nand g2858 (n_2668, n_978, n_977);
  nand g2859 (n_2669, n_976, n_978);
  nand g2860 (n_996, n_2667, n_2668, n_2669);
  xor g2861 (n_2670, n_979, n_980);
  xor g2862 (n_984, n_2670, n_981);
  nand g2863 (n_2671, n_979, n_980);
  nand g2864 (n_2672, n_981, n_980);
  nand g2865 (n_2673, n_979, n_981);
  nand g2866 (n_997, n_2671, n_2672, n_2673);
  xor g2867 (n_2674, n_982, n_983);
  xor g2868 (n_986, n_2674, n_984);
  nand g2869 (n_2675, n_982, n_983);
  nand g2870 (n_2676, n_984, n_983);
  nand g2871 (n_2677, n_982, n_984);
  nand g2872 (n_1000, n_2675, n_2676, n_2677);
  xor g2873 (n_2678, n_985, n_986);
  xor g2874 (n_154, n_2678, n_987);
  nand g2875 (n_2679, n_985, n_986);
  nand g2876 (n_2680, n_987, n_986);
  nand g2877 (n_2681, n_985, n_987);
  nand g2878 (n_75, n_2679, n_2680, n_2681);
  xor g2885 (n_2686, A[44], A[50]);
  xor g2886 (n_992, n_2686, A[54]);
  nand g2889 (n_2689, A[44], A[54]);
  nand g2890 (n_1004, n_2305, n_2496, n_2689);
  xor g2891 (n_2690, A[48], A[46]);
  xor g2892 (n_993, n_2690, A[57]);
  nand g2893 (n_2691, A[48], A[46]);
  nand g2894 (n_2692, A[57], A[46]);
  nand g2895 (n_2693, A[48], A[57]);
  nand g2896 (n_1007, n_2691, n_2692, n_2693);
  xor g2897 (n_2694, n_989, n_990);
  xor g2898 (n_995, n_2694, n_963);
  nand g2899 (n_2695, n_989, n_990);
  nand g2900 (n_2696, n_963, n_990);
  nand g2901 (n_2697, n_989, n_963);
  nand g2902 (n_1009, n_2695, n_2696, n_2697);
  xor g2903 (n_2698, n_992, n_993);
  xor g2904 (n_998, n_2698, n_994);
  nand g2905 (n_2699, n_992, n_993);
  nand g2906 (n_2700, n_994, n_993);
  nand g2907 (n_2701, n_992, n_994);
  nand g2908 (n_1011, n_2699, n_2700, n_2701);
  xor g2909 (n_2702, n_995, n_996);
  xor g2910 (n_999, n_2702, n_997);
  nand g2911 (n_2703, n_995, n_996);
  nand g2912 (n_2704, n_997, n_996);
  nand g2913 (n_2705, n_995, n_997);
  nand g2914 (n_1013, n_2703, n_2704, n_2705);
  xor g2915 (n_2706, n_998, n_999);
  xor g2916 (n_153, n_2706, n_1000);
  nand g2917 (n_2707, n_998, n_999);
  nand g2918 (n_2708, n_1000, n_999);
  nand g2919 (n_2709, n_998, n_1000);
  nand g2920 (n_152, n_2707, n_2708, n_2709);
  xor g2923 (n_2710, A[55], A[51]);
  xor g2924 (n_1006, n_2710, A[49]);
  nand g2928 (n_1015, n_2528, n_2335, n_2465);
  xor g2929 (n_2714, A[53], A[47]);
  xor g2930 (n_1005, n_2714, A[45]);
  nand g2932 (n_2716, A[45], A[47]);
  nand g2933 (n_2717, A[53], A[45]);
  nand g2934 (n_1016, n_2401, n_2716, n_2717);
  xor g2936 (n_1008, n_2718, n_1004);
  nand g2938 (n_2720, n_1004, n_975);
  nand g2940 (n_1020, n_2664, n_2720, n_2721);
  xor g2941 (n_2722, n_1005, n_1006);
  xor g2942 (n_1010, n_2722, n_1007);
  nand g2943 (n_2723, n_1005, n_1006);
  nand g2944 (n_2724, n_1007, n_1006);
  nand g2945 (n_2725, n_1005, n_1007);
  nand g2946 (n_1021, n_2723, n_2724, n_2725);
  xor g2947 (n_2726, n_1008, n_1009);
  xor g2948 (n_1012, n_2726, n_1010);
  nand g2949 (n_2727, n_1008, n_1009);
  nand g2950 (n_2728, n_1010, n_1009);
  nand g2951 (n_2729, n_1008, n_1010);
  nand g2952 (n_1024, n_2727, n_2728, n_2729);
  xor g2953 (n_2730, n_1011, n_1012);
  xor g2954 (n_74, n_2730, n_1013);
  nand g2955 (n_2731, n_1011, n_1012);
  nand g2956 (n_2732, n_1013, n_1012);
  nand g2957 (n_2733, n_1011, n_1013);
  nand g2958 (n_73, n_2731, n_2732, n_2733);
  xor g2971 (n_2742, A[46], A[57]);
  xor g2972 (n_1019, n_2742, n_1015);
  nand g2974 (n_2744, n_1015, A[57]);
  nand g2975 (n_2745, A[46], n_1015);
  nand g2976 (n_1031, n_2692, n_2744, n_2745);
  xor g2977 (n_2746, n_1016, n_930);
  xor g2978 (n_1022, n_2746, n_963);
  nand g2979 (n_2747, n_1016, n_930);
  nand g2980 (n_2748, n_963, n_930);
  nand g2981 (n_2749, n_1016, n_963);
  nand g2982 (n_1032, n_2747, n_2748, n_2749);
  xor g2983 (n_2750, n_1019, n_1020);
  xor g2984 (n_1023, n_2750, n_1021);
  nand g2985 (n_2751, n_1019, n_1020);
  nand g2986 (n_2752, n_1021, n_1020);
  nand g2987 (n_2753, n_1019, n_1021);
  nand g2988 (n_1035, n_2751, n_2752, n_2753);
  xor g2989 (n_2754, n_1022, n_1023);
  xor g2990 (n_151, n_2754, n_1024);
  nand g2991 (n_2755, n_1022, n_1023);
  nand g2992 (n_2756, n_1024, n_1023);
  nand g2993 (n_2757, n_1022, n_1024);
  nand g2994 (n_72, n_2755, n_2756, n_2757);
  xor g2998 (n_1029, n_2334, A[57]);
  nand g3002 (n_1037, n_2335, n_2596, n_2529);
  nand g3008 (n_1040, n_2401, n_2764, n_2765);
  xor g3009 (n_2766, n_944, n_975);
  xor g3010 (n_1033, n_2766, n_1029);
  nand g3011 (n_2767, n_944, n_975);
  nand g3012 (n_2768, n_1029, n_975);
  nand g3013 (n_2769, n_944, n_1029);
  nand g3014 (n_1042, n_2767, n_2768, n_2769);
  xor g3015 (n_2770, n_1030, n_1031);
  xor g3016 (n_1034, n_2770, n_1032);
  nand g3017 (n_2771, n_1030, n_1031);
  nand g3018 (n_2772, n_1032, n_1031);
  nand g3019 (n_2773, n_1030, n_1032);
  nand g3020 (n_1044, n_2771, n_2772, n_2773);
  xor g3021 (n_2774, n_1033, n_1034);
  xor g3022 (n_150, n_2774, n_1035);
  nand g3023 (n_2775, n_1033, n_1034);
  nand g3024 (n_2776, n_1035, n_1034);
  nand g3025 (n_2777, n_1033, n_1035);
  nand g3026 (n_71, n_2775, n_2776, n_2777);
  xor g3039 (n_2786, A[55], n_1037);
  xor g3040 (n_1041, n_2786, n_930);
  nand g3041 (n_2787, A[55], n_1037);
  nand g3042 (n_2788, n_930, n_1037);
  nand g3043 (n_2789, A[55], n_930);
  nand g3044 (n_1051, n_2787, n_2788, n_2789);
  xor g3045 (n_2790, n_963, n_1040);
  xor g3046 (n_1043, n_2790, n_1041);
  nand g3047 (n_2791, n_963, n_1040);
  nand g3048 (n_2792, n_1041, n_1040);
  nand g3049 (n_2793, n_963, n_1041);
  nand g3050 (n_1053, n_2791, n_2792, n_2793);
  xor g3051 (n_2794, n_1042, n_1043);
  xor g3052 (n_149, n_2794, n_1044);
  nand g3053 (n_2795, n_1042, n_1043);
  nand g3054 (n_2796, n_1044, n_1043);
  nand g3055 (n_2797, n_1042, n_1044);
  nand g3056 (n_70, n_2795, n_2796, n_2797);
  nand g3069 (n_2805, A[53], n_944);
  nand g3070 (n_1058, n_2764, n_2804, n_2805);
  xor g3071 (n_2806, n_975, n_1029);
  xor g3072 (n_1052, n_2806, n_1050);
  nand g3074 (n_2808, n_1050, n_1029);
  nand g3075 (n_2809, n_975, n_1050);
  nand g3076 (n_1060, n_2768, n_2808, n_2809);
  xor g3077 (n_2810, n_1051, n_1052);
  xor g3078 (n_148, n_2810, n_1053);
  nand g3079 (n_2811, n_1051, n_1052);
  nand g3080 (n_2812, n_1053, n_1052);
  nand g3081 (n_2813, n_1051, n_1053);
  nand g3082 (n_147, n_2811, n_2812, n_2813);
  xor g3090 (n_1057, n_2566, A[55]);
  nand g3092 (n_2820, A[55], A[54]);
  nand g3093 (n_2821, A[50], A[55]);
  nand g3094 (n_1065, n_2496, n_2820, n_2821);
  xor g3095 (n_2822, n_1037, n_963);
  xor g3096 (n_1059, n_2822, n_1057);
  nand g3097 (n_2823, n_1037, n_963);
  nand g3098 (n_2824, n_1057, n_963);
  nand g3099 (n_2825, n_1037, n_1057);
  nand g3100 (n_1067, n_2823, n_2824, n_2825);
  xor g3101 (n_2826, n_1058, n_1059);
  xor g3102 (n_69, n_2826, n_1060);
  nand g3103 (n_2827, n_1058, n_1059);
  nand g3104 (n_2828, n_1060, n_1059);
  nand g3105 (n_2829, n_1058, n_1060);
  nand g3106 (n_146, n_2827, n_2828, n_2829);
  xor g3110 (n_1064, n_2710, A[53]);
  nand g3114 (n_1069, n_2528, n_2463, n_2399);
  xor g3116 (n_1066, n_2718, n_1064);
  nand g3118 (n_2836, n_1064, n_975);
  nand g3120 (n_1072, n_2664, n_2836, n_2837);
  xor g3121 (n_2838, n_1065, n_1066);
  xor g3122 (n_68, n_2838, n_1067);
  nand g3123 (n_2839, n_1065, n_1066);
  nand g3124 (n_2840, n_1067, n_1066);
  nand g3125 (n_2841, n_1065, n_1067);
  nand g3126 (n_145, n_2839, n_2840, n_2841);
  xor g3133 (n_2846, A[54], A[57]);
  xor g3134 (n_1071, n_2846, n_1069);
  nand g3135 (n_2847, A[54], A[57]);
  nand g3136 (n_2848, n_1069, A[57]);
  nand g3137 (n_2849, A[54], n_1069);
  nand g3138 (n_1077, n_2847, n_2848, n_2849);
  xor g3139 (n_2850, n_963, n_1071);
  xor g3140 (n_67, n_2850, n_1072);
  nand g3141 (n_2851, n_963, n_1071);
  nand g3142 (n_2852, n_1072, n_1071);
  nand g3143 (n_2853, n_963, n_1072);
  nand g3144 (n_144, n_2851, n_2852, n_2853);
  nand g3152 (n_1080, n_2463, n_2856, n_2857);
  xor g3153 (n_2858, n_975, n_1076);
  xor g3154 (n_66, n_2858, n_1077);
  nand g3155 (n_2859, n_975, n_1076);
  nand g3156 (n_2860, n_1077, n_1076);
  nand g3157 (n_2861, n_975, n_1077);
  nand g3158 (n_143, n_2859, n_2860, n_2861);
  xor g3160 (n_1079, n_2622, A[54]);
  nand g3164 (n_1083, n_2623, n_2495, n_2631);
  xor g3165 (n_2866, A[57], n_1079);
  xor g3166 (n_65, n_2866, n_1080);
  nand g3167 (n_2867, A[57], n_1079);
  nand g3168 (n_2868, n_1080, n_1079);
  nand g3169 (n_2869, A[57], n_1080);
  nand g3170 (n_142, n_2867, n_2868, n_2869);
  nand g3177 (n_2873, A[57], n_1083);
  nand g3178 (n_141, n_2871, n_2872, n_2873);
  xor g3180 (n_63, n_2622, A[55]);
  nand g3182 (n_2876, A[55], A[56]);
  nand g3184 (n_140, n_2623, n_2876, n_2877);
  nor g11 (n_2893, A[2], A[0]);
  nor g13 (n_2889, A[1], A[3]);
  nor g15 (n_2899, A[2], n_211);
  nand g16 (n_2894, A[2], n_211);
  nor g17 (n_2895, n_132, n_210);
  nand g18 (n_2896, n_132, n_210);
  nor g19 (n_2905, n_131, n_209);
  nand g20 (n_2900, n_131, n_209);
  nor g21 (n_2901, n_130, n_208);
  nand g22 (n_2902, n_130, n_208);
  nor g23 (n_2911, n_129, n_207);
  nand g24 (n_2906, n_129, n_207);
  nor g25 (n_2907, n_128, n_206);
  nand g26 (n_2908, n_128, n_206);
  nor g27 (n_2917, n_127, n_205);
  nand g28 (n_2912, n_127, n_205);
  nor g29 (n_2913, n_126, n_204);
  nand g30 (n_2914, n_126, n_204);
  nor g31 (n_2923, n_125, n_203);
  nand g32 (n_2918, n_125, n_203);
  nor g33 (n_2919, n_124, n_202);
  nand g34 (n_2920, n_124, n_202);
  nor g35 (n_2929, n_123, n_201);
  nand g36 (n_2924, n_123, n_201);
  nor g37 (n_2925, n_122, n_200);
  nand g38 (n_2926, n_122, n_200);
  nor g39 (n_2935, n_121, n_199);
  nand g40 (n_2930, n_121, n_199);
  nor g41 (n_2931, n_120, n_198);
  nand g42 (n_2932, n_120, n_198);
  nor g43 (n_2941, n_119, n_197);
  nand g44 (n_2936, n_119, n_197);
  nor g45 (n_2937, n_118, n_196);
  nand g46 (n_2938, n_118, n_196);
  nor g47 (n_2947, n_117, n_195);
  nand g48 (n_2942, n_117, n_195);
  nor g49 (n_2943, n_116, n_194);
  nand g50 (n_2944, n_116, n_194);
  nor g51 (n_2953, n_115, n_193);
  nand g52 (n_2948, n_115, n_193);
  nor g53 (n_2949, n_114, n_192);
  nand g54 (n_2950, n_114, n_192);
  nor g55 (n_2959, n_113, n_191);
  nand g56 (n_2954, n_113, n_191);
  nor g57 (n_2955, n_112, n_190);
  nand g58 (n_2956, n_112, n_190);
  nor g59 (n_2965, n_111, n_189);
  nand g60 (n_2960, n_111, n_189);
  nor g61 (n_2961, n_110, n_188);
  nand g62 (n_2962, n_110, n_188);
  nor g63 (n_2971, n_109, n_187);
  nand g64 (n_2966, n_109, n_187);
  nor g65 (n_2967, n_108, n_186);
  nand g66 (n_2968, n_108, n_186);
  nor g67 (n_2977, n_107, n_185);
  nand g68 (n_2972, n_107, n_185);
  nor g69 (n_2973, n_106, n_184);
  nand g70 (n_2974, n_106, n_184);
  nor g71 (n_2983, n_105, n_183);
  nand g72 (n_2978, n_105, n_183);
  nor g73 (n_2979, n_104, n_182);
  nand g74 (n_2980, n_104, n_182);
  nor g75 (n_2989, n_103, n_181);
  nand g76 (n_2984, n_103, n_181);
  nor g77 (n_2985, n_102, n_180);
  nand g78 (n_2986, n_102, n_180);
  nor g79 (n_2995, n_101, n_179);
  nand g80 (n_2990, n_101, n_179);
  nor g81 (n_2991, n_100, n_178);
  nand g82 (n_2992, n_100, n_178);
  nor g83 (n_3001, n_99, n_177);
  nand g84 (n_2996, n_99, n_177);
  nor g85 (n_2997, n_98, n_176);
  nand g86 (n_2998, n_98, n_176);
  nor g87 (n_3007, n_97, n_175);
  nand g88 (n_3002, n_97, n_175);
  nor g89 (n_3003, n_96, n_174);
  nand g90 (n_3004, n_96, n_174);
  nor g91 (n_3013, n_95, n_173);
  nand g92 (n_3008, n_95, n_173);
  nor g93 (n_3009, n_94, n_172);
  nand g94 (n_3010, n_94, n_172);
  nor g95 (n_3019, n_93, n_171);
  nand g96 (n_3014, n_93, n_171);
  nor g97 (n_3015, n_92, n_170);
  nand g98 (n_3016, n_92, n_170);
  nor g99 (n_3025, n_91, n_169);
  nand g100 (n_3020, n_91, n_169);
  nor g101 (n_3021, n_90, n_168);
  nand g102 (n_3022, n_90, n_168);
  nor g103 (n_3031, n_89, n_167);
  nand g104 (n_3026, n_89, n_167);
  nor g105 (n_3027, n_88, n_166);
  nand g106 (n_3028, n_88, n_166);
  nor g107 (n_3037, n_87, n_165);
  nand g108 (n_3032, n_87, n_165);
  nor g109 (n_3033, n_86, n_164);
  nand g110 (n_3034, n_86, n_164);
  nor g111 (n_3043, n_85, n_163);
  nand g112 (n_3038, n_85, n_163);
  nor g113 (n_3039, n_84, n_162);
  nand g114 (n_3040, n_84, n_162);
  nor g115 (n_3049, n_83, n_161);
  nand g116 (n_3044, n_83, n_161);
  nor g117 (n_3045, n_82, n_160);
  nand g118 (n_3046, n_82, n_160);
  nor g119 (n_3055, n_81, n_159);
  nand g120 (n_3050, n_81, n_159);
  nor g121 (n_3051, n_80, n_158);
  nand g122 (n_3052, n_80, n_158);
  nor g123 (n_3061, n_79, n_157);
  nand g124 (n_3056, n_79, n_157);
  nor g125 (n_3057, n_78, n_156);
  nand g126 (n_3058, n_78, n_156);
  nor g127 (n_3067, n_77, n_155);
  nand g128 (n_3062, n_77, n_155);
  nor g129 (n_3063, n_76, n_154);
  nand g130 (n_3064, n_76, n_154);
  nor g131 (n_3073, n_75, n_153);
  nand g132 (n_3068, n_75, n_153);
  nor g133 (n_3069, n_74, n_152);
  nand g134 (n_3070, n_74, n_152);
  nor g135 (n_3079, n_73, n_151);
  nand g136 (n_3074, n_73, n_151);
  nor g137 (n_3075, n_72, n_150);
  nand g138 (n_3076, n_72, n_150);
  nor g139 (n_3085, n_71, n_149);
  nand g140 (n_3080, n_71, n_149);
  nor g141 (n_3081, n_70, n_148);
  nand g142 (n_3082, n_70, n_148);
  nor g143 (n_3091, n_69, n_147);
  nand g144 (n_3086, n_69, n_147);
  nor g145 (n_3087, n_68, n_146);
  nand g146 (n_3088, n_68, n_146);
  nor g147 (n_3097, n_67, n_145);
  nand g148 (n_3092, n_67, n_145);
  nor g149 (n_3093, n_66, n_144);
  nand g150 (n_3094, n_66, n_144);
  nor g151 (n_3103, n_65, n_143);
  nand g152 (n_3098, n_65, n_143);
  nor g153 (n_3099, n_64, n_142);
  nand g154 (n_3100, n_64, n_142);
  nor g155 (n_3109, n_63, n_141);
  nand g156 (n_3104, n_63, n_141);
  nor g166 (n_2891, n_1091, n_2889);
  nor g170 (n_2897, n_2894, n_2895);
  nor g173 (n_3123, n_2899, n_2895);
  nor g174 (n_2903, n_2900, n_2901);
  nor g177 (n_3125, n_2905, n_2901);
  nor g178 (n_2909, n_2906, n_2907);
  nor g181 (n_3133, n_2911, n_2907);
  nor g182 (n_2915, n_2912, n_2913);
  nor g185 (n_3135, n_2917, n_2913);
  nor g186 (n_2921, n_2918, n_2919);
  nor g189 (n_3143, n_2923, n_2919);
  nor g190 (n_2927, n_2924, n_2925);
  nor g193 (n_3145, n_2929, n_2925);
  nor g194 (n_2933, n_2930, n_2931);
  nor g197 (n_3153, n_2935, n_2931);
  nor g198 (n_2939, n_2936, n_2937);
  nor g201 (n_3155, n_2941, n_2937);
  nor g202 (n_2945, n_2942, n_2943);
  nor g205 (n_3163, n_2947, n_2943);
  nor g206 (n_2951, n_2948, n_2949);
  nor g209 (n_3165, n_2953, n_2949);
  nor g210 (n_2957, n_2954, n_2955);
  nor g213 (n_3173, n_2959, n_2955);
  nor g214 (n_2963, n_2960, n_2961);
  nor g217 (n_3175, n_2965, n_2961);
  nor g218 (n_2969, n_2966, n_2967);
  nor g221 (n_3183, n_2971, n_2967);
  nor g222 (n_2975, n_2972, n_2973);
  nor g225 (n_3185, n_2977, n_2973);
  nor g226 (n_2981, n_2978, n_2979);
  nor g229 (n_3193, n_2983, n_2979);
  nor g230 (n_2987, n_2984, n_2985);
  nor g233 (n_3195, n_2989, n_2985);
  nor g234 (n_2993, n_2990, n_2991);
  nor g237 (n_3203, n_2995, n_2991);
  nor g238 (n_2999, n_2996, n_2997);
  nor g241 (n_3205, n_3001, n_2997);
  nor g242 (n_3005, n_3002, n_3003);
  nor g245 (n_3213, n_3007, n_3003);
  nor g246 (n_3011, n_3008, n_3009);
  nor g249 (n_3215, n_3013, n_3009);
  nor g250 (n_3017, n_3014, n_3015);
  nor g253 (n_3223, n_3019, n_3015);
  nor g254 (n_3023, n_3020, n_3021);
  nor g257 (n_3225, n_3025, n_3021);
  nor g258 (n_3029, n_3026, n_3027);
  nor g261 (n_3233, n_3031, n_3027);
  nor g262 (n_3035, n_3032, n_3033);
  nor g265 (n_3235, n_3037, n_3033);
  nor g266 (n_3041, n_3038, n_3039);
  nor g269 (n_3243, n_3043, n_3039);
  nor g270 (n_3047, n_3044, n_3045);
  nor g273 (n_3245, n_3049, n_3045);
  nor g274 (n_3053, n_3050, n_3051);
  nor g277 (n_3253, n_3055, n_3051);
  nor g278 (n_3059, n_3056, n_3057);
  nor g281 (n_3255, n_3061, n_3057);
  nor g282 (n_3065, n_3062, n_3063);
  nor g285 (n_3263, n_3067, n_3063);
  nor g286 (n_3071, n_3068, n_3069);
  nor g289 (n_3265, n_3073, n_3069);
  nor g290 (n_3077, n_3074, n_3075);
  nor g293 (n_3273, n_3079, n_3075);
  nor g294 (n_3083, n_3080, n_3081);
  nor g297 (n_3275, n_3085, n_3081);
  nor g298 (n_3089, n_3086, n_3087);
  nor g301 (n_3283, n_3091, n_3087);
  nor g302 (n_3095, n_3092, n_3093);
  nor g305 (n_3285, n_3097, n_3093);
  nor g306 (n_3101, n_3098, n_3099);
  nor g309 (n_3293, n_3103, n_3099);
  nor g310 (n_3107, n_3104, n_3105);
  nor g313 (n_3295, n_3109, n_3105);
  nor g323 (n_3121, n_2905, n_3120);
  nand g332 (n_3308, n_3123, n_3125);
  nor g333 (n_3131, n_2917, n_3130);
  nand g342 (n_3315, n_3133, n_3135);
  nor g343 (n_3141, n_2929, n_3140);
  nand g352 (n_3323, n_3143, n_3145);
  nor g353 (n_3151, n_2941, n_3150);
  nand g362 (n_3330, n_3153, n_3155);
  nor g363 (n_3161, n_2953, n_3160);
  nand g372 (n_3338, n_3163, n_3165);
  nor g373 (n_3171, n_2965, n_3170);
  nand g382 (n_3345, n_3173, n_3175);
  nor g383 (n_3181, n_2977, n_3180);
  nand g392 (n_3353, n_3183, n_3185);
  nor g393 (n_3191, n_2989, n_3190);
  nand g402 (n_3360, n_3193, n_3195);
  nor g403 (n_3201, n_3001, n_3200);
  nand g412 (n_3368, n_3203, n_3205);
  nor g413 (n_3211, n_3013, n_3210);
  nand g422 (n_3375, n_3213, n_3215);
  nor g423 (n_3221, n_3025, n_3220);
  nand g432 (n_3383, n_3223, n_3225);
  nor g433 (n_3231, n_3037, n_3230);
  nand g442 (n_3390, n_3233, n_3235);
  nor g443 (n_3241, n_3049, n_3240);
  nand g452 (n_3398, n_3243, n_3245);
  nor g453 (n_3251, n_3061, n_3250);
  nand g462 (n_3405, n_3253, n_3255);
  nor g463 (n_3261, n_3073, n_3260);
  nand g3196 (n_3413, n_3263, n_3265);
  nor g3197 (n_3271, n_3085, n_3270);
  nand g3206 (n_3420, n_3273, n_3275);
  nor g3207 (n_3281, n_3097, n_3280);
  nand g3216 (n_3428, n_3283, n_3285);
  nor g3217 (n_3291, n_3109, n_3290);
  nand g3226 (n_3435, n_3293, n_3295);
  nand g3229 (n_3847, n_2894, n_3302);
  nand g3231 (n_3849, n_3120, n_3303);
  nand g3234 (n_3852, n_3306, n_3307);
  nand g3237 (n_3436, n_3310, n_3311);
  nor g3238 (n_3313, n_2923, n_3312);
  nor g3241 (n_3446, n_2923, n_3315);
  nor g3247 (n_3321, n_3319, n_3312);
  nor g3250 (n_3452, n_3315, n_3319);
  nor g3251 (n_3325, n_3323, n_3312);
  nor g3254 (n_3455, n_3315, n_3323);
  nor g3255 (n_3328, n_2947, n_3327);
  nor g3258 (n_3597, n_2947, n_3330);
  nor g3264 (n_3336, n_3334, n_3327);
  nor g3267 (n_3603, n_3330, n_3334);
  nor g3268 (n_3340, n_3338, n_3327);
  nor g3271 (n_3461, n_3330, n_3338);
  nor g3272 (n_3343, n_2971, n_3342);
  nor g3275 (n_3474, n_2971, n_3345);
  nor g3281 (n_3351, n_3349, n_3342);
  nor g3284 (n_3484, n_3345, n_3349);
  nor g3285 (n_3355, n_3353, n_3342);
  nor g3288 (n_3489, n_3345, n_3353);
  nor g3289 (n_3358, n_2995, n_3357);
  nor g3292 (n_3712, n_2995, n_3360);
  nor g3298 (n_3366, n_3364, n_3357);
  nor g3301 (n_3718, n_3360, n_3364);
  nor g3302 (n_3370, n_3368, n_3357);
  nor g3305 (n_3497, n_3360, n_3368);
  nor g3306 (n_3373, n_3019, n_3372);
  nor g3309 (n_3510, n_3019, n_3375);
  nor g3315 (n_3381, n_3379, n_3372);
  nor g3318 (n_3520, n_3375, n_3379);
  nor g3319 (n_3385, n_3383, n_3372);
  nor g3322 (n_3525, n_3375, n_3383);
  nor g3323 (n_3388, n_3043, n_3387);
  nor g3326 (n_3652, n_3043, n_3390);
  nor g3332 (n_3396, n_3394, n_3387);
  nor g3335 (n_3662, n_3390, n_3394);
  nor g3336 (n_3400, n_3398, n_3387);
  nor g3339 (n_3533, n_3390, n_3398);
  nor g3340 (n_3403, n_3067, n_3402);
  nor g3343 (n_3546, n_3067, n_3405);
  nor g3349 (n_3411, n_3409, n_3402);
  nor g3352 (n_3556, n_3405, n_3409);
  nor g3353 (n_3415, n_3413, n_3402);
  nor g3356 (n_3561, n_3405, n_3413);
  nor g3357 (n_3418, n_3091, n_3417);
  nor g3360 (n_3810, n_3091, n_3420);
  nor g3366 (n_3426, n_3424, n_3417);
  nor g3369 (n_3816, n_3420, n_3424);
  nor g3370 (n_3430, n_3428, n_3417);
  nor g3373 (n_3569, n_3420, n_3428);
  nor g3374 (n_3433, n_3113, n_3432);
  nor g3377 (n_3582, n_3113, n_3435);
  nand g3380 (n_3856, n_2906, n_3438);
  nand g3381 (n_3439, n_3133, n_3436);
  nand g3382 (n_3858, n_3130, n_3439);
  nand g3385 (n_3861, n_3442, n_3443);
  nand g3388 (n_3864, n_3312, n_3445);
  nand g3389 (n_3448, n_3446, n_3436);
  nand g3390 (n_3867, n_3447, n_3448);
  nand g3391 (n_3451, n_3449, n_3436);
  nand g3392 (n_3869, n_3450, n_3451);
  nand g3393 (n_3454, n_3452, n_3436);
  nand g3394 (n_3872, n_3453, n_3454);
  nand g3395 (n_3457, n_3455, n_3436);
  nand g3396 (n_3587, n_3456, n_3457);
  nor g3397 (n_3459, n_2959, n_3458);
  nand g3406 (n_3611, n_3173, n_3461);
  nor g3407 (n_3468, n_3466, n_3458);
  nor g3412 (n_3471, n_3345, n_3458);
  nand g3421 (n_3623, n_3461, n_3474);
  nand g3426 (n_3627, n_3461, n_3479);
  nand g3431 (n_3631, n_3461, n_3484);
  nand g3436 (n_3635, n_3461, n_3489);
  nor g3437 (n_3495, n_3007, n_3494);
  nand g3446 (n_3726, n_3213, n_3497);
  nor g3447 (n_3504, n_3502, n_3494);
  nor g3452 (n_3507, n_3375, n_3494);
  nand g3461 (n_3738, n_3497, n_3510);
  nand g3466 (n_3742, n_3497, n_3515);
  nand g3471 (n_3746, n_3497, n_3520);
  nand g3476 (n_3642, n_3497, n_3525);
  nor g3477 (n_3531, n_3055, n_3530);
  nand g3486 (n_3674, n_3253, n_3533);
  nor g3487 (n_3540, n_3538, n_3530);
  nor g3492 (n_3543, n_3405, n_3530);
  nand g3501 (n_3686, n_3533, n_3546);
  nand g3506 (n_3690, n_3533, n_3551);
  nand g3511 (n_3694, n_3533, n_3556);
  nand g3516 (n_3698, n_3533, n_3561);
  nor g3517 (n_3567, n_3103, n_3566);
  nand g3526 (n_3824, n_3293, n_3569);
  nor g3527 (n_3576, n_3574, n_3566);
  nor g3532 (n_3579, n_3435, n_3566);
  nand g3541 (n_3836, n_3569, n_3582);
  nand g3544 (n_3876, n_2930, n_3589);
  nand g3545 (n_3590, n_3153, n_3587);
  nand g3546 (n_3878, n_3150, n_3590);
  nand g3549 (n_3881, n_3593, n_3594);
  nand g3552 (n_3884, n_3327, n_3596);
  nand g3553 (n_3599, n_3597, n_3587);
  nand g3554 (n_3887, n_3598, n_3599);
  nand g3555 (n_3602, n_3600, n_3587);
  nand g3556 (n_3889, n_3601, n_3602);
  nand g3557 (n_3605, n_3603, n_3587);
  nand g3558 (n_3892, n_3604, n_3605);
  nand g3559 (n_3606, n_3461, n_3587);
  nand g3560 (n_3894, n_3458, n_3606);
  nand g3563 (n_3897, n_3609, n_3610);
  nand g3566 (n_3899, n_3613, n_3614);
  nand g3569 (n_3902, n_3617, n_3618);
  nand g3572 (n_3905, n_3621, n_3622);
  nand g3575 (n_3908, n_3625, n_3626);
  nand g3578 (n_3910, n_3629, n_3630);
  nand g3581 (n_3913, n_3633, n_3634);
  nand g3584 (n_3702, n_3637, n_3638);
  nor g3585 (n_3640, n_3031, n_3639);
  nor g3588 (n_3752, n_3031, n_3642);
  nor g3594 (n_3648, n_3646, n_3639);
  nor g3597 (n_3758, n_3646, n_3642);
  nor g3598 (n_3650, n_3390, n_3639);
  nor g3601 (n_3761, n_3390, n_3642);
  nor g3622 (n_3672, n_3670, n_3639);
  nor g3625 (n_3776, n_3642, n_3670);
  nor g3626 (n_3676, n_3674, n_3639);
  nor g3629 (n_3779, n_3642, n_3674);
  nor g3630 (n_3680, n_3678, n_3639);
  nor g3633 (n_3782, n_3642, n_3678);
  nor g3634 (n_3684, n_3682, n_3639);
  nor g3637 (n_3785, n_3642, n_3682);
  nor g3638 (n_3688, n_3686, n_3639);
  nor g3641 (n_3788, n_3642, n_3686);
  nor g3642 (n_3692, n_3690, n_3639);
  nor g3645 (n_3791, n_3642, n_3690);
  nor g3646 (n_3696, n_3694, n_3639);
  nor g3649 (n_3794, n_3642, n_3694);
  nor g3650 (n_3700, n_3698, n_3639);
  nor g3653 (n_3797, n_3642, n_3698);
  nand g3656 (n_3917, n_2978, n_3704);
  nand g3657 (n_3705, n_3193, n_3702);
  nand g3658 (n_3919, n_3190, n_3705);
  nand g3661 (n_3922, n_3708, n_3709);
  nand g3664 (n_3925, n_3357, n_3711);
  nand g3665 (n_3714, n_3712, n_3702);
  nand g3666 (n_3928, n_3713, n_3714);
  nand g3667 (n_3717, n_3715, n_3702);
  nand g3668 (n_3930, n_3716, n_3717);
  nand g3669 (n_3720, n_3718, n_3702);
  nand g3670 (n_3933, n_3719, n_3720);
  nand g3671 (n_3721, n_3497, n_3702);
  nand g3672 (n_3935, n_3494, n_3721);
  nand g3675 (n_3938, n_3724, n_3725);
  nand g3678 (n_3940, n_3728, n_3729);
  nand g3681 (n_3943, n_3732, n_3733);
  nand g3684 (n_3946, n_3736, n_3737);
  nand g3687 (n_3949, n_3740, n_3741);
  nand g3690 (n_3951, n_3744, n_3745);
  nand g3693 (n_3954, n_3748, n_3749);
  nand g3696 (n_3957, n_3639, n_3751);
  nand g3697 (n_3754, n_3752, n_3702);
  nand g3698 (n_3960, n_3753, n_3754);
  nand g3699 (n_3757, n_3755, n_3702);
  nand g3700 (n_3962, n_3756, n_3757);
  nand g3701 (n_3760, n_3758, n_3702);
  nand g3702 (n_3965, n_3759, n_3760);
  nand g3703 (n_3763, n_3761, n_3702);
  nand g3704 (n_3968, n_3762, n_3763);
  nand g3705 (n_3766, n_3764, n_3702);
  nand g3706 (n_3971, n_3765, n_3766);
  nand g3707 (n_3769, n_3767, n_3702);
  nand g3708 (n_3973, n_3768, n_3769);
  nand g3709 (n_3772, n_3770, n_3702);
  nand g3710 (n_3976, n_3771, n_3772);
  nand g3711 (n_3775, n_3773, n_3702);
  nand g3712 (n_3978, n_3774, n_3775);
  nand g3713 (n_3778, n_3776, n_3702);
  nand g3714 (n_3981, n_3777, n_3778);
  nand g3715 (n_3781, n_3779, n_3702);
  nand g3716 (n_3983, n_3780, n_3781);
  nand g3717 (n_3784, n_3782, n_3702);
  nand g3718 (n_3986, n_3783, n_3784);
  nand g3719 (n_3787, n_3785, n_3702);
  nand g3720 (n_3989, n_3786, n_3787);
  nand g3721 (n_3790, n_3788, n_3702);
  nand g3722 (n_3992, n_3789, n_3790);
  nand g3723 (n_3793, n_3791, n_3702);
  nand g3724 (n_3994, n_3792, n_3793);
  nand g3725 (n_3796, n_3794, n_3702);
  nand g3726 (n_3997, n_3795, n_3796);
  nand g3727 (n_3799, n_3797, n_3702);
  nand g3728 (n_3800, n_3798, n_3799);
  nand g3731 (n_4001, n_3074, n_3802);
  nand g3732 (n_3803, n_3273, n_3800);
  nand g3733 (n_4003, n_3270, n_3803);
  nand g3736 (n_4006, n_3806, n_3807);
  nand g3739 (n_4009, n_3417, n_3809);
  nand g3740 (n_3812, n_3810, n_3800);
  nand g3741 (n_4012, n_3811, n_3812);
  nand g3742 (n_3815, n_3813, n_3800);
  nand g3743 (n_4014, n_3814, n_3815);
  nand g3744 (n_3818, n_3816, n_3800);
  nand g3745 (n_4017, n_3817, n_3818);
  nand g3746 (n_3819, n_3569, n_3800);
  nand g3747 (n_4019, n_3566, n_3819);
  nand g3750 (n_4022, n_3822, n_3823);
  nand g3753 (n_4024, n_3826, n_3827);
  nand g3756 (n_4027, n_3830, n_3831);
  nand g3759 (n_4030, n_3834, n_3835);
  nand g3762 (n_4033, n_3838, n_3839);
  xnor g3774 (Z[5], n_3847, n_3848);
  xnor g3776 (Z[6], n_3849, n_3850);
  xnor g3779 (Z[7], n_3852, n_3853);
  xnor g3781 (Z[8], n_3436, n_3854);
  xnor g3784 (Z[9], n_3856, n_3857);
  xnor g3786 (Z[10], n_3858, n_3859);
  xnor g3789 (Z[11], n_3861, n_3862);
  xnor g3792 (Z[12], n_3864, n_3865);
  xnor g3795 (Z[13], n_3867, n_3868);
  xnor g3797 (Z[14], n_3869, n_3870);
  xnor g3800 (Z[15], n_3872, n_3873);
  xnor g3802 (Z[16], n_3587, n_3874);
  xnor g3805 (Z[17], n_3876, n_3877);
  xnor g3807 (Z[18], n_3878, n_3879);
  xnor g3810 (Z[19], n_3881, n_3882);
  xnor g3813 (Z[20], n_3884, n_3885);
  xnor g3816 (Z[21], n_3887, n_3888);
  xnor g3818 (Z[22], n_3889, n_3890);
  xnor g3821 (Z[23], n_3892, n_3893);
  xnor g3823 (Z[24], n_3894, n_3895);
  xnor g3826 (Z[25], n_3897, n_3898);
  xnor g3828 (Z[26], n_3899, n_3900);
  xnor g3831 (Z[27], n_3902, n_3903);
  xnor g3834 (Z[28], n_3905, n_3906);
  xnor g3837 (Z[29], n_3908, n_3909);
  xnor g3839 (Z[30], n_3910, n_3911);
  xnor g3842 (Z[31], n_3913, n_3914);
  xnor g3844 (Z[32], n_3702, n_3915);
  xnor g3847 (Z[33], n_3917, n_3918);
  xnor g3849 (Z[34], n_3919, n_3920);
  xnor g3852 (Z[35], n_3922, n_3923);
  xnor g3855 (Z[36], n_3925, n_3926);
  xnor g3858 (Z[37], n_3928, n_3929);
  xnor g3860 (Z[38], n_3930, n_3931);
  xnor g3863 (Z[39], n_3933, n_3934);
  xnor g3865 (Z[40], n_3935, n_3936);
  xnor g3868 (Z[41], n_3938, n_3939);
  xnor g3870 (Z[42], n_3940, n_3941);
  xnor g3873 (Z[43], n_3943, n_3944);
  xnor g3876 (Z[44], n_3946, n_3947);
  xnor g3879 (Z[45], n_3949, n_3950);
  xnor g3881 (Z[46], n_3951, n_3952);
  xnor g3884 (Z[47], n_3954, n_3955);
  xnor g3887 (Z[48], n_3957, n_3958);
  xnor g3890 (Z[49], n_3960, n_3961);
  xnor g3892 (Z[50], n_3962, n_3963);
  xnor g3895 (Z[51], n_3965, n_3966);
  xnor g3898 (Z[52], n_3968, n_3969);
  xnor g3901 (Z[53], n_3971, n_3972);
  xnor g3903 (Z[54], n_3973, n_3974);
  xnor g3906 (Z[55], n_3976, n_3977);
  xnor g3908 (Z[56], n_3978, n_3979);
  xnor g3911 (Z[57], n_3981, n_3982);
  xnor g3913 (Z[58], n_3983, n_3984);
  xnor g3916 (Z[59], n_3986, n_3987);
  xnor g3919 (Z[60], n_3989, n_3990);
  xnor g3922 (Z[61], n_3992, n_3993);
  xnor g3924 (Z[62], n_3994, n_3995);
  xnor g3927 (Z[63], n_3997, n_3998);
  xnor g3929 (Z[64], n_3800, n_3999);
  xnor g3932 (Z[65], n_4001, n_4002);
  xnor g3934 (Z[66], n_4003, n_4004);
  xnor g3937 (Z[67], n_4006, n_4007);
  xnor g3940 (Z[68], n_4009, n_4010);
  xnor g3943 (Z[69], n_4012, n_4013);
  xnor g3945 (Z[70], n_4014, n_4015);
  xnor g3948 (Z[71], n_4017, n_4018);
  xnor g3950 (Z[72], n_4019, n_4020);
  xnor g3953 (Z[73], n_4022, n_4023);
  xnor g3955 (Z[74], n_4024, n_4025);
  xnor g3958 (Z[75], n_4027, n_4028);
  xnor g3961 (Z[76], n_4030, n_4031);
  or g3975 (n_302, wc, wc0, n_132);
  not gc0 (wc0, n_1091);
  not gc (wc, n_1105);
  or g3976 (n_311, wc1, wc2, n_296);
  not gc2 (wc2, n_1105);
  not gc1 (wc1, n_1124);
  or g3977 (n_324, wc3, n_301, n_296);
  not gc3 (wc3, n_1152);
  or g3978 (n_342, wc4, wc5, n_301);
  not gc5 (wc5, n_1187);
  not gc4 (wc4, n_1188);
  or g3979 (n_364, wc6, wc7, n_301);
  not gc7 (wc7, n_1235);
  not gc6 (wc6, n_1236);
  or g3980 (n_410, wc8, wc9, n_361);
  not gc9 (wc9, n_1344);
  not gc8 (wc8, n_1345);
  or g3981 (n_411, wc10, wc11, n_296);
  not gc11 (wc11, n_1236);
  not gc10 (wc10, n_1284);
  or g3982 (n_438, wc12, wc13, n_361);
  not gc13 (wc13, n_1408);
  not gc12 (wc12, n_1409);
  or g3983 (n_439, wc14, wc15, n_301);
  not gc15 (wc15, n_1412);
  not gc14 (wc14, n_1413);
  or g3984 (n_466, wc16, wc17, n_361);
  not gc17 (wc17, n_1472);
  not gc16 (wc16, n_1473);
  or g3985 (n_467, wc18, wc19, n_310);
  not gc19 (wc19, n_1475);
  not gc18 (wc18, n_1477);
  or g3986 (n_493, wc20, wc21, n_323);
  not gc21 (wc21, n_1352);
  not gc20 (wc20, n_1539);
  or g3987 (n_519, wc22, wc23, n_361);
  not gc23 (wc23, n_1599);
  not gc22 (wc22, n_1601);
  or g3988 (n_575, wc24, wc25, n_361);
  not gc25 (wc25, n_1665);
  not gc24 (wc24, n_1729);
  xnor g3989 (n_2622, A[58], A[56]);
  or g3990 (n_2623, wc26, A[58]);
  not gc26 (wc26, A[56]);
  or g3991 (n_2625, wc27, A[58]);
  not gc27 (wc27, A[52]);
  xnor g3992 (n_2662, A[57], A[45]);
  or g3993 (n_2663, wc28, A[57]);
  not gc28 (wc28, A[45]);
  xnor g3994 (n_1030, n_2714, A[55]);
  or g3995 (n_2764, wc29, A[55]);
  not gc29 (wc29, A[53]);
  or g3996 (n_2765, wc30, A[55]);
  not gc30 (wc30, A[47]);
  xnor g3998 (n_1076, n_2462, A[57]);
  or g3999 (n_2856, wc31, A[57]);
  not gc31 (wc31, A[53]);
  or g4000 (n_2857, wc32, A[57]);
  not gc32 (wc32, A[55]);
  or g4001 (n_2631, wc33, A[58]);
  not gc33 (wc33, A[54]);
  or g4003 (n_2871, A[55], wc34);
  not gc34 (wc34, A[57]);
  or g4004 (n_2877, wc35, A[58]);
  not gc35 (wc35, A[55]);
  and g4005 (n_3113, wc36, A[58]);
  not gc36 (wc36, A[57]);
  or g4006 (n_3110, wc37, A[58]);
  not gc37 (wc37, A[57]);
  or g4007 (n_390, wc38, wc39, n_301);
  not gc39 (wc39, n_1292);
  not gc38 (wc38, n_1293);
  or g4008 (n_2721, A[57], wc40);
  not gc40 (wc40, n_1004);
  xnor g4009 (n_1050, n_2462, n_944);
  or g4010 (n_2804, A[55], wc41);
  not gc41 (wc41, n_944);
  or g4011 (n_2837, A[57], wc42);
  not gc42 (wc42, n_1064);
  and g4012 (n_3118, wc43, n_1087);
  not gc43 (wc43, n_2891);
  or g4014 (n_3841, n_2893, wc44);
  not gc44 (wc44, n_1091);
  or g4015 (n_3844, n_2889, wc45);
  not gc45 (wc45, n_1087);
  xnor g4016 (n_2630, A[58], A[54]);
  or g4017 (n_2633, wc46, A[58]);
  not gc46 (wc46, A[48]);
  or g4018 (n_2664, A[57], wc47);
  not gc47 (wc47, n_975);
  xnor g4019 (n_2718, n_975, A[57]);
  xnor g4020 (n_64, n_2526, n_1083);
  or g4021 (n_2872, A[55], wc48);
  not gc48 (wc48, n_1083);
  and g4022 (n_3105, A[57], wc49);
  not gc49 (wc49, n_140);
  or g4023 (n_3106, A[57], wc50);
  not gc50 (wc50, n_140);
  or g4024 (n_3845, wc51, n_2899);
  not gc51 (wc51, n_2894);
  or g4025 (n_4031, wc52, n_3113);
  not gc52 (wc52, n_3110);
  and g4026 (n_3120, wc53, n_2896);
  not gc53 (wc53, n_2897);
  or g4027 (n_3304, wc54, n_2905);
  not gc54 (wc54, n_3123);
  not g4028 (Z[2], n_3841);
  or g4029 (n_3848, wc55, n_2895);
  not gc55 (wc55, n_2896);
  or g4030 (n_3850, wc56, n_2905);
  not gc56 (wc56, n_2900);
  and g4031 (n_3127, wc57, n_2902);
  not gc57 (wc57, n_2903);
  or g4034 (n_3853, wc58, n_2901);
  not gc58 (wc58, n_2902);
  or g4035 (n_4028, wc59, n_3105);
  not gc59 (wc59, n_3106);
  and g4036 (n_3130, wc60, n_2908);
  not gc60 (wc60, n_2909);
  and g4037 (n_3306, wc61, n_2900);
  not gc61 (wc61, n_3121);
  and g4038 (n_3128, wc62, n_3125);
  not gc62 (wc62, n_3120);
  or g4039 (n_3302, n_2899, n_3118);
  or g4040 (n_3303, n_3118, wc63);
  not gc63 (wc63, n_3123);
  or g4041 (n_3307, n_3118, n_3304);
  xor g4042 (Z[3], n_1091, n_3844);
  xor g4043 (Z[4], n_3118, n_3845);
  or g4044 (n_3854, wc64, n_2911);
  not gc64 (wc64, n_2906);
  or g4045 (n_3857, wc65, n_2907);
  not gc65 (wc65, n_2908);
  and g4046 (n_3297, n_3106, wc66);
  not gc66 (wc66, n_3107);
  and g4047 (n_3310, wc67, n_3127);
  not gc67 (wc67, n_3128);
  or g4048 (n_3440, wc68, n_2917);
  not gc68 (wc68, n_3133);
  or g4049 (n_3311, n_3308, n_3118);
  or g4050 (n_3859, wc69, n_2917);
  not gc69 (wc69, n_2912);
  or g4051 (n_4023, wc70, n_3099);
  not gc70 (wc70, n_3100);
  or g4052 (n_4025, wc71, n_3109);
  not gc71 (wc71, n_3104);
  and g4053 (n_3137, wc72, n_2914);
  not gc72 (wc72, n_2915);
  and g4054 (n_3140, wc73, n_2920);
  not gc73 (wc73, n_2921);
  and g4055 (n_3290, wc74, n_3100);
  not gc74 (wc74, n_3101);
  and g4056 (n_3442, wc75, n_2912);
  not gc75 (wc75, n_3131);
  or g4057 (n_3574, wc76, n_3109);
  not gc76 (wc76, n_3293);
  or g4058 (n_3862, wc77, n_2913);
  not gc77 (wc77, n_2914);
  or g4059 (n_3865, wc78, n_2923);
  not gc78 (wc78, n_2918);
  or g4060 (n_3868, wc79, n_2919);
  not gc79 (wc79, n_2920);
  or g4061 (n_4020, wc80, n_3103);
  not gc80 (wc80, n_3098);
  and g4062 (n_3147, wc81, n_2926);
  not gc81 (wc81, n_2927);
  and g4063 (n_3287, wc82, n_3094);
  not gc82 (wc82, n_3095);
  and g4064 (n_3138, wc83, n_3135);
  not gc83 (wc83, n_3130);
  or g4065 (n_3319, wc84, n_2929);
  not gc84 (wc84, n_3143);
  and g4066 (n_3298, wc85, n_3295);
  not gc85 (wc85, n_3290);
  and g4067 (n_3449, wc86, n_3143);
  not gc86 (wc86, n_3315);
  or g4068 (n_3438, wc87, n_2911);
  not gc87 (wc87, n_3436);
  or g4069 (n_3443, n_3440, wc88);
  not gc88 (wc88, n_3436);
  or g4070 (n_3870, wc89, n_2929);
  not gc89 (wc89, n_2924);
  or g4071 (n_3873, wc90, n_2925);
  not gc90 (wc90, n_2926);
  or g4072 (n_4013, wc91, n_3087);
  not gc91 (wc91, n_3088);
  or g4073 (n_4015, wc92, n_3097);
  not gc92 (wc92, n_3092);
  or g4074 (n_4018, wc93, n_3093);
  not gc93 (wc93, n_3094);
  and g4075 (n_3150, wc94, n_2932);
  not gc94 (wc94, n_2933);
  and g4076 (n_3157, wc95, n_2938);
  not gc95 (wc95, n_2939);
  and g4077 (n_3280, wc96, n_3088);
  not gc96 (wc96, n_3089);
  and g4078 (n_3312, wc97, n_3137);
  not gc97 (wc97, n_3138);
  and g4079 (n_3320, wc98, n_2924);
  not gc98 (wc98, n_3141);
  and g4080 (n_3148, wc99, n_3145);
  not gc99 (wc99, n_3140);
  or g4081 (n_3591, wc100, n_2941);
  not gc100 (wc100, n_3153);
  or g4082 (n_3424, wc101, n_3097);
  not gc101 (wc101, n_3283);
  and g4083 (n_3575, wc102, n_3104);
  not gc102 (wc102, n_3291);
  and g4084 (n_3432, wc103, n_3297);
  not gc103 (wc103, n_3298);
  or g4085 (n_3445, wc104, n_3315);
  not gc104 (wc104, n_3436);
  or g4086 (n_3874, wc105, n_2935);
  not gc105 (wc105, n_2930);
  or g4087 (n_3877, wc106, n_2931);
  not gc106 (wc106, n_2932);
  or g4088 (n_3879, wc107, n_2941);
  not gc107 (wc107, n_2936);
  or g4089 (n_3882, wc108, n_2937);
  not gc108 (wc108, n_2938);
  or g4090 (n_3885, wc109, n_2947);
  not gc109 (wc109, n_2942);
  or g4091 (n_4010, wc110, n_3091);
  not gc110 (wc110, n_3086);
  and g4092 (n_3160, wc111, n_2944);
  not gc111 (wc111, n_2945);
  and g4093 (n_3277, wc112, n_3082);
  not gc112 (wc112, n_3083);
  and g4094 (n_3324, wc113, n_3147);
  not gc113 (wc113, n_3148);
  and g4095 (n_3158, wc114, n_3155);
  not gc114 (wc114, n_3150);
  and g4096 (n_3288, wc115, n_3285);
  not gc115 (wc115, n_3280);
  and g4097 (n_3317, wc116, n_3143);
  not gc116 (wc116, n_3312);
  or g4098 (n_3888, wc117, n_2943);
  not gc117 (wc117, n_2944);
  or g4099 (n_4002, wc118, n_3075);
  not gc118 (wc118, n_3076);
  or g4100 (n_4004, wc119, n_3085);
  not gc119 (wc119, n_3080);
  or g4101 (n_4007, wc120, n_3081);
  not gc120 (wc120, n_3082);
  and g4102 (n_3167, wc121, n_2950);
  not gc121 (wc121, n_2951);
  and g4103 (n_3170, wc122, n_2956);
  not gc122 (wc122, n_2957);
  and g4104 (n_3177, wc123, n_2962);
  not gc123 (wc123, n_2963);
  and g4105 (n_3180, wc124, n_2968);
  not gc124 (wc124, n_2969);
  and g4106 (n_3187, wc125, n_2974);
  not gc125 (wc125, n_2975);
  and g4107 (n_3190, wc126, n_2980);
  not gc126 (wc126, n_2981);
  and g4108 (n_3197, wc127, n_2986);
  not gc127 (wc127, n_2987);
  and g4109 (n_3200, wc128, n_2992);
  not gc128 (wc128, n_2993);
  and g4110 (n_3207, wc129, n_2998);
  not gc129 (wc129, n_2999);
  and g4111 (n_3210, wc130, n_3004);
  not gc130 (wc130, n_3005);
  and g4112 (n_3217, wc131, n_3010);
  not gc131 (wc131, n_3011);
  and g4113 (n_3220, wc132, n_3016);
  not gc132 (wc132, n_3017);
  and g4114 (n_3227, wc133, n_3022);
  not gc133 (wc133, n_3023);
  and g4115 (n_3230, wc134, n_3028);
  not gc134 (wc134, n_3029);
  and g4116 (n_3237, wc135, n_3034);
  not gc135 (wc135, n_3035);
  and g4117 (n_3240, wc136, n_3040);
  not gc136 (wc136, n_3041);
  and g4118 (n_3247, wc137, n_3046);
  not gc137 (wc137, n_3047);
  and g4119 (n_3250, wc138, n_3052);
  not gc138 (wc138, n_3053);
  and g4120 (n_3257, wc139, n_3058);
  not gc139 (wc139, n_3059);
  and g4121 (n_3593, wc140, n_2936);
  not gc140 (wc140, n_3151);
  and g4122 (n_3327, wc141, n_3157);
  not gc141 (wc141, n_3158);
  or g4123 (n_3334, wc142, n_2953);
  not gc142 (wc142, n_3163);
  or g4124 (n_3466, wc143, n_2965);
  not gc143 (wc143, n_3173);
  or g4125 (n_3349, wc144, n_2977);
  not gc144 (wc144, n_3183);
  or g4126 (n_3706, wc145, n_2989);
  not gc145 (wc145, n_3193);
  or g4127 (n_3364, wc146, n_3001);
  not gc146 (wc146, n_3203);
  or g4128 (n_3502, wc147, n_3013);
  not gc147 (wc147, n_3213);
  or g4129 (n_3379, wc148, n_3025);
  not gc148 (wc148, n_3223);
  or g4130 (n_3646, wc149, n_3037);
  not gc149 (wc149, n_3233);
  or g4131 (n_3394, wc150, n_3049);
  not gc150 (wc150, n_3243);
  or g4132 (n_3538, wc151, n_3061);
  not gc151 (wc151, n_3253);
  and g4133 (n_3425, wc152, n_3092);
  not gc152 (wc152, n_3281);
  and g4134 (n_3429, wc153, n_3287);
  not gc153 (wc153, n_3288);
  and g4135 (n_3447, wc154, n_2918);
  not gc154 (wc154, n_3313);
  and g4136 (n_3450, wc155, n_3140);
  not gc155 (wc155, n_3317);
  and g4137 (n_3453, n_3320, wc156);
  not gc156 (wc156, n_3321);
  and g4138 (n_3600, wc157, n_3163);
  not gc157 (wc157, n_3330);
  and g4139 (n_3584, n_3110, wc158);
  not gc158 (wc158, n_3433);
  or g4140 (n_3890, wc159, n_2953);
  not gc159 (wc159, n_2948);
  or g4141 (n_3893, wc160, n_2949);
  not gc160 (wc160, n_2950);
  or g4142 (n_3895, wc161, n_2959);
  not gc161 (wc161, n_2954);
  or g4143 (n_3898, wc162, n_2955);
  not gc162 (wc162, n_2956);
  or g4144 (n_3900, wc163, n_2965);
  not gc163 (wc163, n_2960);
  or g4145 (n_3903, wc164, n_2961);
  not gc164 (wc164, n_2962);
  or g4146 (n_3906, wc165, n_2971);
  not gc165 (wc165, n_2966);
  or g4147 (n_3909, wc166, n_2967);
  not gc166 (wc166, n_2968);
  or g4148 (n_3911, wc167, n_2977);
  not gc167 (wc167, n_2972);
  or g4149 (n_3914, wc168, n_2973);
  not gc168 (wc168, n_2974);
  or g4150 (n_3915, wc169, n_2983);
  not gc169 (wc169, n_2978);
  or g4151 (n_3918, wc170, n_2979);
  not gc170 (wc170, n_2980);
  or g4152 (n_3920, wc171, n_2989);
  not gc171 (wc171, n_2984);
  or g4153 (n_3923, wc172, n_2985);
  not gc172 (wc172, n_2986);
  or g4154 (n_3926, wc173, n_2995);
  not gc173 (wc173, n_2990);
  or g4155 (n_3929, wc174, n_2991);
  not gc174 (wc174, n_2992);
  or g4156 (n_3931, wc175, n_3001);
  not gc175 (wc175, n_2996);
  or g4157 (n_3934, wc176, n_2997);
  not gc176 (wc176, n_2998);
  or g4158 (n_3936, wc177, n_3007);
  not gc177 (wc177, n_3002);
  or g4159 (n_3939, wc178, n_3003);
  not gc178 (wc178, n_3004);
  or g4160 (n_3941, wc179, n_3013);
  not gc179 (wc179, n_3008);
  or g4161 (n_3944, wc180, n_3009);
  not gc180 (wc180, n_3010);
  or g4162 (n_3947, wc181, n_3019);
  not gc181 (wc181, n_3014);
  or g4163 (n_3950, wc182, n_3015);
  not gc182 (wc182, n_3016);
  or g4164 (n_3952, wc183, n_3025);
  not gc183 (wc183, n_3020);
  or g4165 (n_3955, wc184, n_3021);
  not gc184 (wc184, n_3022);
  or g4166 (n_3958, wc185, n_3031);
  not gc185 (wc185, n_3026);
  or g4167 (n_3961, wc186, n_3027);
  not gc186 (wc186, n_3028);
  or g4168 (n_3963, wc187, n_3037);
  not gc187 (wc187, n_3032);
  or g4169 (n_3966, wc188, n_3033);
  not gc188 (wc188, n_3034);
  or g4170 (n_3969, wc189, n_3043);
  not gc189 (wc189, n_3038);
  or g4171 (n_3972, wc190, n_3039);
  not gc190 (wc190, n_3040);
  or g4172 (n_3974, wc191, n_3049);
  not gc191 (wc191, n_3044);
  or g4173 (n_3977, wc192, n_3045);
  not gc192 (wc192, n_3046);
  or g4174 (n_3979, wc193, n_3055);
  not gc193 (wc193, n_3050);
  or g4175 (n_3982, wc194, n_3051);
  not gc194 (wc194, n_3052);
  or g4176 (n_3984, wc195, n_3061);
  not gc195 (wc195, n_3056);
  or g4177 (n_3987, wc196, n_3057);
  not gc196 (wc196, n_3058);
  and g4178 (n_3260, wc197, n_3064);
  not gc197 (wc197, n_3065);
  and g4179 (n_3335, wc198, n_2948);
  not gc198 (wc198, n_3161);
  and g4180 (n_3168, wc199, n_3165);
  not gc199 (wc199, n_3160);
  and g4181 (n_3178, wc200, n_3175);
  not gc200 (wc200, n_3170);
  and g4182 (n_3188, wc201, n_3185);
  not gc201 (wc201, n_3180);
  and g4183 (n_3198, wc202, n_3195);
  not gc202 (wc202, n_3190);
  and g4184 (n_3208, wc203, n_3205);
  not gc203 (wc203, n_3200);
  and g4185 (n_3218, wc204, n_3215);
  not gc204 (wc204, n_3210);
  and g4186 (n_3228, wc205, n_3225);
  not gc205 (wc205, n_3220);
  and g4187 (n_3238, wc206, n_3235);
  not gc206 (wc206, n_3230);
  and g4188 (n_3248, wc207, n_3245);
  not gc207 (wc207, n_3240);
  and g4189 (n_3258, wc208, n_3255);
  not gc208 (wc208, n_3250);
  and g4190 (n_3456, n_3324, wc209);
  not gc209 (wc209, n_3325);
  and g4191 (n_3332, wc210, n_3163);
  not gc210 (wc210, n_3327);
  and g4192 (n_3479, wc211, n_3183);
  not gc211 (wc211, n_3345);
  and g4193 (n_3715, wc212, n_3203);
  not gc212 (wc212, n_3360);
  and g4194 (n_3515, wc213, n_3223);
  not gc213 (wc213, n_3375);
  and g4195 (n_3657, wc214, n_3243);
  not gc214 (wc214, n_3390);
  or g4196 (n_3990, wc215, n_3067);
  not gc215 (wc215, n_3062);
  or g4197 (n_3993, wc216, n_3063);
  not gc216 (wc216, n_3064);
  and g4198 (n_3267, wc217, n_3070);
  not gc217 (wc217, n_3071);
  and g4199 (n_3339, wc218, n_3167);
  not gc218 (wc218, n_3168);
  and g4200 (n_3467, wc219, n_2960);
  not gc219 (wc219, n_3171);
  and g4201 (n_3342, wc220, n_3177);
  not gc220 (wc220, n_3178);
  and g4202 (n_3350, wc221, n_2972);
  not gc221 (wc221, n_3181);
  and g4203 (n_3354, wc222, n_3187);
  not gc222 (wc222, n_3188);
  and g4204 (n_3708, wc223, n_2984);
  not gc223 (wc223, n_3191);
  and g4205 (n_3357, wc224, n_3197);
  not gc224 (wc224, n_3198);
  and g4206 (n_3365, wc225, n_2996);
  not gc225 (wc225, n_3201);
  and g4207 (n_3369, wc226, n_3207);
  not gc226 (wc226, n_3208);
  and g4208 (n_3503, wc227, n_3008);
  not gc227 (wc227, n_3211);
  and g4209 (n_3372, wc228, n_3217);
  not gc228 (wc228, n_3218);
  and g4210 (n_3380, wc229, n_3020);
  not gc229 (wc229, n_3221);
  and g4211 (n_3384, wc230, n_3227);
  not gc230 (wc230, n_3228);
  and g4212 (n_3647, wc231, n_3032);
  not gc231 (wc231, n_3231);
  and g4213 (n_3387, wc232, n_3237);
  not gc232 (wc232, n_3238);
  and g4214 (n_3395, wc233, n_3044);
  not gc233 (wc233, n_3241);
  and g4215 (n_3399, wc234, n_3247);
  not gc234 (wc234, n_3248);
  and g4216 (n_3539, wc235, n_3056);
  not gc235 (wc235, n_3251);
  and g4217 (n_3402, wc236, n_3257);
  not gc236 (wc236, n_3258);
  or g4218 (n_3409, wc237, n_3073);
  not gc237 (wc237, n_3263);
  and g4219 (n_3598, wc238, n_2942);
  not gc238 (wc238, n_3328);
  and g4220 (n_3601, wc239, n_3160);
  not gc239 (wc239, n_3332);
  and g4221 (n_3551, wc240, n_3263);
  not gc240 (wc240, n_3405);
  or g4222 (n_3607, wc241, n_2959);
  not gc241 (wc241, n_3461);
  or g4223 (n_3615, n_3466, wc242);
  not gc242 (wc242, n_3461);
  or g4224 (n_3619, wc243, n_3345);
  not gc243 (wc243, n_3461);
  or g4225 (n_3722, wc244, n_3007);
  not gc244 (wc244, n_3497);
  or g4226 (n_3730, n_3502, wc245);
  not gc245 (wc245, n_3497);
  or g4227 (n_3734, wc246, n_3375);
  not gc246 (wc246, n_3497);
  or g4228 (n_3670, wc247, n_3055);
  not gc247 (wc247, n_3533);
  or g4229 (n_3678, n_3538, wc248);
  not gc248 (wc248, n_3533);
  or g4230 (n_3682, wc249, n_3405);
  not gc249 (wc249, n_3533);
  or g4231 (n_3995, wc250, n_3073);
  not gc250 (wc250, n_3068);
  or g4232 (n_3998, wc251, n_3069);
  not gc251 (wc251, n_3070);
  and g4233 (n_3270, wc252, n_3076);
  not gc252 (wc252, n_3077);
  and g4234 (n_3410, wc253, n_3068);
  not gc253 (wc253, n_3261);
  and g4235 (n_3268, wc254, n_3265);
  not gc254 (wc254, n_3260);
  or g4236 (n_3804, wc255, n_3085);
  not gc255 (wc255, n_3273);
  and g4237 (n_3604, n_3335, wc256);
  not gc256 (wc256, n_3336);
  and g4238 (n_3347, wc257, n_3183);
  not gc257 (wc257, n_3342);
  and g4239 (n_3362, wc258, n_3203);
  not gc258 (wc258, n_3357);
  and g4240 (n_3377, wc259, n_3223);
  not gc259 (wc259, n_3372);
  and g4241 (n_3392, wc260, n_3243);
  not gc260 (wc260, n_3387);
  and g4242 (n_3407, wc261, n_3263);
  not gc261 (wc261, n_3402);
  or g4243 (n_3589, wc262, n_2935);
  not gc262 (wc262, n_3587);
  or g4244 (n_3594, n_3591, wc263);
  not gc263 (wc263, n_3587);
  or g4245 (n_3596, wc264, n_3330);
  not gc264 (wc264, n_3587);
  and g4246 (n_3755, wc265, n_3233);
  not gc265 (wc265, n_3642);
  and g4247 (n_3764, wc266, n_3652);
  not gc266 (wc266, n_3642);
  and g4248 (n_3767, n_3657, wc267);
  not gc267 (wc267, n_3642);
  and g4249 (n_3770, wc268, n_3662);
  not gc268 (wc268, n_3642);
  and g4250 (n_3773, wc269, n_3533);
  not gc269 (wc269, n_3642);
  or g4251 (n_3999, wc270, n_3079);
  not gc270 (wc270, n_3074);
  and g4252 (n_3414, wc271, n_3267);
  not gc271 (wc271, n_3268);
  and g4253 (n_3278, wc272, n_3275);
  not gc272 (wc272, n_3270);
  and g4254 (n_3458, n_3339, wc273);
  not gc273 (wc273, n_3340);
  and g4255 (n_3476, wc274, n_2966);
  not gc274 (wc274, n_3343);
  and g4256 (n_3481, wc275, n_3180);
  not gc275 (wc275, n_3347);
  and g4257 (n_3486, n_3350, wc276);
  not gc276 (wc276, n_3351);
  and g4258 (n_3491, n_3354, wc277);
  not gc277 (wc277, n_3355);
  and g4259 (n_3713, wc278, n_2990);
  not gc278 (wc278, n_3358);
  and g4260 (n_3716, wc279, n_3200);
  not gc279 (wc279, n_3362);
  and g4261 (n_3719, n_3365, wc280);
  not gc280 (wc280, n_3366);
  and g4262 (n_3494, n_3369, wc281);
  not gc281 (wc281, n_3370);
  and g4263 (n_3512, wc282, n_3014);
  not gc282 (wc282, n_3373);
  and g4264 (n_3517, wc283, n_3220);
  not gc283 (wc283, n_3377);
  and g4265 (n_3522, n_3380, wc284);
  not gc284 (wc284, n_3381);
  and g4266 (n_3527, n_3384, wc285);
  not gc285 (wc285, n_3385);
  and g4267 (n_3654, wc286, n_3038);
  not gc286 (wc286, n_3388);
  and g4268 (n_3659, wc287, n_3240);
  not gc287 (wc287, n_3392);
  and g4269 (n_3664, n_3395, wc288);
  not gc288 (wc288, n_3396);
  and g4270 (n_3530, n_3399, wc289);
  not gc289 (wc289, n_3400);
  and g4271 (n_3548, wc290, n_3062);
  not gc290 (wc290, n_3403);
  and g4272 (n_3553, wc291, n_3260);
  not gc291 (wc291, n_3407);
  and g4273 (n_3813, wc292, n_3283);
  not gc292 (wc292, n_3420);
  or g4274 (n_3610, n_3607, wc293);
  not gc293 (wc293, n_3587);
  or g4275 (n_3614, n_3611, wc294);
  not gc294 (wc294, n_3587);
  or g4276 (n_3618, n_3615, wc295);
  not gc295 (wc295, n_3587);
  or g4277 (n_3622, n_3619, wc296);
  not gc296 (wc296, n_3587);
  or g4278 (n_3626, n_3623, wc297);
  not gc297 (wc297, n_3587);
  or g4279 (n_3630, n_3627, wc298);
  not gc298 (wc298, n_3587);
  or g4280 (n_3634, n_3631, wc299);
  not gc299 (wc299, n_3587);
  or g4281 (n_3638, n_3635, wc300);
  not gc300 (wc300, n_3587);
  and g4282 (n_3806, wc301, n_3080);
  not gc301 (wc301, n_3271);
  and g4283 (n_3417, wc302, n_3277);
  not gc302 (wc302, n_3278);
  and g4284 (n_3558, n_3410, wc303);
  not gc303 (wc303, n_3411);
  and g4285 (n_3464, wc304, n_3173);
  not gc304 (wc304, n_3458);
  and g4286 (n_3477, wc305, n_3474);
  not gc305 (wc305, n_3458);
  and g4287 (n_3482, wc306, n_3479);
  not gc306 (wc306, n_3458);
  and g4288 (n_3487, wc307, n_3484);
  not gc307 (wc307, n_3458);
  and g4289 (n_3492, wc308, n_3489);
  not gc308 (wc308, n_3458);
  and g4290 (n_3500, wc309, n_3213);
  not gc309 (wc309, n_3494);
  and g4291 (n_3513, wc310, n_3510);
  not gc310 (wc310, n_3494);
  and g4292 (n_3518, wc311, n_3515);
  not gc311 (wc311, n_3494);
  and g4293 (n_3523, wc312, n_3520);
  not gc312 (wc312, n_3494);
  and g4294 (n_3528, wc313, n_3525);
  not gc313 (wc313, n_3494);
  and g4295 (n_3536, wc314, n_3253);
  not gc314 (wc314, n_3530);
  and g4296 (n_3549, wc315, n_3546);
  not gc315 (wc315, n_3530);
  and g4297 (n_3554, wc316, n_3551);
  not gc316 (wc316, n_3530);
  and g4298 (n_3559, wc317, n_3556);
  not gc317 (wc317, n_3530);
  and g4299 (n_3564, wc318, n_3561);
  not gc318 (wc318, n_3530);
  or g4300 (n_3820, wc319, n_3103);
  not gc319 (wc319, n_3569);
  or g4301 (n_3828, n_3574, wc320);
  not gc320 (wc320, n_3569);
  or g4302 (n_3832, wc321, n_3435);
  not gc321 (wc321, n_3569);
  and g4303 (n_3563, n_3414, wc322);
  not gc322 (wc322, n_3415);
  and g4304 (n_3422, wc323, n_3283);
  not gc323 (wc323, n_3417);
  and g4305 (n_3609, wc324, n_2954);
  not gc324 (wc324, n_3459);
  and g4306 (n_3613, wc325, n_3170);
  not gc325 (wc325, n_3464);
  and g4307 (n_3617, n_3467, wc326);
  not gc326 (wc326, n_3468);
  and g4308 (n_3621, n_3342, wc327);
  not gc327 (wc327, n_3471);
  and g4309 (n_3625, wc328, n_3476);
  not gc328 (wc328, n_3477);
  and g4310 (n_3629, wc329, n_3481);
  not gc329 (wc329, n_3482);
  and g4311 (n_3633, wc330, n_3486);
  not gc330 (wc330, n_3487);
  and g4312 (n_3637, wc331, n_3491);
  not gc331 (wc331, n_3492);
  and g4313 (n_3724, wc332, n_3002);
  not gc332 (wc332, n_3495);
  and g4314 (n_3728, wc333, n_3210);
  not gc333 (wc333, n_3500);
  and g4315 (n_3732, n_3503, wc334);
  not gc334 (wc334, n_3504);
  and g4316 (n_3736, n_3372, wc335);
  not gc335 (wc335, n_3507);
  and g4317 (n_3740, wc336, n_3512);
  not gc336 (wc336, n_3513);
  and g4318 (n_3744, wc337, n_3517);
  not gc337 (wc337, n_3518);
  and g4319 (n_3748, wc338, n_3522);
  not gc338 (wc338, n_3523);
  and g4320 (n_3639, wc339, n_3527);
  not gc339 (wc339, n_3528);
  and g4321 (n_3671, wc340, n_3050);
  not gc340 (wc340, n_3531);
  and g4322 (n_3675, wc341, n_3250);
  not gc341 (wc341, n_3536);
  and g4323 (n_3679, n_3539, wc342);
  not gc342 (wc342, n_3540);
  and g4324 (n_3683, n_3402, wc343);
  not gc343 (wc343, n_3543);
  and g4325 (n_3687, wc344, n_3548);
  not gc344 (wc344, n_3549);
  and g4326 (n_3691, wc345, n_3553);
  not gc345 (wc345, n_3554);
  and g4327 (n_3811, wc346, n_3086);
  not gc346 (wc346, n_3418);
  and g4328 (n_3814, wc347, n_3280);
  not gc347 (wc347, n_3422);
  and g4329 (n_3817, n_3425, wc348);
  not gc348 (wc348, n_3426);
  and g4330 (n_3566, n_3429, wc349);
  not gc349 (wc349, n_3430);
  and g4331 (n_3695, wc350, n_3558);
  not gc350 (wc350, n_3559);
  and g4332 (n_3644, wc351, n_3233);
  not gc351 (wc351, n_3639);
  and g4333 (n_3655, wc352, n_3652);
  not gc352 (wc352, n_3639);
  and g4334 (n_3660, wc353, n_3657);
  not gc353 (wc353, n_3639);
  and g4335 (n_3665, wc354, n_3662);
  not gc354 (wc354, n_3639);
  and g4336 (n_3668, wc355, n_3533);
  not gc355 (wc355, n_3639);
  and g4337 (n_3699, n_3563, wc356);
  not gc356 (wc356, n_3564);
  and g4338 (n_3572, wc357, n_3293);
  not gc357 (wc357, n_3566);
  and g4339 (n_3585, wc358, n_3582);
  not gc358 (wc358, n_3566);
  and g4340 (n_3753, wc359, n_3026);
  not gc359 (wc359, n_3640);
  and g4341 (n_3756, wc360, n_3230);
  not gc360 (wc360, n_3644);
  and g4342 (n_3759, n_3647, wc361);
  not gc361 (wc361, n_3648);
  and g4343 (n_3762, n_3387, wc362);
  not gc362 (wc362, n_3650);
  and g4344 (n_3765, wc363, n_3654);
  not gc363 (wc363, n_3655);
  and g4345 (n_3768, wc364, n_3659);
  not gc364 (wc364, n_3660);
  and g4346 (n_3771, wc365, n_3664);
  not gc365 (wc365, n_3665);
  and g4347 (n_3774, wc366, n_3530);
  not gc366 (wc366, n_3668);
  and g4348 (n_3777, n_3671, wc367);
  not gc367 (wc367, n_3672);
  and g4349 (n_3780, n_3675, wc368);
  not gc368 (wc368, n_3676);
  and g4350 (n_3783, n_3679, wc369);
  not gc369 (wc369, n_3680);
  and g4351 (n_3786, n_3683, wc370);
  not gc370 (wc370, n_3684);
  and g4352 (n_3789, n_3687, wc371);
  not gc371 (wc371, n_3688);
  and g4353 (n_3792, n_3691, wc372);
  not gc372 (wc372, n_3692);
  or g4354 (n_3704, wc373, n_2983);
  not gc373 (wc373, n_3702);
  or g4355 (n_3709, n_3706, wc374);
  not gc374 (wc374, n_3702);
  or g4356 (n_3711, wc375, n_3360);
  not gc375 (wc375, n_3702);
  or g4357 (n_3725, n_3722, wc376);
  not gc376 (wc376, n_3702);
  or g4358 (n_3729, wc377, n_3726);
  not gc377 (wc377, n_3702);
  or g4359 (n_3733, n_3730, wc378);
  not gc378 (wc378, n_3702);
  or g4360 (n_3737, n_3734, wc379);
  not gc379 (wc379, n_3702);
  or g4361 (n_3741, wc380, n_3738);
  not gc380 (wc380, n_3702);
  or g4362 (n_3745, wc381, n_3742);
  not gc381 (wc381, n_3702);
  or g4363 (n_3749, wc382, n_3746);
  not gc382 (wc382, n_3702);
  or g4364 (n_3751, wc383, n_3642);
  not gc383 (wc383, n_3702);
  and g4365 (n_3822, wc384, n_3098);
  not gc384 (wc384, n_3567);
  and g4366 (n_3826, wc385, n_3290);
  not gc385 (wc385, n_3572);
  and g4367 (n_3830, n_3575, wc386);
  not gc386 (wc386, n_3576);
  and g4368 (n_3834, n_3432, wc387);
  not gc387 (wc387, n_3579);
  and g4369 (n_3838, wc388, n_3584);
  not gc388 (wc388, n_3585);
  and g4370 (n_3795, n_3695, wc389);
  not gc389 (wc389, n_3696);
  and g4371 (n_3798, n_3699, wc390);
  not gc390 (wc390, n_3700);
  or g4372 (n_3802, wc391, n_3079);
  not gc391 (wc391, n_3800);
  or g4373 (n_3807, n_3804, wc392);
  not gc392 (wc392, n_3800);
  or g4374 (n_3809, wc393, n_3420);
  not gc393 (wc393, n_3800);
  or g4375 (n_3823, n_3820, wc394);
  not gc394 (wc394, n_3800);
  or g4376 (n_3827, wc395, n_3824);
  not gc395 (wc395, n_3800);
  or g4377 (n_3831, n_3828, wc396);
  not gc396 (wc396, n_3800);
  or g4378 (n_3835, n_3832, wc397);
  not gc397 (wc397, n_3800);
  or g4379 (n_3839, wc398, n_3836);
  not gc398 (wc398, n_3800);
  not g4380 (Z[77], n_4033);
endmodule

module mult_signed_const_13291_GENERIC(A, Z);
  input [58:0] A;
  output [77:0] Z;
  wire [58:0] A;
  wire [77:0] Z;
  mult_signed_const_13291_GENERIC_REAL g1(.A ({A[58:2], A[0], A[0]}),
       .Z (Z));
endmodule

module mult_signed_const_13758_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [58:0] A;
  output [77:0] Z;
  wire [58:0] A;
  wire [77:0] Z;
  wire n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78;
  wire n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_295, n_296, n_297;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_310, n_311, n_312, n_313;
  wire n_314, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538;
  wire n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562;
  wire n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578;
  wire n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586;
  wire n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594;
  wire n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602;
  wire n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610;
  wire n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618;
  wire n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626;
  wire n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634;
  wire n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642;
  wire n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650;
  wire n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658;
  wire n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666;
  wire n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674;
  wire n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682;
  wire n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690;
  wire n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698;
  wire n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706;
  wire n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714;
  wire n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722;
  wire n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730;
  wire n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738;
  wire n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746;
  wire n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754;
  wire n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762;
  wire n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770;
  wire n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778;
  wire n_779, n_780, n_781, n_782, n_783, n_784, n_785, n_786;
  wire n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794;
  wire n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802;
  wire n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810;
  wire n_811, n_812, n_813, n_814, n_815, n_816, n_817, n_818;
  wire n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826;
  wire n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834;
  wire n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842;
  wire n_843, n_844, n_845, n_846, n_847, n_848, n_849, n_850;
  wire n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858;
  wire n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866;
  wire n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874;
  wire n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882;
  wire n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890;
  wire n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898;
  wire n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906;
  wire n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914;
  wire n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922;
  wire n_923, n_924, n_927, n_928, n_929, n_930, n_931, n_932;
  wire n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940;
  wire n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951;
  wire n_952, n_953, n_954, n_955, n_956, n_957, n_959, n_960;
  wire n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968;
  wire n_969, n_970, n_971, n_972, n_975, n_976, n_977, n_978;
  wire n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986;
  wire n_987, n_989, n_990, n_992, n_993, n_994, n_995, n_996;
  wire n_997, n_998, n_999, n_1000, n_1004, n_1006, n_1007, n_1008;
  wire n_1009, n_1010, n_1011, n_1012, n_1013, n_1015, n_1019, n_1020;
  wire n_1021, n_1022, n_1023, n_1024, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1037, n_1040, n_1041, n_1042, n_1043;
  wire n_1044, n_1050, n_1051, n_1052, n_1053, n_1057, n_1058, n_1059;
  wire n_1060, n_1064, n_1065, n_1066, n_1067, n_1069, n_1071, n_1072;
  wire n_1076, n_1077, n_1079, n_1080, n_1083, n_1086, n_1087, n_1088;
  wire n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1097;
  wire n_1098, n_1099, n_1100, n_1101, n_1105, n_1106, n_1107, n_1108;
  wire n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1116, n_1117;
  wire n_1118, n_1119, n_1120, n_1121, n_1122, n_1124, n_1126, n_1127;
  wire n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135;
  wire n_1136, n_1137, n_1138, n_1142, n_1143, n_1144, n_1145, n_1146;
  wire n_1147, n_1148, n_1149, n_1152, n_1156, n_1157, n_1158, n_1159;
  wire n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167;
  wire n_1168, n_1169, n_1170, n_1174, n_1175, n_1176, n_1177, n_1178;
  wire n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186;
  wire n_1187, n_1188, n_1190, n_1191, n_1193, n_1194, n_1195, n_1196;
  wire n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204;
  wire n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1213, n_1216;
  wire n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224;
  wire n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1233, n_1234;
  wire n_1235, n_1236, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243;
  wire n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251;
  wire n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1260;
  wire n_1262, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271;
  wire n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279;
  wire n_1280, n_1281, n_1282, n_1283, n_1285, n_1286, n_1288, n_1289;
  wire n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299;
  wire n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307;
  wire n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1316, n_1318;
  wire n_1319, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328;
  wire n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336;
  wire n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344;
  wire n_1345, n_1350, n_1351, n_1352, n_1354, n_1355, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1382, n_1383, n_1386, n_1387;
  wire n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395;
  wire n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403;
  wire n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1412, n_1413;
  wire n_1414, n_1415, n_1416, n_1418, n_1419, n_1420, n_1421, n_1422;
  wire n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430;
  wire n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438;
  wire n_1439, n_1440, n_1441, n_1444, n_1446, n_1447, n_1450, n_1451;
  wire n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467;
  wire n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1476, n_1478;
  wire n_1479, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488;
  wire n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496;
  wire n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504;
  wire n_1505, n_1508, n_1510, n_1511, n_1514, n_1515, n_1516, n_1517;
  wire n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525;
  wire n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533;
  wire n_1534, n_1535, n_1536, n_1537, n_1540, n_1542, n_1543, n_1546;
  wire n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554;
  wire n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562;
  wire n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1572;
  wire n_1574, n_1575, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583;
  wire n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591;
  wire n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599;
  wire n_1600, n_1601, n_1604, n_1606, n_1607, n_1610, n_1611, n_1612;
  wire n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620;
  wire n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628;
  wire n_1629, n_1630, n_1631, n_1632, n_1633, n_1636, n_1638, n_1639;
  wire n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649;
  wire n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657;
  wire n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665;
  wire n_1668, n_1670, n_1671, n_1674, n_1675, n_1676, n_1677, n_1678;
  wire n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686;
  wire n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694;
  wire n_1695, n_1696, n_1697, n_1700, n_1702, n_1703, n_1706, n_1707;
  wire n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715;
  wire n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723;
  wire n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1732, n_1734;
  wire n_1735, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744;
  wire n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752;
  wire n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760;
  wire n_1761, n_1764, n_1766, n_1767, n_1770, n_1771, n_1772, n_1773;
  wire n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781;
  wire n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789;
  wire n_1790, n_1791, n_1792, n_1793, n_1796, n_1798, n_1799, n_1802;
  wire n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810;
  wire n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818;
  wire n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1828;
  wire n_1830, n_1831, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839;
  wire n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847;
  wire n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855;
  wire n_1856, n_1857, n_1860, n_1862, n_1863, n_1866, n_1867, n_1868;
  wire n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876;
  wire n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884;
  wire n_1885, n_1886, n_1887, n_1888, n_1889, n_1892, n_1894, n_1895;
  wire n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905;
  wire n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913;
  wire n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921;
  wire n_1924, n_1926, n_1927, n_1930, n_1931, n_1932, n_1933, n_1934;
  wire n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942;
  wire n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950;
  wire n_1951, n_1952, n_1953, n_1956, n_1958, n_1959, n_1962, n_1963;
  wire n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971;
  wire n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979;
  wire n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1988, n_1990;
  wire n_1991, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000;
  wire n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008;
  wire n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016;
  wire n_2017, n_2020, n_2022, n_2023, n_2026, n_2027, n_2028, n_2029;
  wire n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037;
  wire n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045;
  wire n_2046, n_2047, n_2048, n_2049, n_2052, n_2054, n_2055, n_2058;
  wire n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066;
  wire n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074;
  wire n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2084;
  wire n_2086, n_2087, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095;
  wire n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103;
  wire n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111;
  wire n_2112, n_2113, n_2116, n_2118, n_2119, n_2122, n_2123, n_2124;
  wire n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132;
  wire n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140;
  wire n_2141, n_2142, n_2143, n_2144, n_2145, n_2148, n_2150, n_2151;
  wire n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161;
  wire n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169;
  wire n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177;
  wire n_2180, n_2182, n_2183, n_2186, n_2187, n_2188, n_2189, n_2190;
  wire n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198;
  wire n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206;
  wire n_2207, n_2208, n_2209, n_2212, n_2214, n_2215, n_2218, n_2219;
  wire n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227;
  wire n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235;
  wire n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2244, n_2246;
  wire n_2247, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256;
  wire n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264;
  wire n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272;
  wire n_2273, n_2276, n_2278, n_2279, n_2282, n_2283, n_2284, n_2285;
  wire n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293;
  wire n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301;
  wire n_2302, n_2303, n_2304, n_2305, n_2308, n_2310, n_2311, n_2314;
  wire n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322;
  wire n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330;
  wire n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2340;
  wire n_2342, n_2343, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351;
  wire n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359;
  wire n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367;
  wire n_2368, n_2369, n_2372, n_2374, n_2375, n_2378, n_2379, n_2380;
  wire n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388;
  wire n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396;
  wire n_2397, n_2398, n_2399, n_2400, n_2401, n_2404, n_2406, n_2407;
  wire n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417;
  wire n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425;
  wire n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433;
  wire n_2436, n_2438, n_2439, n_2442, n_2443, n_2444, n_2445, n_2446;
  wire n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454;
  wire n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462;
  wire n_2463, n_2464, n_2465, n_2468, n_2470, n_2471, n_2474, n_2475;
  wire n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483;
  wire n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491;
  wire n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2500, n_2502;
  wire n_2503, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512;
  wire n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520;
  wire n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528;
  wire n_2529, n_2532, n_2534, n_2535, n_2538, n_2539, n_2540, n_2541;
  wire n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549;
  wire n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557;
  wire n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2566;
  wire n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577;
  wire n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585;
  wire n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2593, n_2594;
  wire n_2595, n_2598, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606;
  wire n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614;
  wire n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622;
  wire n_2623, n_2624, n_2625, n_2628, n_2630, n_2633, n_2634, n_2635;
  wire n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643;
  wire n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651;
  wire n_2652, n_2653, n_2654, n_2655, n_2658, n_2662, n_2663, n_2664;
  wire n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672;
  wire n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680;
  wire n_2681, n_2686, n_2689, n_2692, n_2693, n_2694, n_2695, n_2696;
  wire n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704;
  wire n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2718, n_2720;
  wire n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728;
  wire n_2729, n_2730, n_2731, n_2732, n_2733, n_2742, n_2744, n_2745;
  wire n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753;
  wire n_2754, n_2755, n_2756, n_2757, n_2764, n_2765, n_2766, n_2767;
  wire n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775;
  wire n_2776, n_2777, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791;
  wire n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2804, n_2805;
  wire n_2806, n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2820;
  wire n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828;
  wire n_2829, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2846;
  wire n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2856;
  wire n_2857, n_2858, n_2859, n_2860, n_2861, n_2865, n_2866, n_2867;
  wire n_2868, n_2869, n_2871, n_2872, n_2873, n_2876, n_2877, n_2889;
  wire n_2891, n_2893, n_2894, n_2895, n_2896, n_2897, n_2899, n_2900;
  wire n_2901, n_2902, n_2903, n_2905, n_2906, n_2907, n_2908, n_2909;
  wire n_2911, n_2912, n_2913, n_2914, n_2915, n_2917, n_2918, n_2919;
  wire n_2920, n_2921, n_2923, n_2924, n_2925, n_2926, n_2927, n_2929;
  wire n_2930, n_2931, n_2932, n_2933, n_2935, n_2936, n_2937, n_2938;
  wire n_2939, n_2941, n_2942, n_2943, n_2944, n_2945, n_2947, n_2948;
  wire n_2949, n_2950, n_2951, n_2953, n_2954, n_2955, n_2956, n_2957;
  wire n_2959, n_2960, n_2961, n_2962, n_2963, n_2965, n_2966, n_2967;
  wire n_2968, n_2969, n_2971, n_2972, n_2973, n_2974, n_2975, n_2977;
  wire n_2978, n_2979, n_2980, n_2981, n_2983, n_2984, n_2985, n_2986;
  wire n_2987, n_2989, n_2990, n_2991, n_2992, n_2993, n_2995, n_2996;
  wire n_2997, n_2998, n_2999, n_3001, n_3002, n_3003, n_3004, n_3005;
  wire n_3007, n_3008, n_3009, n_3010, n_3011, n_3013, n_3014, n_3015;
  wire n_3016, n_3017, n_3019, n_3020, n_3021, n_3022, n_3023, n_3025;
  wire n_3026, n_3027, n_3028, n_3029, n_3031, n_3032, n_3033, n_3034;
  wire n_3035, n_3037, n_3038, n_3039, n_3040, n_3041, n_3043, n_3044;
  wire n_3045, n_3046, n_3047, n_3049, n_3050, n_3051, n_3052, n_3053;
  wire n_3055, n_3056, n_3057, n_3058, n_3059, n_3061, n_3062, n_3063;
  wire n_3064, n_3065, n_3067, n_3068, n_3069, n_3070, n_3071, n_3073;
  wire n_3074, n_3075, n_3076, n_3077, n_3079, n_3080, n_3081, n_3082;
  wire n_3083, n_3085, n_3086, n_3087, n_3088, n_3089, n_3091, n_3092;
  wire n_3093, n_3094, n_3095, n_3097, n_3098, n_3099, n_3100, n_3101;
  wire n_3103, n_3104, n_3105, n_3106, n_3107, n_3109, n_3110, n_3113;
  wire n_3116, n_3118, n_3119, n_3121, n_3122, n_3124, n_3125, n_3126;
  wire n_3128, n_3129, n_3131, n_3132, n_3133, n_3135, n_3136, n_3138;
  wire n_3139, n_3140, n_3142, n_3143, n_3145, n_3146, n_3147, n_3149;
  wire n_3150, n_3152, n_3153, n_3154, n_3156, n_3157, n_3159, n_3160;
  wire n_3161, n_3163, n_3164, n_3166, n_3167, n_3168, n_3170, n_3171;
  wire n_3173, n_3174, n_3175, n_3177, n_3178, n_3180, n_3181, n_3182;
  wire n_3184, n_3185, n_3187, n_3188, n_3189, n_3191, n_3192, n_3194;
  wire n_3195, n_3196, n_3198, n_3199, n_3201, n_3202, n_3203, n_3205;
  wire n_3206, n_3208, n_3209, n_3210, n_3212, n_3213, n_3215, n_3216;
  wire n_3217, n_3219, n_3220, n_3222, n_3223, n_3224, n_3226, n_3227;
  wire n_3229, n_3230, n_3231, n_3233, n_3234, n_3236, n_3237, n_3238;
  wire n_3240, n_3241, n_3243, n_3244, n_3247, n_3248, n_3249, n_3250;
  wire n_3251, n_3252, n_3254, n_3255, n_3256, n_3257, n_3258, n_3260;
  wire n_3261, n_3262, n_3263, n_3264, n_3266, n_3267, n_3268, n_3269;
  wire n_3270, n_3272, n_3273, n_3274, n_3275, n_3276, n_3278, n_3279;
  wire n_3280, n_3281, n_3282, n_3284, n_3285, n_3286, n_3287, n_3288;
  wire n_3290, n_3291, n_3292, n_3293, n_3294, n_3296, n_3297, n_3298;
  wire n_3299, n_3300, n_3301, n_3302, n_3304, n_3305, n_3307, n_3308;
  wire n_3309, n_3311, n_3312, n_3314, n_3315, n_3316, n_3318, n_3319;
  wire n_3321, n_3322, n_3323, n_3325, n_3326, n_3327, n_3328, n_3329;
  wire n_3330, n_3332, n_3333, n_3334, n_3335, n_3336, n_3338, n_3339;
  wire n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3348;
  wire n_3350, n_3351, n_3353, n_3355, n_3356, n_3358, n_3360, n_3361;
  wire n_3363, n_3365, n_3366, n_3367, n_3369, n_3370, n_3371, n_3372;
  wire n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, n_3380;
  wire n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388;
  wire n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396;
  wire n_3397, n_3401, n_3402, n_3404, n_3406, n_3407, n_3409, n_3411;
  wire n_3412, n_3414, n_3416, n_3417, n_3419, n_3421, n_3422, n_3424;
  wire n_3426, n_3427, n_3429, n_3431, n_3432, n_3434, n_3436, n_3437;
  wire n_3439, n_3441, n_3442, n_3444, n_3446, n_3447, n_3449, n_3451;
  wire n_3452, n_3454, n_3456, n_3457, n_3459, n_3461, n_3462, n_3464;
  wire n_3466, n_3467, n_3469, n_3471, n_3472, n_3474, n_3476, n_3477;
  wire n_3479, n_3481, n_3482, n_3484, n_3486, n_3487, n_3489, n_3491;
  wire n_3493, n_3496, n_3497, n_3499, n_3500, n_3501, n_3503, n_3504;
  wire n_3505, n_3507, n_3508, n_3509, n_3511, n_3512, n_3513, n_3515;
  wire n_3516, n_3517, n_3519, n_3520, n_3521, n_3523, n_3524, n_3525;
  wire n_3527, n_3528, n_3529, n_3531, n_3532, n_3533, n_3535, n_3536;
  wire n_3537, n_3539, n_3540, n_3541, n_3543, n_3544, n_3545, n_3547;
  wire n_3548, n_3549, n_3551, n_3552, n_3553, n_3555, n_3556, n_3557;
  wire n_3559, n_3560, n_3561, n_3563, n_3564, n_3565, n_3567, n_3568;
  wire n_3569, n_3571, n_3572, n_3573, n_3575, n_3576, n_3577, n_3579;
  wire n_3580, n_3581, n_3583, n_3584, n_3585, n_3587, n_3588, n_3589;
  wire n_3591, n_3592, n_3593, n_3595, n_3596, n_3597, n_3599, n_3600;
  wire n_3601, n_3603, n_3604, n_3605, n_3607, n_3608, n_3609, n_3611;
  wire n_3612, n_3613, n_3615, n_3616, n_3617, n_3619, n_3620, n_3621;
  wire n_3623, n_3624, n_3625, n_3627, n_3628, n_3629, n_3631, n_3632;
  wire n_3633, n_3635, n_3636, n_3637, n_3639, n_3640, n_3641, n_3643;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g468 (n_211, A[4], A[0]);
  and g2 (n_132, A[4], A[0]);
  xor g469 (n_1086, A[5], A[3]);
  xor g470 (n_210, n_1086, A[1]);
  nand g3 (n_1087, A[5], A[3]);
  nand g471 (n_1088, A[1], A[3]);
  nand g472 (n_1089, A[5], A[1]);
  nand g473 (n_131, n_1087, n_1088, n_1089);
  xor g474 (n_295, A[6], A[4]);
  and g475 (n_296, A[6], A[4]);
  xor g476 (n_1090, A[0], A[2]);
  xor g477 (n_209, n_1090, n_295);
  nand g478 (n_1091, A[0], A[2]);
  nand g4 (n_1092, n_295, A[2]);
  nand g5 (n_1093, A[0], n_295);
  nand g479 (n_130, n_1091, n_1092, n_1093);
  xor g480 (n_1094, A[7], A[5]);
  xor g481 (n_297, n_1094, A[1]);
  nand g482 (n_1095, A[7], A[5]);
  nand g484 (n_1097, A[7], A[1]);
  nand g6 (n_299, n_1095, n_1089, n_1097);
  xor g485 (n_1098, A[3], n_296);
  xor g486 (n_208, n_1098, n_297);
  nand g487 (n_1099, A[3], n_296);
  nand g488 (n_1100, n_297, n_296);
  nand g489 (n_1101, A[3], n_297);
  nand g490 (n_129, n_1099, n_1100, n_1101);
  xor g491 (n_298, A[8], A[6]);
  and g492 (n_301, A[8], A[6]);
  xor g494 (n_300, n_1090, A[4]);
  nand g497 (n_1105, A[2], A[4]);
  xor g499 (n_1106, n_298, n_299);
  xor g500 (n_207, n_1106, n_300);
  nand g501 (n_1107, n_298, n_299);
  nand g502 (n_1108, n_300, n_299);
  nand g503 (n_1109, n_298, n_300);
  nand g504 (n_128, n_1107, n_1108, n_1109);
  xor g505 (n_1110, A[9], A[7]);
  xor g506 (n_303, n_1110, A[3]);
  nand g507 (n_1111, A[9], A[7]);
  nand g508 (n_1112, A[3], A[7]);
  nand g509 (n_1113, A[9], A[3]);
  nand g510 (n_306, n_1111, n_1112, n_1113);
  xor g511 (n_1114, A[1], A[5]);
  xor g512 (n_304, n_1114, n_301);
  nand g514 (n_1116, n_301, A[5]);
  nand g515 (n_1117, A[1], n_301);
  nand g516 (n_308, n_1089, n_1116, n_1117);
  xor g517 (n_1118, n_302, n_303);
  xor g518 (n_206, n_1118, n_304);
  nand g519 (n_1119, n_302, n_303);
  nand g520 (n_1120, n_304, n_303);
  nand g521 (n_1121, n_302, n_304);
  nand g522 (n_127, n_1119, n_1120, n_1121);
  xor g523 (n_305, A[10], A[8]);
  and g524 (n_310, A[10], A[8]);
  xor g525 (n_1122, A[4], A[2]);
  xor g526 (n_307, n_1122, A[6]);
  nand g528 (n_1124, A[6], A[2]);
  xor g531 (n_1126, A[0], n_305);
  xor g532 (n_309, n_1126, n_306);
  nand g533 (n_1127, A[0], n_305);
  nand g534 (n_1128, n_306, n_305);
  nand g535 (n_1129, A[0], n_306);
  nand g536 (n_314, n_1127, n_1128, n_1129);
  xor g537 (n_1130, n_307, n_308);
  xor g538 (n_205, n_1130, n_309);
  nand g539 (n_1131, n_307, n_308);
  nand g540 (n_1132, n_309, n_308);
  nand g541 (n_1133, n_307, n_309);
  nand g542 (n_126, n_1131, n_1132, n_1133);
  xor g543 (n_1134, A[11], A[9]);
  xor g544 (n_312, n_1134, A[5]);
  nand g545 (n_1135, A[11], A[9]);
  nand g546 (n_1136, A[5], A[9]);
  nand g547 (n_1137, A[11], A[5]);
  nand g548 (n_317, n_1135, n_1136, n_1137);
  xor g549 (n_1138, A[3], A[7]);
  xor g550 (n_313, n_1138, A[1]);
  nand g554 (n_318, n_1112, n_1097, n_1088);
  xor g555 (n_1142, n_310, n_311);
  xor g556 (n_315, n_1142, n_312);
  nand g557 (n_1143, n_310, n_311);
  nand g558 (n_1144, n_312, n_311);
  nand g559 (n_1145, n_310, n_312);
  nand g560 (n_322, n_1143, n_1144, n_1145);
  xor g561 (n_1146, n_313, n_314);
  xor g562 (n_204, n_1146, n_315);
  nand g563 (n_1147, n_313, n_314);
  nand g564 (n_1148, n_315, n_314);
  nand g565 (n_1149, n_313, n_315);
  nand g566 (n_125, n_1147, n_1148, n_1149);
  xor g567 (n_316, A[12], A[10]);
  and g568 (n_323, A[12], A[10]);
  xor g570 (n_319, n_295, A[8]);
  nand g572 (n_1152, A[8], A[4]);
  xor g576 (n_320, n_1090, n_316);
  nand g578 (n_1156, n_316, A[0]);
  nand g579 (n_1157, A[2], n_316);
  nand g580 (n_327, n_1091, n_1156, n_1157);
  xor g581 (n_1158, n_317, n_318);
  xor g582 (n_321, n_1158, n_319);
  nand g583 (n_1159, n_317, n_318);
  nand g584 (n_1160, n_319, n_318);
  nand g585 (n_1161, n_317, n_319);
  nand g586 (n_329, n_1159, n_1160, n_1161);
  xor g587 (n_1162, n_320, n_321);
  xor g588 (n_203, n_1162, n_322);
  nand g589 (n_1163, n_320, n_321);
  nand g590 (n_1164, n_322, n_321);
  nand g591 (n_1165, n_320, n_322);
  nand g592 (n_124, n_1163, n_1164, n_1165);
  xor g593 (n_1166, A[13], A[11]);
  xor g594 (n_326, n_1166, A[7]);
  nand g595 (n_1167, A[13], A[11]);
  nand g596 (n_1168, A[7], A[11]);
  nand g597 (n_1169, A[13], A[7]);
  nand g598 (n_332, n_1167, n_1168, n_1169);
  xor g599 (n_1170, A[5], A[9]);
  xor g600 (n_325, n_1170, A[3]);
  nand g604 (n_333, n_1136, n_1113, n_1087);
  xor g605 (n_1174, A[1], n_323);
  xor g606 (n_328, n_1174, n_324);
  nand g607 (n_1175, A[1], n_323);
  nand g608 (n_1176, n_324, n_323);
  nand g609 (n_1177, A[1], n_324);
  nand g610 (n_336, n_1175, n_1176, n_1177);
  xor g611 (n_1178, n_325, n_326);
  xor g612 (n_330, n_1178, n_327);
  nand g613 (n_1179, n_325, n_326);
  nand g614 (n_1180, n_327, n_326);
  nand g615 (n_1181, n_325, n_327);
  nand g616 (n_338, n_1179, n_1180, n_1181);
  xor g617 (n_1182, n_328, n_329);
  xor g618 (n_202, n_1182, n_330);
  nand g619 (n_1183, n_328, n_329);
  nand g620 (n_1184, n_330, n_329);
  nand g621 (n_1185, n_328, n_330);
  nand g622 (n_123, n_1183, n_1184, n_1185);
  xor g623 (n_331, A[14], A[12]);
  and g624 (n_340, A[14], A[12]);
  xor g625 (n_1186, A[8], A[0]);
  xor g626 (n_335, n_1186, A[6]);
  nand g627 (n_1187, A[8], A[0]);
  nand g628 (n_1188, A[6], A[0]);
  xor g631 (n_1190, A[10], A[4]);
  xor g632 (n_334, n_1190, A[2]);
  nand g633 (n_1191, A[10], A[4]);
  nand g635 (n_1193, A[10], A[2]);
  nand g636 (n_342, n_1191, n_1105, n_1193);
  xor g637 (n_1194, n_331, n_332);
  xor g638 (n_337, n_1194, n_333);
  nand g639 (n_1195, n_331, n_332);
  nand g640 (n_1196, n_333, n_332);
  nand g641 (n_1197, n_331, n_333);
  nand g642 (n_346, n_1195, n_1196, n_1197);
  xor g643 (n_1198, n_334, n_335);
  xor g644 (n_339, n_1198, n_336);
  nand g645 (n_1199, n_334, n_335);
  nand g646 (n_1200, n_336, n_335);
  nand g647 (n_1201, n_334, n_336);
  nand g648 (n_349, n_1199, n_1200, n_1201);
  xor g649 (n_1202, n_337, n_338);
  xor g650 (n_201, n_1202, n_339);
  nand g651 (n_1203, n_337, n_338);
  nand g652 (n_1204, n_339, n_338);
  nand g653 (n_1205, n_337, n_339);
  nand g654 (n_122, n_1203, n_1204, n_1205);
  xor g655 (n_1206, A[15], A[13]);
  xor g656 (n_343, n_1206, A[9]);
  nand g657 (n_1207, A[15], A[13]);
  nand g658 (n_1208, A[9], A[13]);
  nand g659 (n_1209, A[15], A[9]);
  nand g660 (n_351, n_1207, n_1208, n_1209);
  xor g661 (n_1210, A[1], A[7]);
  xor g662 (n_344, n_1210, A[11]);
  nand g665 (n_1213, A[1], A[11]);
  nand g666 (n_352, n_1097, n_1168, n_1213);
  xor g668 (n_345, n_1086, n_340);
  nand g670 (n_1216, n_340, A[3]);
  nand g671 (n_1217, A[5], n_340);
  nand g672 (n_355, n_1087, n_1216, n_1217);
  xor g673 (n_1218, n_341, n_342);
  xor g674 (n_347, n_1218, n_343);
  nand g675 (n_1219, n_341, n_342);
  nand g676 (n_1220, n_343, n_342);
  nand g677 (n_1221, n_341, n_343);
  nand g678 (n_357, n_1219, n_1220, n_1221);
  xor g679 (n_1222, n_344, n_345);
  xor g680 (n_348, n_1222, n_346);
  nand g681 (n_1223, n_344, n_345);
  nand g682 (n_1224, n_346, n_345);
  nand g683 (n_1225, n_344, n_346);
  nand g684 (n_359, n_1223, n_1224, n_1225);
  xor g685 (n_1226, n_347, n_348);
  xor g686 (n_200, n_1226, n_349);
  nand g687 (n_1227, n_347, n_348);
  nand g688 (n_1228, n_349, n_348);
  nand g689 (n_1229, n_347, n_349);
  nand g690 (n_121, n_1227, n_1228, n_1229);
  xor g691 (n_350, A[16], A[14]);
  and g692 (n_361, A[16], A[14]);
  xor g693 (n_1230, A[10], A[2]);
  xor g694 (n_354, n_1230, A[0]);
  nand g697 (n_1233, A[10], A[0]);
  nand g698 (n_362, n_1193, n_1091, n_1233);
  xor g699 (n_1234, A[8], A[12]);
  xor g700 (n_353, n_1234, A[6]);
  nand g701 (n_1235, A[8], A[12]);
  nand g702 (n_1236, A[6], A[12]);
  xor g705 (n_1238, A[4], n_350);
  xor g706 (n_356, n_1238, n_351);
  nand g707 (n_1239, A[4], n_350);
  nand g708 (n_1240, n_351, n_350);
  nand g709 (n_1241, A[4], n_351);
  nand g710 (n_367, n_1239, n_1240, n_1241);
  xor g711 (n_1242, n_352, n_353);
  xor g712 (n_358, n_1242, n_354);
  nand g713 (n_1243, n_352, n_353);
  nand g714 (n_1244, n_354, n_353);
  nand g715 (n_1245, n_352, n_354);
  nand g716 (n_369, n_1243, n_1244, n_1245);
  xor g717 (n_1246, n_355, n_356);
  xor g718 (n_360, n_1246, n_357);
  nand g719 (n_1247, n_355, n_356);
  nand g720 (n_1248, n_357, n_356);
  nand g721 (n_1249, n_355, n_357);
  nand g722 (n_371, n_1247, n_1248, n_1249);
  xor g723 (n_1250, n_358, n_359);
  xor g724 (n_199, n_1250, n_360);
  nand g725 (n_1251, n_358, n_359);
  nand g726 (n_1252, n_360, n_359);
  nand g727 (n_1253, n_358, n_360);
  nand g728 (n_120, n_1251, n_1252, n_1253);
  xor g729 (n_1254, A[17], A[15]);
  xor g730 (n_365, n_1254, A[11]);
  nand g731 (n_1255, A[17], A[15]);
  nand g732 (n_1256, A[11], A[15]);
  nand g733 (n_1257, A[17], A[11]);
  nand g734 (n_374, n_1255, n_1256, n_1257);
  xor g735 (n_1258, A[3], A[1]);
  xor g736 (n_366, n_1258, A[9]);
  nand g738 (n_1260, A[9], A[1]);
  nand g740 (n_376, n_1088, n_1260, n_1113);
  xor g741 (n_1262, A[13], A[7]);
  xor g742 (n_364, n_1262, A[5]);
  nand g745 (n_1265, A[13], A[5]);
  nand g746 (n_375, n_1169, n_1095, n_1265);
  xor g747 (n_1266, n_361, n_362);
  xor g748 (n_368, n_1266, n_363);
  nand g749 (n_1267, n_361, n_362);
  nand g750 (n_1268, n_363, n_362);
  nand g751 (n_1269, n_361, n_363);
  nand g752 (n_380, n_1267, n_1268, n_1269);
  xor g753 (n_1270, n_364, n_365);
  xor g754 (n_370, n_1270, n_366);
  nand g755 (n_1271, n_364, n_365);
  nand g756 (n_1272, n_366, n_365);
  nand g757 (n_1273, n_364, n_366);
  nand g758 (n_382, n_1271, n_1272, n_1273);
  xor g759 (n_1274, n_367, n_368);
  xor g760 (n_372, n_1274, n_369);
  nand g761 (n_1275, n_367, n_368);
  nand g762 (n_1276, n_369, n_368);
  nand g763 (n_1277, n_367, n_369);
  nand g764 (n_384, n_1275, n_1276, n_1277);
  xor g765 (n_1278, n_370, n_371);
  xor g766 (n_198, n_1278, n_372);
  nand g767 (n_1279, n_370, n_371);
  nand g768 (n_1280, n_372, n_371);
  nand g769 (n_1281, n_370, n_372);
  nand g770 (n_119, n_1279, n_1280, n_1281);
  xor g771 (n_373, A[18], A[16]);
  and g772 (n_386, A[18], A[16]);
  xor g773 (n_1282, A[12], A[4]);
  xor g774 (n_377, n_1282, A[2]);
  nand g775 (n_1283, A[12], A[4]);
  nand g777 (n_1285, A[12], A[2]);
  nand g778 (n_387, n_1283, n_1105, n_1285);
  xor g779 (n_1286, A[10], A[0]);
  xor g780 (n_378, n_1286, A[14]);
  nand g782 (n_1288, A[14], A[0]);
  nand g783 (n_1289, A[10], A[14]);
  nand g784 (n_388, n_1233, n_1288, n_1289);
  xor g786 (n_379, n_298, n_373);
  nand g788 (n_1292, n_373, A[6]);
  nand g789 (n_1293, A[8], n_373);
  xor g791 (n_1294, n_374, n_375);
  xor g792 (n_381, n_1294, n_376);
  nand g793 (n_1295, n_374, n_375);
  nand g794 (n_1296, n_376, n_375);
  nand g795 (n_1297, n_374, n_376);
  nand g796 (n_394, n_1295, n_1296, n_1297);
  xor g797 (n_1298, n_377, n_378);
  xor g798 (n_383, n_1298, n_379);
  nand g799 (n_1299, n_377, n_378);
  nand g800 (n_1300, n_379, n_378);
  nand g801 (n_1301, n_377, n_379);
  nand g802 (n_395, n_1299, n_1300, n_1301);
  xor g803 (n_1302, n_380, n_381);
  xor g804 (n_385, n_1302, n_382);
  nand g805 (n_1303, n_380, n_381);
  nand g806 (n_1304, n_382, n_381);
  nand g807 (n_1305, n_380, n_382);
  nand g808 (n_398, n_1303, n_1304, n_1305);
  xor g809 (n_1306, n_383, n_384);
  xor g810 (n_197, n_1306, n_385);
  nand g811 (n_1307, n_383, n_384);
  nand g812 (n_1308, n_385, n_384);
  nand g813 (n_1309, n_383, n_385);
  nand g814 (n_118, n_1307, n_1308, n_1309);
  xor g815 (n_1310, A[19], A[17]);
  xor g816 (n_390, n_1310, A[13]);
  nand g817 (n_1311, A[19], A[17]);
  nand g818 (n_1312, A[13], A[17]);
  nand g819 (n_1313, A[19], A[13]);
  nand g820 (n_400, n_1311, n_1312, n_1313);
  xor g822 (n_391, n_1086, A[11]);
  nand g824 (n_1316, A[11], A[3]);
  nand g826 (n_401, n_1087, n_1316, n_1137);
  xor g827 (n_1318, A[1], A[15]);
  xor g828 (n_389, n_1318, A[9]);
  nand g829 (n_1319, A[1], A[15]);
  nand g832 (n_402, n_1319, n_1209, n_1260);
  xor g833 (n_1322, A[7], n_386);
  xor g834 (n_393, n_1322, n_387);
  nand g835 (n_1323, A[7], n_386);
  nand g836 (n_1324, n_387, n_386);
  nand g837 (n_1325, A[7], n_387);
  nand g838 (n_134, n_1323, n_1324, n_1325);
  xor g839 (n_1326, n_388, n_389);
  xor g840 (n_396, n_1326, n_390);
  nand g841 (n_1327, n_388, n_389);
  nand g842 (n_1328, n_390, n_389);
  nand g843 (n_1329, n_388, n_390);
  nand g844 (n_136, n_1327, n_1328, n_1329);
  xor g845 (n_1330, n_391, n_392);
  xor g846 (n_397, n_1330, n_393);
  nand g847 (n_1331, n_391, n_392);
  nand g848 (n_1332, n_393, n_392);
  nand g849 (n_1333, n_391, n_393);
  nand g850 (n_405, n_1331, n_1332, n_1333);
  xor g851 (n_1334, n_394, n_395);
  xor g852 (n_399, n_1334, n_396);
  nand g853 (n_1335, n_394, n_395);
  nand g854 (n_1336, n_396, n_395);
  nand g855 (n_1337, n_394, n_396);
  nand g856 (n_407, n_1335, n_1336, n_1337);
  xor g857 (n_1338, n_397, n_398);
  xor g858 (n_196, n_1338, n_399);
  nand g859 (n_1339, n_397, n_398);
  nand g860 (n_1340, n_399, n_398);
  nand g861 (n_1341, n_397, n_399);
  nand g862 (n_117, n_1339, n_1340, n_1341);
  xor g863 (n_1342, A[20], A[18]);
  xor g864 (n_404, n_1342, A[14]);
  nand g865 (n_1343, A[20], A[18]);
  nand g866 (n_1344, A[14], A[18]);
  nand g867 (n_1345, A[20], A[14]);
  nand g868 (n_409, n_1343, n_1344, n_1345);
  xor g870 (n_133, n_295, A[12]);
  xor g875 (n_1350, A[2], A[16]);
  xor g876 (n_403, n_1350, A[10]);
  nand g877 (n_1351, A[2], A[16]);
  nand g878 (n_1352, A[10], A[16]);
  nand g880 (n_411, n_1351, n_1352, n_1193);
  xor g881 (n_1354, A[8], n_400);
  xor g882 (n_135, n_1354, n_401);
  nand g883 (n_1355, A[8], n_400);
  nand g884 (n_1356, n_401, n_400);
  nand g885 (n_1357, A[8], n_401);
  nand g886 (n_415, n_1355, n_1356, n_1357);
  xor g887 (n_1358, n_402, n_403);
  xor g888 (n_137, n_1358, n_404);
  nand g889 (n_1359, n_402, n_403);
  nand g890 (n_1360, n_404, n_403);
  nand g891 (n_1361, n_402, n_404);
  nand g892 (n_417, n_1359, n_1360, n_1361);
  xor g893 (n_1362, n_133, n_134);
  xor g894 (n_406, n_1362, n_135);
  nand g895 (n_1363, n_133, n_134);
  nand g896 (n_1364, n_135, n_134);
  nand g897 (n_1365, n_133, n_135);
  nand g898 (n_419, n_1363, n_1364, n_1365);
  xor g899 (n_1366, n_136, n_137);
  xor g900 (n_408, n_1366, n_405);
  nand g901 (n_1367, n_136, n_137);
  nand g902 (n_1368, n_405, n_137);
  nand g903 (n_1369, n_136, n_405);
  nand g904 (n_421, n_1367, n_1368, n_1369);
  xor g905 (n_1370, n_406, n_407);
  xor g906 (n_195, n_1370, n_408);
  nand g907 (n_1371, n_406, n_407);
  nand g908 (n_1372, n_408, n_407);
  nand g909 (n_1373, n_406, n_408);
  nand g910 (n_116, n_1371, n_1372, n_1373);
  xor g911 (n_1374, A[21], A[19]);
  xor g912 (n_413, n_1374, A[15]);
  nand g913 (n_1375, A[21], A[19]);
  nand g914 (n_1376, A[15], A[19]);
  nand g915 (n_1377, A[21], A[15]);
  nand g916 (n_423, n_1375, n_1376, n_1377);
  xor g918 (n_414, n_1094, A[13]);
  xor g923 (n_1382, A[3], A[17]);
  xor g924 (n_412, n_1382, A[11]);
  nand g925 (n_1383, A[3], A[17]);
  nand g928 (n_425, n_1383, n_1257, n_1316);
  xor g929 (n_1386, A[9], n_409);
  xor g930 (n_416, n_1386, n_410);
  nand g931 (n_1387, A[9], n_409);
  nand g932 (n_1388, n_410, n_409);
  nand g933 (n_1389, A[9], n_410);
  nand g934 (n_429, n_1387, n_1388, n_1389);
  xor g935 (n_1390, n_411, n_412);
  xor g936 (n_418, n_1390, n_413);
  nand g937 (n_1391, n_411, n_412);
  nand g938 (n_1392, n_413, n_412);
  nand g939 (n_1393, n_411, n_413);
  nand g940 (n_431, n_1391, n_1392, n_1393);
  xor g941 (n_1394, n_414, n_415);
  xor g942 (n_420, n_1394, n_416);
  nand g943 (n_1395, n_414, n_415);
  nand g944 (n_1396, n_416, n_415);
  nand g945 (n_1397, n_414, n_416);
  nand g946 (n_433, n_1395, n_1396, n_1397);
  xor g947 (n_1398, n_417, n_418);
  xor g948 (n_422, n_1398, n_419);
  nand g949 (n_1399, n_417, n_418);
  nand g950 (n_1400, n_419, n_418);
  nand g951 (n_1401, n_417, n_419);
  nand g952 (n_436, n_1399, n_1400, n_1401);
  xor g953 (n_1402, n_420, n_421);
  xor g954 (n_194, n_1402, n_422);
  nand g955 (n_1403, n_420, n_421);
  nand g956 (n_1404, n_422, n_421);
  nand g957 (n_1405, n_420, n_422);
  nand g958 (n_115, n_1403, n_1404, n_1405);
  xor g959 (n_1406, A[22], A[20]);
  xor g960 (n_427, n_1406, A[16]);
  nand g961 (n_1407, A[22], A[20]);
  nand g962 (n_1408, A[16], A[20]);
  nand g963 (n_1409, A[22], A[16]);
  nand g964 (n_437, n_1407, n_1408, n_1409);
  xor g966 (n_428, n_298, A[14]);
  nand g968 (n_1412, A[14], A[6]);
  nand g969 (n_1413, A[8], A[14]);
  xor g971 (n_1414, A[4], A[18]);
  xor g972 (n_426, n_1414, A[12]);
  nand g973 (n_1415, A[4], A[18]);
  nand g974 (n_1416, A[12], A[18]);
  nand g976 (n_439, n_1415, n_1416, n_1283);
  xor g977 (n_1418, A[10], n_423);
  xor g978 (n_430, n_1418, n_375);
  nand g979 (n_1419, A[10], n_423);
  nand g980 (n_1420, n_375, n_423);
  nand g981 (n_1421, A[10], n_375);
  nand g982 (n_443, n_1419, n_1420, n_1421);
  xor g983 (n_1422, n_425, n_426);
  xor g984 (n_432, n_1422, n_427);
  nand g985 (n_1423, n_425, n_426);
  nand g986 (n_1424, n_427, n_426);
  nand g987 (n_1425, n_425, n_427);
  nand g988 (n_445, n_1423, n_1424, n_1425);
  xor g989 (n_1426, n_428, n_429);
  xor g990 (n_434, n_1426, n_430);
  nand g991 (n_1427, n_428, n_429);
  nand g992 (n_1428, n_430, n_429);
  nand g993 (n_1429, n_428, n_430);
  nand g994 (n_447, n_1427, n_1428, n_1429);
  xor g995 (n_1430, n_431, n_432);
  xor g996 (n_435, n_1430, n_433);
  nand g997 (n_1431, n_431, n_432);
  nand g998 (n_1432, n_433, n_432);
  nand g999 (n_1433, n_431, n_433);
  nand g1000 (n_450, n_1431, n_1432, n_1433);
  xor g1001 (n_1434, n_434, n_435);
  xor g1002 (n_193, n_1434, n_436);
  nand g1003 (n_1435, n_434, n_435);
  nand g1004 (n_1436, n_436, n_435);
  nand g1005 (n_1437, n_434, n_436);
  nand g1006 (n_114, n_1435, n_1436, n_1437);
  xor g1007 (n_1438, A[23], A[21]);
  xor g1008 (n_441, n_1438, A[17]);
  nand g1009 (n_1439, A[23], A[21]);
  nand g1010 (n_1440, A[17], A[21]);
  nand g1011 (n_1441, A[23], A[17]);
  nand g1012 (n_451, n_1439, n_1440, n_1441);
  xor g1014 (n_442, n_1110, A[15]);
  nand g1016 (n_1444, A[15], A[7]);
  nand g1018 (n_452, n_1111, n_1444, n_1209);
  xor g1019 (n_1446, A[5], A[19]);
  xor g1020 (n_440, n_1446, A[13]);
  nand g1021 (n_1447, A[5], A[19]);
  nand g1024 (n_453, n_1447, n_1313, n_1265);
  xor g1025 (n_1450, A[11], n_437);
  xor g1026 (n_444, n_1450, n_438);
  nand g1027 (n_1451, A[11], n_437);
  nand g1028 (n_1452, n_438, n_437);
  nand g1029 (n_1453, A[11], n_438);
  nand g1030 (n_457, n_1451, n_1452, n_1453);
  xor g1031 (n_1454, n_439, n_440);
  xor g1032 (n_446, n_1454, n_441);
  nand g1033 (n_1455, n_439, n_440);
  nand g1034 (n_1456, n_441, n_440);
  nand g1035 (n_1457, n_439, n_441);
  nand g1036 (n_459, n_1455, n_1456, n_1457);
  xor g1037 (n_1458, n_442, n_443);
  xor g1038 (n_448, n_1458, n_444);
  nand g1039 (n_1459, n_442, n_443);
  nand g1040 (n_1460, n_444, n_443);
  nand g1041 (n_1461, n_442, n_444);
  nand g1042 (n_461, n_1459, n_1460, n_1461);
  xor g1043 (n_1462, n_445, n_446);
  xor g1044 (n_449, n_1462, n_447);
  nand g1045 (n_1463, n_445, n_446);
  nand g1046 (n_1464, n_447, n_446);
  nand g1047 (n_1465, n_445, n_447);
  nand g1048 (n_464, n_1463, n_1464, n_1465);
  xor g1049 (n_1466, n_448, n_449);
  xor g1050 (n_192, n_1466, n_450);
  nand g1051 (n_1467, n_448, n_449);
  nand g1052 (n_1468, n_450, n_449);
  nand g1053 (n_1469, n_448, n_450);
  nand g1054 (n_113, n_1467, n_1468, n_1469);
  xor g1055 (n_1470, A[24], A[22]);
  xor g1056 (n_455, n_1470, A[18]);
  nand g1057 (n_1471, A[24], A[22]);
  nand g1058 (n_1472, A[18], A[22]);
  nand g1059 (n_1473, A[24], A[18]);
  nand g1060 (n_465, n_1471, n_1472, n_1473);
  xor g1062 (n_456, n_305, A[16]);
  nand g1064 (n_1476, A[16], A[8]);
  xor g1067 (n_1478, A[6], A[20]);
  xor g1068 (n_454, n_1478, A[14]);
  nand g1069 (n_1479, A[6], A[20]);
  nand g1072 (n_467, n_1479, n_1345, n_1412);
  xor g1073 (n_1482, A[12], n_451);
  xor g1074 (n_458, n_1482, n_452);
  nand g1075 (n_1483, A[12], n_451);
  nand g1076 (n_1484, n_452, n_451);
  nand g1077 (n_1485, A[12], n_452);
  nand g1078 (n_471, n_1483, n_1484, n_1485);
  xor g1079 (n_1486, n_453, n_454);
  xor g1080 (n_460, n_1486, n_455);
  nand g1081 (n_1487, n_453, n_454);
  nand g1082 (n_1488, n_455, n_454);
  nand g1083 (n_1489, n_453, n_455);
  nand g1084 (n_473, n_1487, n_1488, n_1489);
  xor g1085 (n_1490, n_456, n_457);
  xor g1086 (n_462, n_1490, n_458);
  nand g1087 (n_1491, n_456, n_457);
  nand g1088 (n_1492, n_458, n_457);
  nand g1089 (n_1493, n_456, n_458);
  nand g1090 (n_213, n_1491, n_1492, n_1493);
  xor g1091 (n_1494, n_459, n_460);
  xor g1092 (n_463, n_1494, n_461);
  nand g1093 (n_1495, n_459, n_460);
  nand g1094 (n_1496, n_461, n_460);
  nand g1095 (n_1497, n_459, n_461);
  nand g1096 (n_476, n_1495, n_1496, n_1497);
  xor g1097 (n_1498, n_462, n_463);
  xor g1098 (n_191, n_1498, n_464);
  nand g1099 (n_1499, n_462, n_463);
  nand g1100 (n_1500, n_464, n_463);
  nand g1101 (n_1501, n_462, n_464);
  nand g1102 (n_112, n_1499, n_1500, n_1501);
  xor g1103 (n_1502, A[25], A[23]);
  xor g1104 (n_469, n_1502, A[19]);
  nand g1105 (n_1503, A[25], A[23]);
  nand g1106 (n_1504, A[19], A[23]);
  nand g1107 (n_1505, A[25], A[19]);
  nand g1108 (n_477, n_1503, n_1504, n_1505);
  xor g1110 (n_470, n_1134, A[17]);
  nand g1112 (n_1508, A[17], A[9]);
  nand g1114 (n_478, n_1135, n_1508, n_1257);
  xor g1115 (n_1510, A[7], A[21]);
  xor g1116 (n_468, n_1510, A[15]);
  nand g1117 (n_1511, A[7], A[21]);
  nand g1120 (n_479, n_1511, n_1377, n_1444);
  xor g1121 (n_1514, A[13], n_465);
  xor g1122 (n_472, n_1514, n_466);
  nand g1123 (n_1515, A[13], n_465);
  nand g1124 (n_1516, n_466, n_465);
  nand g1125 (n_1517, A[13], n_466);
  nand g1126 (n_483, n_1515, n_1516, n_1517);
  xor g1127 (n_1518, n_467, n_468);
  xor g1128 (n_212, n_1518, n_469);
  nand g1129 (n_1519, n_467, n_468);
  nand g1130 (n_1520, n_469, n_468);
  nand g1131 (n_1521, n_467, n_469);
  nand g1132 (n_485, n_1519, n_1520, n_1521);
  xor g1133 (n_1522, n_470, n_471);
  xor g1134 (n_474, n_1522, n_472);
  nand g1135 (n_1523, n_470, n_471);
  nand g1136 (n_1524, n_472, n_471);
  nand g1137 (n_1525, n_470, n_472);
  nand g1138 (n_487, n_1523, n_1524, n_1525);
  xor g1139 (n_1526, n_473, n_212);
  xor g1140 (n_475, n_1526, n_213);
  nand g1141 (n_1527, n_473, n_212);
  nand g1142 (n_1528, n_213, n_212);
  nand g1143 (n_1529, n_473, n_213);
  nand g1144 (n_490, n_1527, n_1528, n_1529);
  xor g1145 (n_1530, n_474, n_475);
  xor g1146 (n_190, n_1530, n_476);
  nand g1147 (n_1531, n_474, n_475);
  nand g1148 (n_1532, n_476, n_475);
  nand g1149 (n_1533, n_474, n_476);
  nand g1150 (n_111, n_1531, n_1532, n_1533);
  xor g1151 (n_1534, A[26], A[24]);
  xor g1152 (n_481, n_1534, A[20]);
  nand g1153 (n_1535, A[26], A[24]);
  nand g1154 (n_1536, A[20], A[24]);
  nand g1155 (n_1537, A[26], A[20]);
  nand g1156 (n_491, n_1535, n_1536, n_1537);
  xor g1158 (n_482, n_316, A[18]);
  nand g1160 (n_1540, A[18], A[10]);
  xor g1163 (n_1542, A[8], A[22]);
  xor g1164 (n_480, n_1542, A[16]);
  nand g1165 (n_1543, A[8], A[22]);
  nand g1168 (n_493, n_1543, n_1409, n_1476);
  xor g1169 (n_1546, A[14], n_477);
  xor g1170 (n_484, n_1546, n_478);
  nand g1171 (n_1547, A[14], n_477);
  nand g1172 (n_1548, n_478, n_477);
  nand g1173 (n_1549, A[14], n_478);
  nand g1174 (n_497, n_1547, n_1548, n_1549);
  xor g1175 (n_1550, n_479, n_480);
  xor g1176 (n_486, n_1550, n_481);
  nand g1177 (n_1551, n_479, n_480);
  nand g1178 (n_1552, n_481, n_480);
  nand g1179 (n_1553, n_479, n_481);
  nand g1180 (n_499, n_1551, n_1552, n_1553);
  xor g1181 (n_1554, n_482, n_483);
  xor g1182 (n_488, n_1554, n_484);
  nand g1183 (n_1555, n_482, n_483);
  nand g1184 (n_1556, n_484, n_483);
  nand g1185 (n_1557, n_482, n_484);
  nand g1186 (n_501, n_1555, n_1556, n_1557);
  xor g1187 (n_1558, n_485, n_486);
  xor g1188 (n_489, n_1558, n_487);
  nand g1189 (n_1559, n_485, n_486);
  nand g1190 (n_1560, n_487, n_486);
  nand g1191 (n_1561, n_485, n_487);
  nand g1192 (n_504, n_1559, n_1560, n_1561);
  xor g1193 (n_1562, n_488, n_489);
  xor g1194 (n_189, n_1562, n_490);
  nand g1195 (n_1563, n_488, n_489);
  nand g1196 (n_1564, n_490, n_489);
  nand g1197 (n_1565, n_488, n_490);
  nand g1198 (n_110, n_1563, n_1564, n_1565);
  xor g1199 (n_1566, A[27], A[25]);
  xor g1200 (n_495, n_1566, A[21]);
  nand g1201 (n_1567, A[27], A[25]);
  nand g1202 (n_1568, A[21], A[25]);
  nand g1203 (n_1569, A[27], A[21]);
  nand g1204 (n_505, n_1567, n_1568, n_1569);
  xor g1206 (n_496, n_1166, A[19]);
  nand g1208 (n_1572, A[19], A[11]);
  nand g1210 (n_506, n_1167, n_1572, n_1313);
  xor g1211 (n_1574, A[9], A[23]);
  xor g1212 (n_494, n_1574, A[17]);
  nand g1213 (n_1575, A[9], A[23]);
  nand g1216 (n_507, n_1575, n_1441, n_1508);
  xor g1217 (n_1578, A[15], n_491);
  xor g1218 (n_498, n_1578, n_492);
  nand g1219 (n_1579, A[15], n_491);
  nand g1220 (n_1580, n_492, n_491);
  nand g1221 (n_1581, A[15], n_492);
  nand g1222 (n_511, n_1579, n_1580, n_1581);
  xor g1223 (n_1582, n_493, n_494);
  xor g1224 (n_500, n_1582, n_495);
  nand g1225 (n_1583, n_493, n_494);
  nand g1226 (n_1584, n_495, n_494);
  nand g1227 (n_1585, n_493, n_495);
  nand g1228 (n_513, n_1583, n_1584, n_1585);
  xor g1229 (n_1586, n_496, n_497);
  xor g1230 (n_502, n_1586, n_498);
  nand g1231 (n_1587, n_496, n_497);
  nand g1232 (n_1588, n_498, n_497);
  nand g1233 (n_1589, n_496, n_498);
  nand g1234 (n_515, n_1587, n_1588, n_1589);
  xor g1235 (n_1590, n_499, n_500);
  xor g1236 (n_503, n_1590, n_501);
  nand g1237 (n_1591, n_499, n_500);
  nand g1238 (n_1592, n_501, n_500);
  nand g1239 (n_1593, n_499, n_501);
  nand g1240 (n_518, n_1591, n_1592, n_1593);
  xor g1241 (n_1594, n_502, n_503);
  xor g1242 (n_188, n_1594, n_504);
  nand g1243 (n_1595, n_502, n_503);
  nand g1244 (n_1596, n_504, n_503);
  nand g1245 (n_1597, n_502, n_504);
  nand g1246 (n_109, n_1595, n_1596, n_1597);
  xor g1247 (n_1598, A[28], A[26]);
  xor g1248 (n_509, n_1598, A[22]);
  nand g1249 (n_1599, A[28], A[26]);
  nand g1250 (n_1600, A[22], A[26]);
  nand g1251 (n_1601, A[28], A[22]);
  nand g1252 (n_519, n_1599, n_1600, n_1601);
  xor g1254 (n_510, n_331, A[20]);
  nand g1256 (n_1604, A[20], A[12]);
  xor g1259 (n_1606, A[10], A[24]);
  xor g1260 (n_508, n_1606, A[18]);
  nand g1261 (n_1607, A[10], A[24]);
  nand g1264 (n_521, n_1607, n_1473, n_1540);
  xor g1265 (n_1610, A[16], n_505);
  xor g1266 (n_512, n_1610, n_506);
  nand g1267 (n_1611, A[16], n_505);
  nand g1268 (n_1612, n_506, n_505);
  nand g1269 (n_1613, A[16], n_506);
  nand g1270 (n_525, n_1611, n_1612, n_1613);
  xor g1271 (n_1614, n_507, n_508);
  xor g1272 (n_514, n_1614, n_509);
  nand g1273 (n_1615, n_507, n_508);
  nand g1274 (n_1616, n_509, n_508);
  nand g1275 (n_1617, n_507, n_509);
  nand g1276 (n_527, n_1615, n_1616, n_1617);
  xor g1277 (n_1618, n_510, n_511);
  xor g1278 (n_516, n_1618, n_512);
  nand g1279 (n_1619, n_510, n_511);
  nand g1280 (n_1620, n_512, n_511);
  nand g1281 (n_1621, n_510, n_512);
  nand g1282 (n_529, n_1619, n_1620, n_1621);
  xor g1283 (n_1622, n_513, n_514);
  xor g1284 (n_517, n_1622, n_515);
  nand g1285 (n_1623, n_513, n_514);
  nand g1286 (n_1624, n_515, n_514);
  nand g1287 (n_1625, n_513, n_515);
  nand g1288 (n_532, n_1623, n_1624, n_1625);
  xor g1289 (n_1626, n_516, n_517);
  xor g1290 (n_187, n_1626, n_518);
  nand g1291 (n_1627, n_516, n_517);
  nand g1292 (n_1628, n_518, n_517);
  nand g1293 (n_1629, n_516, n_518);
  nand g1294 (n_108, n_1627, n_1628, n_1629);
  xor g1295 (n_1630, A[29], A[27]);
  xor g1296 (n_523, n_1630, A[23]);
  nand g1297 (n_1631, A[29], A[27]);
  nand g1298 (n_1632, A[23], A[27]);
  nand g1299 (n_1633, A[29], A[23]);
  nand g1300 (n_533, n_1631, n_1632, n_1633);
  xor g1302 (n_524, n_1206, A[21]);
  nand g1304 (n_1636, A[21], A[13]);
  nand g1306 (n_534, n_1207, n_1636, n_1377);
  xor g1307 (n_1638, A[11], A[25]);
  xor g1308 (n_522, n_1638, A[19]);
  nand g1309 (n_1639, A[11], A[25]);
  nand g1312 (n_535, n_1639, n_1505, n_1572);
  xor g1313 (n_1642, A[17], n_519);
  xor g1314 (n_526, n_1642, n_520);
  nand g1315 (n_1643, A[17], n_519);
  nand g1316 (n_1644, n_520, n_519);
  nand g1317 (n_1645, A[17], n_520);
  nand g1318 (n_539, n_1643, n_1644, n_1645);
  xor g1319 (n_1646, n_521, n_522);
  xor g1320 (n_528, n_1646, n_523);
  nand g1321 (n_1647, n_521, n_522);
  nand g1322 (n_1648, n_523, n_522);
  nand g1323 (n_1649, n_521, n_523);
  nand g1324 (n_541, n_1647, n_1648, n_1649);
  xor g1325 (n_1650, n_524, n_525);
  xor g1326 (n_530, n_1650, n_526);
  nand g1327 (n_1651, n_524, n_525);
  nand g1328 (n_1652, n_526, n_525);
  nand g1329 (n_1653, n_524, n_526);
  nand g1330 (n_543, n_1651, n_1652, n_1653);
  xor g1331 (n_1654, n_527, n_528);
  xor g1332 (n_531, n_1654, n_529);
  nand g1333 (n_1655, n_527, n_528);
  nand g1334 (n_1656, n_529, n_528);
  nand g1335 (n_1657, n_527, n_529);
  nand g1336 (n_546, n_1655, n_1656, n_1657);
  xor g1337 (n_1658, n_530, n_531);
  xor g1338 (n_186, n_1658, n_532);
  nand g1339 (n_1659, n_530, n_531);
  nand g1340 (n_1660, n_532, n_531);
  nand g1341 (n_1661, n_530, n_532);
  nand g1342 (n_107, n_1659, n_1660, n_1661);
  xor g1343 (n_1662, A[30], A[28]);
  xor g1344 (n_537, n_1662, A[24]);
  nand g1345 (n_1663, A[30], A[28]);
  nand g1346 (n_1664, A[24], A[28]);
  nand g1347 (n_1665, A[30], A[24]);
  nand g1348 (n_547, n_1663, n_1664, n_1665);
  xor g1350 (n_538, n_350, A[22]);
  nand g1352 (n_1668, A[22], A[14]);
  xor g1355 (n_1670, A[12], A[26]);
  xor g1356 (n_536, n_1670, A[20]);
  nand g1357 (n_1671, A[12], A[26]);
  nand g1360 (n_549, n_1671, n_1537, n_1604);
  xor g1361 (n_1674, A[18], n_533);
  xor g1362 (n_540, n_1674, n_534);
  nand g1363 (n_1675, A[18], n_533);
  nand g1364 (n_1676, n_534, n_533);
  nand g1365 (n_1677, A[18], n_534);
  nand g1366 (n_553, n_1675, n_1676, n_1677);
  xor g1367 (n_1678, n_535, n_536);
  xor g1368 (n_542, n_1678, n_537);
  nand g1369 (n_1679, n_535, n_536);
  nand g1370 (n_1680, n_537, n_536);
  nand g1371 (n_1681, n_535, n_537);
  nand g1372 (n_555, n_1679, n_1680, n_1681);
  xor g1373 (n_1682, n_538, n_539);
  xor g1374 (n_544, n_1682, n_540);
  nand g1375 (n_1683, n_538, n_539);
  nand g1376 (n_1684, n_540, n_539);
  nand g1377 (n_1685, n_538, n_540);
  nand g1378 (n_557, n_1683, n_1684, n_1685);
  xor g1379 (n_1686, n_541, n_542);
  xor g1380 (n_545, n_1686, n_543);
  nand g1381 (n_1687, n_541, n_542);
  nand g1382 (n_1688, n_543, n_542);
  nand g1383 (n_1689, n_541, n_543);
  nand g1384 (n_560, n_1687, n_1688, n_1689);
  xor g1385 (n_1690, n_544, n_545);
  xor g1386 (n_185, n_1690, n_546);
  nand g1387 (n_1691, n_544, n_545);
  nand g1388 (n_1692, n_546, n_545);
  nand g1389 (n_1693, n_544, n_546);
  nand g1390 (n_106, n_1691, n_1692, n_1693);
  xor g1391 (n_1694, A[31], A[29]);
  xor g1392 (n_551, n_1694, A[25]);
  nand g1393 (n_1695, A[31], A[29]);
  nand g1394 (n_1696, A[25], A[29]);
  nand g1395 (n_1697, A[31], A[25]);
  nand g1396 (n_561, n_1695, n_1696, n_1697);
  xor g1398 (n_552, n_1254, A[23]);
  nand g1400 (n_1700, A[23], A[15]);
  nand g1402 (n_562, n_1255, n_1700, n_1441);
  xor g1403 (n_1702, A[13], A[27]);
  xor g1404 (n_550, n_1702, A[21]);
  nand g1405 (n_1703, A[13], A[27]);
  nand g1408 (n_563, n_1703, n_1569, n_1636);
  xor g1409 (n_1706, A[19], n_547);
  xor g1410 (n_554, n_1706, n_548);
  nand g1411 (n_1707, A[19], n_547);
  nand g1412 (n_1708, n_548, n_547);
  nand g1413 (n_1709, A[19], n_548);
  nand g1414 (n_567, n_1707, n_1708, n_1709);
  xor g1415 (n_1710, n_549, n_550);
  xor g1416 (n_556, n_1710, n_551);
  nand g1417 (n_1711, n_549, n_550);
  nand g1418 (n_1712, n_551, n_550);
  nand g1419 (n_1713, n_549, n_551);
  nand g1420 (n_569, n_1711, n_1712, n_1713);
  xor g1421 (n_1714, n_552, n_553);
  xor g1422 (n_558, n_1714, n_554);
  nand g1423 (n_1715, n_552, n_553);
  nand g1424 (n_1716, n_554, n_553);
  nand g1425 (n_1717, n_552, n_554);
  nand g1426 (n_571, n_1715, n_1716, n_1717);
  xor g1427 (n_1718, n_555, n_556);
  xor g1428 (n_559, n_1718, n_557);
  nand g1429 (n_1719, n_555, n_556);
  nand g1430 (n_1720, n_557, n_556);
  nand g1431 (n_1721, n_555, n_557);
  nand g1432 (n_574, n_1719, n_1720, n_1721);
  xor g1433 (n_1722, n_558, n_559);
  xor g1434 (n_184, n_1722, n_560);
  nand g1435 (n_1723, n_558, n_559);
  nand g1436 (n_1724, n_560, n_559);
  nand g1437 (n_1725, n_558, n_560);
  nand g1438 (n_105, n_1723, n_1724, n_1725);
  xor g1439 (n_1726, A[32], A[30]);
  xor g1440 (n_565, n_1726, A[26]);
  nand g1441 (n_1727, A[32], A[30]);
  nand g1442 (n_1728, A[26], A[30]);
  nand g1443 (n_1729, A[32], A[26]);
  nand g1444 (n_575, n_1727, n_1728, n_1729);
  xor g1446 (n_566, n_373, A[24]);
  nand g1448 (n_1732, A[24], A[16]);
  xor g1451 (n_1734, A[14], A[28]);
  xor g1452 (n_564, n_1734, A[22]);
  nand g1453 (n_1735, A[14], A[28]);
  nand g1456 (n_577, n_1735, n_1601, n_1668);
  xor g1457 (n_1738, A[20], n_561);
  xor g1458 (n_568, n_1738, n_562);
  nand g1459 (n_1739, A[20], n_561);
  nand g1460 (n_1740, n_562, n_561);
  nand g1461 (n_1741, A[20], n_562);
  nand g1462 (n_581, n_1739, n_1740, n_1741);
  xor g1463 (n_1742, n_563, n_564);
  xor g1464 (n_570, n_1742, n_565);
  nand g1465 (n_1743, n_563, n_564);
  nand g1466 (n_1744, n_565, n_564);
  nand g1467 (n_1745, n_563, n_565);
  nand g1468 (n_583, n_1743, n_1744, n_1745);
  xor g1469 (n_1746, n_566, n_567);
  xor g1470 (n_572, n_1746, n_568);
  nand g1471 (n_1747, n_566, n_567);
  nand g1472 (n_1748, n_568, n_567);
  nand g1473 (n_1749, n_566, n_568);
  nand g1474 (n_585, n_1747, n_1748, n_1749);
  xor g1475 (n_1750, n_569, n_570);
  xor g1476 (n_573, n_1750, n_571);
  nand g1477 (n_1751, n_569, n_570);
  nand g1478 (n_1752, n_571, n_570);
  nand g1479 (n_1753, n_569, n_571);
  nand g1480 (n_588, n_1751, n_1752, n_1753);
  xor g1481 (n_1754, n_572, n_573);
  xor g1482 (n_183, n_1754, n_574);
  nand g1483 (n_1755, n_572, n_573);
  nand g1484 (n_1756, n_574, n_573);
  nand g1485 (n_1757, n_572, n_574);
  nand g1486 (n_104, n_1755, n_1756, n_1757);
  xor g1487 (n_1758, A[33], A[31]);
  xor g1488 (n_579, n_1758, A[27]);
  nand g1489 (n_1759, A[33], A[31]);
  nand g1490 (n_1760, A[27], A[31]);
  nand g1491 (n_1761, A[33], A[27]);
  nand g1492 (n_589, n_1759, n_1760, n_1761);
  xor g1494 (n_580, n_1310, A[25]);
  nand g1496 (n_1764, A[25], A[17]);
  nand g1498 (n_590, n_1311, n_1764, n_1505);
  xor g1499 (n_1766, A[15], A[29]);
  xor g1500 (n_578, n_1766, A[23]);
  nand g1501 (n_1767, A[15], A[29]);
  nand g1504 (n_591, n_1767, n_1633, n_1700);
  xor g1505 (n_1770, A[21], n_575);
  xor g1506 (n_582, n_1770, n_576);
  nand g1507 (n_1771, A[21], n_575);
  nand g1508 (n_1772, n_576, n_575);
  nand g1509 (n_1773, A[21], n_576);
  nand g1510 (n_595, n_1771, n_1772, n_1773);
  xor g1511 (n_1774, n_577, n_578);
  xor g1512 (n_584, n_1774, n_579);
  nand g1513 (n_1775, n_577, n_578);
  nand g1514 (n_1776, n_579, n_578);
  nand g1515 (n_1777, n_577, n_579);
  nand g1516 (n_597, n_1775, n_1776, n_1777);
  xor g1517 (n_1778, n_580, n_581);
  xor g1518 (n_586, n_1778, n_582);
  nand g1519 (n_1779, n_580, n_581);
  nand g1520 (n_1780, n_582, n_581);
  nand g1521 (n_1781, n_580, n_582);
  nand g1522 (n_599, n_1779, n_1780, n_1781);
  xor g1523 (n_1782, n_583, n_584);
  xor g1524 (n_587, n_1782, n_585);
  nand g1525 (n_1783, n_583, n_584);
  nand g1526 (n_1784, n_585, n_584);
  nand g1527 (n_1785, n_583, n_585);
  nand g1528 (n_602, n_1783, n_1784, n_1785);
  xor g1529 (n_1786, n_586, n_587);
  xor g1530 (n_182, n_1786, n_588);
  nand g1531 (n_1787, n_586, n_587);
  nand g1532 (n_1788, n_588, n_587);
  nand g1533 (n_1789, n_586, n_588);
  nand g1534 (n_103, n_1787, n_1788, n_1789);
  xor g1535 (n_1790, A[34], A[32]);
  xor g1536 (n_593, n_1790, A[28]);
  nand g1537 (n_1791, A[34], A[32]);
  nand g1538 (n_1792, A[28], A[32]);
  nand g1539 (n_1793, A[34], A[28]);
  nand g1540 (n_603, n_1791, n_1792, n_1793);
  xor g1542 (n_594, n_1342, A[26]);
  nand g1544 (n_1796, A[26], A[18]);
  nand g1546 (n_604, n_1343, n_1796, n_1537);
  xor g1547 (n_1798, A[16], A[30]);
  xor g1548 (n_592, n_1798, A[24]);
  nand g1549 (n_1799, A[16], A[30]);
  nand g1552 (n_605, n_1799, n_1665, n_1732);
  xor g1553 (n_1802, A[22], n_589);
  xor g1554 (n_596, n_1802, n_590);
  nand g1555 (n_1803, A[22], n_589);
  nand g1556 (n_1804, n_590, n_589);
  nand g1557 (n_1805, A[22], n_590);
  nand g1558 (n_609, n_1803, n_1804, n_1805);
  xor g1559 (n_1806, n_591, n_592);
  xor g1560 (n_598, n_1806, n_593);
  nand g1561 (n_1807, n_591, n_592);
  nand g1562 (n_1808, n_593, n_592);
  nand g1563 (n_1809, n_591, n_593);
  nand g1564 (n_611, n_1807, n_1808, n_1809);
  xor g1565 (n_1810, n_594, n_595);
  xor g1566 (n_600, n_1810, n_596);
  nand g1567 (n_1811, n_594, n_595);
  nand g1568 (n_1812, n_596, n_595);
  nand g1569 (n_1813, n_594, n_596);
  nand g1570 (n_613, n_1811, n_1812, n_1813);
  xor g1571 (n_1814, n_597, n_598);
  xor g1572 (n_601, n_1814, n_599);
  nand g1573 (n_1815, n_597, n_598);
  nand g1574 (n_1816, n_599, n_598);
  nand g1575 (n_1817, n_597, n_599);
  nand g1576 (n_616, n_1815, n_1816, n_1817);
  xor g1577 (n_1818, n_600, n_601);
  xor g1578 (n_181, n_1818, n_602);
  nand g1579 (n_1819, n_600, n_601);
  nand g1580 (n_1820, n_602, n_601);
  nand g1581 (n_1821, n_600, n_602);
  nand g1582 (n_102, n_1819, n_1820, n_1821);
  xor g1583 (n_1822, A[35], A[33]);
  xor g1584 (n_607, n_1822, A[29]);
  nand g1585 (n_1823, A[35], A[33]);
  nand g1586 (n_1824, A[29], A[33]);
  nand g1587 (n_1825, A[35], A[29]);
  nand g1588 (n_617, n_1823, n_1824, n_1825);
  xor g1590 (n_608, n_1374, A[27]);
  nand g1592 (n_1828, A[27], A[19]);
  nand g1594 (n_618, n_1375, n_1828, n_1569);
  xor g1595 (n_1830, A[17], A[31]);
  xor g1596 (n_606, n_1830, A[25]);
  nand g1597 (n_1831, A[17], A[31]);
  nand g1600 (n_619, n_1831, n_1697, n_1764);
  xor g1601 (n_1834, A[23], n_603);
  xor g1602 (n_610, n_1834, n_604);
  nand g1603 (n_1835, A[23], n_603);
  nand g1604 (n_1836, n_604, n_603);
  nand g1605 (n_1837, A[23], n_604);
  nand g1606 (n_623, n_1835, n_1836, n_1837);
  xor g1607 (n_1838, n_605, n_606);
  xor g1608 (n_612, n_1838, n_607);
  nand g1609 (n_1839, n_605, n_606);
  nand g1610 (n_1840, n_607, n_606);
  nand g1611 (n_1841, n_605, n_607);
  nand g1612 (n_625, n_1839, n_1840, n_1841);
  xor g1613 (n_1842, n_608, n_609);
  xor g1614 (n_614, n_1842, n_610);
  nand g1615 (n_1843, n_608, n_609);
  nand g1616 (n_1844, n_610, n_609);
  nand g1617 (n_1845, n_608, n_610);
  nand g1618 (n_627, n_1843, n_1844, n_1845);
  xor g1619 (n_1846, n_611, n_612);
  xor g1620 (n_615, n_1846, n_613);
  nand g1621 (n_1847, n_611, n_612);
  nand g1622 (n_1848, n_613, n_612);
  nand g1623 (n_1849, n_611, n_613);
  nand g1624 (n_630, n_1847, n_1848, n_1849);
  xor g1625 (n_1850, n_614, n_615);
  xor g1626 (n_180, n_1850, n_616);
  nand g1627 (n_1851, n_614, n_615);
  nand g1628 (n_1852, n_616, n_615);
  nand g1629 (n_1853, n_614, n_616);
  nand g1630 (n_101, n_1851, n_1852, n_1853);
  xor g1631 (n_1854, A[36], A[34]);
  xor g1632 (n_621, n_1854, A[30]);
  nand g1633 (n_1855, A[36], A[34]);
  nand g1634 (n_1856, A[30], A[34]);
  nand g1635 (n_1857, A[36], A[30]);
  nand g1636 (n_631, n_1855, n_1856, n_1857);
  xor g1638 (n_622, n_1406, A[28]);
  nand g1640 (n_1860, A[28], A[20]);
  nand g1642 (n_632, n_1407, n_1860, n_1601);
  xor g1643 (n_1862, A[18], A[32]);
  xor g1644 (n_620, n_1862, A[26]);
  nand g1645 (n_1863, A[18], A[32]);
  nand g1648 (n_633, n_1863, n_1729, n_1796);
  xor g1649 (n_1866, A[24], n_617);
  xor g1650 (n_624, n_1866, n_618);
  nand g1651 (n_1867, A[24], n_617);
  nand g1652 (n_1868, n_618, n_617);
  nand g1653 (n_1869, A[24], n_618);
  nand g1654 (n_637, n_1867, n_1868, n_1869);
  xor g1655 (n_1870, n_619, n_620);
  xor g1656 (n_626, n_1870, n_621);
  nand g1657 (n_1871, n_619, n_620);
  nand g1658 (n_1872, n_621, n_620);
  nand g1659 (n_1873, n_619, n_621);
  nand g1660 (n_639, n_1871, n_1872, n_1873);
  xor g1661 (n_1874, n_622, n_623);
  xor g1662 (n_628, n_1874, n_624);
  nand g1663 (n_1875, n_622, n_623);
  nand g1664 (n_1876, n_624, n_623);
  nand g1665 (n_1877, n_622, n_624);
  nand g1666 (n_641, n_1875, n_1876, n_1877);
  xor g1667 (n_1878, n_625, n_626);
  xor g1668 (n_629, n_1878, n_627);
  nand g1669 (n_1879, n_625, n_626);
  nand g1670 (n_1880, n_627, n_626);
  nand g1671 (n_1881, n_625, n_627);
  nand g1672 (n_644, n_1879, n_1880, n_1881);
  xor g1673 (n_1882, n_628, n_629);
  xor g1674 (n_179, n_1882, n_630);
  nand g1675 (n_1883, n_628, n_629);
  nand g1676 (n_1884, n_630, n_629);
  nand g1677 (n_1885, n_628, n_630);
  nand g1678 (n_100, n_1883, n_1884, n_1885);
  xor g1679 (n_1886, A[37], A[35]);
  xor g1680 (n_635, n_1886, A[31]);
  nand g1681 (n_1887, A[37], A[35]);
  nand g1682 (n_1888, A[31], A[35]);
  nand g1683 (n_1889, A[37], A[31]);
  nand g1684 (n_645, n_1887, n_1888, n_1889);
  xor g1686 (n_636, n_1438, A[29]);
  nand g1688 (n_1892, A[29], A[21]);
  nand g1690 (n_646, n_1439, n_1892, n_1633);
  xor g1691 (n_1894, A[19], A[33]);
  xor g1692 (n_634, n_1894, A[27]);
  nand g1693 (n_1895, A[19], A[33]);
  nand g1696 (n_647, n_1895, n_1761, n_1828);
  xor g1697 (n_1898, A[25], n_631);
  xor g1698 (n_638, n_1898, n_632);
  nand g1699 (n_1899, A[25], n_631);
  nand g1700 (n_1900, n_632, n_631);
  nand g1701 (n_1901, A[25], n_632);
  nand g1702 (n_651, n_1899, n_1900, n_1901);
  xor g1703 (n_1902, n_633, n_634);
  xor g1704 (n_640, n_1902, n_635);
  nand g1705 (n_1903, n_633, n_634);
  nand g1706 (n_1904, n_635, n_634);
  nand g1707 (n_1905, n_633, n_635);
  nand g1708 (n_653, n_1903, n_1904, n_1905);
  xor g1709 (n_1906, n_636, n_637);
  xor g1710 (n_642, n_1906, n_638);
  nand g1711 (n_1907, n_636, n_637);
  nand g1712 (n_1908, n_638, n_637);
  nand g1713 (n_1909, n_636, n_638);
  nand g1714 (n_655, n_1907, n_1908, n_1909);
  xor g1715 (n_1910, n_639, n_640);
  xor g1716 (n_643, n_1910, n_641);
  nand g1717 (n_1911, n_639, n_640);
  nand g1718 (n_1912, n_641, n_640);
  nand g1719 (n_1913, n_639, n_641);
  nand g1720 (n_658, n_1911, n_1912, n_1913);
  xor g1721 (n_1914, n_642, n_643);
  xor g1722 (n_178, n_1914, n_644);
  nand g1723 (n_1915, n_642, n_643);
  nand g1724 (n_1916, n_644, n_643);
  nand g1725 (n_1917, n_642, n_644);
  nand g1726 (n_99, n_1915, n_1916, n_1917);
  xor g1727 (n_1918, A[38], A[36]);
  xor g1728 (n_649, n_1918, A[32]);
  nand g1729 (n_1919, A[38], A[36]);
  nand g1730 (n_1920, A[32], A[36]);
  nand g1731 (n_1921, A[38], A[32]);
  nand g1732 (n_659, n_1919, n_1920, n_1921);
  xor g1734 (n_650, n_1470, A[30]);
  nand g1736 (n_1924, A[30], A[22]);
  nand g1738 (n_660, n_1471, n_1924, n_1665);
  xor g1739 (n_1926, A[20], A[34]);
  xor g1740 (n_648, n_1926, A[28]);
  nand g1741 (n_1927, A[20], A[34]);
  nand g1744 (n_661, n_1927, n_1793, n_1860);
  xor g1745 (n_1930, A[26], n_645);
  xor g1746 (n_652, n_1930, n_646);
  nand g1747 (n_1931, A[26], n_645);
  nand g1748 (n_1932, n_646, n_645);
  nand g1749 (n_1933, A[26], n_646);
  nand g1750 (n_665, n_1931, n_1932, n_1933);
  xor g1751 (n_1934, n_647, n_648);
  xor g1752 (n_654, n_1934, n_649);
  nand g1753 (n_1935, n_647, n_648);
  nand g1754 (n_1936, n_649, n_648);
  nand g1755 (n_1937, n_647, n_649);
  nand g1756 (n_667, n_1935, n_1936, n_1937);
  xor g1757 (n_1938, n_650, n_651);
  xor g1758 (n_656, n_1938, n_652);
  nand g1759 (n_1939, n_650, n_651);
  nand g1760 (n_1940, n_652, n_651);
  nand g1761 (n_1941, n_650, n_652);
  nand g1762 (n_669, n_1939, n_1940, n_1941);
  xor g1763 (n_1942, n_653, n_654);
  xor g1764 (n_657, n_1942, n_655);
  nand g1765 (n_1943, n_653, n_654);
  nand g1766 (n_1944, n_655, n_654);
  nand g1767 (n_1945, n_653, n_655);
  nand g1768 (n_672, n_1943, n_1944, n_1945);
  xor g1769 (n_1946, n_656, n_657);
  xor g1770 (n_177, n_1946, n_658);
  nand g1771 (n_1947, n_656, n_657);
  nand g1772 (n_1948, n_658, n_657);
  nand g1773 (n_1949, n_656, n_658);
  nand g1774 (n_98, n_1947, n_1948, n_1949);
  xor g1775 (n_1950, A[39], A[37]);
  xor g1776 (n_663, n_1950, A[33]);
  nand g1777 (n_1951, A[39], A[37]);
  nand g1778 (n_1952, A[33], A[37]);
  nand g1779 (n_1953, A[39], A[33]);
  nand g1780 (n_673, n_1951, n_1952, n_1953);
  xor g1782 (n_664, n_1502, A[31]);
  nand g1784 (n_1956, A[31], A[23]);
  nand g1786 (n_674, n_1503, n_1956, n_1697);
  xor g1787 (n_1958, A[21], A[35]);
  xor g1788 (n_662, n_1958, A[29]);
  nand g1789 (n_1959, A[21], A[35]);
  nand g1792 (n_675, n_1959, n_1825, n_1892);
  xor g1793 (n_1962, A[27], n_659);
  xor g1794 (n_666, n_1962, n_660);
  nand g1795 (n_1963, A[27], n_659);
  nand g1796 (n_1964, n_660, n_659);
  nand g1797 (n_1965, A[27], n_660);
  nand g1798 (n_679, n_1963, n_1964, n_1965);
  xor g1799 (n_1966, n_661, n_662);
  xor g1800 (n_668, n_1966, n_663);
  nand g1801 (n_1967, n_661, n_662);
  nand g1802 (n_1968, n_663, n_662);
  nand g1803 (n_1969, n_661, n_663);
  nand g1804 (n_681, n_1967, n_1968, n_1969);
  xor g1805 (n_1970, n_664, n_665);
  xor g1806 (n_670, n_1970, n_666);
  nand g1807 (n_1971, n_664, n_665);
  nand g1808 (n_1972, n_666, n_665);
  nand g1809 (n_1973, n_664, n_666);
  nand g1810 (n_683, n_1971, n_1972, n_1973);
  xor g1811 (n_1974, n_667, n_668);
  xor g1812 (n_671, n_1974, n_669);
  nand g1813 (n_1975, n_667, n_668);
  nand g1814 (n_1976, n_669, n_668);
  nand g1815 (n_1977, n_667, n_669);
  nand g1816 (n_686, n_1975, n_1976, n_1977);
  xor g1817 (n_1978, n_670, n_671);
  xor g1818 (n_176, n_1978, n_672);
  nand g1819 (n_1979, n_670, n_671);
  nand g1820 (n_1980, n_672, n_671);
  nand g1821 (n_1981, n_670, n_672);
  nand g1822 (n_97, n_1979, n_1980, n_1981);
  xor g1823 (n_1982, A[40], A[38]);
  xor g1824 (n_677, n_1982, A[34]);
  nand g1825 (n_1983, A[40], A[38]);
  nand g1826 (n_1984, A[34], A[38]);
  nand g1827 (n_1985, A[40], A[34]);
  nand g1828 (n_687, n_1983, n_1984, n_1985);
  xor g1830 (n_678, n_1534, A[32]);
  nand g1832 (n_1988, A[32], A[24]);
  nand g1834 (n_688, n_1535, n_1988, n_1729);
  xor g1835 (n_1990, A[22], A[36]);
  xor g1836 (n_676, n_1990, A[30]);
  nand g1837 (n_1991, A[22], A[36]);
  nand g1840 (n_689, n_1991, n_1857, n_1924);
  xor g1841 (n_1994, A[28], n_673);
  xor g1842 (n_680, n_1994, n_674);
  nand g1843 (n_1995, A[28], n_673);
  nand g1844 (n_1996, n_674, n_673);
  nand g1845 (n_1997, A[28], n_674);
  nand g1846 (n_693, n_1995, n_1996, n_1997);
  xor g1847 (n_1998, n_675, n_676);
  xor g1848 (n_682, n_1998, n_677);
  nand g1849 (n_1999, n_675, n_676);
  nand g1850 (n_2000, n_677, n_676);
  nand g1851 (n_2001, n_675, n_677);
  nand g1852 (n_695, n_1999, n_2000, n_2001);
  xor g1853 (n_2002, n_678, n_679);
  xor g1854 (n_684, n_2002, n_680);
  nand g1855 (n_2003, n_678, n_679);
  nand g1856 (n_2004, n_680, n_679);
  nand g1857 (n_2005, n_678, n_680);
  nand g1858 (n_697, n_2003, n_2004, n_2005);
  xor g1859 (n_2006, n_681, n_682);
  xor g1860 (n_685, n_2006, n_683);
  nand g1861 (n_2007, n_681, n_682);
  nand g1862 (n_2008, n_683, n_682);
  nand g1863 (n_2009, n_681, n_683);
  nand g1864 (n_700, n_2007, n_2008, n_2009);
  xor g1865 (n_2010, n_684, n_685);
  xor g1866 (n_175, n_2010, n_686);
  nand g1867 (n_2011, n_684, n_685);
  nand g1868 (n_2012, n_686, n_685);
  nand g1869 (n_2013, n_684, n_686);
  nand g1870 (n_96, n_2011, n_2012, n_2013);
  xor g1871 (n_2014, A[41], A[39]);
  xor g1872 (n_691, n_2014, A[35]);
  nand g1873 (n_2015, A[41], A[39]);
  nand g1874 (n_2016, A[35], A[39]);
  nand g1875 (n_2017, A[41], A[35]);
  nand g1876 (n_701, n_2015, n_2016, n_2017);
  xor g1878 (n_692, n_1566, A[33]);
  nand g1880 (n_2020, A[33], A[25]);
  nand g1882 (n_702, n_1567, n_2020, n_1761);
  xor g1883 (n_2022, A[23], A[37]);
  xor g1884 (n_690, n_2022, A[31]);
  nand g1885 (n_2023, A[23], A[37]);
  nand g1888 (n_703, n_2023, n_1889, n_1956);
  xor g1889 (n_2026, A[29], n_687);
  xor g1890 (n_694, n_2026, n_688);
  nand g1891 (n_2027, A[29], n_687);
  nand g1892 (n_2028, n_688, n_687);
  nand g1893 (n_2029, A[29], n_688);
  nand g1894 (n_707, n_2027, n_2028, n_2029);
  xor g1895 (n_2030, n_689, n_690);
  xor g1896 (n_696, n_2030, n_691);
  nand g1897 (n_2031, n_689, n_690);
  nand g1898 (n_2032, n_691, n_690);
  nand g1899 (n_2033, n_689, n_691);
  nand g1900 (n_709, n_2031, n_2032, n_2033);
  xor g1901 (n_2034, n_692, n_693);
  xor g1902 (n_698, n_2034, n_694);
  nand g1903 (n_2035, n_692, n_693);
  nand g1904 (n_2036, n_694, n_693);
  nand g1905 (n_2037, n_692, n_694);
  nand g1906 (n_711, n_2035, n_2036, n_2037);
  xor g1907 (n_2038, n_695, n_696);
  xor g1908 (n_699, n_2038, n_697);
  nand g1909 (n_2039, n_695, n_696);
  nand g1910 (n_2040, n_697, n_696);
  nand g1911 (n_2041, n_695, n_697);
  nand g1912 (n_714, n_2039, n_2040, n_2041);
  xor g1913 (n_2042, n_698, n_699);
  xor g1914 (n_174, n_2042, n_700);
  nand g1915 (n_2043, n_698, n_699);
  nand g1916 (n_2044, n_700, n_699);
  nand g1917 (n_2045, n_698, n_700);
  nand g1918 (n_95, n_2043, n_2044, n_2045);
  xor g1919 (n_2046, A[42], A[40]);
  xor g1920 (n_705, n_2046, A[36]);
  nand g1921 (n_2047, A[42], A[40]);
  nand g1922 (n_2048, A[36], A[40]);
  nand g1923 (n_2049, A[42], A[36]);
  nand g1924 (n_715, n_2047, n_2048, n_2049);
  xor g1926 (n_706, n_1598, A[34]);
  nand g1928 (n_2052, A[34], A[26]);
  nand g1930 (n_716, n_1599, n_2052, n_1793);
  xor g1931 (n_2054, A[24], A[38]);
  xor g1932 (n_704, n_2054, A[32]);
  nand g1933 (n_2055, A[24], A[38]);
  nand g1936 (n_717, n_2055, n_1921, n_1988);
  xor g1937 (n_2058, A[30], n_701);
  xor g1938 (n_708, n_2058, n_702);
  nand g1939 (n_2059, A[30], n_701);
  nand g1940 (n_2060, n_702, n_701);
  nand g1941 (n_2061, A[30], n_702);
  nand g1942 (n_721, n_2059, n_2060, n_2061);
  xor g1943 (n_2062, n_703, n_704);
  xor g1944 (n_710, n_2062, n_705);
  nand g1945 (n_2063, n_703, n_704);
  nand g1946 (n_2064, n_705, n_704);
  nand g1947 (n_2065, n_703, n_705);
  nand g1948 (n_723, n_2063, n_2064, n_2065);
  xor g1949 (n_2066, n_706, n_707);
  xor g1950 (n_712, n_2066, n_708);
  nand g1951 (n_2067, n_706, n_707);
  nand g1952 (n_2068, n_708, n_707);
  nand g1953 (n_2069, n_706, n_708);
  nand g1954 (n_725, n_2067, n_2068, n_2069);
  xor g1955 (n_2070, n_709, n_710);
  xor g1956 (n_713, n_2070, n_711);
  nand g1957 (n_2071, n_709, n_710);
  nand g1958 (n_2072, n_711, n_710);
  nand g1959 (n_2073, n_709, n_711);
  nand g1960 (n_728, n_2071, n_2072, n_2073);
  xor g1961 (n_2074, n_712, n_713);
  xor g1962 (n_173, n_2074, n_714);
  nand g1963 (n_2075, n_712, n_713);
  nand g1964 (n_2076, n_714, n_713);
  nand g1965 (n_2077, n_712, n_714);
  nand g1966 (n_94, n_2075, n_2076, n_2077);
  xor g1967 (n_2078, A[43], A[41]);
  xor g1968 (n_719, n_2078, A[37]);
  nand g1969 (n_2079, A[43], A[41]);
  nand g1970 (n_2080, A[37], A[41]);
  nand g1971 (n_2081, A[43], A[37]);
  nand g1972 (n_729, n_2079, n_2080, n_2081);
  xor g1974 (n_720, n_1630, A[35]);
  nand g1976 (n_2084, A[35], A[27]);
  nand g1978 (n_730, n_1631, n_2084, n_1825);
  xor g1979 (n_2086, A[25], A[39]);
  xor g1980 (n_718, n_2086, A[33]);
  nand g1981 (n_2087, A[25], A[39]);
  nand g1984 (n_731, n_2087, n_1953, n_2020);
  xor g1985 (n_2090, A[31], n_715);
  xor g1986 (n_722, n_2090, n_716);
  nand g1987 (n_2091, A[31], n_715);
  nand g1988 (n_2092, n_716, n_715);
  nand g1989 (n_2093, A[31], n_716);
  nand g1990 (n_735, n_2091, n_2092, n_2093);
  xor g1991 (n_2094, n_717, n_718);
  xor g1992 (n_724, n_2094, n_719);
  nand g1993 (n_2095, n_717, n_718);
  nand g1994 (n_2096, n_719, n_718);
  nand g1995 (n_2097, n_717, n_719);
  nand g1996 (n_737, n_2095, n_2096, n_2097);
  xor g1997 (n_2098, n_720, n_721);
  xor g1998 (n_726, n_2098, n_722);
  nand g1999 (n_2099, n_720, n_721);
  nand g2000 (n_2100, n_722, n_721);
  nand g2001 (n_2101, n_720, n_722);
  nand g2002 (n_739, n_2099, n_2100, n_2101);
  xor g2003 (n_2102, n_723, n_724);
  xor g2004 (n_727, n_2102, n_725);
  nand g2005 (n_2103, n_723, n_724);
  nand g2006 (n_2104, n_725, n_724);
  nand g2007 (n_2105, n_723, n_725);
  nand g2008 (n_742, n_2103, n_2104, n_2105);
  xor g2009 (n_2106, n_726, n_727);
  xor g2010 (n_172, n_2106, n_728);
  nand g2011 (n_2107, n_726, n_727);
  nand g2012 (n_2108, n_728, n_727);
  nand g2013 (n_2109, n_726, n_728);
  nand g2014 (n_93, n_2107, n_2108, n_2109);
  xor g2015 (n_2110, A[44], A[42]);
  xor g2016 (n_733, n_2110, A[38]);
  nand g2017 (n_2111, A[44], A[42]);
  nand g2018 (n_2112, A[38], A[42]);
  nand g2019 (n_2113, A[44], A[38]);
  nand g2020 (n_743, n_2111, n_2112, n_2113);
  xor g2022 (n_734, n_1662, A[36]);
  nand g2024 (n_2116, A[36], A[28]);
  nand g2026 (n_744, n_1663, n_2116, n_1857);
  xor g2027 (n_2118, A[26], A[40]);
  xor g2028 (n_732, n_2118, A[34]);
  nand g2029 (n_2119, A[26], A[40]);
  nand g2032 (n_745, n_2119, n_1985, n_2052);
  xor g2033 (n_2122, A[32], n_729);
  xor g2034 (n_736, n_2122, n_730);
  nand g2035 (n_2123, A[32], n_729);
  nand g2036 (n_2124, n_730, n_729);
  nand g2037 (n_2125, A[32], n_730);
  nand g2038 (n_749, n_2123, n_2124, n_2125);
  xor g2039 (n_2126, n_731, n_732);
  xor g2040 (n_738, n_2126, n_733);
  nand g2041 (n_2127, n_731, n_732);
  nand g2042 (n_2128, n_733, n_732);
  nand g2043 (n_2129, n_731, n_733);
  nand g2044 (n_751, n_2127, n_2128, n_2129);
  xor g2045 (n_2130, n_734, n_735);
  xor g2046 (n_740, n_2130, n_736);
  nand g2047 (n_2131, n_734, n_735);
  nand g2048 (n_2132, n_736, n_735);
  nand g2049 (n_2133, n_734, n_736);
  nand g2050 (n_753, n_2131, n_2132, n_2133);
  xor g2051 (n_2134, n_737, n_738);
  xor g2052 (n_741, n_2134, n_739);
  nand g2053 (n_2135, n_737, n_738);
  nand g2054 (n_2136, n_739, n_738);
  nand g2055 (n_2137, n_737, n_739);
  nand g2056 (n_756, n_2135, n_2136, n_2137);
  xor g2057 (n_2138, n_740, n_741);
  xor g2058 (n_171, n_2138, n_742);
  nand g2059 (n_2139, n_740, n_741);
  nand g2060 (n_2140, n_742, n_741);
  nand g2061 (n_2141, n_740, n_742);
  nand g2062 (n_92, n_2139, n_2140, n_2141);
  xor g2063 (n_2142, A[45], A[43]);
  xor g2064 (n_747, n_2142, A[39]);
  nand g2065 (n_2143, A[45], A[43]);
  nand g2066 (n_2144, A[39], A[43]);
  nand g2067 (n_2145, A[45], A[39]);
  nand g2068 (n_757, n_2143, n_2144, n_2145);
  xor g2070 (n_748, n_1694, A[37]);
  nand g2072 (n_2148, A[37], A[29]);
  nand g2074 (n_758, n_1695, n_2148, n_1889);
  xor g2075 (n_2150, A[27], A[41]);
  xor g2076 (n_746, n_2150, A[35]);
  nand g2077 (n_2151, A[27], A[41]);
  nand g2080 (n_759, n_2151, n_2017, n_2084);
  xor g2081 (n_2154, A[33], n_743);
  xor g2082 (n_750, n_2154, n_744);
  nand g2083 (n_2155, A[33], n_743);
  nand g2084 (n_2156, n_744, n_743);
  nand g2085 (n_2157, A[33], n_744);
  nand g2086 (n_763, n_2155, n_2156, n_2157);
  xor g2087 (n_2158, n_745, n_746);
  xor g2088 (n_752, n_2158, n_747);
  nand g2089 (n_2159, n_745, n_746);
  nand g2090 (n_2160, n_747, n_746);
  nand g2091 (n_2161, n_745, n_747);
  nand g2092 (n_765, n_2159, n_2160, n_2161);
  xor g2093 (n_2162, n_748, n_749);
  xor g2094 (n_754, n_2162, n_750);
  nand g2095 (n_2163, n_748, n_749);
  nand g2096 (n_2164, n_750, n_749);
  nand g2097 (n_2165, n_748, n_750);
  nand g2098 (n_767, n_2163, n_2164, n_2165);
  xor g2099 (n_2166, n_751, n_752);
  xor g2100 (n_755, n_2166, n_753);
  nand g2101 (n_2167, n_751, n_752);
  nand g2102 (n_2168, n_753, n_752);
  nand g2103 (n_2169, n_751, n_753);
  nand g2104 (n_770, n_2167, n_2168, n_2169);
  xor g2105 (n_2170, n_754, n_755);
  xor g2106 (n_170, n_2170, n_756);
  nand g2107 (n_2171, n_754, n_755);
  nand g2108 (n_2172, n_756, n_755);
  nand g2109 (n_2173, n_754, n_756);
  nand g2110 (n_91, n_2171, n_2172, n_2173);
  xor g2111 (n_2174, A[46], A[44]);
  xor g2112 (n_761, n_2174, A[40]);
  nand g2113 (n_2175, A[46], A[44]);
  nand g2114 (n_2176, A[40], A[44]);
  nand g2115 (n_2177, A[46], A[40]);
  nand g2116 (n_771, n_2175, n_2176, n_2177);
  xor g2118 (n_762, n_1726, A[38]);
  nand g2120 (n_2180, A[38], A[30]);
  nand g2122 (n_772, n_1727, n_2180, n_1921);
  xor g2123 (n_2182, A[28], A[42]);
  xor g2124 (n_760, n_2182, A[36]);
  nand g2125 (n_2183, A[28], A[42]);
  nand g2128 (n_773, n_2183, n_2049, n_2116);
  xor g2129 (n_2186, A[34], n_757);
  xor g2130 (n_764, n_2186, n_758);
  nand g2131 (n_2187, A[34], n_757);
  nand g2132 (n_2188, n_758, n_757);
  nand g2133 (n_2189, A[34], n_758);
  nand g2134 (n_777, n_2187, n_2188, n_2189);
  xor g2135 (n_2190, n_759, n_760);
  xor g2136 (n_766, n_2190, n_761);
  nand g2137 (n_2191, n_759, n_760);
  nand g2138 (n_2192, n_761, n_760);
  nand g2139 (n_2193, n_759, n_761);
  nand g2140 (n_779, n_2191, n_2192, n_2193);
  xor g2141 (n_2194, n_762, n_763);
  xor g2142 (n_768, n_2194, n_764);
  nand g2143 (n_2195, n_762, n_763);
  nand g2144 (n_2196, n_764, n_763);
  nand g2145 (n_2197, n_762, n_764);
  nand g2146 (n_781, n_2195, n_2196, n_2197);
  xor g2147 (n_2198, n_765, n_766);
  xor g2148 (n_769, n_2198, n_767);
  nand g2149 (n_2199, n_765, n_766);
  nand g2150 (n_2200, n_767, n_766);
  nand g2151 (n_2201, n_765, n_767);
  nand g2152 (n_784, n_2199, n_2200, n_2201);
  xor g2153 (n_2202, n_768, n_769);
  xor g2154 (n_169, n_2202, n_770);
  nand g2155 (n_2203, n_768, n_769);
  nand g2156 (n_2204, n_770, n_769);
  nand g2157 (n_2205, n_768, n_770);
  nand g2158 (n_90, n_2203, n_2204, n_2205);
  xor g2159 (n_2206, A[47], A[45]);
  xor g2160 (n_775, n_2206, A[41]);
  nand g2161 (n_2207, A[47], A[45]);
  nand g2162 (n_2208, A[41], A[45]);
  nand g2163 (n_2209, A[47], A[41]);
  nand g2164 (n_785, n_2207, n_2208, n_2209);
  xor g2166 (n_776, n_1758, A[39]);
  nand g2168 (n_2212, A[39], A[31]);
  nand g2170 (n_786, n_1759, n_2212, n_1953);
  xor g2171 (n_2214, A[29], A[43]);
  xor g2172 (n_774, n_2214, A[37]);
  nand g2173 (n_2215, A[29], A[43]);
  nand g2176 (n_787, n_2215, n_2081, n_2148);
  xor g2177 (n_2218, A[35], n_771);
  xor g2178 (n_778, n_2218, n_772);
  nand g2179 (n_2219, A[35], n_771);
  nand g2180 (n_2220, n_772, n_771);
  nand g2181 (n_2221, A[35], n_772);
  nand g2182 (n_791, n_2219, n_2220, n_2221);
  xor g2183 (n_2222, n_773, n_774);
  xor g2184 (n_780, n_2222, n_775);
  nand g2185 (n_2223, n_773, n_774);
  nand g2186 (n_2224, n_775, n_774);
  nand g2187 (n_2225, n_773, n_775);
  nand g2188 (n_793, n_2223, n_2224, n_2225);
  xor g2189 (n_2226, n_776, n_777);
  xor g2190 (n_782, n_2226, n_778);
  nand g2191 (n_2227, n_776, n_777);
  nand g2192 (n_2228, n_778, n_777);
  nand g2193 (n_2229, n_776, n_778);
  nand g2194 (n_795, n_2227, n_2228, n_2229);
  xor g2195 (n_2230, n_779, n_780);
  xor g2196 (n_783, n_2230, n_781);
  nand g2197 (n_2231, n_779, n_780);
  nand g2198 (n_2232, n_781, n_780);
  nand g2199 (n_2233, n_779, n_781);
  nand g2200 (n_798, n_2231, n_2232, n_2233);
  xor g2201 (n_2234, n_782, n_783);
  xor g2202 (n_168, n_2234, n_784);
  nand g2203 (n_2235, n_782, n_783);
  nand g2204 (n_2236, n_784, n_783);
  nand g2205 (n_2237, n_782, n_784);
  nand g2206 (n_89, n_2235, n_2236, n_2237);
  xor g2207 (n_2238, A[48], A[46]);
  xor g2208 (n_789, n_2238, A[42]);
  nand g2209 (n_2239, A[48], A[46]);
  nand g2210 (n_2240, A[42], A[46]);
  nand g2211 (n_2241, A[48], A[42]);
  nand g2212 (n_799, n_2239, n_2240, n_2241);
  xor g2214 (n_790, n_1790, A[40]);
  nand g2216 (n_2244, A[40], A[32]);
  nand g2218 (n_800, n_1791, n_2244, n_1985);
  xor g2219 (n_2246, A[30], A[44]);
  xor g2220 (n_788, n_2246, A[38]);
  nand g2221 (n_2247, A[30], A[44]);
  nand g2224 (n_801, n_2247, n_2113, n_2180);
  xor g2225 (n_2250, A[36], n_785);
  xor g2226 (n_792, n_2250, n_786);
  nand g2227 (n_2251, A[36], n_785);
  nand g2228 (n_2252, n_786, n_785);
  nand g2229 (n_2253, A[36], n_786);
  nand g2230 (n_805, n_2251, n_2252, n_2253);
  xor g2231 (n_2254, n_787, n_788);
  xor g2232 (n_794, n_2254, n_789);
  nand g2233 (n_2255, n_787, n_788);
  nand g2234 (n_2256, n_789, n_788);
  nand g2235 (n_2257, n_787, n_789);
  nand g2236 (n_807, n_2255, n_2256, n_2257);
  xor g2237 (n_2258, n_790, n_791);
  xor g2238 (n_796, n_2258, n_792);
  nand g2239 (n_2259, n_790, n_791);
  nand g2240 (n_2260, n_792, n_791);
  nand g2241 (n_2261, n_790, n_792);
  nand g2242 (n_809, n_2259, n_2260, n_2261);
  xor g2243 (n_2262, n_793, n_794);
  xor g2244 (n_797, n_2262, n_795);
  nand g2245 (n_2263, n_793, n_794);
  nand g2246 (n_2264, n_795, n_794);
  nand g2247 (n_2265, n_793, n_795);
  nand g2248 (n_812, n_2263, n_2264, n_2265);
  xor g2249 (n_2266, n_796, n_797);
  xor g2250 (n_167, n_2266, n_798);
  nand g2251 (n_2267, n_796, n_797);
  nand g2252 (n_2268, n_798, n_797);
  nand g2253 (n_2269, n_796, n_798);
  nand g2254 (n_88, n_2267, n_2268, n_2269);
  xor g2255 (n_2270, A[49], A[47]);
  xor g2256 (n_803, n_2270, A[43]);
  nand g2257 (n_2271, A[49], A[47]);
  nand g2258 (n_2272, A[43], A[47]);
  nand g2259 (n_2273, A[49], A[43]);
  nand g2260 (n_813, n_2271, n_2272, n_2273);
  xor g2262 (n_804, n_1822, A[41]);
  nand g2264 (n_2276, A[41], A[33]);
  nand g2266 (n_814, n_1823, n_2276, n_2017);
  xor g2267 (n_2278, A[31], A[45]);
  xor g2268 (n_802, n_2278, A[39]);
  nand g2269 (n_2279, A[31], A[45]);
  nand g2272 (n_815, n_2279, n_2145, n_2212);
  xor g2273 (n_2282, A[37], n_799);
  xor g2274 (n_806, n_2282, n_800);
  nand g2275 (n_2283, A[37], n_799);
  nand g2276 (n_2284, n_800, n_799);
  nand g2277 (n_2285, A[37], n_800);
  nand g2278 (n_819, n_2283, n_2284, n_2285);
  xor g2279 (n_2286, n_801, n_802);
  xor g2280 (n_808, n_2286, n_803);
  nand g2281 (n_2287, n_801, n_802);
  nand g2282 (n_2288, n_803, n_802);
  nand g2283 (n_2289, n_801, n_803);
  nand g2284 (n_821, n_2287, n_2288, n_2289);
  xor g2285 (n_2290, n_804, n_805);
  xor g2286 (n_810, n_2290, n_806);
  nand g2287 (n_2291, n_804, n_805);
  nand g2288 (n_2292, n_806, n_805);
  nand g2289 (n_2293, n_804, n_806);
  nand g2290 (n_823, n_2291, n_2292, n_2293);
  xor g2291 (n_2294, n_807, n_808);
  xor g2292 (n_811, n_2294, n_809);
  nand g2293 (n_2295, n_807, n_808);
  nand g2294 (n_2296, n_809, n_808);
  nand g2295 (n_2297, n_807, n_809);
  nand g2296 (n_826, n_2295, n_2296, n_2297);
  xor g2297 (n_2298, n_810, n_811);
  xor g2298 (n_166, n_2298, n_812);
  nand g2299 (n_2299, n_810, n_811);
  nand g2300 (n_2300, n_812, n_811);
  nand g2301 (n_2301, n_810, n_812);
  nand g2302 (n_87, n_2299, n_2300, n_2301);
  xor g2303 (n_2302, A[50], A[48]);
  xor g2304 (n_817, n_2302, A[44]);
  nand g2305 (n_2303, A[50], A[48]);
  nand g2306 (n_2304, A[44], A[48]);
  nand g2307 (n_2305, A[50], A[44]);
  nand g2308 (n_827, n_2303, n_2304, n_2305);
  xor g2310 (n_818, n_1854, A[42]);
  nand g2312 (n_2308, A[42], A[34]);
  nand g2314 (n_828, n_1855, n_2308, n_2049);
  xor g2315 (n_2310, A[32], A[46]);
  xor g2316 (n_816, n_2310, A[40]);
  nand g2317 (n_2311, A[32], A[46]);
  nand g2320 (n_829, n_2311, n_2177, n_2244);
  xor g2321 (n_2314, A[38], n_813);
  xor g2322 (n_820, n_2314, n_814);
  nand g2323 (n_2315, A[38], n_813);
  nand g2324 (n_2316, n_814, n_813);
  nand g2325 (n_2317, A[38], n_814);
  nand g2326 (n_833, n_2315, n_2316, n_2317);
  xor g2327 (n_2318, n_815, n_816);
  xor g2328 (n_822, n_2318, n_817);
  nand g2329 (n_2319, n_815, n_816);
  nand g2330 (n_2320, n_817, n_816);
  nand g2331 (n_2321, n_815, n_817);
  nand g2332 (n_835, n_2319, n_2320, n_2321);
  xor g2333 (n_2322, n_818, n_819);
  xor g2334 (n_824, n_2322, n_820);
  nand g2335 (n_2323, n_818, n_819);
  nand g2336 (n_2324, n_820, n_819);
  nand g2337 (n_2325, n_818, n_820);
  nand g2338 (n_837, n_2323, n_2324, n_2325);
  xor g2339 (n_2326, n_821, n_822);
  xor g2340 (n_825, n_2326, n_823);
  nand g2341 (n_2327, n_821, n_822);
  nand g2342 (n_2328, n_823, n_822);
  nand g2343 (n_2329, n_821, n_823);
  nand g2344 (n_840, n_2327, n_2328, n_2329);
  xor g2345 (n_2330, n_824, n_825);
  xor g2346 (n_165, n_2330, n_826);
  nand g2347 (n_2331, n_824, n_825);
  nand g2348 (n_2332, n_826, n_825);
  nand g2349 (n_2333, n_824, n_826);
  nand g2350 (n_86, n_2331, n_2332, n_2333);
  xor g2351 (n_2334, A[51], A[49]);
  xor g2352 (n_831, n_2334, A[45]);
  nand g2353 (n_2335, A[51], A[49]);
  nand g2354 (n_2336, A[45], A[49]);
  nand g2355 (n_2337, A[51], A[45]);
  nand g2356 (n_841, n_2335, n_2336, n_2337);
  xor g2358 (n_832, n_1886, A[43]);
  nand g2360 (n_2340, A[43], A[35]);
  nand g2362 (n_842, n_1887, n_2340, n_2081);
  xor g2363 (n_2342, A[33], A[47]);
  xor g2364 (n_830, n_2342, A[41]);
  nand g2365 (n_2343, A[33], A[47]);
  nand g2368 (n_843, n_2343, n_2209, n_2276);
  xor g2369 (n_2346, A[39], n_827);
  xor g2370 (n_834, n_2346, n_828);
  nand g2371 (n_2347, A[39], n_827);
  nand g2372 (n_2348, n_828, n_827);
  nand g2373 (n_2349, A[39], n_828);
  nand g2374 (n_847, n_2347, n_2348, n_2349);
  xor g2375 (n_2350, n_829, n_830);
  xor g2376 (n_836, n_2350, n_831);
  nand g2377 (n_2351, n_829, n_830);
  nand g2378 (n_2352, n_831, n_830);
  nand g2379 (n_2353, n_829, n_831);
  nand g2380 (n_849, n_2351, n_2352, n_2353);
  xor g2381 (n_2354, n_832, n_833);
  xor g2382 (n_838, n_2354, n_834);
  nand g2383 (n_2355, n_832, n_833);
  nand g2384 (n_2356, n_834, n_833);
  nand g2385 (n_2357, n_832, n_834);
  nand g2386 (n_851, n_2355, n_2356, n_2357);
  xor g2387 (n_2358, n_835, n_836);
  xor g2388 (n_839, n_2358, n_837);
  nand g2389 (n_2359, n_835, n_836);
  nand g2390 (n_2360, n_837, n_836);
  nand g2391 (n_2361, n_835, n_837);
  nand g2392 (n_854, n_2359, n_2360, n_2361);
  xor g2393 (n_2362, n_838, n_839);
  xor g2394 (n_164, n_2362, n_840);
  nand g2395 (n_2363, n_838, n_839);
  nand g2396 (n_2364, n_840, n_839);
  nand g2397 (n_2365, n_838, n_840);
  nand g2398 (n_85, n_2363, n_2364, n_2365);
  xor g2399 (n_2366, A[52], A[50]);
  xor g2400 (n_845, n_2366, A[46]);
  nand g2401 (n_2367, A[52], A[50]);
  nand g2402 (n_2368, A[46], A[50]);
  nand g2403 (n_2369, A[52], A[46]);
  nand g2404 (n_855, n_2367, n_2368, n_2369);
  xor g2406 (n_846, n_1918, A[44]);
  nand g2408 (n_2372, A[44], A[36]);
  nand g2410 (n_856, n_1919, n_2372, n_2113);
  xor g2411 (n_2374, A[34], A[48]);
  xor g2412 (n_844, n_2374, A[42]);
  nand g2413 (n_2375, A[34], A[48]);
  nand g2416 (n_857, n_2375, n_2241, n_2308);
  xor g2417 (n_2378, A[40], n_841);
  xor g2418 (n_848, n_2378, n_842);
  nand g2419 (n_2379, A[40], n_841);
  nand g2420 (n_2380, n_842, n_841);
  nand g2421 (n_2381, A[40], n_842);
  nand g2422 (n_861, n_2379, n_2380, n_2381);
  xor g2423 (n_2382, n_843, n_844);
  xor g2424 (n_850, n_2382, n_845);
  nand g2425 (n_2383, n_843, n_844);
  nand g2426 (n_2384, n_845, n_844);
  nand g2427 (n_2385, n_843, n_845);
  nand g2428 (n_863, n_2383, n_2384, n_2385);
  xor g2429 (n_2386, n_846, n_847);
  xor g2430 (n_852, n_2386, n_848);
  nand g2431 (n_2387, n_846, n_847);
  nand g2432 (n_2388, n_848, n_847);
  nand g2433 (n_2389, n_846, n_848);
  nand g2434 (n_865, n_2387, n_2388, n_2389);
  xor g2435 (n_2390, n_849, n_850);
  xor g2436 (n_853, n_2390, n_851);
  nand g2437 (n_2391, n_849, n_850);
  nand g2438 (n_2392, n_851, n_850);
  nand g2439 (n_2393, n_849, n_851);
  nand g2440 (n_868, n_2391, n_2392, n_2393);
  xor g2441 (n_2394, n_852, n_853);
  xor g2442 (n_163, n_2394, n_854);
  nand g2443 (n_2395, n_852, n_853);
  nand g2444 (n_2396, n_854, n_853);
  nand g2445 (n_2397, n_852, n_854);
  nand g2446 (n_84, n_2395, n_2396, n_2397);
  xor g2447 (n_2398, A[53], A[51]);
  xor g2448 (n_859, n_2398, A[47]);
  nand g2449 (n_2399, A[53], A[51]);
  nand g2450 (n_2400, A[47], A[51]);
  nand g2451 (n_2401, A[53], A[47]);
  nand g2452 (n_869, n_2399, n_2400, n_2401);
  xor g2454 (n_860, n_1950, A[45]);
  nand g2456 (n_2404, A[45], A[37]);
  nand g2458 (n_870, n_1951, n_2404, n_2145);
  xor g2459 (n_2406, A[35], A[49]);
  xor g2460 (n_858, n_2406, A[43]);
  nand g2461 (n_2407, A[35], A[49]);
  nand g2464 (n_871, n_2407, n_2273, n_2340);
  xor g2465 (n_2410, A[41], n_855);
  xor g2466 (n_862, n_2410, n_856);
  nand g2467 (n_2411, A[41], n_855);
  nand g2468 (n_2412, n_856, n_855);
  nand g2469 (n_2413, A[41], n_856);
  nand g2470 (n_875, n_2411, n_2412, n_2413);
  xor g2471 (n_2414, n_857, n_858);
  xor g2472 (n_864, n_2414, n_859);
  nand g2473 (n_2415, n_857, n_858);
  nand g2474 (n_2416, n_859, n_858);
  nand g2475 (n_2417, n_857, n_859);
  nand g2476 (n_877, n_2415, n_2416, n_2417);
  xor g2477 (n_2418, n_860, n_861);
  xor g2478 (n_866, n_2418, n_862);
  nand g2479 (n_2419, n_860, n_861);
  nand g2480 (n_2420, n_862, n_861);
  nand g2481 (n_2421, n_860, n_862);
  nand g2482 (n_879, n_2419, n_2420, n_2421);
  xor g2483 (n_2422, n_863, n_864);
  xor g2484 (n_867, n_2422, n_865);
  nand g2485 (n_2423, n_863, n_864);
  nand g2486 (n_2424, n_865, n_864);
  nand g2487 (n_2425, n_863, n_865);
  nand g2488 (n_882, n_2423, n_2424, n_2425);
  xor g2489 (n_2426, n_866, n_867);
  xor g2490 (n_162, n_2426, n_868);
  nand g2491 (n_2427, n_866, n_867);
  nand g2492 (n_2428, n_868, n_867);
  nand g2493 (n_2429, n_866, n_868);
  nand g2494 (n_83, n_2427, n_2428, n_2429);
  xor g2495 (n_2430, A[54], A[52]);
  xor g2496 (n_873, n_2430, A[48]);
  nand g2497 (n_2431, A[54], A[52]);
  nand g2498 (n_2432, A[48], A[52]);
  nand g2499 (n_2433, A[54], A[48]);
  nand g2500 (n_883, n_2431, n_2432, n_2433);
  xor g2502 (n_874, n_1982, A[46]);
  nand g2504 (n_2436, A[46], A[38]);
  nand g2506 (n_884, n_1983, n_2436, n_2177);
  xor g2507 (n_2438, A[36], A[50]);
  xor g2508 (n_872, n_2438, A[44]);
  nand g2509 (n_2439, A[36], A[50]);
  nand g2512 (n_885, n_2439, n_2305, n_2372);
  xor g2513 (n_2442, A[42], n_869);
  xor g2514 (n_876, n_2442, n_870);
  nand g2515 (n_2443, A[42], n_869);
  nand g2516 (n_2444, n_870, n_869);
  nand g2517 (n_2445, A[42], n_870);
  nand g2518 (n_889, n_2443, n_2444, n_2445);
  xor g2519 (n_2446, n_871, n_872);
  xor g2520 (n_878, n_2446, n_873);
  nand g2521 (n_2447, n_871, n_872);
  nand g2522 (n_2448, n_873, n_872);
  nand g2523 (n_2449, n_871, n_873);
  nand g2524 (n_891, n_2447, n_2448, n_2449);
  xor g2525 (n_2450, n_874, n_875);
  xor g2526 (n_880, n_2450, n_876);
  nand g2527 (n_2451, n_874, n_875);
  nand g2528 (n_2452, n_876, n_875);
  nand g2529 (n_2453, n_874, n_876);
  nand g2530 (n_893, n_2451, n_2452, n_2453);
  xor g2531 (n_2454, n_877, n_878);
  xor g2532 (n_881, n_2454, n_879);
  nand g2533 (n_2455, n_877, n_878);
  nand g2534 (n_2456, n_879, n_878);
  nand g2535 (n_2457, n_877, n_879);
  nand g2536 (n_896, n_2455, n_2456, n_2457);
  xor g2537 (n_2458, n_880, n_881);
  xor g2538 (n_161, n_2458, n_882);
  nand g2539 (n_2459, n_880, n_881);
  nand g2540 (n_2460, n_882, n_881);
  nand g2541 (n_2461, n_880, n_882);
  nand g2542 (n_82, n_2459, n_2460, n_2461);
  xor g2543 (n_2462, A[55], A[53]);
  xor g2544 (n_887, n_2462, A[49]);
  nand g2545 (n_2463, A[55], A[53]);
  nand g2546 (n_2464, A[49], A[53]);
  nand g2547 (n_2465, A[55], A[49]);
  nand g2548 (n_897, n_2463, n_2464, n_2465);
  xor g2550 (n_888, n_2014, A[47]);
  nand g2552 (n_2468, A[47], A[39]);
  nand g2554 (n_898, n_2015, n_2468, n_2209);
  xor g2555 (n_2470, A[37], A[51]);
  xor g2556 (n_886, n_2470, A[45]);
  nand g2557 (n_2471, A[37], A[51]);
  nand g2560 (n_899, n_2471, n_2337, n_2404);
  xor g2561 (n_2474, A[43], n_883);
  xor g2562 (n_890, n_2474, n_884);
  nand g2563 (n_2475, A[43], n_883);
  nand g2564 (n_2476, n_884, n_883);
  nand g2565 (n_2477, A[43], n_884);
  nand g2566 (n_903, n_2475, n_2476, n_2477);
  xor g2567 (n_2478, n_885, n_886);
  xor g2568 (n_892, n_2478, n_887);
  nand g2569 (n_2479, n_885, n_886);
  nand g2570 (n_2480, n_887, n_886);
  nand g2571 (n_2481, n_885, n_887);
  nand g2572 (n_905, n_2479, n_2480, n_2481);
  xor g2573 (n_2482, n_888, n_889);
  xor g2574 (n_894, n_2482, n_890);
  nand g2575 (n_2483, n_888, n_889);
  nand g2576 (n_2484, n_890, n_889);
  nand g2577 (n_2485, n_888, n_890);
  nand g2578 (n_907, n_2483, n_2484, n_2485);
  xor g2579 (n_2486, n_891, n_892);
  xor g2580 (n_895, n_2486, n_893);
  nand g2581 (n_2487, n_891, n_892);
  nand g2582 (n_2488, n_893, n_892);
  nand g2583 (n_2489, n_891, n_893);
  nand g2584 (n_910, n_2487, n_2488, n_2489);
  xor g2585 (n_2490, n_894, n_895);
  xor g2586 (n_160, n_2490, n_896);
  nand g2587 (n_2491, n_894, n_895);
  nand g2588 (n_2492, n_896, n_895);
  nand g2589 (n_2493, n_894, n_896);
  nand g2590 (n_81, n_2491, n_2492, n_2493);
  xor g2591 (n_2494, A[56], A[54]);
  xor g2592 (n_901, n_2494, A[50]);
  nand g2593 (n_2495, A[56], A[54]);
  nand g2594 (n_2496, A[50], A[54]);
  nand g2595 (n_2497, A[56], A[50]);
  nand g2596 (n_911, n_2495, n_2496, n_2497);
  xor g2598 (n_902, n_2046, A[48]);
  nand g2600 (n_2500, A[48], A[40]);
  nand g2602 (n_912, n_2047, n_2500, n_2241);
  xor g2603 (n_2502, A[38], A[52]);
  xor g2604 (n_900, n_2502, A[46]);
  nand g2605 (n_2503, A[38], A[52]);
  nand g2608 (n_913, n_2503, n_2369, n_2436);
  xor g2609 (n_2506, A[44], n_897);
  xor g2610 (n_904, n_2506, n_898);
  nand g2611 (n_2507, A[44], n_897);
  nand g2612 (n_2508, n_898, n_897);
  nand g2613 (n_2509, A[44], n_898);
  nand g2614 (n_917, n_2507, n_2508, n_2509);
  xor g2615 (n_2510, n_899, n_900);
  xor g2616 (n_906, n_2510, n_901);
  nand g2617 (n_2511, n_899, n_900);
  nand g2618 (n_2512, n_901, n_900);
  nand g2619 (n_2513, n_899, n_901);
  nand g2620 (n_919, n_2511, n_2512, n_2513);
  xor g2621 (n_2514, n_902, n_903);
  xor g2622 (n_908, n_2514, n_904);
  nand g2623 (n_2515, n_902, n_903);
  nand g2624 (n_2516, n_904, n_903);
  nand g2625 (n_2517, n_902, n_904);
  nand g2626 (n_921, n_2515, n_2516, n_2517);
  xor g2627 (n_2518, n_905, n_906);
  xor g2628 (n_909, n_2518, n_907);
  nand g2629 (n_2519, n_905, n_906);
  nand g2630 (n_2520, n_907, n_906);
  nand g2631 (n_2521, n_905, n_907);
  nand g2632 (n_924, n_2519, n_2520, n_2521);
  xor g2633 (n_2522, n_908, n_909);
  xor g2634 (n_159, n_2522, n_910);
  nand g2635 (n_2523, n_908, n_909);
  nand g2636 (n_2524, n_910, n_909);
  nand g2637 (n_2525, n_908, n_910);
  nand g2638 (n_80, n_2523, n_2524, n_2525);
  xor g2639 (n_2526, A[57], A[55]);
  xor g2640 (n_915, n_2526, A[51]);
  nand g2641 (n_2527, A[57], A[55]);
  nand g2642 (n_2528, A[51], A[55]);
  nand g2643 (n_2529, A[57], A[51]);
  nand g2644 (n_928, n_2527, n_2528, n_2529);
  xor g2646 (n_916, n_2078, A[49]);
  nand g2648 (n_2532, A[49], A[41]);
  nand g2650 (n_929, n_2079, n_2532, n_2273);
  xor g2651 (n_2534, A[39], A[53]);
  xor g2652 (n_914, n_2534, A[47]);
  nand g2653 (n_2535, A[39], A[53]);
  nand g2656 (n_927, n_2535, n_2401, n_2468);
  xor g2657 (n_2538, A[45], n_911);
  xor g2658 (n_918, n_2538, n_912);
  nand g2659 (n_2539, A[45], n_911);
  nand g2660 (n_2540, n_912, n_911);
  nand g2661 (n_2541, A[45], n_912);
  nand g2662 (n_933, n_2539, n_2540, n_2541);
  xor g2663 (n_2542, n_913, n_914);
  xor g2664 (n_920, n_2542, n_915);
  nand g2665 (n_2543, n_913, n_914);
  nand g2666 (n_2544, n_915, n_914);
  nand g2667 (n_2545, n_913, n_915);
  nand g2668 (n_935, n_2543, n_2544, n_2545);
  xor g2669 (n_2546, n_916, n_917);
  xor g2670 (n_922, n_2546, n_918);
  nand g2671 (n_2547, n_916, n_917);
  nand g2672 (n_2548, n_918, n_917);
  nand g2673 (n_2549, n_916, n_918);
  nand g2674 (n_937, n_2547, n_2548, n_2549);
  xor g2675 (n_2550, n_919, n_920);
  xor g2676 (n_923, n_2550, n_921);
  nand g2677 (n_2551, n_919, n_920);
  nand g2678 (n_2552, n_921, n_920);
  nand g2679 (n_2553, n_919, n_921);
  nand g2680 (n_940, n_2551, n_2552, n_2553);
  xor g2681 (n_2554, n_922, n_923);
  xor g2682 (n_158, n_2554, n_924);
  nand g2683 (n_2555, n_922, n_923);
  nand g2684 (n_2556, n_924, n_923);
  nand g2685 (n_2557, n_922, n_924);
  nand g2686 (n_79, n_2555, n_2556, n_2557);
  xor g2689 (n_2558, A[58], A[52]);
  xor g2690 (n_931, n_2558, A[44]);
  nand g2691 (n_2559, A[58], A[52]);
  nand g2692 (n_2560, A[44], A[52]);
  nand g2693 (n_2561, A[58], A[44]);
  nand g2694 (n_944, n_2559, n_2560, n_2561);
  xor g2695 (n_2562, A[42], A[56]);
  xor g2696 (n_932, n_2562, A[40]);
  nand g2697 (n_2563, A[42], A[56]);
  nand g2698 (n_2564, A[40], A[56]);
  nand g2700 (n_945, n_2563, n_2564, n_2047);
  xor g2701 (n_2566, A[50], A[54]);
  xor g2702 (n_930, n_2566, A[48]);
  nand g2706 (n_946, n_2496, n_2433, n_2303);
  xor g2707 (n_2570, A[46], n_927);
  xor g2708 (n_934, n_2570, n_928);
  nand g2709 (n_2571, A[46], n_927);
  nand g2710 (n_2572, n_928, n_927);
  nand g2711 (n_2573, A[46], n_928);
  nand g2712 (n_950, n_2571, n_2572, n_2573);
  xor g2713 (n_2574, n_929, n_930);
  xor g2714 (n_936, n_2574, n_931);
  nand g2715 (n_2575, n_929, n_930);
  nand g2716 (n_2576, n_931, n_930);
  nand g2717 (n_2577, n_929, n_931);
  nand g2718 (n_952, n_2575, n_2576, n_2577);
  xor g2719 (n_2578, n_932, n_933);
  xor g2720 (n_938, n_2578, n_934);
  nand g2721 (n_2579, n_932, n_933);
  nand g2722 (n_2580, n_934, n_933);
  nand g2723 (n_2581, n_932, n_934);
  nand g2724 (n_955, n_2579, n_2580, n_2581);
  xor g2725 (n_2582, n_935, n_936);
  xor g2726 (n_939, n_2582, n_937);
  nand g2727 (n_2583, n_935, n_936);
  nand g2728 (n_2584, n_937, n_936);
  nand g2729 (n_2585, n_935, n_937);
  nand g2730 (n_957, n_2583, n_2584, n_2585);
  xor g2731 (n_2586, n_938, n_939);
  xor g2732 (n_157, n_2586, n_940);
  nand g2733 (n_2587, n_938, n_939);
  nand g2734 (n_2588, n_940, n_939);
  nand g2735 (n_2589, n_938, n_940);
  nand g2736 (n_78, n_2587, n_2588, n_2589);
  xor g2739 (n_2590, A[51], A[43]);
  xor g2740 (n_948, n_2590, A[41]);
  nand g2741 (n_2591, A[51], A[43]);
  nand g2743 (n_2593, A[51], A[41]);
  nand g2744 (n_959, n_2591, n_2079, n_2593);
  xor g2745 (n_2594, A[57], A[49]);
  xor g2746 (n_949, n_2594, A[55]);
  nand g2747 (n_2595, A[57], A[49]);
  nand g2750 (n_961, n_2595, n_2465, n_2527);
  xor g2751 (n_2598, A[53], A[47]);
  xor g2752 (n_947, n_2598, A[45]);
  nand g2755 (n_2601, A[53], A[45]);
  nand g2756 (n_960, n_2401, n_2207, n_2601);
  xor g2757 (n_2602, A[58], n_944);
  xor g2758 (n_951, n_2602, n_945);
  nand g2759 (n_2603, A[58], n_944);
  nand g2760 (n_2604, n_945, n_944);
  nand g2761 (n_2605, A[58], n_945);
  nand g2762 (n_965, n_2603, n_2604, n_2605);
  xor g2763 (n_2606, n_946, n_947);
  xor g2764 (n_953, n_2606, n_948);
  nand g2765 (n_2607, n_946, n_947);
  nand g2766 (n_2608, n_948, n_947);
  nand g2767 (n_2609, n_946, n_948);
  nand g2768 (n_967, n_2607, n_2608, n_2609);
  xor g2769 (n_2610, n_949, n_950);
  xor g2770 (n_954, n_2610, n_951);
  nand g2771 (n_2611, n_949, n_950);
  nand g2772 (n_2612, n_951, n_950);
  nand g2773 (n_2613, n_949, n_951);
  nand g2774 (n_970, n_2611, n_2612, n_2613);
  xor g2775 (n_2614, n_952, n_953);
  xor g2776 (n_956, n_2614, n_954);
  nand g2777 (n_2615, n_952, n_953);
  nand g2778 (n_2616, n_954, n_953);
  nand g2779 (n_2617, n_952, n_954);
  nand g2780 (n_972, n_2615, n_2616, n_2617);
  xor g2781 (n_2618, n_955, n_956);
  xor g2782 (n_156, n_2618, n_957);
  nand g2783 (n_2619, n_955, n_956);
  nand g2784 (n_2620, n_957, n_956);
  nand g2785 (n_2621, n_955, n_957);
  nand g2786 (n_77, n_2619, n_2620, n_2621);
  xor g2788 (n_963, n_2622, A[52]);
  nand g2790 (n_2624, A[52], A[56]);
  nand g2792 (n_975, n_2623, n_2624, n_2625);
  xor g2794 (n_964, n_2110, A[50]);
  nand g2796 (n_2628, A[50], A[42]);
  nand g2798 (n_976, n_2111, n_2628, n_2305);
  xor g2799 (n_2630, A[54], A[48]);
  xor g2800 (n_962, n_2630, A[46]);
  nand g2803 (n_2633, A[54], A[46]);
  nand g2804 (n_977, n_2433, n_2239, n_2633);
  xor g2806 (n_966, n_2634, n_960);
  nand g2808 (n_2636, n_960, n_959);
  nand g2810 (n_981, n_2635, n_2636, n_2637);
  xor g2811 (n_2638, n_961, n_962);
  xor g2812 (n_968, n_2638, n_963);
  nand g2813 (n_2639, n_961, n_962);
  nand g2814 (n_2640, n_963, n_962);
  nand g2815 (n_2641, n_961, n_963);
  nand g2816 (n_983, n_2639, n_2640, n_2641);
  xor g2817 (n_2642, n_964, n_965);
  xor g2818 (n_969, n_2642, n_966);
  nand g2819 (n_2643, n_964, n_965);
  nand g2820 (n_2644, n_966, n_965);
  nand g2821 (n_2645, n_964, n_966);
  nand g2822 (n_985, n_2643, n_2644, n_2645);
  xor g2823 (n_2646, n_967, n_968);
  xor g2824 (n_971, n_2646, n_969);
  nand g2825 (n_2647, n_967, n_968);
  nand g2826 (n_2648, n_969, n_968);
  nand g2827 (n_2649, n_967, n_969);
  nand g2828 (n_987, n_2647, n_2648, n_2649);
  xor g2829 (n_2650, n_970, n_971);
  xor g2830 (n_155, n_2650, n_972);
  nand g2831 (n_2651, n_970, n_971);
  nand g2832 (n_2652, n_972, n_971);
  nand g2833 (n_2653, n_970, n_972);
  nand g2834 (n_76, n_2651, n_2652, n_2653);
  xor g2837 (n_2654, A[55], A[43]);
  xor g2838 (n_979, n_2654, A[51]);
  nand g2839 (n_2655, A[55], A[43]);
  nand g2842 (n_990, n_2655, n_2591, n_2528);
  xor g2843 (n_2658, A[49], A[53]);
  xor g2844 (n_978, n_2658, A[47]);
  nand g2848 (n_989, n_2464, n_2401, n_2271);
  xor g2850 (n_980, n_2662, n_975);
  nand g2853 (n_2665, A[45], n_975);
  nand g2854 (n_994, n_2663, n_2664, n_2665);
  xor g2855 (n_2666, n_976, n_977);
  xor g2856 (n_982, n_2666, n_978);
  nand g2857 (n_2667, n_976, n_977);
  nand g2858 (n_2668, n_978, n_977);
  nand g2859 (n_2669, n_976, n_978);
  nand g2860 (n_996, n_2667, n_2668, n_2669);
  xor g2861 (n_2670, n_979, n_980);
  xor g2862 (n_984, n_2670, n_981);
  nand g2863 (n_2671, n_979, n_980);
  nand g2864 (n_2672, n_981, n_980);
  nand g2865 (n_2673, n_979, n_981);
  nand g2866 (n_997, n_2671, n_2672, n_2673);
  xor g2867 (n_2674, n_982, n_983);
  xor g2868 (n_986, n_2674, n_984);
  nand g2869 (n_2675, n_982, n_983);
  nand g2870 (n_2676, n_984, n_983);
  nand g2871 (n_2677, n_982, n_984);
  nand g2872 (n_1000, n_2675, n_2676, n_2677);
  xor g2873 (n_2678, n_985, n_986);
  xor g2874 (n_154, n_2678, n_987);
  nand g2875 (n_2679, n_985, n_986);
  nand g2876 (n_2680, n_987, n_986);
  nand g2877 (n_2681, n_985, n_987);
  nand g2878 (n_75, n_2679, n_2680, n_2681);
  xor g2885 (n_2686, A[44], A[50]);
  xor g2886 (n_992, n_2686, A[54]);
  nand g2889 (n_2689, A[44], A[54]);
  nand g2890 (n_1004, n_2305, n_2496, n_2689);
  xor g2892 (n_993, n_2238, A[57]);
  nand g2894 (n_2692, A[57], A[46]);
  nand g2895 (n_2693, A[48], A[57]);
  nand g2896 (n_1007, n_2239, n_2692, n_2693);
  xor g2897 (n_2694, n_989, n_990);
  xor g2898 (n_995, n_2694, n_963);
  nand g2899 (n_2695, n_989, n_990);
  nand g2900 (n_2696, n_963, n_990);
  nand g2901 (n_2697, n_989, n_963);
  nand g2902 (n_1009, n_2695, n_2696, n_2697);
  xor g2903 (n_2698, n_992, n_993);
  xor g2904 (n_998, n_2698, n_994);
  nand g2905 (n_2699, n_992, n_993);
  nand g2906 (n_2700, n_994, n_993);
  nand g2907 (n_2701, n_992, n_994);
  nand g2908 (n_1011, n_2699, n_2700, n_2701);
  xor g2909 (n_2702, n_995, n_996);
  xor g2910 (n_999, n_2702, n_997);
  nand g2911 (n_2703, n_995, n_996);
  nand g2912 (n_2704, n_997, n_996);
  nand g2913 (n_2705, n_995, n_997);
  nand g2914 (n_1013, n_2703, n_2704, n_2705);
  xor g2915 (n_2706, n_998, n_999);
  xor g2916 (n_153, n_2706, n_1000);
  nand g2917 (n_2707, n_998, n_999);
  nand g2918 (n_2708, n_1000, n_999);
  nand g2919 (n_2709, n_998, n_1000);
  nand g2920 (n_152, n_2707, n_2708, n_2709);
  xor g2923 (n_2710, A[55], A[51]);
  xor g2924 (n_1006, n_2710, A[49]);
  nand g2928 (n_1015, n_2528, n_2335, n_2465);
  xor g2936 (n_1008, n_2718, n_1004);
  nand g2938 (n_2720, n_1004, n_975);
  nand g2940 (n_1020, n_2664, n_2720, n_2721);
  xor g2941 (n_2722, n_947, n_1006);
  xor g2942 (n_1010, n_2722, n_1007);
  nand g2943 (n_2723, n_947, n_1006);
  nand g2944 (n_2724, n_1007, n_1006);
  nand g2945 (n_2725, n_947, n_1007);
  nand g2946 (n_1021, n_2723, n_2724, n_2725);
  xor g2947 (n_2726, n_1008, n_1009);
  xor g2948 (n_1012, n_2726, n_1010);
  nand g2949 (n_2727, n_1008, n_1009);
  nand g2950 (n_2728, n_1010, n_1009);
  nand g2951 (n_2729, n_1008, n_1010);
  nand g2952 (n_1024, n_2727, n_2728, n_2729);
  xor g2953 (n_2730, n_1011, n_1012);
  xor g2954 (n_74, n_2730, n_1013);
  nand g2955 (n_2731, n_1011, n_1012);
  nand g2956 (n_2732, n_1013, n_1012);
  nand g2957 (n_2733, n_1011, n_1013);
  nand g2958 (n_73, n_2731, n_2732, n_2733);
  xor g2971 (n_2742, A[46], A[57]);
  xor g2972 (n_1019, n_2742, n_1015);
  nand g2974 (n_2744, n_1015, A[57]);
  nand g2975 (n_2745, A[46], n_1015);
  nand g2976 (n_1031, n_2692, n_2744, n_2745);
  xor g2977 (n_2746, n_960, n_930);
  xor g2978 (n_1022, n_2746, n_963);
  nand g2979 (n_2747, n_960, n_930);
  nand g2980 (n_2748, n_963, n_930);
  nand g2981 (n_2749, n_960, n_963);
  nand g2982 (n_1032, n_2747, n_2748, n_2749);
  xor g2983 (n_2750, n_1019, n_1020);
  xor g2984 (n_1023, n_2750, n_1021);
  nand g2985 (n_2751, n_1019, n_1020);
  nand g2986 (n_2752, n_1021, n_1020);
  nand g2987 (n_2753, n_1019, n_1021);
  nand g2988 (n_1035, n_2751, n_2752, n_2753);
  xor g2989 (n_2754, n_1022, n_1023);
  xor g2990 (n_151, n_2754, n_1024);
  nand g2991 (n_2755, n_1022, n_1023);
  nand g2992 (n_2756, n_1024, n_1023);
  nand g2993 (n_2757, n_1022, n_1024);
  nand g2994 (n_72, n_2755, n_2756, n_2757);
  xor g2998 (n_1029, n_2334, A[57]);
  nand g3002 (n_1037, n_2335, n_2595, n_2529);
  nand g3008 (n_1040, n_2401, n_2764, n_2765);
  xor g3009 (n_2766, n_946, n_975);
  xor g3010 (n_1033, n_2766, n_1029);
  nand g3011 (n_2767, n_946, n_975);
  nand g3012 (n_2768, n_1029, n_975);
  nand g3013 (n_2769, n_946, n_1029);
  nand g3014 (n_1042, n_2767, n_2768, n_2769);
  xor g3015 (n_2770, n_1030, n_1031);
  xor g3016 (n_1034, n_2770, n_1032);
  nand g3017 (n_2771, n_1030, n_1031);
  nand g3018 (n_2772, n_1032, n_1031);
  nand g3019 (n_2773, n_1030, n_1032);
  nand g3020 (n_1044, n_2771, n_2772, n_2773);
  xor g3021 (n_2774, n_1033, n_1034);
  xor g3022 (n_150, n_2774, n_1035);
  nand g3023 (n_2775, n_1033, n_1034);
  nand g3024 (n_2776, n_1035, n_1034);
  nand g3025 (n_2777, n_1033, n_1035);
  nand g3026 (n_71, n_2775, n_2776, n_2777);
  xor g3039 (n_2786, A[55], n_1037);
  xor g3040 (n_1041, n_2786, n_930);
  nand g3041 (n_2787, A[55], n_1037);
  nand g3042 (n_2788, n_930, n_1037);
  nand g3043 (n_2789, A[55], n_930);
  nand g3044 (n_1051, n_2787, n_2788, n_2789);
  xor g3045 (n_2790, n_963, n_1040);
  xor g3046 (n_1043, n_2790, n_1041);
  nand g3047 (n_2791, n_963, n_1040);
  nand g3048 (n_2792, n_1041, n_1040);
  nand g3049 (n_2793, n_963, n_1041);
  nand g3050 (n_1053, n_2791, n_2792, n_2793);
  xor g3051 (n_2794, n_1042, n_1043);
  xor g3052 (n_149, n_2794, n_1044);
  nand g3053 (n_2795, n_1042, n_1043);
  nand g3054 (n_2796, n_1044, n_1043);
  nand g3055 (n_2797, n_1042, n_1044);
  nand g3056 (n_70, n_2795, n_2796, n_2797);
  nand g3069 (n_2805, A[53], n_946);
  nand g3070 (n_1058, n_2764, n_2804, n_2805);
  xor g3071 (n_2806, n_975, n_1029);
  xor g3072 (n_1052, n_2806, n_1050);
  nand g3074 (n_2808, n_1050, n_1029);
  nand g3075 (n_2809, n_975, n_1050);
  nand g3076 (n_1060, n_2768, n_2808, n_2809);
  xor g3077 (n_2810, n_1051, n_1052);
  xor g3078 (n_148, n_2810, n_1053);
  nand g3079 (n_2811, n_1051, n_1052);
  nand g3080 (n_2812, n_1053, n_1052);
  nand g3081 (n_2813, n_1051, n_1053);
  nand g3082 (n_147, n_2811, n_2812, n_2813);
  xor g3090 (n_1057, n_2566, A[55]);
  nand g3092 (n_2820, A[55], A[54]);
  nand g3093 (n_2821, A[50], A[55]);
  nand g3094 (n_1065, n_2496, n_2820, n_2821);
  xor g3095 (n_2822, n_1037, n_963);
  xor g3096 (n_1059, n_2822, n_1057);
  nand g3097 (n_2823, n_1037, n_963);
  nand g3098 (n_2824, n_1057, n_963);
  nand g3099 (n_2825, n_1037, n_1057);
  nand g3100 (n_1067, n_2823, n_2824, n_2825);
  xor g3101 (n_2826, n_1058, n_1059);
  xor g3102 (n_69, n_2826, n_1060);
  nand g3103 (n_2827, n_1058, n_1059);
  nand g3104 (n_2828, n_1060, n_1059);
  nand g3105 (n_2829, n_1058, n_1060);
  nand g3106 (n_146, n_2827, n_2828, n_2829);
  xor g3110 (n_1064, n_2710, A[53]);
  nand g3114 (n_1069, n_2528, n_2463, n_2399);
  xor g3116 (n_1066, n_2718, n_1064);
  nand g3118 (n_2836, n_1064, n_975);
  nand g3120 (n_1072, n_2664, n_2836, n_2837);
  xor g3121 (n_2838, n_1065, n_1066);
  xor g3122 (n_68, n_2838, n_1067);
  nand g3123 (n_2839, n_1065, n_1066);
  nand g3124 (n_2840, n_1067, n_1066);
  nand g3125 (n_2841, n_1065, n_1067);
  nand g3126 (n_145, n_2839, n_2840, n_2841);
  xor g3133 (n_2846, A[54], A[57]);
  xor g3134 (n_1071, n_2846, n_1069);
  nand g3135 (n_2847, A[54], A[57]);
  nand g3136 (n_2848, n_1069, A[57]);
  nand g3137 (n_2849, A[54], n_1069);
  nand g3138 (n_1077, n_2847, n_2848, n_2849);
  xor g3139 (n_2850, n_963, n_1071);
  xor g3140 (n_67, n_2850, n_1072);
  nand g3141 (n_2851, n_963, n_1071);
  nand g3142 (n_2852, n_1072, n_1071);
  nand g3143 (n_2853, n_963, n_1072);
  nand g3144 (n_144, n_2851, n_2852, n_2853);
  nand g3152 (n_1080, n_2463, n_2856, n_2857);
  xor g3153 (n_2858, n_975, n_1076);
  xor g3154 (n_66, n_2858, n_1077);
  nand g3155 (n_2859, n_975, n_1076);
  nand g3156 (n_2860, n_1077, n_1076);
  nand g3157 (n_2861, n_975, n_1077);
  nand g3158 (n_143, n_2859, n_2860, n_2861);
  xor g3160 (n_1079, n_2622, A[54]);
  nand g3164 (n_1083, n_2623, n_2495, n_2865);
  xor g3165 (n_2866, A[57], n_1079);
  xor g3166 (n_65, n_2866, n_1080);
  nand g3167 (n_2867, A[57], n_1079);
  nand g3168 (n_2868, n_1080, n_1079);
  nand g3169 (n_2869, A[57], n_1080);
  nand g3170 (n_142, n_2867, n_2868, n_2869);
  nand g3177 (n_2873, A[57], n_1083);
  nand g3178 (n_141, n_2871, n_2872, n_2873);
  xor g3180 (n_63, n_2622, A[55]);
  nand g3182 (n_2876, A[55], A[56]);
  nand g3184 (n_140, n_2623, n_2876, n_2877);
  nor g11 (n_2893, A[2], A[0]);
  nor g13 (n_2889, A[3], A[1]);
  nor g15 (n_2899, A[2], n_211);
  nand g16 (n_2894, A[2], n_211);
  nor g17 (n_2895, n_132, n_210);
  nand g18 (n_2896, n_132, n_210);
  nor g19 (n_2905, n_131, n_209);
  nand g20 (n_2900, n_131, n_209);
  nor g21 (n_2901, n_130, n_208);
  nand g22 (n_2902, n_130, n_208);
  nor g23 (n_2911, n_129, n_207);
  nand g24 (n_2906, n_129, n_207);
  nor g25 (n_2907, n_128, n_206);
  nand g26 (n_2908, n_128, n_206);
  nor g27 (n_2917, n_127, n_205);
  nand g28 (n_2912, n_127, n_205);
  nor g29 (n_2913, n_126, n_204);
  nand g30 (n_2914, n_126, n_204);
  nor g31 (n_2923, n_125, n_203);
  nand g32 (n_2918, n_125, n_203);
  nor g33 (n_2919, n_124, n_202);
  nand g34 (n_2920, n_124, n_202);
  nor g35 (n_2929, n_123, n_201);
  nand g36 (n_2924, n_123, n_201);
  nor g37 (n_2925, n_122, n_200);
  nand g38 (n_2926, n_122, n_200);
  nor g39 (n_2935, n_121, n_199);
  nand g40 (n_2930, n_121, n_199);
  nor g41 (n_2931, n_120, n_198);
  nand g42 (n_2932, n_120, n_198);
  nor g43 (n_2941, n_119, n_197);
  nand g44 (n_2936, n_119, n_197);
  nor g45 (n_2937, n_118, n_196);
  nand g46 (n_2938, n_118, n_196);
  nor g47 (n_2947, n_117, n_195);
  nand g48 (n_2942, n_117, n_195);
  nor g49 (n_2943, n_116, n_194);
  nand g50 (n_2944, n_116, n_194);
  nor g51 (n_2953, n_115, n_193);
  nand g52 (n_2948, n_115, n_193);
  nor g53 (n_2949, n_114, n_192);
  nand g54 (n_2950, n_114, n_192);
  nor g55 (n_2959, n_113, n_191);
  nand g56 (n_2954, n_113, n_191);
  nor g57 (n_2955, n_112, n_190);
  nand g58 (n_2956, n_112, n_190);
  nor g59 (n_2965, n_111, n_189);
  nand g60 (n_2960, n_111, n_189);
  nor g61 (n_2961, n_110, n_188);
  nand g62 (n_2962, n_110, n_188);
  nor g63 (n_2971, n_109, n_187);
  nand g64 (n_2966, n_109, n_187);
  nor g65 (n_2967, n_108, n_186);
  nand g66 (n_2968, n_108, n_186);
  nor g67 (n_2977, n_107, n_185);
  nand g68 (n_2972, n_107, n_185);
  nor g69 (n_2973, n_106, n_184);
  nand g70 (n_2974, n_106, n_184);
  nor g71 (n_2983, n_105, n_183);
  nand g72 (n_2978, n_105, n_183);
  nor g73 (n_2979, n_104, n_182);
  nand g74 (n_2980, n_104, n_182);
  nor g75 (n_2989, n_103, n_181);
  nand g76 (n_2984, n_103, n_181);
  nor g77 (n_2985, n_102, n_180);
  nand g78 (n_2986, n_102, n_180);
  nor g79 (n_2995, n_101, n_179);
  nand g80 (n_2990, n_101, n_179);
  nor g81 (n_2991, n_100, n_178);
  nand g82 (n_2992, n_100, n_178);
  nor g83 (n_3001, n_99, n_177);
  nand g84 (n_2996, n_99, n_177);
  nor g85 (n_2997, n_98, n_176);
  nand g86 (n_2998, n_98, n_176);
  nor g87 (n_3007, n_97, n_175);
  nand g88 (n_3002, n_97, n_175);
  nor g89 (n_3003, n_96, n_174);
  nand g90 (n_3004, n_96, n_174);
  nor g91 (n_3013, n_95, n_173);
  nand g92 (n_3008, n_95, n_173);
  nor g93 (n_3009, n_94, n_172);
  nand g94 (n_3010, n_94, n_172);
  nor g95 (n_3019, n_93, n_171);
  nand g96 (n_3014, n_93, n_171);
  nor g97 (n_3015, n_92, n_170);
  nand g98 (n_3016, n_92, n_170);
  nor g99 (n_3025, n_91, n_169);
  nand g100 (n_3020, n_91, n_169);
  nor g101 (n_3021, n_90, n_168);
  nand g102 (n_3022, n_90, n_168);
  nor g103 (n_3031, n_89, n_167);
  nand g104 (n_3026, n_89, n_167);
  nor g105 (n_3027, n_88, n_166);
  nand g106 (n_3028, n_88, n_166);
  nor g107 (n_3037, n_87, n_165);
  nand g108 (n_3032, n_87, n_165);
  nor g109 (n_3033, n_86, n_164);
  nand g110 (n_3034, n_86, n_164);
  nor g111 (n_3043, n_85, n_163);
  nand g112 (n_3038, n_85, n_163);
  nor g113 (n_3039, n_84, n_162);
  nand g114 (n_3040, n_84, n_162);
  nor g115 (n_3049, n_83, n_161);
  nand g116 (n_3044, n_83, n_161);
  nor g117 (n_3045, n_82, n_160);
  nand g118 (n_3046, n_82, n_160);
  nor g119 (n_3055, n_81, n_159);
  nand g120 (n_3050, n_81, n_159);
  nor g121 (n_3051, n_80, n_158);
  nand g122 (n_3052, n_80, n_158);
  nor g123 (n_3061, n_79, n_157);
  nand g124 (n_3056, n_79, n_157);
  nor g125 (n_3057, n_78, n_156);
  nand g126 (n_3058, n_78, n_156);
  nor g127 (n_3067, n_77, n_155);
  nand g128 (n_3062, n_77, n_155);
  nor g129 (n_3063, n_76, n_154);
  nand g130 (n_3064, n_76, n_154);
  nor g131 (n_3073, n_75, n_153);
  nand g132 (n_3068, n_75, n_153);
  nor g133 (n_3069, n_74, n_152);
  nand g134 (n_3070, n_74, n_152);
  nor g135 (n_3079, n_73, n_151);
  nand g136 (n_3074, n_73, n_151);
  nor g137 (n_3075, n_72, n_150);
  nand g138 (n_3076, n_72, n_150);
  nor g139 (n_3085, n_71, n_149);
  nand g140 (n_3080, n_71, n_149);
  nor g141 (n_3081, n_70, n_148);
  nand g142 (n_3082, n_70, n_148);
  nor g143 (n_3091, n_69, n_147);
  nand g144 (n_3086, n_69, n_147);
  nor g145 (n_3087, n_68, n_146);
  nand g146 (n_3088, n_68, n_146);
  nor g147 (n_3097, n_67, n_145);
  nand g148 (n_3092, n_67, n_145);
  nor g149 (n_3093, n_66, n_144);
  nand g150 (n_3094, n_66, n_144);
  nor g151 (n_3103, n_65, n_143);
  nand g152 (n_3098, n_65, n_143);
  nor g153 (n_3099, n_64, n_142);
  nand g154 (n_3100, n_64, n_142);
  nor g155 (n_3109, n_63, n_141);
  nand g156 (n_3104, n_63, n_141);
  nor g166 (n_2891, n_1091, n_2889);
  nor g170 (n_2897, n_2894, n_2895);
  nor g173 (n_3124, n_2899, n_2895);
  nor g174 (n_2903, n_2900, n_2901);
  nor g177 (n_3118, n_2905, n_2901);
  nor g178 (n_2909, n_2906, n_2907);
  nor g181 (n_3131, n_2911, n_2907);
  nor g182 (n_2915, n_2912, n_2913);
  nor g185 (n_3125, n_2917, n_2913);
  nor g186 (n_2921, n_2918, n_2919);
  nor g189 (n_3138, n_2923, n_2919);
  nor g190 (n_2927, n_2924, n_2925);
  nor g193 (n_3132, n_2929, n_2925);
  nor g194 (n_2933, n_2930, n_2931);
  nor g197 (n_3145, n_2935, n_2931);
  nor g198 (n_2939, n_2936, n_2937);
  nor g201 (n_3139, n_2941, n_2937);
  nor g202 (n_2945, n_2942, n_2943);
  nor g205 (n_3152, n_2947, n_2943);
  nor g206 (n_2951, n_2948, n_2949);
  nor g209 (n_3146, n_2953, n_2949);
  nor g210 (n_2957, n_2954, n_2955);
  nor g213 (n_3159, n_2959, n_2955);
  nor g214 (n_2963, n_2960, n_2961);
  nor g217 (n_3153, n_2965, n_2961);
  nor g218 (n_2969, n_2966, n_2967);
  nor g221 (n_3166, n_2971, n_2967);
  nor g222 (n_2975, n_2972, n_2973);
  nor g225 (n_3160, n_2977, n_2973);
  nor g226 (n_2981, n_2978, n_2979);
  nor g229 (n_3173, n_2983, n_2979);
  nor g230 (n_2987, n_2984, n_2985);
  nor g233 (n_3167, n_2989, n_2985);
  nor g234 (n_2993, n_2990, n_2991);
  nor g237 (n_3180, n_2995, n_2991);
  nor g238 (n_2999, n_2996, n_2997);
  nor g241 (n_3174, n_3001, n_2997);
  nor g242 (n_3005, n_3002, n_3003);
  nor g245 (n_3187, n_3007, n_3003);
  nor g246 (n_3011, n_3008, n_3009);
  nor g249 (n_3181, n_3013, n_3009);
  nor g250 (n_3017, n_3014, n_3015);
  nor g253 (n_3194, n_3019, n_3015);
  nor g254 (n_3023, n_3020, n_3021);
  nor g257 (n_3188, n_3025, n_3021);
  nor g258 (n_3029, n_3026, n_3027);
  nor g261 (n_3201, n_3031, n_3027);
  nor g262 (n_3035, n_3032, n_3033);
  nor g265 (n_3195, n_3037, n_3033);
  nor g266 (n_3041, n_3038, n_3039);
  nor g269 (n_3208, n_3043, n_3039);
  nor g270 (n_3047, n_3044, n_3045);
  nor g273 (n_3202, n_3049, n_3045);
  nor g274 (n_3053, n_3050, n_3051);
  nor g277 (n_3215, n_3055, n_3051);
  nor g278 (n_3059, n_3056, n_3057);
  nor g281 (n_3209, n_3061, n_3057);
  nor g282 (n_3065, n_3062, n_3063);
  nor g285 (n_3222, n_3067, n_3063);
  nor g286 (n_3071, n_3068, n_3069);
  nor g289 (n_3216, n_3073, n_3069);
  nor g290 (n_3077, n_3074, n_3075);
  nor g293 (n_3229, n_3079, n_3075);
  nor g294 (n_3083, n_3080, n_3081);
  nor g297 (n_3223, n_3085, n_3081);
  nor g298 (n_3089, n_3086, n_3087);
  nor g301 (n_3236, n_3091, n_3087);
  nor g302 (n_3095, n_3092, n_3093);
  nor g305 (n_3230, n_3097, n_3093);
  nor g306 (n_3101, n_3098, n_3099);
  nor g309 (n_3243, n_3103, n_3099);
  nor g310 (n_3107, n_3104, n_3105);
  nor g313 (n_3237, n_3109, n_3105);
  nand g324 (n_3244, n_3124, n_3118);
  nand g329 (n_3254, n_3131, n_3125);
  nand g334 (n_3249, n_3138, n_3132);
  nand g339 (n_3260, n_3145, n_3139);
  nand g344 (n_3255, n_3152, n_3146);
  nand g349 (n_3266, n_3159, n_3153);
  nand g354 (n_3261, n_3166, n_3160);
  nand g359 (n_3272, n_3173, n_3167);
  nand g364 (n_3267, n_3180, n_3174);
  nand g369 (n_3278, n_3187, n_3181);
  nand g374 (n_3273, n_3194, n_3188);
  nand g379 (n_3284, n_3201, n_3195);
  nand g384 (n_3279, n_3208, n_3202);
  nand g389 (n_3290, n_3215, n_3209);
  nand g394 (n_3285, n_3222, n_3216);
  nand g399 (n_3296, n_3229, n_3223);
  nand g404 (n_3291, n_3236, n_3230);
  nand g409 (n_3366, n_3243, n_3237);
  nand g412 (n_3298, n_3247, n_3248);
  nor g413 (n_3252, n_3249, n_3250);
  nor g416 (n_3297, n_3254, n_3249);
  nor g417 (n_3258, n_3255, n_3256);
  nor g420 (n_3307, n_3260, n_3255);
  nor g421 (n_3264, n_3261, n_3262);
  nor g424 (n_3301, n_3266, n_3261);
  nor g425 (n_3270, n_3267, n_3268);
  nor g428 (n_3314, n_3272, n_3267);
  nor g429 (n_3276, n_3273, n_3274);
  nor g432 (n_3308, n_3278, n_3273);
  nor g433 (n_3282, n_3279, n_3280);
  nor g436 (n_3321, n_3284, n_3279);
  nor g437 (n_3288, n_3285, n_3286);
  nor g440 (n_3315, n_3290, n_3285);
  nor g441 (n_3294, n_3291, n_3292);
  nor g444 (n_3343, n_3296, n_3291);
  nand g445 (n_3300, n_3297, n_3298);
  nand g446 (n_3323, n_3299, n_3300);
  nand g451 (n_3322, n_3307, n_3301);
  nand g456 (n_3332, n_3314, n_3308);
  nand g461 (n_3327, n_3321, n_3315);
  nand g464 (n_3334, n_3325, n_3326);
  nor g465 (n_3330, n_3327, n_3328);
  nor g3192 (n_3333, n_3332, n_3327);
  nand g3193 (n_3336, n_3333, n_3334);
  nand g3194 (n_3344, n_3335, n_3336);
  nand g3197 (n_3341, n_3328, n_3338);
  nand g3198 (n_3339, n_3307, n_3323);
  nand g3199 (n_3351, n_3302, n_3339);
  nand g3200 (n_3340, n_3314, n_3334);
  nand g3201 (n_3356, n_3309, n_3340);
  nand g3202 (n_3342, n_3321, n_3341);
  nand g3203 (n_3361, n_3316, n_3342);
  nand g3204 (n_3346, n_3343, n_3344);
  nand g3205 (n_3367, n_3345, n_3346);
  nand g3208 (n_3373, n_3250, n_3348);
  nand g3211 (n_3376, n_3256, n_3350);
  nand g3214 (n_3379, n_3262, n_3353);
  nand g3217 (n_3382, n_3268, n_3355);
  nand g3220 (n_3385, n_3274, n_3358);
  nand g3223 (n_3388, n_3280, n_3360);
  nand g3226 (n_3391, n_3286, n_3363);
  nand g3229 (n_3394, n_3292, n_3365);
  nand g3232 (n_3397, n_3369, n_3370);
  nand g3234 (n_3402, n_3119, n_3371);
  nand g3235 (n_3372, n_3131, n_3298);
  nand g3236 (n_3407, n_3126, n_3372);
  nand g3237 (n_3374, n_3138, n_3373);
  nand g3238 (n_3412, n_3133, n_3374);
  nand g3239 (n_3375, n_3145, n_3323);
  nand g3240 (n_3417, n_3140, n_3375);
  nand g3241 (n_3377, n_3152, n_3376);
  nand g3242 (n_3422, n_3147, n_3377);
  nand g3243 (n_3378, n_3159, n_3351);
  nand g3244 (n_3427, n_3154, n_3378);
  nand g3245 (n_3380, n_3166, n_3379);
  nand g3246 (n_3432, n_3161, n_3380);
  nand g3247 (n_3381, n_3173, n_3334);
  nand g3248 (n_3437, n_3168, n_3381);
  nand g3249 (n_3383, n_3180, n_3382);
  nand g3250 (n_3442, n_3175, n_3383);
  nand g3251 (n_3384, n_3187, n_3356);
  nand g3252 (n_3447, n_3182, n_3384);
  nand g3253 (n_3386, n_3194, n_3385);
  nand g3254 (n_3452, n_3189, n_3386);
  nand g3255 (n_3387, n_3201, n_3341);
  nand g3256 (n_3457, n_3196, n_3387);
  nand g3257 (n_3389, n_3208, n_3388);
  nand g3258 (n_3462, n_3203, n_3389);
  nand g3259 (n_3390, n_3215, n_3361);
  nand g3260 (n_3467, n_3210, n_3390);
  nand g3261 (n_3392, n_3222, n_3391);
  nand g3262 (n_3472, n_3217, n_3392);
  nand g3263 (n_3393, n_3229, n_3344);
  nand g3264 (n_3477, n_3224, n_3393);
  nand g3265 (n_3395, n_3236, n_3394);
  nand g3266 (n_3482, n_3231, n_3395);
  nand g3267 (n_3396, n_3243, n_3367);
  nand g3268 (n_3487, n_3238, n_3396);
  nand g3274 (n_3499, n_2894, n_3401);
  nand g3277 (n_3503, n_2900, n_3404);
  nand g3280 (n_3507, n_2906, n_3406);
  nand g3283 (n_3511, n_2912, n_3409);
  nand g3286 (n_3515, n_2918, n_3411);
  nand g3289 (n_3519, n_2924, n_3414);
  nand g3292 (n_3523, n_2930, n_3416);
  nand g3295 (n_3527, n_2936, n_3419);
  nand g3298 (n_3531, n_2942, n_3421);
  nand g3301 (n_3535, n_2948, n_3424);
  nand g3304 (n_3539, n_2954, n_3426);
  nand g3307 (n_3543, n_2960, n_3429);
  nand g3310 (n_3547, n_2966, n_3431);
  nand g3313 (n_3551, n_2972, n_3434);
  nand g3316 (n_3555, n_2978, n_3436);
  nand g3319 (n_3559, n_2984, n_3439);
  nand g3322 (n_3563, n_2990, n_3441);
  nand g3325 (n_3567, n_2996, n_3444);
  nand g3328 (n_3571, n_3002, n_3446);
  nand g3331 (n_3575, n_3008, n_3449);
  nand g3334 (n_3579, n_3014, n_3451);
  nand g3337 (n_3583, n_3020, n_3454);
  nand g3340 (n_3587, n_3026, n_3456);
  nand g3343 (n_3591, n_3032, n_3459);
  nand g3346 (n_3595, n_3038, n_3461);
  nand g3349 (n_3599, n_3044, n_3464);
  nand g3352 (n_3603, n_3050, n_3466);
  nand g3355 (n_3607, n_3056, n_3469);
  nand g3358 (n_3611, n_3062, n_3471);
  nand g3361 (n_3615, n_3068, n_3474);
  nand g3364 (n_3619, n_3074, n_3476);
  nand g3367 (n_3623, n_3080, n_3479);
  nand g3370 (n_3627, n_3086, n_3481);
  nand g3373 (n_3631, n_3092, n_3484);
  nand g3376 (n_3635, n_3098, n_3486);
  nand g3379 (n_3639, n_3104, n_3489);
  nand g3382 (n_3643, n_3110, n_3491);
  xnor g3394 (Z[5], n_3499, n_3500);
  xnor g3396 (Z[6], n_3402, n_3501);
  xnor g3399 (Z[7], n_3503, n_3504);
  xnor g3401 (Z[8], n_3298, n_3505);
  xnor g3404 (Z[9], n_3507, n_3508);
  xnor g3406 (Z[10], n_3407, n_3509);
  xnor g3409 (Z[11], n_3511, n_3512);
  xnor g3411 (Z[12], n_3373, n_3513);
  xnor g3414 (Z[13], n_3515, n_3516);
  xnor g3416 (Z[14], n_3412, n_3517);
  xnor g3419 (Z[15], n_3519, n_3520);
  xnor g3421 (Z[16], n_3323, n_3521);
  xnor g3424 (Z[17], n_3523, n_3524);
  xnor g3426 (Z[18], n_3417, n_3525);
  xnor g3429 (Z[19], n_3527, n_3528);
  xnor g3431 (Z[20], n_3376, n_3529);
  xnor g3434 (Z[21], n_3531, n_3532);
  xnor g3436 (Z[22], n_3422, n_3533);
  xnor g3439 (Z[23], n_3535, n_3536);
  xnor g3441 (Z[24], n_3351, n_3537);
  xnor g3444 (Z[25], n_3539, n_3540);
  xnor g3446 (Z[26], n_3427, n_3541);
  xnor g3449 (Z[27], n_3543, n_3544);
  xnor g3451 (Z[28], n_3379, n_3545);
  xnor g3454 (Z[29], n_3547, n_3548);
  xnor g3456 (Z[30], n_3432, n_3549);
  xnor g3459 (Z[31], n_3551, n_3552);
  xnor g3461 (Z[32], n_3334, n_3553);
  xnor g3464 (Z[33], n_3555, n_3556);
  xnor g3466 (Z[34], n_3437, n_3557);
  xnor g3469 (Z[35], n_3559, n_3560);
  xnor g3471 (Z[36], n_3382, n_3561);
  xnor g3474 (Z[37], n_3563, n_3564);
  xnor g3476 (Z[38], n_3442, n_3565);
  xnor g3479 (Z[39], n_3567, n_3568);
  xnor g3481 (Z[40], n_3356, n_3569);
  xnor g3484 (Z[41], n_3571, n_3572);
  xnor g3486 (Z[42], n_3447, n_3573);
  xnor g3489 (Z[43], n_3575, n_3576);
  xnor g3491 (Z[44], n_3385, n_3577);
  xnor g3494 (Z[45], n_3579, n_3580);
  xnor g3496 (Z[46], n_3452, n_3581);
  xnor g3499 (Z[47], n_3583, n_3584);
  xnor g3501 (Z[48], n_3341, n_3585);
  xnor g3504 (Z[49], n_3587, n_3588);
  xnor g3506 (Z[50], n_3457, n_3589);
  xnor g3509 (Z[51], n_3591, n_3592);
  xnor g3511 (Z[52], n_3388, n_3593);
  xnor g3514 (Z[53], n_3595, n_3596);
  xnor g3516 (Z[54], n_3462, n_3597);
  xnor g3519 (Z[55], n_3599, n_3600);
  xnor g3521 (Z[56], n_3361, n_3601);
  xnor g3524 (Z[57], n_3603, n_3604);
  xnor g3526 (Z[58], n_3467, n_3605);
  xnor g3529 (Z[59], n_3607, n_3608);
  xnor g3531 (Z[60], n_3391, n_3609);
  xnor g3534 (Z[61], n_3611, n_3612);
  xnor g3536 (Z[62], n_3472, n_3613);
  xnor g3539 (Z[63], n_3615, n_3616);
  xnor g3541 (Z[64], n_3344, n_3617);
  xnor g3544 (Z[65], n_3619, n_3620);
  xnor g3546 (Z[66], n_3477, n_3621);
  xnor g3549 (Z[67], n_3623, n_3624);
  xnor g3551 (Z[68], n_3394, n_3625);
  xnor g3554 (Z[69], n_3627, n_3628);
  xnor g3556 (Z[70], n_3482, n_3629);
  xnor g3559 (Z[71], n_3631, n_3632);
  xnor g3561 (Z[72], n_3367, n_3633);
  xnor g3564 (Z[73], n_3635, n_3636);
  xnor g3566 (Z[74], n_3487, n_3637);
  xnor g3569 (Z[75], n_3639, n_3640);
  xnor g3571 (Z[76], n_3397, n_3641);
  or g3587 (n_302, wc, wc0, n_132);
  not gc0 (wc0, n_1091);
  not gc (wc, n_1105);
  or g3588 (n_311, wc1, wc2, n_296);
  not gc2 (wc2, n_1105);
  not gc1 (wc1, n_1124);
  or g3589 (n_324, wc3, n_301, n_296);
  not gc3 (wc3, n_1152);
  or g3590 (n_341, wc4, wc5, n_301);
  not gc5 (wc5, n_1187);
  not gc4 (wc4, n_1188);
  or g3591 (n_363, wc6, wc7, n_301);
  not gc7 (wc7, n_1235);
  not gc6 (wc6, n_1236);
  or g3592 (n_410, wc8, wc9, n_296);
  not gc9 (wc9, n_1236);
  not gc8 (wc8, n_1283);
  or g3593 (n_438, wc10, wc11, n_301);
  not gc11 (wc11, n_1412);
  not gc10 (wc10, n_1413);
  or g3594 (n_466, wc12, wc13, n_310);
  not gc13 (wc13, n_1352);
  not gc12 (wc12, n_1476);
  or g3595 (n_492, wc14, wc15, n_323);
  not gc15 (wc15, n_1416);
  not gc14 (wc14, n_1540);
  or g3596 (n_520, wc16, wc17, n_340);
  not gc17 (wc17, n_1345);
  not gc16 (wc16, n_1604);
  or g3597 (n_548, wc18, wc19, n_361);
  not gc19 (wc19, n_1409);
  not gc18 (wc18, n_1668);
  or g3598 (n_576, wc20, wc21, n_386);
  not gc21 (wc21, n_1473);
  not gc20 (wc20, n_1732);
  xnor g3599 (n_2622, A[58], A[56]);
  or g3600 (n_2623, wc22, A[58]);
  not gc22 (wc22, A[56]);
  or g3601 (n_2625, wc23, A[58]);
  not gc23 (wc23, A[52]);
  xnor g3602 (n_2662, A[57], A[45]);
  or g3603 (n_2663, wc24, A[57]);
  not gc24 (wc24, A[45]);
  xnor g3604 (n_1030, n_2598, A[55]);
  or g3605 (n_2764, wc25, A[55]);
  not gc25 (wc25, A[53]);
  or g3606 (n_2765, wc26, A[55]);
  not gc26 (wc26, A[47]);
  xnor g3608 (n_1076, n_2462, A[57]);
  or g3609 (n_2856, wc27, A[57]);
  not gc27 (wc27, A[53]);
  or g3610 (n_2857, wc28, A[57]);
  not gc28 (wc28, A[55]);
  or g3611 (n_2865, wc29, A[58]);
  not gc29 (wc29, A[54]);
  or g3613 (n_2871, A[55], wc30);
  not gc30 (wc30, A[57]);
  or g3614 (n_2877, wc31, A[58]);
  not gc31 (wc31, A[55]);
  and g3615 (n_3113, wc32, A[58]);
  not gc32 (wc32, A[57]);
  or g3616 (n_3110, wc33, A[58]);
  not gc33 (wc33, A[57]);
  or g3617 (n_392, wc34, wc35, n_301);
  not gc35 (wc35, n_1292);
  not gc34 (wc34, n_1293);
  or g3618 (n_2721, A[57], wc36);
  not gc36 (wc36, n_1004);
  xnor g3619 (n_1050, n_2462, n_946);
  or g3620 (n_2804, A[55], wc37);
  not gc37 (wc37, n_946);
  or g3621 (n_2837, A[57], wc38);
  not gc38 (wc38, n_1064);
  and g3622 (n_3116, wc39, n_1088);
  not gc39 (wc39, n_2891);
  or g3624 (n_3493, n_2893, wc40);
  not gc40 (wc40, n_1091);
  or g3625 (n_3496, n_2889, wc41);
  not gc41 (wc41, n_1088);
  xnor g3626 (n_2634, n_959, A[58]);
  or g3627 (n_2635, A[58], wc42);
  not gc42 (wc42, n_959);
  or g3628 (n_2637, A[58], wc43);
  not gc43 (wc43, n_960);
  or g3629 (n_2664, A[57], wc44);
  not gc44 (wc44, n_975);
  xnor g3630 (n_2718, n_975, A[57]);
  xnor g3631 (n_64, n_2526, n_1083);
  or g3632 (n_2872, A[55], wc45);
  not gc45 (wc45, n_1083);
  and g3633 (n_3105, A[57], wc46);
  not gc46 (wc46, n_140);
  or g3634 (n_3106, A[57], wc47);
  not gc47 (wc47, n_140);
  or g3635 (n_3497, wc48, n_2899);
  not gc48 (wc48, n_2894);
  or g3636 (n_3641, wc49, n_3113);
  not gc49 (wc49, n_3110);
  and g3637 (n_3119, wc50, n_2896);
  not gc50 (wc50, n_2897);
  not g3638 (Z[2], n_3493);
  or g3639 (n_3500, wc51, n_2895);
  not gc51 (wc51, n_2896);
  or g3640 (n_3501, wc52, n_2905);
  not gc52 (wc52, n_2900);
  and g3641 (n_3121, wc53, n_2902);
  not gc53 (wc53, n_2903);
  or g3644 (n_3504, wc54, n_2901);
  not gc54 (wc54, n_2902);
  or g3645 (n_3640, wc55, n_3105);
  not gc55 (wc55, n_3106);
  and g3646 (n_3126, wc56, n_2908);
  not gc56 (wc56, n_2909);
  and g3647 (n_3122, wc57, n_3118);
  not gc57 (wc57, n_3119);
  or g3648 (n_3371, n_3116, wc58);
  not gc58 (wc58, n_3124);
  or g3649 (n_3401, n_2899, n_3116);
  xor g3650 (Z[3], n_1091, n_3496);
  xor g3651 (Z[4], n_3116, n_3497);
  or g3652 (n_3505, wc59, n_2911);
  not gc59 (wc59, n_2906);
  or g3653 (n_3508, wc60, n_2907);
  not gc60 (wc60, n_2908);
  and g3654 (n_3240, n_3106, wc61);
  not gc61 (wc61, n_3107);
  and g3655 (n_3247, wc62, n_3121);
  not gc62 (wc62, n_3122);
  or g3656 (n_3248, n_3244, n_3116);
  or g3657 (n_3509, wc63, n_2917);
  not gc63 (wc63, n_2912);
  or g3658 (n_3636, wc64, n_3099);
  not gc64 (wc64, n_3100);
  or g3659 (n_3637, wc65, n_3109);
  not gc65 (wc65, n_3104);
  and g3660 (n_3128, wc66, n_2914);
  not gc66 (wc66, n_2915);
  and g3661 (n_3133, wc67, n_2920);
  not gc67 (wc67, n_2921);
  and g3662 (n_3238, wc68, n_3100);
  not gc68 (wc68, n_3101);
  or g3663 (n_3404, wc69, n_2905);
  not gc69 (wc69, n_3402);
  or g3664 (n_3512, wc70, n_2913);
  not gc70 (wc70, n_2914);
  or g3665 (n_3513, wc71, n_2923);
  not gc71 (wc71, n_2918);
  or g3666 (n_3516, wc72, n_2919);
  not gc72 (wc72, n_2920);
  or g3667 (n_3633, wc73, n_3103);
  not gc73 (wc73, n_3098);
  and g3668 (n_3135, wc74, n_2926);
  not gc74 (wc74, n_2927);
  and g3669 (n_3233, wc75, n_3094);
  not gc75 (wc75, n_3095);
  and g3670 (n_3129, wc76, n_3125);
  not gc76 (wc76, n_3126);
  and g3671 (n_3241, wc77, n_3237);
  not gc77 (wc77, n_3238);
  or g3672 (n_3406, wc78, n_2911);
  not gc78 (wc78, n_3298);
  or g3673 (n_3517, wc79, n_2929);
  not gc79 (wc79, n_2924);
  or g3674 (n_3520, wc80, n_2925);
  not gc80 (wc80, n_2926);
  or g3675 (n_3628, wc81, n_3087);
  not gc81 (wc81, n_3088);
  or g3676 (n_3629, wc82, n_3097);
  not gc82 (wc82, n_3092);
  or g3677 (n_3632, wc83, n_3093);
  not gc83 (wc83, n_3094);
  and g3678 (n_3140, wc84, n_2932);
  not gc84 (wc84, n_2933);
  and g3679 (n_3142, wc85, n_2938);
  not gc85 (wc85, n_2939);
  and g3680 (n_3231, wc86, n_3088);
  not gc86 (wc86, n_3089);
  and g3681 (n_3250, wc87, n_3128);
  not gc87 (wc87, n_3129);
  and g3682 (n_3136, wc88, n_3132);
  not gc88 (wc88, n_3133);
  and g3683 (n_3369, wc89, n_3240);
  not gc89 (wc89, n_3241);
  or g3684 (n_3348, wc90, n_3254);
  not gc90 (wc90, n_3298);
  or g3685 (n_3521, wc91, n_2935);
  not gc91 (wc91, n_2930);
  or g3686 (n_3524, wc92, n_2931);
  not gc92 (wc92, n_2932);
  or g3687 (n_3525, wc93, n_2941);
  not gc93 (wc93, n_2936);
  or g3688 (n_3528, wc94, n_2937);
  not gc94 (wc94, n_2938);
  or g3689 (n_3529, wc95, n_2947);
  not gc95 (wc95, n_2942);
  or g3690 (n_3625, wc96, n_3091);
  not gc96 (wc96, n_3086);
  and g3691 (n_3147, wc97, n_2944);
  not gc97 (wc97, n_2945);
  and g3692 (n_3226, wc98, n_3082);
  not gc98 (wc98, n_3083);
  and g3693 (n_3251, wc99, n_3135);
  not gc99 (wc99, n_3136);
  and g3694 (n_3143, wc100, n_3139);
  not gc100 (wc100, n_3140);
  and g3695 (n_3234, wc101, n_3230);
  not gc101 (wc101, n_3231);
  or g3696 (n_3409, wc102, n_2917);
  not gc102 (wc102, n_3407);
  or g3697 (n_3532, wc103, n_2943);
  not gc103 (wc103, n_2944);
  or g3698 (n_3533, wc104, n_2953);
  not gc104 (wc104, n_2948);
  or g3699 (n_3620, wc105, n_3075);
  not gc105 (wc105, n_3076);
  or g3700 (n_3621, wc106, n_3085);
  not gc106 (wc106, n_3080);
  or g3701 (n_3624, wc107, n_3081);
  not gc107 (wc107, n_3082);
  and g3702 (n_3149, wc108, n_2950);
  not gc108 (wc108, n_2951);
  and g3703 (n_3154, wc109, n_2956);
  not gc109 (wc109, n_2957);
  and g3704 (n_3156, wc110, n_2962);
  not gc110 (wc110, n_2963);
  and g3705 (n_3161, wc111, n_2968);
  not gc111 (wc111, n_2969);
  and g3706 (n_3163, wc112, n_2974);
  not gc112 (wc112, n_2975);
  and g3707 (n_3168, wc113, n_2980);
  not gc113 (wc113, n_2981);
  and g3708 (n_3170, wc114, n_2986);
  not gc114 (wc114, n_2987);
  and g3709 (n_3175, wc115, n_2992);
  not gc115 (wc115, n_2993);
  and g3710 (n_3177, wc116, n_2998);
  not gc116 (wc116, n_2999);
  and g3711 (n_3182, wc117, n_3004);
  not gc117 (wc117, n_3005);
  and g3712 (n_3184, wc118, n_3010);
  not gc118 (wc118, n_3011);
  and g3713 (n_3189, wc119, n_3016);
  not gc119 (wc119, n_3017);
  and g3714 (n_3191, wc120, n_3022);
  not gc120 (wc120, n_3023);
  and g3715 (n_3196, wc121, n_3028);
  not gc121 (wc121, n_3029);
  and g3716 (n_3198, wc122, n_3034);
  not gc122 (wc122, n_3035);
  and g3717 (n_3203, wc123, n_3040);
  not gc123 (wc123, n_3041);
  and g3718 (n_3205, wc124, n_3046);
  not gc124 (wc124, n_3047);
  and g3719 (n_3210, wc125, n_3052);
  not gc125 (wc125, n_3053);
  and g3720 (n_3212, wc126, n_3058);
  not gc126 (wc126, n_3059);
  and g3721 (n_3256, wc127, n_3142);
  not gc127 (wc127, n_3143);
  and g3722 (n_3293, wc128, n_3233);
  not gc128 (wc128, n_3234);
  or g3723 (n_3411, wc129, n_2923);
  not gc129 (wc129, n_3373);
  or g3724 (n_3536, wc130, n_2949);
  not gc130 (wc130, n_2950);
  or g3725 (n_3537, wc131, n_2959);
  not gc131 (wc131, n_2954);
  or g3726 (n_3540, wc132, n_2955);
  not gc132 (wc132, n_2956);
  or g3727 (n_3541, wc133, n_2965);
  not gc133 (wc133, n_2960);
  or g3728 (n_3544, wc134, n_2961);
  not gc134 (wc134, n_2962);
  or g3729 (n_3545, wc135, n_2971);
  not gc135 (wc135, n_2966);
  or g3730 (n_3548, wc136, n_2967);
  not gc136 (wc136, n_2968);
  or g3731 (n_3549, wc137, n_2977);
  not gc137 (wc137, n_2972);
  or g3732 (n_3552, wc138, n_2973);
  not gc138 (wc138, n_2974);
  or g3733 (n_3553, wc139, n_2983);
  not gc139 (wc139, n_2978);
  or g3734 (n_3556, wc140, n_2979);
  not gc140 (wc140, n_2980);
  or g3735 (n_3557, wc141, n_2989);
  not gc141 (wc141, n_2984);
  or g3736 (n_3560, wc142, n_2985);
  not gc142 (wc142, n_2986);
  or g3737 (n_3561, wc143, n_2995);
  not gc143 (wc143, n_2990);
  or g3738 (n_3564, wc144, n_2991);
  not gc144 (wc144, n_2992);
  or g3739 (n_3565, wc145, n_3001);
  not gc145 (wc145, n_2996);
  or g3740 (n_3568, wc146, n_2997);
  not gc146 (wc146, n_2998);
  or g3741 (n_3569, wc147, n_3007);
  not gc147 (wc147, n_3002);
  or g3742 (n_3572, wc148, n_3003);
  not gc148 (wc148, n_3004);
  or g3743 (n_3573, wc149, n_3013);
  not gc149 (wc149, n_3008);
  or g3744 (n_3576, wc150, n_3009);
  not gc150 (wc150, n_3010);
  or g3745 (n_3577, wc151, n_3019);
  not gc151 (wc151, n_3014);
  or g3746 (n_3580, wc152, n_3015);
  not gc152 (wc152, n_3016);
  or g3747 (n_3581, wc153, n_3025);
  not gc153 (wc153, n_3020);
  or g3748 (n_3584, wc154, n_3021);
  not gc154 (wc154, n_3022);
  or g3749 (n_3585, wc155, n_3031);
  not gc155 (wc155, n_3026);
  or g3750 (n_3588, wc156, n_3027);
  not gc156 (wc156, n_3028);
  or g3751 (n_3589, wc157, n_3037);
  not gc157 (wc157, n_3032);
  or g3752 (n_3592, wc158, n_3033);
  not gc158 (wc158, n_3034);
  or g3753 (n_3593, wc159, n_3043);
  not gc159 (wc159, n_3038);
  or g3754 (n_3596, wc160, n_3039);
  not gc160 (wc160, n_3040);
  or g3755 (n_3597, wc161, n_3049);
  not gc161 (wc161, n_3044);
  or g3756 (n_3600, wc162, n_3045);
  not gc162 (wc162, n_3046);
  or g3757 (n_3601, wc163, n_3055);
  not gc163 (wc163, n_3050);
  or g3758 (n_3604, wc164, n_3051);
  not gc164 (wc164, n_3052);
  or g3759 (n_3605, wc165, n_3061);
  not gc165 (wc165, n_3056);
  or g3760 (n_3608, wc166, n_3057);
  not gc166 (wc166, n_3058);
  or g3761 (n_3616, wc167, n_3069);
  not gc167 (wc167, n_3070);
  and g3762 (n_3217, wc168, n_3064);
  not gc168 (wc168, n_3065);
  and g3763 (n_3224, wc169, n_3076);
  not gc169 (wc169, n_3077);
  and g3764 (n_3150, wc170, n_3146);
  not gc170 (wc170, n_3147);
  and g3765 (n_3157, wc171, n_3153);
  not gc171 (wc171, n_3154);
  and g3766 (n_3164, wc172, n_3160);
  not gc172 (wc172, n_3161);
  and g3767 (n_3171, wc173, n_3167);
  not gc173 (wc173, n_3168);
  and g3768 (n_3178, wc174, n_3174);
  not gc174 (wc174, n_3175);
  and g3769 (n_3185, wc175, n_3181);
  not gc175 (wc175, n_3182);
  and g3770 (n_3192, wc176, n_3188);
  not gc176 (wc176, n_3189);
  and g3771 (n_3199, wc177, n_3195);
  not gc177 (wc177, n_3196);
  and g3772 (n_3206, wc178, n_3202);
  not gc178 (wc178, n_3203);
  and g3773 (n_3213, wc179, n_3209);
  not gc179 (wc179, n_3210);
  and g3774 (n_3299, n_3251, wc180);
  not gc180 (wc180, n_3252);
  or g3775 (n_3609, wc181, n_3067);
  not gc181 (wc181, n_3062);
  or g3776 (n_3612, wc182, n_3063);
  not gc182 (wc182, n_3064);
  or g3777 (n_3617, wc183, n_3079);
  not gc183 (wc183, n_3074);
  and g3778 (n_3219, wc184, n_3070);
  not gc184 (wc184, n_3071);
  and g3779 (n_3257, wc185, n_3149);
  not gc185 (wc185, n_3150);
  and g3780 (n_3262, wc186, n_3156);
  not gc186 (wc186, n_3157);
  and g3781 (n_3263, wc187, n_3163);
  not gc187 (wc187, n_3164);
  and g3782 (n_3268, wc188, n_3170);
  not gc188 (wc188, n_3171);
  and g3783 (n_3269, wc189, n_3177);
  not gc189 (wc189, n_3178);
  and g3784 (n_3274, wc190, n_3184);
  not gc190 (wc190, n_3185);
  and g3785 (n_3275, wc191, n_3191);
  not gc191 (wc191, n_3192);
  and g3786 (n_3280, wc192, n_3198);
  not gc192 (wc192, n_3199);
  and g3787 (n_3281, wc193, n_3205);
  not gc193 (wc193, n_3206);
  and g3788 (n_3286, wc194, n_3212);
  not gc194 (wc194, n_3213);
  and g3789 (n_3227, wc195, n_3223);
  not gc195 (wc195, n_3224);
  or g3790 (n_3414, wc196, n_2929);
  not gc196 (wc196, n_3412);
  or g3791 (n_3613, wc197, n_3073);
  not gc197 (wc197, n_3068);
  and g3792 (n_3220, wc198, n_3216);
  not gc198 (wc198, n_3217);
  and g3793 (n_3292, wc199, n_3226);
  not gc199 (wc199, n_3227);
  or g3794 (n_3350, wc200, n_3260);
  not gc200 (wc200, n_3323);
  or g3795 (n_3416, wc201, n_2935);
  not gc201 (wc201, n_3323);
  and g3796 (n_3287, wc202, n_3219);
  not gc202 (wc202, n_3220);
  and g3797 (n_3302, n_3257, wc203);
  not gc203 (wc203, n_3258);
  and g3798 (n_3304, n_3263, wc204);
  not gc204 (wc204, n_3264);
  and g3799 (n_3309, n_3269, wc205);
  not gc205 (wc205, n_3270);
  and g3800 (n_3311, n_3275, wc206);
  not gc206 (wc206, n_3276);
  and g3801 (n_3316, n_3281, wc207);
  not gc207 (wc207, n_3282);
  or g3802 (n_3326, n_3322, wc208);
  not gc208 (wc208, n_3323);
  and g3803 (n_3345, n_3293, wc209);
  not gc209 (wc209, n_3294);
  and g3804 (n_3305, wc210, n_3301);
  not gc210 (wc210, n_3302);
  and g3805 (n_3312, wc211, n_3308);
  not gc211 (wc211, n_3309);
  and g3806 (n_3319, wc212, n_3315);
  not gc212 (wc212, n_3316);
  or g3807 (n_3419, wc213, n_2941);
  not gc213 (wc213, n_3417);
  or g3808 (n_3421, wc214, n_2947);
  not gc214 (wc214, n_3376);
  and g3809 (n_3318, n_3287, wc215);
  not gc215 (wc215, n_3288);
  and g3810 (n_3325, wc216, n_3304);
  not gc216 (wc216, n_3305);
  and g3811 (n_3328, wc217, n_3311);
  not gc217 (wc217, n_3312);
  or g3812 (n_3353, wc218, n_3266);
  not gc218 (wc218, n_3351);
  or g3813 (n_3426, wc219, n_2959);
  not gc219 (wc219, n_3351);
  or g3814 (n_3424, wc220, n_2953);
  not gc220 (wc220, n_3422);
  and g3815 (n_3329, n_3318, wc221);
  not gc221 (wc221, n_3319);
  or g3816 (n_3338, wc222, n_3332);
  not gc222 (wc222, n_3334);
  or g3817 (n_3355, wc223, n_3272);
  not gc223 (wc223, n_3334);
  or g3818 (n_3429, wc224, n_2965);
  not gc224 (wc224, n_3427);
  or g3819 (n_3431, wc225, n_2971);
  not gc225 (wc225, n_3379);
  or g3820 (n_3436, wc226, n_2983);
  not gc226 (wc226, n_3334);
  and g3821 (n_3335, n_3329, wc227);
  not gc227 (wc227, n_3330);
  or g3822 (n_3358, wc228, n_3278);
  not gc228 (wc228, n_3356);
  or g3823 (n_3360, wc229, n_3284);
  not gc229 (wc229, n_3341);
  or g3824 (n_3434, wc230, n_2977);
  not gc230 (wc230, n_3432);
  or g3825 (n_3439, wc231, n_2989);
  not gc231 (wc231, n_3437);
  or g3826 (n_3441, wc232, n_2995);
  not gc232 (wc232, n_3382);
  or g3827 (n_3446, wc233, n_3007);
  not gc233 (wc233, n_3356);
  or g3828 (n_3456, wc234, n_3031);
  not gc234 (wc234, n_3341);
  or g3829 (n_3363, wc235, n_3290);
  not gc235 (wc235, n_3361);
  or g3830 (n_3365, wc236, n_3296);
  not gc236 (wc236, n_3344);
  or g3831 (n_3444, wc237, n_3001);
  not gc237 (wc237, n_3442);
  or g3832 (n_3449, wc238, n_3013);
  not gc238 (wc238, n_3447);
  or g3833 (n_3451, wc239, n_3019);
  not gc239 (wc239, n_3385);
  or g3834 (n_3459, wc240, n_3037);
  not gc240 (wc240, n_3457);
  or g3835 (n_3461, wc241, n_3043);
  not gc241 (wc241, n_3388);
  or g3836 (n_3466, wc242, n_3055);
  not gc242 (wc242, n_3361);
  or g3837 (n_3476, wc243, n_3079);
  not gc243 (wc243, n_3344);
  or g3838 (n_3370, wc244, n_3366);
  not gc244 (wc244, n_3367);
  or g3839 (n_3454, wc245, n_3025);
  not gc245 (wc245, n_3452);
  or g3840 (n_3464, wc246, n_3049);
  not gc246 (wc246, n_3462);
  or g3841 (n_3469, wc247, n_3061);
  not gc247 (wc247, n_3467);
  or g3842 (n_3471, wc248, n_3067);
  not gc248 (wc248, n_3391);
  or g3843 (n_3479, wc249, n_3085);
  not gc249 (wc249, n_3477);
  or g3844 (n_3481, wc250, n_3091);
  not gc250 (wc250, n_3394);
  or g3845 (n_3486, wc251, n_3103);
  not gc251 (wc251, n_3367);
  or g3846 (n_3474, wc252, n_3073);
  not gc252 (wc252, n_3472);
  or g3847 (n_3484, wc253, n_3097);
  not gc253 (wc253, n_3482);
  or g3848 (n_3489, wc254, n_3109);
  not gc254 (wc254, n_3487);
  or g3849 (n_3491, n_3113, wc255);
  not gc255 (wc255, n_3397);
  not g3850 (Z[77], n_3643);
endmodule

module mult_signed_const_13758_GENERIC(A, Z);
  input [58:0] A;
  output [77:0] Z;
  wire [58:0] A;
  wire [77:0] Z;
  mult_signed_const_13758_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_14241_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [60:0] A;
  output [79:0] Z;
  wire [60:0] A;
  wire [79:0] Z;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112;
  wire n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120;
  wire n_121, n_122, n_123, n_124, n_125, n_126, n_127, n_128;
  wire n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136;
  wire n_137, n_138, n_139, n_140, n_141, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381;
  wire n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389;
  wire n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397;
  wire n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405;
  wire n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413;
  wire n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421;
  wire n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429;
  wire n_430, n_431, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502;
  wire n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510;
  wire n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518;
  wire n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526;
  wire n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550;
  wire n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558;
  wire n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566;
  wire n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574;
  wire n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582;
  wire n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590;
  wire n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598;
  wire n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606;
  wire n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614;
  wire n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622;
  wire n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630;
  wire n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638;
  wire n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646;
  wire n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654;
  wire n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662;
  wire n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670;
  wire n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678;
  wire n_679, n_680, n_681, n_682, n_683, n_684, n_685, n_686;
  wire n_687, n_688, n_689, n_690, n_691, n_692, n_693, n_694;
  wire n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702;
  wire n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710;
  wire n_711, n_712, n_713, n_714, n_715, n_716, n_717, n_718;
  wire n_719, n_720, n_721, n_722, n_723, n_724, n_725, n_726;
  wire n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734;
  wire n_735, n_736, n_737, n_738, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758;
  wire n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766;
  wire n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774;
  wire n_775, n_776, n_777, n_778, n_779, n_780, n_781, n_782;
  wire n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790;
  wire n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798;
  wire n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806;
  wire n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_814;
  wire n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822;
  wire n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830;
  wire n_831, n_832, n_833, n_834, n_835, n_836, n_837, n_838;
  wire n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846;
  wire n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854;
  wire n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862;
  wire n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870;
  wire n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878;
  wire n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886;
  wire n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894;
  wire n_895, n_896, n_897, n_898, n_899, n_900, n_901, n_902;
  wire n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_911;
  wire n_912, n_913, n_914, n_915, n_916, n_917, n_918, n_919;
  wire n_920, n_921, n_922, n_925, n_926, n_927, n_928, n_929;
  wire n_930, n_931, n_932, n_933, n_934, n_935, n_937, n_938;
  wire n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946;
  wire n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954;
  wire n_955, n_956, n_957, n_958, n_959, n_960, n_963, n_964;
  wire n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972;
  wire n_973, n_974, n_975, n_976, n_980, n_981, n_982, n_983;
  wire n_984, n_986, n_987, n_988, n_989, n_990, n_991, n_992;
  wire n_993, n_995, n_996, n_997, n_1000, n_1001, n_1002, n_1003;
  wire n_1004, n_1005, n_1006, n_1007, n_1008, n_1011, n_1012, n_1015;
  wire n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023;
  wire n_1026, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034;
  wire n_1035, n_1036, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044;
  wire n_1045, n_1046, n_1047, n_1048, n_1049, n_1051, n_1052, n_1054;
  wire n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1065, n_1066;
  wire n_1067, n_1068, n_1069, n_1070, n_1071, n_1073, n_1076, n_1077;
  wire n_1078, n_1079, n_1080, n_1086, n_1087, n_1088, n_1089, n_1093;
  wire n_1094, n_1095, n_1096, n_1100, n_1101, n_1102, n_1103, n_1105;
  wire n_1107, n_1108, n_1112, n_1113, n_1115, n_1116, n_1119, n_1122;
  wire n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130;
  wire n_1131, n_1132, n_1134, n_1135, n_1136, n_1137, n_1141, n_1142;
  wire n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1150, n_1152;
  wire n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1160, n_1162;
  wire n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1172;
  wire n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181;
  wire n_1182, n_1183, n_1184, n_1185, n_1188, n_1192, n_1193, n_1194;
  wire n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202;
  wire n_1203, n_1206, n_1207, n_1208, n_1210, n_1211, n_1212, n_1213;
  wire n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221;
  wire n_1222, n_1223, n_1224, n_1226, n_1227, n_1229, n_1230, n_1231;
  wire n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239;
  wire n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247;
  wire n_1249, n_1250, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257;
  wire n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265;
  wire n_1266, n_1269, n_1270, n_1271, n_1272, n_1274, n_1275, n_1276;
  wire n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284;
  wire n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292;
  wire n_1298, n_1299, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307;
  wire n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315;
  wire n_1316, n_1317, n_1318, n_1319, n_1321, n_1322, n_1324, n_1325;
  wire n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335;
  wire n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343;
  wire n_1344, n_1345, n_1346, n_1347, n_1348, n_1352, n_1353, n_1354;
  wire n_1355, n_1356, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363;
  wire n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371;
  wire n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379;
  wire n_1380, n_1381, n_1386, n_1387, n_1388, n_1390, n_1391, n_1392;
  wire n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400;
  wire n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408;
  wire n_1409, n_1410, n_1411, n_1412, n_1413, n_1418, n_1420, n_1422;
  wire n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430;
  wire n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438;
  wire n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1448;
  wire n_1449, n_1450, n_1451, n_1452, n_1454, n_1455, n_1456, n_1457;
  wire n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465;
  wire n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473;
  wire n_1474, n_1475, n_1476, n_1477, n_1480, n_1482, n_1483, n_1486;
  wire n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494;
  wire n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502;
  wire n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1512;
  wire n_1514, n_1515, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523;
  wire n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531;
  wire n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539;
  wire n_1540, n_1541, n_1542, n_1544, n_1546, n_1547, n_1550, n_1551;
  wire n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559;
  wire n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567;
  wire n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1576, n_1578;
  wire n_1579, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588;
  wire n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596;
  wire n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604;
  wire n_1605, n_1606, n_1607, n_1608, n_1610, n_1611, n_1614, n_1615;
  wire n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623;
  wire n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631;
  wire n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1640, n_1642;
  wire n_1643, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652;
  wire n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660;
  wire n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668;
  wire n_1669, n_1670, n_1672, n_1674, n_1675, n_1678, n_1679, n_1680;
  wire n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688;
  wire n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696;
  wire n_1697, n_1698, n_1699, n_1700, n_1701, n_1704, n_1706, n_1707;
  wire n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717;
  wire n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725;
  wire n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733;
  wire n_1734, n_1736, n_1738, n_1739, n_1742, n_1743, n_1744, n_1745;
  wire n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753;
  wire n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761;
  wire n_1762, n_1763, n_1764, n_1765, n_1768, n_1770, n_1771, n_1774;
  wire n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782;
  wire n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790;
  wire n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798;
  wire n_1799, n_1800, n_1802, n_1803, n_1806, n_1807, n_1808, n_1809;
  wire n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817;
  wire n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825;
  wire n_1826, n_1827, n_1828, n_1829, n_1832, n_1834, n_1835, n_1838;
  wire n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846;
  wire n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854;
  wire n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1864;
  wire n_1866, n_1867, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875;
  wire n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883;
  wire n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891;
  wire n_1892, n_1893, n_1896, n_1898, n_1899, n_1902, n_1903, n_1904;
  wire n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912;
  wire n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920;
  wire n_1921, n_1922, n_1923, n_1924, n_1925, n_1928, n_1930, n_1931;
  wire n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941;
  wire n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949;
  wire n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957;
  wire n_1960, n_1962, n_1963, n_1966, n_1967, n_1968, n_1969, n_1970;
  wire n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978;
  wire n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986;
  wire n_1987, n_1988, n_1989, n_1992, n_1994, n_1995, n_1998, n_1999;
  wire n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007;
  wire n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015;
  wire n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2024, n_2026;
  wire n_2027, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036;
  wire n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044;
  wire n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052;
  wire n_2053, n_2056, n_2058, n_2059, n_2062, n_2063, n_2064, n_2065;
  wire n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073;
  wire n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081;
  wire n_2082, n_2083, n_2084, n_2085, n_2088, n_2090, n_2091, n_2094;
  wire n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102;
  wire n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110;
  wire n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2120;
  wire n_2122, n_2123, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131;
  wire n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139;
  wire n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147;
  wire n_2148, n_2149, n_2152, n_2154, n_2155, n_2158, n_2159, n_2160;
  wire n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168;
  wire n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176;
  wire n_2177, n_2178, n_2179, n_2180, n_2181, n_2184, n_2186, n_2187;
  wire n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197;
  wire n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205;
  wire n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213;
  wire n_2216, n_2218, n_2219, n_2222, n_2223, n_2224, n_2225, n_2226;
  wire n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234;
  wire n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242;
  wire n_2243, n_2244, n_2245, n_2248, n_2250, n_2251, n_2254, n_2255;
  wire n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263;
  wire n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271;
  wire n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279;
  wire n_2280, n_2282, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290;
  wire n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298;
  wire n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306;
  wire n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2314, n_2317;
  wire n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325;
  wire n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333;
  wire n_2334, n_2335, n_2336, n_2337, n_2341, n_2342, n_2344, n_2348;
  wire n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356;
  wire n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364;
  wire n_2365, n_2366, n_2367, n_2368, n_2369, n_2373, n_2374, n_2376;
  wire n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387;
  wire n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395;
  wire n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2405, n_2410;
  wire n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418;
  wire n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426;
  wire n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2437;
  wire n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449;
  wire n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457;
  wire n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465;
  wire n_2466, n_2470, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479;
  wire n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487;
  wire n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495;
  wire n_2496, n_2497, n_2498, n_2502, n_2506, n_2507, n_2508, n_2509;
  wire n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517;
  wire n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525;
  wire n_2526, n_2527, n_2528, n_2529, n_2536, n_2537, n_2542, n_2543;
  wire n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551;
  wire n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559;
  wire n_2560, n_2561, n_2568, n_2569, n_2574, n_2575, n_2576, n_2577;
  wire n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585;
  wire n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593;
  wire n_2598, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606;
  wire n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614;
  wire n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622;
  wire n_2623, n_2624, n_2625, n_2630, n_2632, n_2633, n_2634, n_2635;
  wire n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643;
  wire n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, n_2651;
  wire n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659;
  wire n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2668, n_2670;
  wire n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678;
  wire n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686;
  wire n_2687, n_2688, n_2689, n_2692, n_2693, n_2694, n_2695, n_2697;
  wire n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709;
  wire n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717;
  wire n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2725, n_2726;
  wire n_2727, n_2729, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739;
  wire n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747;
  wire n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2762;
  wire n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770;
  wire n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778;
  wire n_2779, n_2780, n_2781, n_2784, n_2786, n_2789, n_2790, n_2792;
  wire n_2793, n_2794, n_2795, n_2796, n_2798, n_2799, n_2800, n_2801;
  wire n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809;
  wire n_2810, n_2813, n_2814, n_2817, n_2818, n_2819, n_2820, n_2821;
  wire n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829;
  wire n_2830, n_2831, n_2832, n_2833, n_2834, n_2842, n_2844, n_2845;
  wire n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853;
  wire n_2854, n_2855, n_2856, n_2857, n_2858, n_2861, n_2864, n_2865;
  wire n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875;
  wire n_2876, n_2877, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891;
  wire n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2904, n_2906;
  wire n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2920, n_2921;
  wire n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929;
  wire n_2932, n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940;
  wire n_2941, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952;
  wire n_2953, n_2954, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961;
  wire n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971;
  wire n_2972, n_2973, n_2976, n_2977, n_2989, n_2991, n_2993, n_2994;
  wire n_2995, n_2996, n_2997, n_2999, n_3000, n_3001, n_3002, n_3003;
  wire n_3005, n_3006, n_3007, n_3008, n_3009, n_3011, n_3012, n_3013;
  wire n_3014, n_3015, n_3017, n_3018, n_3019, n_3020, n_3021, n_3023;
  wire n_3024, n_3025, n_3026, n_3027, n_3029, n_3030, n_3031, n_3032;
  wire n_3033, n_3035, n_3036, n_3037, n_3038, n_3039, n_3041, n_3042;
  wire n_3043, n_3044, n_3045, n_3047, n_3048, n_3049, n_3050, n_3051;
  wire n_3053, n_3054, n_3055, n_3056, n_3057, n_3059, n_3060, n_3061;
  wire n_3062, n_3063, n_3065, n_3066, n_3067, n_3068, n_3069, n_3071;
  wire n_3072, n_3073, n_3074, n_3075, n_3077, n_3078, n_3079, n_3080;
  wire n_3081, n_3083, n_3084, n_3085, n_3086, n_3087, n_3089, n_3090;
  wire n_3091, n_3092, n_3093, n_3095, n_3096, n_3097, n_3098, n_3099;
  wire n_3101, n_3102, n_3103, n_3104, n_3105, n_3107, n_3108, n_3109;
  wire n_3110, n_3111, n_3113, n_3114, n_3115, n_3116, n_3117, n_3119;
  wire n_3120, n_3121, n_3122, n_3123, n_3125, n_3126, n_3127, n_3128;
  wire n_3129, n_3131, n_3132, n_3133, n_3134, n_3135, n_3137, n_3138;
  wire n_3139, n_3140, n_3141, n_3143, n_3144, n_3145, n_3146, n_3147;
  wire n_3149, n_3150, n_3151, n_3152, n_3153, n_3155, n_3156, n_3157;
  wire n_3158, n_3159, n_3161, n_3162, n_3163, n_3164, n_3165, n_3167;
  wire n_3168, n_3169, n_3170, n_3171, n_3173, n_3174, n_3175, n_3176;
  wire n_3177, n_3179, n_3180, n_3181, n_3182, n_3183, n_3185, n_3186;
  wire n_3187, n_3188, n_3189, n_3191, n_3192, n_3193, n_3194, n_3195;
  wire n_3197, n_3198, n_3199, n_3200, n_3201, n_3203, n_3204, n_3205;
  wire n_3206, n_3207, n_3209, n_3210, n_3211, n_3212, n_3213, n_3215;
  wire n_3216, n_3219, n_3222, n_3224, n_3225, n_3227, n_3228, n_3230;
  wire n_3231, n_3232, n_3234, n_3235, n_3237, n_3238, n_3239, n_3241;
  wire n_3242, n_3244, n_3245, n_3246, n_3248, n_3249, n_3251, n_3252;
  wire n_3253, n_3255, n_3256, n_3258, n_3259, n_3260, n_3262, n_3263;
  wire n_3265, n_3266, n_3267, n_3269, n_3270, n_3272, n_3273, n_3274;
  wire n_3276, n_3277, n_3279, n_3280, n_3281, n_3283, n_3284, n_3286;
  wire n_3287, n_3288, n_3290, n_3291, n_3293, n_3294, n_3295, n_3297;
  wire n_3298, n_3300, n_3301, n_3302, n_3304, n_3305, n_3307, n_3308;
  wire n_3309, n_3311, n_3312, n_3314, n_3315, n_3316, n_3318, n_3319;
  wire n_3321, n_3322, n_3323, n_3325, n_3326, n_3328, n_3329, n_3330;
  wire n_3332, n_3333, n_3335, n_3336, n_3337, n_3339, n_3340, n_3342;
  wire n_3343, n_3344, n_3346, n_3347, n_3349, n_3350, n_3351, n_3352;
  wire n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3362, n_3363;
  wire n_3364, n_3365, n_3366, n_3368, n_3369, n_3370, n_3371, n_3372;
  wire n_3374, n_3375, n_3376, n_3377, n_3378, n_3380, n_3381, n_3382;
  wire n_3383, n_3384, n_3386, n_3387, n_3388, n_3389, n_3390, n_3392;
  wire n_3393, n_3394, n_3395, n_3396, n_3398, n_3399, n_3400, n_3401;
  wire n_3402, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410;
  wire n_3411, n_3412, n_3414, n_3415, n_3417, n_3418, n_3419, n_3421;
  wire n_3422, n_3424, n_3425, n_3426, n_3428, n_3429, n_3431, n_3432;
  wire n_3433, n_3434, n_3435, n_3437, n_3438, n_3439, n_3440, n_3441;
  wire n_3442, n_3444, n_3445, n_3446, n_3447, n_3448, n_3450, n_3451;
  wire n_3452, n_3453, n_3454, n_3455, n_3456, n_3458, n_3460, n_3461;
  wire n_3463, n_3465, n_3466, n_3468, n_3470, n_3471, n_3473, n_3475;
  wire n_3476, n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484;
  wire n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492;
  wire n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500;
  wire n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3510, n_3511;
  wire n_3513, n_3515, n_3516, n_3518, n_3520, n_3521, n_3523, n_3525;
  wire n_3526, n_3528, n_3530, n_3531, n_3533, n_3535, n_3536, n_3538;
  wire n_3540, n_3541, n_3543, n_3545, n_3546, n_3548, n_3550, n_3551;
  wire n_3553, n_3555, n_3556, n_3558, n_3560, n_3561, n_3563, n_3565;
  wire n_3566, n_3568, n_3570, n_3571, n_3573, n_3575, n_3576, n_3578;
  wire n_3580, n_3581, n_3583, n_3585, n_3586, n_3588, n_3590, n_3591;
  wire n_3593, n_3595, n_3596, n_3598, n_3600, n_3601, n_3603, n_3605;
  wire n_3608, n_3609, n_3611, n_3612, n_3613, n_3615, n_3616, n_3617;
  wire n_3619, n_3620, n_3621, n_3623, n_3624, n_3625, n_3627, n_3628;
  wire n_3629, n_3631, n_3632, n_3633, n_3635, n_3636, n_3637, n_3639;
  wire n_3640, n_3641, n_3643, n_3644, n_3645, n_3647, n_3648, n_3649;
  wire n_3651, n_3652, n_3653, n_3655, n_3656, n_3657, n_3659, n_3660;
  wire n_3661, n_3663, n_3664, n_3665, n_3667, n_3668, n_3669, n_3671;
  wire n_3672, n_3673, n_3675, n_3676, n_3677, n_3679, n_3680, n_3681;
  wire n_3683, n_3684, n_3685, n_3687, n_3688, n_3689, n_3691, n_3692;
  wire n_3693, n_3695, n_3696, n_3697, n_3699, n_3700, n_3701, n_3703;
  wire n_3704, n_3705, n_3707, n_3708, n_3709, n_3711, n_3712, n_3713;
  wire n_3715, n_3716, n_3717, n_3719, n_3720, n_3721, n_3723, n_3724;
  wire n_3725, n_3727, n_3728, n_3729, n_3731, n_3732, n_3733, n_3735;
  wire n_3736, n_3737, n_3739, n_3740, n_3741, n_3743, n_3744, n_3745;
  wire n_3747, n_3748, n_3749, n_3751, n_3752, n_3753, n_3755, n_3756;
  wire n_3757, n_3759;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g484 (n_217, A[4], A[0]);
  and g2 (n_136, A[4], A[0]);
  xor g485 (n_1122, A[1], A[3]);
  xor g486 (n_216, n_1122, A[5]);
  nand g3 (n_1123, A[1], A[3]);
  nand g487 (n_1124, A[5], A[3]);
  nand g488 (n_1125, A[1], A[5]);
  nand g489 (n_135, n_1123, n_1124, n_1125);
  xor g490 (n_303, A[6], A[4]);
  and g491 (n_304, A[6], A[4]);
  xor g492 (n_1126, A[0], A[2]);
  xor g493 (n_215, n_1126, n_303);
  nand g494 (n_1127, A[0], A[2]);
  nand g4 (n_1128, n_303, A[2]);
  nand g5 (n_1129, A[0], n_303);
  nand g495 (n_134, n_1127, n_1128, n_1129);
  xor g496 (n_1130, A[1], A[7]);
  xor g497 (n_305, n_1130, A[5]);
  nand g498 (n_1131, A[1], A[7]);
  nand g499 (n_1132, A[5], A[7]);
  nand g6 (n_307, n_1131, n_1132, n_1125);
  xor g501 (n_1134, A[3], n_304);
  xor g502 (n_214, n_1134, n_305);
  nand g503 (n_1135, A[3], n_304);
  nand g504 (n_1136, n_305, n_304);
  nand g505 (n_1137, A[3], n_305);
  nand g506 (n_133, n_1135, n_1136, n_1137);
  xor g507 (n_306, A[8], A[6]);
  and g508 (n_309, A[8], A[6]);
  xor g510 (n_308, n_1126, A[4]);
  nand g513 (n_1141, A[2], A[4]);
  xor g515 (n_1142, n_306, n_307);
  xor g516 (n_213, n_1142, n_308);
  nand g517 (n_1143, n_306, n_307);
  nand g518 (n_1144, n_308, n_307);
  nand g519 (n_1145, n_306, n_308);
  nand g520 (n_132, n_1143, n_1144, n_1145);
  xor g521 (n_1146, A[1], A[9]);
  xor g522 (n_311, n_1146, A[3]);
  nand g523 (n_1147, A[1], A[9]);
  nand g524 (n_1148, A[3], A[9]);
  nand g526 (n_314, n_1147, n_1148, n_1123);
  xor g527 (n_1150, A[7], A[5]);
  xor g528 (n_312, n_1150, n_309);
  nand g530 (n_1152, n_309, A[5]);
  nand g531 (n_1153, A[7], n_309);
  nand g532 (n_316, n_1132, n_1152, n_1153);
  xor g533 (n_1154, n_310, n_311);
  xor g534 (n_212, n_1154, n_312);
  nand g535 (n_1155, n_310, n_311);
  nand g536 (n_1156, n_312, n_311);
  nand g537 (n_1157, n_310, n_312);
  nand g538 (n_131, n_1155, n_1156, n_1157);
  xor g539 (n_313, A[10], A[8]);
  and g540 (n_318, A[10], A[8]);
  xor g541 (n_1158, A[4], A[2]);
  xor g542 (n_315, n_1158, A[6]);
  nand g544 (n_1160, A[6], A[2]);
  xor g547 (n_1162, A[0], n_313);
  xor g548 (n_317, n_1162, n_314);
  nand g549 (n_1163, A[0], n_313);
  nand g550 (n_1164, n_314, n_313);
  nand g551 (n_1165, A[0], n_314);
  nand g552 (n_322, n_1163, n_1164, n_1165);
  xor g553 (n_1166, n_315, n_316);
  xor g554 (n_211, n_1166, n_317);
  nand g555 (n_1167, n_315, n_316);
  nand g556 (n_1168, n_317, n_316);
  nand g557 (n_1169, n_315, n_317);
  nand g558 (n_130, n_1167, n_1168, n_1169);
  xor g560 (n_320, n_1146, A[5]);
  nand g562 (n_1172, A[5], A[9]);
  nand g564 (n_325, n_1147, n_1172, n_1125);
  xor g565 (n_1174, A[3], A[11]);
  xor g566 (n_321, n_1174, A[7]);
  nand g567 (n_1175, A[3], A[11]);
  nand g568 (n_1176, A[7], A[11]);
  nand g569 (n_1177, A[3], A[7]);
  nand g570 (n_326, n_1175, n_1176, n_1177);
  xor g571 (n_1178, n_318, n_319);
  xor g572 (n_323, n_1178, n_320);
  nand g573 (n_1179, n_318, n_319);
  nand g574 (n_1180, n_320, n_319);
  nand g575 (n_1181, n_318, n_320);
  nand g576 (n_330, n_1179, n_1180, n_1181);
  xor g577 (n_1182, n_321, n_322);
  xor g578 (n_210, n_1182, n_323);
  nand g579 (n_1183, n_321, n_322);
  nand g580 (n_1184, n_323, n_322);
  nand g581 (n_1185, n_321, n_323);
  nand g582 (n_129, n_1183, n_1184, n_1185);
  xor g583 (n_324, A[12], A[10]);
  and g584 (n_331, A[12], A[10]);
  xor g586 (n_327, n_303, A[8]);
  nand g588 (n_1188, A[8], A[4]);
  xor g592 (n_328, n_1126, n_324);
  nand g594 (n_1192, n_324, A[0]);
  nand g595 (n_1193, A[2], n_324);
  nand g596 (n_335, n_1127, n_1192, n_1193);
  xor g597 (n_1194, n_325, n_326);
  xor g598 (n_329, n_1194, n_327);
  nand g599 (n_1195, n_325, n_326);
  nand g600 (n_1196, n_327, n_326);
  nand g601 (n_1197, n_325, n_327);
  nand g602 (n_337, n_1195, n_1196, n_1197);
  xor g603 (n_1198, n_328, n_329);
  xor g604 (n_209, n_1198, n_330);
  nand g605 (n_1199, n_328, n_329);
  nand g606 (n_1200, n_330, n_329);
  nand g607 (n_1201, n_328, n_330);
  nand g608 (n_128, n_1199, n_1200, n_1201);
  xor g609 (n_1202, A[1], A[11]);
  xor g610 (n_334, n_1202, A[7]);
  nand g611 (n_1203, A[1], A[11]);
  nand g614 (n_340, n_1203, n_1176, n_1131);
  xor g615 (n_1206, A[5], A[13]);
  xor g616 (n_333, n_1206, A[3]);
  nand g617 (n_1207, A[5], A[13]);
  nand g618 (n_1208, A[3], A[13]);
  nand g620 (n_341, n_1207, n_1208, n_1124);
  xor g621 (n_1210, A[9], n_331);
  xor g622 (n_336, n_1210, n_332);
  nand g623 (n_1211, A[9], n_331);
  nand g624 (n_1212, n_332, n_331);
  nand g625 (n_1213, A[9], n_332);
  nand g626 (n_344, n_1211, n_1212, n_1213);
  xor g627 (n_1214, n_333, n_334);
  xor g628 (n_338, n_1214, n_335);
  nand g629 (n_1215, n_333, n_334);
  nand g630 (n_1216, n_335, n_334);
  nand g631 (n_1217, n_333, n_335);
  nand g632 (n_346, n_1215, n_1216, n_1217);
  xor g633 (n_1218, n_336, n_337);
  xor g634 (n_208, n_1218, n_338);
  nand g635 (n_1219, n_336, n_337);
  nand g636 (n_1220, n_338, n_337);
  nand g637 (n_1221, n_336, n_338);
  nand g638 (n_127, n_1219, n_1220, n_1221);
  xor g639 (n_339, A[14], A[12]);
  and g640 (n_348, A[14], A[12]);
  xor g641 (n_1222, A[8], A[0]);
  xor g642 (n_343, n_1222, A[6]);
  nand g643 (n_1223, A[8], A[0]);
  nand g644 (n_1224, A[6], A[0]);
  xor g647 (n_1226, A[10], A[4]);
  xor g648 (n_342, n_1226, A[2]);
  nand g649 (n_1227, A[10], A[4]);
  nand g651 (n_1229, A[10], A[2]);
  nand g652 (n_350, n_1227, n_1141, n_1229);
  xor g653 (n_1230, n_339, n_340);
  xor g654 (n_345, n_1230, n_341);
  nand g655 (n_1231, n_339, n_340);
  nand g656 (n_1232, n_341, n_340);
  nand g657 (n_1233, n_339, n_341);
  nand g658 (n_354, n_1231, n_1232, n_1233);
  xor g659 (n_1234, n_342, n_343);
  xor g660 (n_347, n_1234, n_344);
  nand g661 (n_1235, n_342, n_343);
  nand g662 (n_1236, n_344, n_343);
  nand g663 (n_1237, n_342, n_344);
  nand g664 (n_357, n_1235, n_1236, n_1237);
  xor g665 (n_1238, n_345, n_346);
  xor g666 (n_207, n_1238, n_347);
  nand g667 (n_1239, n_345, n_346);
  nand g668 (n_1240, n_347, n_346);
  nand g669 (n_1241, n_345, n_347);
  nand g670 (n_126, n_1239, n_1240, n_1241);
  xor g671 (n_1242, A[1], A[15]);
  xor g672 (n_351, n_1242, A[13]);
  nand g673 (n_1243, A[1], A[15]);
  nand g674 (n_1244, A[13], A[15]);
  nand g675 (n_1245, A[1], A[13]);
  nand g676 (n_359, n_1243, n_1244, n_1245);
  xor g677 (n_1246, A[9], A[7]);
  xor g678 (n_352, n_1246, A[11]);
  nand g679 (n_1247, A[9], A[7]);
  nand g681 (n_1249, A[9], A[11]);
  nand g682 (n_360, n_1247, n_1176, n_1249);
  xor g683 (n_1250, A[5], A[3]);
  xor g684 (n_353, n_1250, n_348);
  nand g686 (n_1252, n_348, A[3]);
  nand g687 (n_1253, A[5], n_348);
  nand g688 (n_363, n_1124, n_1252, n_1253);
  xor g689 (n_1254, n_349, n_350);
  xor g690 (n_355, n_1254, n_351);
  nand g691 (n_1255, n_349, n_350);
  nand g692 (n_1256, n_351, n_350);
  nand g693 (n_1257, n_349, n_351);
  nand g694 (n_365, n_1255, n_1256, n_1257);
  xor g695 (n_1258, n_352, n_353);
  xor g696 (n_356, n_1258, n_354);
  nand g697 (n_1259, n_352, n_353);
  nand g698 (n_1260, n_354, n_353);
  nand g699 (n_1261, n_352, n_354);
  nand g700 (n_367, n_1259, n_1260, n_1261);
  xor g701 (n_1262, n_355, n_356);
  xor g702 (n_206, n_1262, n_357);
  nand g703 (n_1263, n_355, n_356);
  nand g704 (n_1264, n_357, n_356);
  nand g705 (n_1265, n_355, n_357);
  nand g706 (n_125, n_1263, n_1264, n_1265);
  xor g707 (n_358, A[16], A[14]);
  and g708 (n_369, A[16], A[14]);
  xor g709 (n_1266, A[10], A[2]);
  xor g710 (n_362, n_1266, A[0]);
  nand g713 (n_1269, A[10], A[0]);
  nand g714 (n_370, n_1229, n_1127, n_1269);
  xor g715 (n_1270, A[8], A[12]);
  xor g716 (n_361, n_1270, A[6]);
  nand g717 (n_1271, A[8], A[12]);
  nand g718 (n_1272, A[6], A[12]);
  xor g721 (n_1274, A[4], n_358);
  xor g722 (n_364, n_1274, n_359);
  nand g723 (n_1275, A[4], n_358);
  nand g724 (n_1276, n_359, n_358);
  nand g725 (n_1277, A[4], n_359);
  nand g726 (n_375, n_1275, n_1276, n_1277);
  xor g727 (n_1278, n_360, n_361);
  xor g728 (n_366, n_1278, n_362);
  nand g729 (n_1279, n_360, n_361);
  nand g730 (n_1280, n_362, n_361);
  nand g731 (n_1281, n_360, n_362);
  nand g732 (n_377, n_1279, n_1280, n_1281);
  xor g733 (n_1282, n_363, n_364);
  xor g734 (n_368, n_1282, n_365);
  nand g735 (n_1283, n_363, n_364);
  nand g736 (n_1284, n_365, n_364);
  nand g737 (n_1285, n_363, n_365);
  nand g738 (n_379, n_1283, n_1284, n_1285);
  xor g739 (n_1286, n_366, n_367);
  xor g740 (n_205, n_1286, n_368);
  nand g741 (n_1287, n_366, n_367);
  nand g742 (n_1288, n_368, n_367);
  nand g743 (n_1289, n_366, n_368);
  nand g744 (n_124, n_1287, n_1288, n_1289);
  xor g745 (n_1290, A[1], A[17]);
  xor g746 (n_373, n_1290, A[15]);
  nand g747 (n_1291, A[1], A[17]);
  nand g748 (n_1292, A[15], A[17]);
  nand g750 (n_382, n_1291, n_1292, n_1243);
  xor g752 (n_374, n_1174, A[9]);
  nand g756 (n_384, n_1175, n_1249, n_1148);
  xor g757 (n_1298, A[13], A[7]);
  xor g758 (n_372, n_1298, A[5]);
  nand g759 (n_1299, A[13], A[7]);
  nand g762 (n_383, n_1299, n_1132, n_1207);
  xor g763 (n_1302, n_369, n_370);
  xor g764 (n_376, n_1302, n_371);
  nand g765 (n_1303, n_369, n_370);
  nand g766 (n_1304, n_371, n_370);
  nand g767 (n_1305, n_369, n_371);
  nand g768 (n_388, n_1303, n_1304, n_1305);
  xor g769 (n_1306, n_372, n_373);
  xor g770 (n_378, n_1306, n_374);
  nand g771 (n_1307, n_372, n_373);
  nand g772 (n_1308, n_374, n_373);
  nand g773 (n_1309, n_372, n_374);
  nand g774 (n_390, n_1307, n_1308, n_1309);
  xor g775 (n_1310, n_375, n_376);
  xor g776 (n_380, n_1310, n_377);
  nand g777 (n_1311, n_375, n_376);
  nand g778 (n_1312, n_377, n_376);
  nand g779 (n_1313, n_375, n_377);
  nand g780 (n_392, n_1311, n_1312, n_1313);
  xor g781 (n_1314, n_378, n_379);
  xor g782 (n_204, n_1314, n_380);
  nand g783 (n_1315, n_378, n_379);
  nand g784 (n_1316, n_380, n_379);
  nand g785 (n_1317, n_378, n_380);
  nand g786 (n_123, n_1315, n_1316, n_1317);
  xor g787 (n_381, A[18], A[16]);
  and g788 (n_394, A[18], A[16]);
  xor g789 (n_1318, A[12], A[4]);
  xor g790 (n_385, n_1318, A[2]);
  nand g791 (n_1319, A[12], A[4]);
  nand g793 (n_1321, A[12], A[2]);
  nand g794 (n_395, n_1319, n_1141, n_1321);
  xor g795 (n_1322, A[10], A[0]);
  xor g796 (n_386, n_1322, A[14]);
  nand g798 (n_1324, A[14], A[0]);
  nand g799 (n_1325, A[10], A[14]);
  nand g800 (n_396, n_1269, n_1324, n_1325);
  xor g802 (n_387, n_306, n_381);
  nand g804 (n_1328, n_381, A[6]);
  nand g805 (n_1329, A[8], n_381);
  xor g807 (n_1330, n_382, n_383);
  xor g808 (n_389, n_1330, n_384);
  nand g809 (n_1331, n_382, n_383);
  nand g810 (n_1332, n_384, n_383);
  nand g811 (n_1333, n_382, n_384);
  nand g812 (n_402, n_1331, n_1332, n_1333);
  xor g813 (n_1334, n_385, n_386);
  xor g814 (n_391, n_1334, n_387);
  nand g815 (n_1335, n_385, n_386);
  nand g816 (n_1336, n_387, n_386);
  nand g817 (n_1337, n_385, n_387);
  nand g818 (n_403, n_1335, n_1336, n_1337);
  xor g819 (n_1338, n_388, n_389);
  xor g820 (n_393, n_1338, n_390);
  nand g821 (n_1339, n_388, n_389);
  nand g822 (n_1340, n_390, n_389);
  nand g823 (n_1341, n_388, n_390);
  nand g824 (n_406, n_1339, n_1340, n_1341);
  xor g825 (n_1342, n_391, n_392);
  xor g826 (n_203, n_1342, n_393);
  nand g827 (n_1343, n_391, n_392);
  nand g828 (n_1344, n_393, n_392);
  nand g829 (n_1345, n_391, n_393);
  nand g830 (n_122, n_1343, n_1344, n_1345);
  xor g831 (n_1346, A[1], A[19]);
  xor g832 (n_398, n_1346, A[13]);
  nand g833 (n_1347, A[1], A[19]);
  nand g834 (n_1348, A[13], A[19]);
  nand g836 (n_408, n_1347, n_1348, n_1245);
  xor g838 (n_399, n_1250, A[17]);
  nand g840 (n_1352, A[17], A[3]);
  nand g841 (n_1353, A[5], A[17]);
  nand g842 (n_409, n_1124, n_1352, n_1353);
  xor g843 (n_1354, A[11], A[15]);
  xor g844 (n_397, n_1354, A[9]);
  nand g845 (n_1355, A[11], A[15]);
  nand g846 (n_1356, A[9], A[15]);
  nand g848 (n_410, n_1355, n_1356, n_1249);
  xor g849 (n_1358, A[7], n_394);
  xor g850 (n_401, n_1358, n_395);
  nand g851 (n_1359, A[7], n_394);
  nand g852 (n_1360, n_395, n_394);
  nand g853 (n_1361, A[7], n_395);
  nand g854 (n_414, n_1359, n_1360, n_1361);
  xor g855 (n_1362, n_396, n_397);
  xor g856 (n_404, n_1362, n_398);
  nand g857 (n_1363, n_396, n_397);
  nand g858 (n_1364, n_398, n_397);
  nand g859 (n_1365, n_396, n_398);
  nand g860 (n_416, n_1363, n_1364, n_1365);
  xor g861 (n_1366, n_399, n_400);
  xor g862 (n_405, n_1366, n_401);
  nand g863 (n_1367, n_399, n_400);
  nand g864 (n_1368, n_401, n_400);
  nand g865 (n_1369, n_399, n_401);
  nand g866 (n_138, n_1367, n_1368, n_1369);
  xor g867 (n_1370, n_402, n_403);
  xor g868 (n_407, n_1370, n_404);
  nand g869 (n_1371, n_402, n_403);
  nand g870 (n_1372, n_404, n_403);
  nand g871 (n_1373, n_402, n_404);
  nand g872 (n_140, n_1371, n_1372, n_1373);
  xor g873 (n_1374, n_405, n_406);
  xor g874 (n_202, n_1374, n_407);
  nand g875 (n_1375, n_405, n_406);
  nand g876 (n_1376, n_407, n_406);
  nand g877 (n_1377, n_405, n_407);
  nand g878 (n_121, n_1375, n_1376, n_1377);
  xor g879 (n_1378, A[20], A[18]);
  xor g880 (n_412, n_1378, A[14]);
  nand g881 (n_1379, A[20], A[18]);
  nand g882 (n_1380, A[14], A[18]);
  nand g883 (n_1381, A[20], A[14]);
  nand g884 (n_417, n_1379, n_1380, n_1381);
  xor g886 (n_413, n_303, A[12]);
  xor g891 (n_1386, A[2], A[16]);
  xor g892 (n_411, n_1386, A[10]);
  nand g893 (n_1387, A[2], A[16]);
  nand g894 (n_1388, A[10], A[16]);
  nand g896 (n_419, n_1387, n_1388, n_1229);
  xor g897 (n_1390, A[8], n_408);
  xor g898 (n_415, n_1390, n_409);
  nand g899 (n_1391, A[8], n_408);
  nand g900 (n_1392, n_409, n_408);
  nand g901 (n_1393, A[8], n_409);
  nand g902 (n_423, n_1391, n_1392, n_1393);
  xor g903 (n_1394, n_410, n_411);
  xor g904 (n_137, n_1394, n_412);
  nand g905 (n_1395, n_410, n_411);
  nand g906 (n_1396, n_412, n_411);
  nand g907 (n_1397, n_410, n_412);
  nand g908 (n_425, n_1395, n_1396, n_1397);
  xor g909 (n_1398, n_413, n_414);
  xor g910 (n_139, n_1398, n_415);
  nand g911 (n_1399, n_413, n_414);
  nand g912 (n_1400, n_415, n_414);
  nand g913 (n_1401, n_413, n_415);
  nand g914 (n_427, n_1399, n_1400, n_1401);
  xor g915 (n_1402, n_416, n_137);
  xor g916 (n_141, n_1402, n_138);
  nand g917 (n_1403, n_416, n_137);
  nand g918 (n_1404, n_138, n_137);
  nand g919 (n_1405, n_416, n_138);
  nand g920 (n_429, n_1403, n_1404, n_1405);
  xor g921 (n_1406, n_139, n_140);
  xor g922 (n_201, n_1406, n_141);
  nand g923 (n_1407, n_139, n_140);
  nand g924 (n_1408, n_141, n_140);
  nand g925 (n_1409, n_139, n_141);
  nand g926 (n_120, n_1407, n_1408, n_1409);
  xor g927 (n_1410, A[21], A[19]);
  xor g928 (n_421, n_1410, A[15]);
  nand g929 (n_1411, A[21], A[19]);
  nand g930 (n_1412, A[15], A[19]);
  nand g931 (n_1413, A[21], A[15]);
  nand g932 (n_431, n_1411, n_1412, n_1413);
  xor g934 (n_422, n_1150, A[13]);
  xor g939 (n_1418, A[3], A[17]);
  xor g940 (n_420, n_1418, A[11]);
  nand g942 (n_1420, A[11], A[17]);
  nand g944 (n_433, n_1352, n_1420, n_1175);
  xor g945 (n_1422, A[9], n_417);
  xor g946 (n_424, n_1422, n_418);
  nand g947 (n_1423, A[9], n_417);
  nand g948 (n_1424, n_418, n_417);
  nand g949 (n_1425, A[9], n_418);
  nand g950 (n_437, n_1423, n_1424, n_1425);
  xor g951 (n_1426, n_419, n_420);
  xor g952 (n_426, n_1426, n_421);
  nand g953 (n_1427, n_419, n_420);
  nand g954 (n_1428, n_421, n_420);
  nand g955 (n_1429, n_419, n_421);
  nand g956 (n_439, n_1427, n_1428, n_1429);
  xor g957 (n_1430, n_422, n_423);
  xor g958 (n_428, n_1430, n_424);
  nand g959 (n_1431, n_422, n_423);
  nand g960 (n_1432, n_424, n_423);
  nand g961 (n_1433, n_422, n_424);
  nand g962 (n_441, n_1431, n_1432, n_1433);
  xor g963 (n_1434, n_425, n_426);
  xor g964 (n_430, n_1434, n_427);
  nand g965 (n_1435, n_425, n_426);
  nand g966 (n_1436, n_427, n_426);
  nand g967 (n_1437, n_425, n_427);
  nand g968 (n_444, n_1435, n_1436, n_1437);
  xor g969 (n_1438, n_428, n_429);
  xor g970 (n_200, n_1438, n_430);
  nand g971 (n_1439, n_428, n_429);
  nand g972 (n_1440, n_430, n_429);
  nand g973 (n_1441, n_428, n_430);
  nand g974 (n_119, n_1439, n_1440, n_1441);
  xor g975 (n_1442, A[22], A[20]);
  xor g976 (n_435, n_1442, A[16]);
  nand g977 (n_1443, A[22], A[20]);
  nand g978 (n_1444, A[16], A[20]);
  nand g979 (n_1445, A[22], A[16]);
  nand g980 (n_445, n_1443, n_1444, n_1445);
  xor g982 (n_436, n_306, A[14]);
  nand g984 (n_1448, A[14], A[6]);
  nand g985 (n_1449, A[8], A[14]);
  xor g987 (n_1450, A[4], A[18]);
  xor g988 (n_434, n_1450, A[12]);
  nand g989 (n_1451, A[4], A[18]);
  nand g990 (n_1452, A[12], A[18]);
  nand g992 (n_447, n_1451, n_1452, n_1319);
  xor g993 (n_1454, A[10], n_431);
  xor g994 (n_438, n_1454, n_383);
  nand g995 (n_1455, A[10], n_431);
  nand g996 (n_1456, n_383, n_431);
  nand g997 (n_1457, A[10], n_383);
  nand g998 (n_451, n_1455, n_1456, n_1457);
  xor g999 (n_1458, n_433, n_434);
  xor g1000 (n_440, n_1458, n_435);
  nand g1001 (n_1459, n_433, n_434);
  nand g1002 (n_1460, n_435, n_434);
  nand g1003 (n_1461, n_433, n_435);
  nand g1004 (n_453, n_1459, n_1460, n_1461);
  xor g1005 (n_1462, n_436, n_437);
  xor g1006 (n_442, n_1462, n_438);
  nand g1007 (n_1463, n_436, n_437);
  nand g1008 (n_1464, n_438, n_437);
  nand g1009 (n_1465, n_436, n_438);
  nand g1010 (n_455, n_1463, n_1464, n_1465);
  xor g1011 (n_1466, n_439, n_440);
  xor g1012 (n_443, n_1466, n_441);
  nand g1013 (n_1467, n_439, n_440);
  nand g1014 (n_1468, n_441, n_440);
  nand g1015 (n_1469, n_439, n_441);
  nand g1016 (n_458, n_1467, n_1468, n_1469);
  xor g1017 (n_1470, n_442, n_443);
  xor g1018 (n_199, n_1470, n_444);
  nand g1019 (n_1471, n_442, n_443);
  nand g1020 (n_1472, n_444, n_443);
  nand g1021 (n_1473, n_442, n_444);
  nand g1022 (n_118, n_1471, n_1472, n_1473);
  xor g1023 (n_1474, A[23], A[21]);
  xor g1024 (n_449, n_1474, A[17]);
  nand g1025 (n_1475, A[23], A[21]);
  nand g1026 (n_1476, A[17], A[21]);
  nand g1027 (n_1477, A[23], A[17]);
  nand g1028 (n_459, n_1475, n_1476, n_1477);
  xor g1030 (n_450, n_1246, A[15]);
  nand g1032 (n_1480, A[15], A[7]);
  nand g1034 (n_460, n_1247, n_1480, n_1356);
  xor g1035 (n_1482, A[5], A[19]);
  xor g1036 (n_448, n_1482, A[13]);
  nand g1037 (n_1483, A[5], A[19]);
  nand g1040 (n_461, n_1483, n_1348, n_1207);
  xor g1041 (n_1486, A[11], n_445);
  xor g1042 (n_452, n_1486, n_446);
  nand g1043 (n_1487, A[11], n_445);
  nand g1044 (n_1488, n_446, n_445);
  nand g1045 (n_1489, A[11], n_446);
  nand g1046 (n_465, n_1487, n_1488, n_1489);
  xor g1047 (n_1490, n_447, n_448);
  xor g1048 (n_454, n_1490, n_449);
  nand g1049 (n_1491, n_447, n_448);
  nand g1050 (n_1492, n_449, n_448);
  nand g1051 (n_1493, n_447, n_449);
  nand g1052 (n_467, n_1491, n_1492, n_1493);
  xor g1053 (n_1494, n_450, n_451);
  xor g1054 (n_456, n_1494, n_452);
  nand g1055 (n_1495, n_450, n_451);
  nand g1056 (n_1496, n_452, n_451);
  nand g1057 (n_1497, n_450, n_452);
  nand g1058 (n_469, n_1495, n_1496, n_1497);
  xor g1059 (n_1498, n_453, n_454);
  xor g1060 (n_457, n_1498, n_455);
  nand g1061 (n_1499, n_453, n_454);
  nand g1062 (n_1500, n_455, n_454);
  nand g1063 (n_1501, n_453, n_455);
  nand g1064 (n_472, n_1499, n_1500, n_1501);
  xor g1065 (n_1502, n_456, n_457);
  xor g1066 (n_198, n_1502, n_458);
  nand g1067 (n_1503, n_456, n_457);
  nand g1068 (n_1504, n_458, n_457);
  nand g1069 (n_1505, n_456, n_458);
  nand g1070 (n_117, n_1503, n_1504, n_1505);
  xor g1071 (n_1506, A[24], A[22]);
  xor g1072 (n_463, n_1506, A[18]);
  nand g1073 (n_1507, A[24], A[22]);
  nand g1074 (n_1508, A[18], A[22]);
  nand g1075 (n_1509, A[24], A[18]);
  nand g1076 (n_473, n_1507, n_1508, n_1509);
  xor g1078 (n_464, n_313, A[16]);
  nand g1080 (n_1512, A[16], A[8]);
  xor g1083 (n_1514, A[6], A[20]);
  xor g1084 (n_462, n_1514, A[14]);
  nand g1085 (n_1515, A[6], A[20]);
  nand g1088 (n_475, n_1515, n_1381, n_1448);
  xor g1089 (n_1518, A[12], n_459);
  xor g1090 (n_466, n_1518, n_460);
  nand g1091 (n_1519, A[12], n_459);
  nand g1092 (n_1520, n_460, n_459);
  nand g1093 (n_1521, A[12], n_460);
  nand g1094 (n_479, n_1519, n_1520, n_1521);
  xor g1095 (n_1522, n_461, n_462);
  xor g1096 (n_468, n_1522, n_463);
  nand g1097 (n_1523, n_461, n_462);
  nand g1098 (n_1524, n_463, n_462);
  nand g1099 (n_1525, n_461, n_463);
  nand g1100 (n_481, n_1523, n_1524, n_1525);
  xor g1101 (n_1526, n_464, n_465);
  xor g1102 (n_470, n_1526, n_466);
  nand g1103 (n_1527, n_464, n_465);
  nand g1104 (n_1528, n_466, n_465);
  nand g1105 (n_1529, n_464, n_466);
  nand g1106 (n_483, n_1527, n_1528, n_1529);
  xor g1107 (n_1530, n_467, n_468);
  xor g1108 (n_471, n_1530, n_469);
  nand g1109 (n_1531, n_467, n_468);
  nand g1110 (n_1532, n_469, n_468);
  nand g1111 (n_1533, n_467, n_469);
  nand g1112 (n_486, n_1531, n_1532, n_1533);
  xor g1113 (n_1534, n_470, n_471);
  xor g1114 (n_197, n_1534, n_472);
  nand g1115 (n_1535, n_470, n_471);
  nand g1116 (n_1536, n_472, n_471);
  nand g1117 (n_1537, n_470, n_472);
  nand g1118 (n_116, n_1535, n_1536, n_1537);
  xor g1119 (n_1538, A[25], A[23]);
  xor g1120 (n_477, n_1538, A[19]);
  nand g1121 (n_1539, A[25], A[23]);
  nand g1122 (n_1540, A[19], A[23]);
  nand g1123 (n_1541, A[25], A[19]);
  nand g1124 (n_218, n_1539, n_1540, n_1541);
  xor g1125 (n_1542, A[11], A[9]);
  xor g1126 (n_478, n_1542, A[17]);
  nand g1128 (n_1544, A[17], A[9]);
  nand g1130 (n_219, n_1249, n_1544, n_1420);
  xor g1131 (n_1546, A[7], A[21]);
  xor g1132 (n_476, n_1546, A[15]);
  nand g1133 (n_1547, A[7], A[21]);
  nand g1136 (n_487, n_1547, n_1413, n_1480);
  xor g1137 (n_1550, A[13], n_473);
  xor g1138 (n_480, n_1550, n_474);
  nand g1139 (n_1551, A[13], n_473);
  nand g1140 (n_1552, n_474, n_473);
  nand g1141 (n_1553, A[13], n_474);
  nand g1142 (n_491, n_1551, n_1552, n_1553);
  xor g1143 (n_1554, n_475, n_476);
  xor g1144 (n_482, n_1554, n_477);
  nand g1145 (n_1555, n_475, n_476);
  nand g1146 (n_1556, n_477, n_476);
  nand g1147 (n_1557, n_475, n_477);
  nand g1148 (n_493, n_1555, n_1556, n_1557);
  xor g1149 (n_1558, n_478, n_479);
  xor g1150 (n_484, n_1558, n_480);
  nand g1151 (n_1559, n_478, n_479);
  nand g1152 (n_1560, n_480, n_479);
  nand g1153 (n_1561, n_478, n_480);
  nand g1154 (n_495, n_1559, n_1560, n_1561);
  xor g1155 (n_1562, n_481, n_482);
  xor g1156 (n_485, n_1562, n_483);
  nand g1157 (n_1563, n_481, n_482);
  nand g1158 (n_1564, n_483, n_482);
  nand g1159 (n_1565, n_481, n_483);
  nand g1160 (n_498, n_1563, n_1564, n_1565);
  xor g1161 (n_1566, n_484, n_485);
  xor g1162 (n_196, n_1566, n_486);
  nand g1163 (n_1567, n_484, n_485);
  nand g1164 (n_1568, n_486, n_485);
  nand g1165 (n_1569, n_484, n_486);
  nand g1166 (n_115, n_1567, n_1568, n_1569);
  xor g1167 (n_1570, A[26], A[24]);
  xor g1168 (n_489, n_1570, A[20]);
  nand g1169 (n_1571, A[26], A[24]);
  nand g1170 (n_1572, A[20], A[24]);
  nand g1171 (n_1573, A[26], A[20]);
  nand g1172 (n_499, n_1571, n_1572, n_1573);
  xor g1174 (n_490, n_324, A[18]);
  nand g1176 (n_1576, A[18], A[10]);
  xor g1179 (n_1578, A[8], A[22]);
  xor g1180 (n_488, n_1578, A[16]);
  nand g1181 (n_1579, A[8], A[22]);
  nand g1184 (n_501, n_1579, n_1445, n_1512);
  xor g1185 (n_1582, A[14], n_218);
  xor g1186 (n_492, n_1582, n_219);
  nand g1187 (n_1583, A[14], n_218);
  nand g1188 (n_1584, n_219, n_218);
  nand g1189 (n_1585, A[14], n_219);
  nand g1190 (n_505, n_1583, n_1584, n_1585);
  xor g1191 (n_1586, n_487, n_488);
  xor g1192 (n_494, n_1586, n_489);
  nand g1193 (n_1587, n_487, n_488);
  nand g1194 (n_1588, n_489, n_488);
  nand g1195 (n_1589, n_487, n_489);
  nand g1196 (n_507, n_1587, n_1588, n_1589);
  xor g1197 (n_1590, n_490, n_491);
  xor g1198 (n_496, n_1590, n_492);
  nand g1199 (n_1591, n_490, n_491);
  nand g1200 (n_1592, n_492, n_491);
  nand g1201 (n_1593, n_490, n_492);
  nand g1202 (n_509, n_1591, n_1592, n_1593);
  xor g1203 (n_1594, n_493, n_494);
  xor g1204 (n_497, n_1594, n_495);
  nand g1205 (n_1595, n_493, n_494);
  nand g1206 (n_1596, n_495, n_494);
  nand g1207 (n_1597, n_493, n_495);
  nand g1208 (n_512, n_1595, n_1596, n_1597);
  xor g1209 (n_1598, n_496, n_497);
  xor g1210 (n_195, n_1598, n_498);
  nand g1211 (n_1599, n_496, n_497);
  nand g1212 (n_1600, n_498, n_497);
  nand g1213 (n_1601, n_496, n_498);
  nand g1214 (n_114, n_1599, n_1600, n_1601);
  xor g1215 (n_1602, A[27], A[25]);
  xor g1216 (n_503, n_1602, A[21]);
  nand g1217 (n_1603, A[27], A[25]);
  nand g1218 (n_1604, A[21], A[25]);
  nand g1219 (n_1605, A[27], A[21]);
  nand g1220 (n_513, n_1603, n_1604, n_1605);
  xor g1221 (n_1606, A[13], A[11]);
  xor g1222 (n_504, n_1606, A[19]);
  nand g1223 (n_1607, A[13], A[11]);
  nand g1224 (n_1608, A[19], A[11]);
  nand g1226 (n_514, n_1607, n_1608, n_1348);
  xor g1227 (n_1610, A[9], A[23]);
  xor g1228 (n_502, n_1610, A[17]);
  nand g1229 (n_1611, A[9], A[23]);
  nand g1232 (n_515, n_1611, n_1477, n_1544);
  xor g1233 (n_1614, A[15], n_499);
  xor g1234 (n_506, n_1614, n_500);
  nand g1235 (n_1615, A[15], n_499);
  nand g1236 (n_1616, n_500, n_499);
  nand g1237 (n_1617, A[15], n_500);
  nand g1238 (n_519, n_1615, n_1616, n_1617);
  xor g1239 (n_1618, n_501, n_502);
  xor g1240 (n_508, n_1618, n_503);
  nand g1241 (n_1619, n_501, n_502);
  nand g1242 (n_1620, n_503, n_502);
  nand g1243 (n_1621, n_501, n_503);
  nand g1244 (n_521, n_1619, n_1620, n_1621);
  xor g1245 (n_1622, n_504, n_505);
  xor g1246 (n_510, n_1622, n_506);
  nand g1247 (n_1623, n_504, n_505);
  nand g1248 (n_1624, n_506, n_505);
  nand g1249 (n_1625, n_504, n_506);
  nand g1250 (n_523, n_1623, n_1624, n_1625);
  xor g1251 (n_1626, n_507, n_508);
  xor g1252 (n_511, n_1626, n_509);
  nand g1253 (n_1627, n_507, n_508);
  nand g1254 (n_1628, n_509, n_508);
  nand g1255 (n_1629, n_507, n_509);
  nand g1256 (n_526, n_1627, n_1628, n_1629);
  xor g1257 (n_1630, n_510, n_511);
  xor g1258 (n_194, n_1630, n_512);
  nand g1259 (n_1631, n_510, n_511);
  nand g1260 (n_1632, n_512, n_511);
  nand g1261 (n_1633, n_510, n_512);
  nand g1262 (n_113, n_1631, n_1632, n_1633);
  xor g1263 (n_1634, A[28], A[26]);
  xor g1264 (n_517, n_1634, A[22]);
  nand g1265 (n_1635, A[28], A[26]);
  nand g1266 (n_1636, A[22], A[26]);
  nand g1267 (n_1637, A[28], A[22]);
  nand g1268 (n_527, n_1635, n_1636, n_1637);
  xor g1270 (n_518, n_339, A[20]);
  nand g1272 (n_1640, A[20], A[12]);
  xor g1275 (n_1642, A[10], A[24]);
  xor g1276 (n_516, n_1642, A[18]);
  nand g1277 (n_1643, A[10], A[24]);
  nand g1280 (n_529, n_1643, n_1509, n_1576);
  xor g1281 (n_1646, A[16], n_513);
  xor g1282 (n_520, n_1646, n_514);
  nand g1283 (n_1647, A[16], n_513);
  nand g1284 (n_1648, n_514, n_513);
  nand g1285 (n_1649, A[16], n_514);
  nand g1286 (n_533, n_1647, n_1648, n_1649);
  xor g1287 (n_1650, n_515, n_516);
  xor g1288 (n_522, n_1650, n_517);
  nand g1289 (n_1651, n_515, n_516);
  nand g1290 (n_1652, n_517, n_516);
  nand g1291 (n_1653, n_515, n_517);
  nand g1292 (n_535, n_1651, n_1652, n_1653);
  xor g1293 (n_1654, n_518, n_519);
  xor g1294 (n_524, n_1654, n_520);
  nand g1295 (n_1655, n_518, n_519);
  nand g1296 (n_1656, n_520, n_519);
  nand g1297 (n_1657, n_518, n_520);
  nand g1298 (n_537, n_1655, n_1656, n_1657);
  xor g1299 (n_1658, n_521, n_522);
  xor g1300 (n_525, n_1658, n_523);
  nand g1301 (n_1659, n_521, n_522);
  nand g1302 (n_1660, n_523, n_522);
  nand g1303 (n_1661, n_521, n_523);
  nand g1304 (n_540, n_1659, n_1660, n_1661);
  xor g1305 (n_1662, n_524, n_525);
  xor g1306 (n_193, n_1662, n_526);
  nand g1307 (n_1663, n_524, n_525);
  nand g1308 (n_1664, n_526, n_525);
  nand g1309 (n_1665, n_524, n_526);
  nand g1310 (n_112, n_1663, n_1664, n_1665);
  xor g1311 (n_1666, A[29], A[27]);
  xor g1312 (n_531, n_1666, A[23]);
  nand g1313 (n_1667, A[29], A[27]);
  nand g1314 (n_1668, A[23], A[27]);
  nand g1315 (n_1669, A[29], A[23]);
  nand g1316 (n_541, n_1667, n_1668, n_1669);
  xor g1317 (n_1670, A[15], A[13]);
  xor g1318 (n_532, n_1670, A[21]);
  nand g1320 (n_1672, A[21], A[13]);
  nand g1322 (n_542, n_1244, n_1672, n_1413);
  xor g1323 (n_1674, A[11], A[25]);
  xor g1324 (n_530, n_1674, A[19]);
  nand g1325 (n_1675, A[11], A[25]);
  nand g1328 (n_543, n_1675, n_1541, n_1608);
  xor g1329 (n_1678, A[17], n_527);
  xor g1330 (n_534, n_1678, n_528);
  nand g1331 (n_1679, A[17], n_527);
  nand g1332 (n_1680, n_528, n_527);
  nand g1333 (n_1681, A[17], n_528);
  nand g1334 (n_547, n_1679, n_1680, n_1681);
  xor g1335 (n_1682, n_529, n_530);
  xor g1336 (n_536, n_1682, n_531);
  nand g1337 (n_1683, n_529, n_530);
  nand g1338 (n_1684, n_531, n_530);
  nand g1339 (n_1685, n_529, n_531);
  nand g1340 (n_549, n_1683, n_1684, n_1685);
  xor g1341 (n_1686, n_532, n_533);
  xor g1342 (n_538, n_1686, n_534);
  nand g1343 (n_1687, n_532, n_533);
  nand g1344 (n_1688, n_534, n_533);
  nand g1345 (n_1689, n_532, n_534);
  nand g1346 (n_551, n_1687, n_1688, n_1689);
  xor g1347 (n_1690, n_535, n_536);
  xor g1348 (n_539, n_1690, n_537);
  nand g1349 (n_1691, n_535, n_536);
  nand g1350 (n_1692, n_537, n_536);
  nand g1351 (n_1693, n_535, n_537);
  nand g1352 (n_554, n_1691, n_1692, n_1693);
  xor g1353 (n_1694, n_538, n_539);
  xor g1354 (n_192, n_1694, n_540);
  nand g1355 (n_1695, n_538, n_539);
  nand g1356 (n_1696, n_540, n_539);
  nand g1357 (n_1697, n_538, n_540);
  nand g1358 (n_111, n_1695, n_1696, n_1697);
  xor g1359 (n_1698, A[30], A[28]);
  xor g1360 (n_545, n_1698, A[24]);
  nand g1361 (n_1699, A[30], A[28]);
  nand g1362 (n_1700, A[24], A[28]);
  nand g1363 (n_1701, A[30], A[24]);
  nand g1364 (n_555, n_1699, n_1700, n_1701);
  xor g1366 (n_546, n_358, A[22]);
  nand g1368 (n_1704, A[22], A[14]);
  xor g1371 (n_1706, A[12], A[26]);
  xor g1372 (n_544, n_1706, A[20]);
  nand g1373 (n_1707, A[12], A[26]);
  nand g1376 (n_557, n_1707, n_1573, n_1640);
  xor g1377 (n_1710, A[18], n_541);
  xor g1378 (n_548, n_1710, n_542);
  nand g1379 (n_1711, A[18], n_541);
  nand g1380 (n_1712, n_542, n_541);
  nand g1381 (n_1713, A[18], n_542);
  nand g1382 (n_561, n_1711, n_1712, n_1713);
  xor g1383 (n_1714, n_543, n_544);
  xor g1384 (n_550, n_1714, n_545);
  nand g1385 (n_1715, n_543, n_544);
  nand g1386 (n_1716, n_545, n_544);
  nand g1387 (n_1717, n_543, n_545);
  nand g1388 (n_563, n_1715, n_1716, n_1717);
  xor g1389 (n_1718, n_546, n_547);
  xor g1390 (n_552, n_1718, n_548);
  nand g1391 (n_1719, n_546, n_547);
  nand g1392 (n_1720, n_548, n_547);
  nand g1393 (n_1721, n_546, n_548);
  nand g1394 (n_565, n_1719, n_1720, n_1721);
  xor g1395 (n_1722, n_549, n_550);
  xor g1396 (n_553, n_1722, n_551);
  nand g1397 (n_1723, n_549, n_550);
  nand g1398 (n_1724, n_551, n_550);
  nand g1399 (n_1725, n_549, n_551);
  nand g1400 (n_568, n_1723, n_1724, n_1725);
  xor g1401 (n_1726, n_552, n_553);
  xor g1402 (n_191, n_1726, n_554);
  nand g1403 (n_1727, n_552, n_553);
  nand g1404 (n_1728, n_554, n_553);
  nand g1405 (n_1729, n_552, n_554);
  nand g1406 (n_110, n_1727, n_1728, n_1729);
  xor g1407 (n_1730, A[31], A[29]);
  xor g1408 (n_559, n_1730, A[25]);
  nand g1409 (n_1731, A[31], A[29]);
  nand g1410 (n_1732, A[25], A[29]);
  nand g1411 (n_1733, A[31], A[25]);
  nand g1412 (n_569, n_1731, n_1732, n_1733);
  xor g1413 (n_1734, A[17], A[15]);
  xor g1414 (n_560, n_1734, A[23]);
  nand g1416 (n_1736, A[23], A[15]);
  nand g1418 (n_570, n_1292, n_1736, n_1477);
  xor g1419 (n_1738, A[13], A[27]);
  xor g1420 (n_558, n_1738, A[21]);
  nand g1421 (n_1739, A[13], A[27]);
  nand g1424 (n_571, n_1739, n_1605, n_1672);
  xor g1425 (n_1742, A[19], n_555);
  xor g1426 (n_562, n_1742, n_556);
  nand g1427 (n_1743, A[19], n_555);
  nand g1428 (n_1744, n_556, n_555);
  nand g1429 (n_1745, A[19], n_556);
  nand g1430 (n_575, n_1743, n_1744, n_1745);
  xor g1431 (n_1746, n_557, n_558);
  xor g1432 (n_564, n_1746, n_559);
  nand g1433 (n_1747, n_557, n_558);
  nand g1434 (n_1748, n_559, n_558);
  nand g1435 (n_1749, n_557, n_559);
  nand g1436 (n_577, n_1747, n_1748, n_1749);
  xor g1437 (n_1750, n_560, n_561);
  xor g1438 (n_566, n_1750, n_562);
  nand g1439 (n_1751, n_560, n_561);
  nand g1440 (n_1752, n_562, n_561);
  nand g1441 (n_1753, n_560, n_562);
  nand g1442 (n_579, n_1751, n_1752, n_1753);
  xor g1443 (n_1754, n_563, n_564);
  xor g1444 (n_567, n_1754, n_565);
  nand g1445 (n_1755, n_563, n_564);
  nand g1446 (n_1756, n_565, n_564);
  nand g1447 (n_1757, n_563, n_565);
  nand g1448 (n_582, n_1755, n_1756, n_1757);
  xor g1449 (n_1758, n_566, n_567);
  xor g1450 (n_190, n_1758, n_568);
  nand g1451 (n_1759, n_566, n_567);
  nand g1452 (n_1760, n_568, n_567);
  nand g1453 (n_1761, n_566, n_568);
  nand g1454 (n_109, n_1759, n_1760, n_1761);
  xor g1455 (n_1762, A[32], A[30]);
  xor g1456 (n_573, n_1762, A[26]);
  nand g1457 (n_1763, A[32], A[30]);
  nand g1458 (n_1764, A[26], A[30]);
  nand g1459 (n_1765, A[32], A[26]);
  nand g1460 (n_583, n_1763, n_1764, n_1765);
  xor g1462 (n_574, n_381, A[24]);
  nand g1464 (n_1768, A[24], A[16]);
  xor g1467 (n_1770, A[14], A[28]);
  xor g1468 (n_572, n_1770, A[22]);
  nand g1469 (n_1771, A[14], A[28]);
  nand g1472 (n_585, n_1771, n_1637, n_1704);
  xor g1473 (n_1774, A[20], n_569);
  xor g1474 (n_576, n_1774, n_570);
  nand g1475 (n_1775, A[20], n_569);
  nand g1476 (n_1776, n_570, n_569);
  nand g1477 (n_1777, A[20], n_570);
  nand g1478 (n_589, n_1775, n_1776, n_1777);
  xor g1479 (n_1778, n_571, n_572);
  xor g1480 (n_578, n_1778, n_573);
  nand g1481 (n_1779, n_571, n_572);
  nand g1482 (n_1780, n_573, n_572);
  nand g1483 (n_1781, n_571, n_573);
  nand g1484 (n_591, n_1779, n_1780, n_1781);
  xor g1485 (n_1782, n_574, n_575);
  xor g1486 (n_580, n_1782, n_576);
  nand g1487 (n_1783, n_574, n_575);
  nand g1488 (n_1784, n_576, n_575);
  nand g1489 (n_1785, n_574, n_576);
  nand g1490 (n_593, n_1783, n_1784, n_1785);
  xor g1491 (n_1786, n_577, n_578);
  xor g1492 (n_581, n_1786, n_579);
  nand g1493 (n_1787, n_577, n_578);
  nand g1494 (n_1788, n_579, n_578);
  nand g1495 (n_1789, n_577, n_579);
  nand g1496 (n_596, n_1787, n_1788, n_1789);
  xor g1497 (n_1790, n_580, n_581);
  xor g1498 (n_189, n_1790, n_582);
  nand g1499 (n_1791, n_580, n_581);
  nand g1500 (n_1792, n_582, n_581);
  nand g1501 (n_1793, n_580, n_582);
  nand g1502 (n_108, n_1791, n_1792, n_1793);
  xor g1503 (n_1794, A[33], A[31]);
  xor g1504 (n_587, n_1794, A[27]);
  nand g1505 (n_1795, A[33], A[31]);
  nand g1506 (n_1796, A[27], A[31]);
  nand g1507 (n_1797, A[33], A[27]);
  nand g1508 (n_597, n_1795, n_1796, n_1797);
  xor g1509 (n_1798, A[19], A[17]);
  xor g1510 (n_588, n_1798, A[25]);
  nand g1511 (n_1799, A[19], A[17]);
  nand g1512 (n_1800, A[25], A[17]);
  nand g1514 (n_598, n_1799, n_1800, n_1541);
  xor g1515 (n_1802, A[15], A[29]);
  xor g1516 (n_586, n_1802, A[23]);
  nand g1517 (n_1803, A[15], A[29]);
  nand g1520 (n_599, n_1803, n_1669, n_1736);
  xor g1521 (n_1806, A[21], n_583);
  xor g1522 (n_590, n_1806, n_584);
  nand g1523 (n_1807, A[21], n_583);
  nand g1524 (n_1808, n_584, n_583);
  nand g1525 (n_1809, A[21], n_584);
  nand g1526 (n_603, n_1807, n_1808, n_1809);
  xor g1527 (n_1810, n_585, n_586);
  xor g1528 (n_592, n_1810, n_587);
  nand g1529 (n_1811, n_585, n_586);
  nand g1530 (n_1812, n_587, n_586);
  nand g1531 (n_1813, n_585, n_587);
  nand g1532 (n_605, n_1811, n_1812, n_1813);
  xor g1533 (n_1814, n_588, n_589);
  xor g1534 (n_594, n_1814, n_590);
  nand g1535 (n_1815, n_588, n_589);
  nand g1536 (n_1816, n_590, n_589);
  nand g1537 (n_1817, n_588, n_590);
  nand g1538 (n_607, n_1815, n_1816, n_1817);
  xor g1539 (n_1818, n_591, n_592);
  xor g1540 (n_595, n_1818, n_593);
  nand g1541 (n_1819, n_591, n_592);
  nand g1542 (n_1820, n_593, n_592);
  nand g1543 (n_1821, n_591, n_593);
  nand g1544 (n_610, n_1819, n_1820, n_1821);
  xor g1545 (n_1822, n_594, n_595);
  xor g1546 (n_188, n_1822, n_596);
  nand g1547 (n_1823, n_594, n_595);
  nand g1548 (n_1824, n_596, n_595);
  nand g1549 (n_1825, n_594, n_596);
  nand g1550 (n_107, n_1823, n_1824, n_1825);
  xor g1551 (n_1826, A[34], A[32]);
  xor g1552 (n_601, n_1826, A[28]);
  nand g1553 (n_1827, A[34], A[32]);
  nand g1554 (n_1828, A[28], A[32]);
  nand g1555 (n_1829, A[34], A[28]);
  nand g1556 (n_611, n_1827, n_1828, n_1829);
  xor g1558 (n_602, n_1378, A[26]);
  nand g1560 (n_1832, A[26], A[18]);
  nand g1562 (n_612, n_1379, n_1832, n_1573);
  xor g1563 (n_1834, A[16], A[30]);
  xor g1564 (n_600, n_1834, A[24]);
  nand g1565 (n_1835, A[16], A[30]);
  nand g1568 (n_613, n_1835, n_1701, n_1768);
  xor g1569 (n_1838, A[22], n_597);
  xor g1570 (n_604, n_1838, n_598);
  nand g1571 (n_1839, A[22], n_597);
  nand g1572 (n_1840, n_598, n_597);
  nand g1573 (n_1841, A[22], n_598);
  nand g1574 (n_617, n_1839, n_1840, n_1841);
  xor g1575 (n_1842, n_599, n_600);
  xor g1576 (n_606, n_1842, n_601);
  nand g1577 (n_1843, n_599, n_600);
  nand g1578 (n_1844, n_601, n_600);
  nand g1579 (n_1845, n_599, n_601);
  nand g1580 (n_619, n_1843, n_1844, n_1845);
  xor g1581 (n_1846, n_602, n_603);
  xor g1582 (n_608, n_1846, n_604);
  nand g1583 (n_1847, n_602, n_603);
  nand g1584 (n_1848, n_604, n_603);
  nand g1585 (n_1849, n_602, n_604);
  nand g1586 (n_621, n_1847, n_1848, n_1849);
  xor g1587 (n_1850, n_605, n_606);
  xor g1588 (n_609, n_1850, n_607);
  nand g1589 (n_1851, n_605, n_606);
  nand g1590 (n_1852, n_607, n_606);
  nand g1591 (n_1853, n_605, n_607);
  nand g1592 (n_624, n_1851, n_1852, n_1853);
  xor g1593 (n_1854, n_608, n_609);
  xor g1594 (n_187, n_1854, n_610);
  nand g1595 (n_1855, n_608, n_609);
  nand g1596 (n_1856, n_610, n_609);
  nand g1597 (n_1857, n_608, n_610);
  nand g1598 (n_106, n_1855, n_1856, n_1857);
  xor g1599 (n_1858, A[35], A[33]);
  xor g1600 (n_615, n_1858, A[29]);
  nand g1601 (n_1859, A[35], A[33]);
  nand g1602 (n_1860, A[29], A[33]);
  nand g1603 (n_1861, A[35], A[29]);
  nand g1604 (n_625, n_1859, n_1860, n_1861);
  xor g1606 (n_616, n_1410, A[27]);
  nand g1608 (n_1864, A[27], A[19]);
  nand g1610 (n_626, n_1411, n_1864, n_1605);
  xor g1611 (n_1866, A[17], A[31]);
  xor g1612 (n_614, n_1866, A[25]);
  nand g1613 (n_1867, A[17], A[31]);
  nand g1616 (n_627, n_1867, n_1733, n_1800);
  xor g1617 (n_1870, A[23], n_611);
  xor g1618 (n_618, n_1870, n_612);
  nand g1619 (n_1871, A[23], n_611);
  nand g1620 (n_1872, n_612, n_611);
  nand g1621 (n_1873, A[23], n_612);
  nand g1622 (n_631, n_1871, n_1872, n_1873);
  xor g1623 (n_1874, n_613, n_614);
  xor g1624 (n_620, n_1874, n_615);
  nand g1625 (n_1875, n_613, n_614);
  nand g1626 (n_1876, n_615, n_614);
  nand g1627 (n_1877, n_613, n_615);
  nand g1628 (n_633, n_1875, n_1876, n_1877);
  xor g1629 (n_1878, n_616, n_617);
  xor g1630 (n_622, n_1878, n_618);
  nand g1631 (n_1879, n_616, n_617);
  nand g1632 (n_1880, n_618, n_617);
  nand g1633 (n_1881, n_616, n_618);
  nand g1634 (n_635, n_1879, n_1880, n_1881);
  xor g1635 (n_1882, n_619, n_620);
  xor g1636 (n_623, n_1882, n_621);
  nand g1637 (n_1883, n_619, n_620);
  nand g1638 (n_1884, n_621, n_620);
  nand g1639 (n_1885, n_619, n_621);
  nand g1640 (n_638, n_1883, n_1884, n_1885);
  xor g1641 (n_1886, n_622, n_623);
  xor g1642 (n_186, n_1886, n_624);
  nand g1643 (n_1887, n_622, n_623);
  nand g1644 (n_1888, n_624, n_623);
  nand g1645 (n_1889, n_622, n_624);
  nand g1646 (n_105, n_1887, n_1888, n_1889);
  xor g1647 (n_1890, A[36], A[34]);
  xor g1648 (n_629, n_1890, A[30]);
  nand g1649 (n_1891, A[36], A[34]);
  nand g1650 (n_1892, A[30], A[34]);
  nand g1651 (n_1893, A[36], A[30]);
  nand g1652 (n_639, n_1891, n_1892, n_1893);
  xor g1654 (n_630, n_1442, A[28]);
  nand g1656 (n_1896, A[28], A[20]);
  nand g1658 (n_640, n_1443, n_1896, n_1637);
  xor g1659 (n_1898, A[18], A[32]);
  xor g1660 (n_628, n_1898, A[26]);
  nand g1661 (n_1899, A[18], A[32]);
  nand g1664 (n_641, n_1899, n_1765, n_1832);
  xor g1665 (n_1902, A[24], n_625);
  xor g1666 (n_632, n_1902, n_626);
  nand g1667 (n_1903, A[24], n_625);
  nand g1668 (n_1904, n_626, n_625);
  nand g1669 (n_1905, A[24], n_626);
  nand g1670 (n_645, n_1903, n_1904, n_1905);
  xor g1671 (n_1906, n_627, n_628);
  xor g1672 (n_634, n_1906, n_629);
  nand g1673 (n_1907, n_627, n_628);
  nand g1674 (n_1908, n_629, n_628);
  nand g1675 (n_1909, n_627, n_629);
  nand g1676 (n_647, n_1907, n_1908, n_1909);
  xor g1677 (n_1910, n_630, n_631);
  xor g1678 (n_636, n_1910, n_632);
  nand g1679 (n_1911, n_630, n_631);
  nand g1680 (n_1912, n_632, n_631);
  nand g1681 (n_1913, n_630, n_632);
  nand g1682 (n_649, n_1911, n_1912, n_1913);
  xor g1683 (n_1914, n_633, n_634);
  xor g1684 (n_637, n_1914, n_635);
  nand g1685 (n_1915, n_633, n_634);
  nand g1686 (n_1916, n_635, n_634);
  nand g1687 (n_1917, n_633, n_635);
  nand g1688 (n_652, n_1915, n_1916, n_1917);
  xor g1689 (n_1918, n_636, n_637);
  xor g1690 (n_185, n_1918, n_638);
  nand g1691 (n_1919, n_636, n_637);
  nand g1692 (n_1920, n_638, n_637);
  nand g1693 (n_1921, n_636, n_638);
  nand g1694 (n_104, n_1919, n_1920, n_1921);
  xor g1695 (n_1922, A[37], A[35]);
  xor g1696 (n_643, n_1922, A[31]);
  nand g1697 (n_1923, A[37], A[35]);
  nand g1698 (n_1924, A[31], A[35]);
  nand g1699 (n_1925, A[37], A[31]);
  nand g1700 (n_653, n_1923, n_1924, n_1925);
  xor g1702 (n_644, n_1474, A[29]);
  nand g1704 (n_1928, A[29], A[21]);
  nand g1706 (n_654, n_1475, n_1928, n_1669);
  xor g1707 (n_1930, A[19], A[33]);
  xor g1708 (n_642, n_1930, A[27]);
  nand g1709 (n_1931, A[19], A[33]);
  nand g1712 (n_655, n_1931, n_1797, n_1864);
  xor g1713 (n_1934, A[25], n_639);
  xor g1714 (n_646, n_1934, n_640);
  nand g1715 (n_1935, A[25], n_639);
  nand g1716 (n_1936, n_640, n_639);
  nand g1717 (n_1937, A[25], n_640);
  nand g1718 (n_659, n_1935, n_1936, n_1937);
  xor g1719 (n_1938, n_641, n_642);
  xor g1720 (n_648, n_1938, n_643);
  nand g1721 (n_1939, n_641, n_642);
  nand g1722 (n_1940, n_643, n_642);
  nand g1723 (n_1941, n_641, n_643);
  nand g1724 (n_661, n_1939, n_1940, n_1941);
  xor g1725 (n_1942, n_644, n_645);
  xor g1726 (n_650, n_1942, n_646);
  nand g1727 (n_1943, n_644, n_645);
  nand g1728 (n_1944, n_646, n_645);
  nand g1729 (n_1945, n_644, n_646);
  nand g1730 (n_663, n_1943, n_1944, n_1945);
  xor g1731 (n_1946, n_647, n_648);
  xor g1732 (n_651, n_1946, n_649);
  nand g1733 (n_1947, n_647, n_648);
  nand g1734 (n_1948, n_649, n_648);
  nand g1735 (n_1949, n_647, n_649);
  nand g1736 (n_666, n_1947, n_1948, n_1949);
  xor g1737 (n_1950, n_650, n_651);
  xor g1738 (n_184, n_1950, n_652);
  nand g1739 (n_1951, n_650, n_651);
  nand g1740 (n_1952, n_652, n_651);
  nand g1741 (n_1953, n_650, n_652);
  nand g1742 (n_103, n_1951, n_1952, n_1953);
  xor g1743 (n_1954, A[38], A[36]);
  xor g1744 (n_657, n_1954, A[32]);
  nand g1745 (n_1955, A[38], A[36]);
  nand g1746 (n_1956, A[32], A[36]);
  nand g1747 (n_1957, A[38], A[32]);
  nand g1748 (n_667, n_1955, n_1956, n_1957);
  xor g1750 (n_658, n_1506, A[30]);
  nand g1752 (n_1960, A[30], A[22]);
  nand g1754 (n_668, n_1507, n_1960, n_1701);
  xor g1755 (n_1962, A[20], A[34]);
  xor g1756 (n_656, n_1962, A[28]);
  nand g1757 (n_1963, A[20], A[34]);
  nand g1760 (n_669, n_1963, n_1829, n_1896);
  xor g1761 (n_1966, A[26], n_653);
  xor g1762 (n_660, n_1966, n_654);
  nand g1763 (n_1967, A[26], n_653);
  nand g1764 (n_1968, n_654, n_653);
  nand g1765 (n_1969, A[26], n_654);
  nand g1766 (n_673, n_1967, n_1968, n_1969);
  xor g1767 (n_1970, n_655, n_656);
  xor g1768 (n_662, n_1970, n_657);
  nand g1769 (n_1971, n_655, n_656);
  nand g1770 (n_1972, n_657, n_656);
  nand g1771 (n_1973, n_655, n_657);
  nand g1772 (n_675, n_1971, n_1972, n_1973);
  xor g1773 (n_1974, n_658, n_659);
  xor g1774 (n_664, n_1974, n_660);
  nand g1775 (n_1975, n_658, n_659);
  nand g1776 (n_1976, n_660, n_659);
  nand g1777 (n_1977, n_658, n_660);
  nand g1778 (n_677, n_1975, n_1976, n_1977);
  xor g1779 (n_1978, n_661, n_662);
  xor g1780 (n_665, n_1978, n_663);
  nand g1781 (n_1979, n_661, n_662);
  nand g1782 (n_1980, n_663, n_662);
  nand g1783 (n_1981, n_661, n_663);
  nand g1784 (n_680, n_1979, n_1980, n_1981);
  xor g1785 (n_1982, n_664, n_665);
  xor g1786 (n_183, n_1982, n_666);
  nand g1787 (n_1983, n_664, n_665);
  nand g1788 (n_1984, n_666, n_665);
  nand g1789 (n_1985, n_664, n_666);
  nand g1790 (n_102, n_1983, n_1984, n_1985);
  xor g1791 (n_1986, A[39], A[37]);
  xor g1792 (n_671, n_1986, A[33]);
  nand g1793 (n_1987, A[39], A[37]);
  nand g1794 (n_1988, A[33], A[37]);
  nand g1795 (n_1989, A[39], A[33]);
  nand g1796 (n_681, n_1987, n_1988, n_1989);
  xor g1798 (n_672, n_1538, A[31]);
  nand g1800 (n_1992, A[31], A[23]);
  nand g1802 (n_682, n_1539, n_1992, n_1733);
  xor g1803 (n_1994, A[21], A[35]);
  xor g1804 (n_670, n_1994, A[29]);
  nand g1805 (n_1995, A[21], A[35]);
  nand g1808 (n_683, n_1995, n_1861, n_1928);
  xor g1809 (n_1998, A[27], n_667);
  xor g1810 (n_674, n_1998, n_668);
  nand g1811 (n_1999, A[27], n_667);
  nand g1812 (n_2000, n_668, n_667);
  nand g1813 (n_2001, A[27], n_668);
  nand g1814 (n_687, n_1999, n_2000, n_2001);
  xor g1815 (n_2002, n_669, n_670);
  xor g1816 (n_676, n_2002, n_671);
  nand g1817 (n_2003, n_669, n_670);
  nand g1818 (n_2004, n_671, n_670);
  nand g1819 (n_2005, n_669, n_671);
  nand g1820 (n_689, n_2003, n_2004, n_2005);
  xor g1821 (n_2006, n_672, n_673);
  xor g1822 (n_678, n_2006, n_674);
  nand g1823 (n_2007, n_672, n_673);
  nand g1824 (n_2008, n_674, n_673);
  nand g1825 (n_2009, n_672, n_674);
  nand g1826 (n_691, n_2007, n_2008, n_2009);
  xor g1827 (n_2010, n_675, n_676);
  xor g1828 (n_679, n_2010, n_677);
  nand g1829 (n_2011, n_675, n_676);
  nand g1830 (n_2012, n_677, n_676);
  nand g1831 (n_2013, n_675, n_677);
  nand g1832 (n_694, n_2011, n_2012, n_2013);
  xor g1833 (n_2014, n_678, n_679);
  xor g1834 (n_182, n_2014, n_680);
  nand g1835 (n_2015, n_678, n_679);
  nand g1836 (n_2016, n_680, n_679);
  nand g1837 (n_2017, n_678, n_680);
  nand g1838 (n_101, n_2015, n_2016, n_2017);
  xor g1839 (n_2018, A[40], A[38]);
  xor g1840 (n_685, n_2018, A[34]);
  nand g1841 (n_2019, A[40], A[38]);
  nand g1842 (n_2020, A[34], A[38]);
  nand g1843 (n_2021, A[40], A[34]);
  nand g1844 (n_695, n_2019, n_2020, n_2021);
  xor g1846 (n_686, n_1570, A[32]);
  nand g1848 (n_2024, A[32], A[24]);
  nand g1850 (n_696, n_1571, n_2024, n_1765);
  xor g1851 (n_2026, A[22], A[36]);
  xor g1852 (n_684, n_2026, A[30]);
  nand g1853 (n_2027, A[22], A[36]);
  nand g1856 (n_697, n_2027, n_1893, n_1960);
  xor g1857 (n_2030, A[28], n_681);
  xor g1858 (n_688, n_2030, n_682);
  nand g1859 (n_2031, A[28], n_681);
  nand g1860 (n_2032, n_682, n_681);
  nand g1861 (n_2033, A[28], n_682);
  nand g1862 (n_701, n_2031, n_2032, n_2033);
  xor g1863 (n_2034, n_683, n_684);
  xor g1864 (n_690, n_2034, n_685);
  nand g1865 (n_2035, n_683, n_684);
  nand g1866 (n_2036, n_685, n_684);
  nand g1867 (n_2037, n_683, n_685);
  nand g1868 (n_703, n_2035, n_2036, n_2037);
  xor g1869 (n_2038, n_686, n_687);
  xor g1870 (n_692, n_2038, n_688);
  nand g1871 (n_2039, n_686, n_687);
  nand g1872 (n_2040, n_688, n_687);
  nand g1873 (n_2041, n_686, n_688);
  nand g1874 (n_705, n_2039, n_2040, n_2041);
  xor g1875 (n_2042, n_689, n_690);
  xor g1876 (n_693, n_2042, n_691);
  nand g1877 (n_2043, n_689, n_690);
  nand g1878 (n_2044, n_691, n_690);
  nand g1879 (n_2045, n_689, n_691);
  nand g1880 (n_708, n_2043, n_2044, n_2045);
  xor g1881 (n_2046, n_692, n_693);
  xor g1882 (n_181, n_2046, n_694);
  nand g1883 (n_2047, n_692, n_693);
  nand g1884 (n_2048, n_694, n_693);
  nand g1885 (n_2049, n_692, n_694);
  nand g1886 (n_100, n_2047, n_2048, n_2049);
  xor g1887 (n_2050, A[41], A[39]);
  xor g1888 (n_699, n_2050, A[35]);
  nand g1889 (n_2051, A[41], A[39]);
  nand g1890 (n_2052, A[35], A[39]);
  nand g1891 (n_2053, A[41], A[35]);
  nand g1892 (n_709, n_2051, n_2052, n_2053);
  xor g1894 (n_700, n_1602, A[33]);
  nand g1896 (n_2056, A[33], A[25]);
  nand g1898 (n_710, n_1603, n_2056, n_1797);
  xor g1899 (n_2058, A[23], A[37]);
  xor g1900 (n_698, n_2058, A[31]);
  nand g1901 (n_2059, A[23], A[37]);
  nand g1904 (n_711, n_2059, n_1925, n_1992);
  xor g1905 (n_2062, A[29], n_695);
  xor g1906 (n_702, n_2062, n_696);
  nand g1907 (n_2063, A[29], n_695);
  nand g1908 (n_2064, n_696, n_695);
  nand g1909 (n_2065, A[29], n_696);
  nand g1910 (n_715, n_2063, n_2064, n_2065);
  xor g1911 (n_2066, n_697, n_698);
  xor g1912 (n_704, n_2066, n_699);
  nand g1913 (n_2067, n_697, n_698);
  nand g1914 (n_2068, n_699, n_698);
  nand g1915 (n_2069, n_697, n_699);
  nand g1916 (n_717, n_2067, n_2068, n_2069);
  xor g1917 (n_2070, n_700, n_701);
  xor g1918 (n_706, n_2070, n_702);
  nand g1919 (n_2071, n_700, n_701);
  nand g1920 (n_2072, n_702, n_701);
  nand g1921 (n_2073, n_700, n_702);
  nand g1922 (n_719, n_2071, n_2072, n_2073);
  xor g1923 (n_2074, n_703, n_704);
  xor g1924 (n_707, n_2074, n_705);
  nand g1925 (n_2075, n_703, n_704);
  nand g1926 (n_2076, n_705, n_704);
  nand g1927 (n_2077, n_703, n_705);
  nand g1928 (n_722, n_2075, n_2076, n_2077);
  xor g1929 (n_2078, n_706, n_707);
  xor g1930 (n_180, n_2078, n_708);
  nand g1931 (n_2079, n_706, n_707);
  nand g1932 (n_2080, n_708, n_707);
  nand g1933 (n_2081, n_706, n_708);
  nand g1934 (n_99, n_2079, n_2080, n_2081);
  xor g1935 (n_2082, A[42], A[40]);
  xor g1936 (n_713, n_2082, A[36]);
  nand g1937 (n_2083, A[42], A[40]);
  nand g1938 (n_2084, A[36], A[40]);
  nand g1939 (n_2085, A[42], A[36]);
  nand g1940 (n_723, n_2083, n_2084, n_2085);
  xor g1942 (n_714, n_1634, A[34]);
  nand g1944 (n_2088, A[34], A[26]);
  nand g1946 (n_724, n_1635, n_2088, n_1829);
  xor g1947 (n_2090, A[24], A[38]);
  xor g1948 (n_712, n_2090, A[32]);
  nand g1949 (n_2091, A[24], A[38]);
  nand g1952 (n_725, n_2091, n_1957, n_2024);
  xor g1953 (n_2094, A[30], n_709);
  xor g1954 (n_716, n_2094, n_710);
  nand g1955 (n_2095, A[30], n_709);
  nand g1956 (n_2096, n_710, n_709);
  nand g1957 (n_2097, A[30], n_710);
  nand g1958 (n_729, n_2095, n_2096, n_2097);
  xor g1959 (n_2098, n_711, n_712);
  xor g1960 (n_718, n_2098, n_713);
  nand g1961 (n_2099, n_711, n_712);
  nand g1962 (n_2100, n_713, n_712);
  nand g1963 (n_2101, n_711, n_713);
  nand g1964 (n_731, n_2099, n_2100, n_2101);
  xor g1965 (n_2102, n_714, n_715);
  xor g1966 (n_720, n_2102, n_716);
  nand g1967 (n_2103, n_714, n_715);
  nand g1968 (n_2104, n_716, n_715);
  nand g1969 (n_2105, n_714, n_716);
  nand g1970 (n_733, n_2103, n_2104, n_2105);
  xor g1971 (n_2106, n_717, n_718);
  xor g1972 (n_721, n_2106, n_719);
  nand g1973 (n_2107, n_717, n_718);
  nand g1974 (n_2108, n_719, n_718);
  nand g1975 (n_2109, n_717, n_719);
  nand g1976 (n_736, n_2107, n_2108, n_2109);
  xor g1977 (n_2110, n_720, n_721);
  xor g1978 (n_179, n_2110, n_722);
  nand g1979 (n_2111, n_720, n_721);
  nand g1980 (n_2112, n_722, n_721);
  nand g1981 (n_2113, n_720, n_722);
  nand g1982 (n_98, n_2111, n_2112, n_2113);
  xor g1983 (n_2114, A[43], A[41]);
  xor g1984 (n_727, n_2114, A[37]);
  nand g1985 (n_2115, A[43], A[41]);
  nand g1986 (n_2116, A[37], A[41]);
  nand g1987 (n_2117, A[43], A[37]);
  nand g1988 (n_737, n_2115, n_2116, n_2117);
  xor g1990 (n_728, n_1666, A[35]);
  nand g1992 (n_2120, A[35], A[27]);
  nand g1994 (n_738, n_1667, n_2120, n_1861);
  xor g1995 (n_2122, A[25], A[39]);
  xor g1996 (n_726, n_2122, A[33]);
  nand g1997 (n_2123, A[25], A[39]);
  nand g2000 (n_739, n_2123, n_1989, n_2056);
  xor g2001 (n_2126, A[31], n_723);
  xor g2002 (n_730, n_2126, n_724);
  nand g2003 (n_2127, A[31], n_723);
  nand g2004 (n_2128, n_724, n_723);
  nand g2005 (n_2129, A[31], n_724);
  nand g2006 (n_743, n_2127, n_2128, n_2129);
  xor g2007 (n_2130, n_725, n_726);
  xor g2008 (n_732, n_2130, n_727);
  nand g2009 (n_2131, n_725, n_726);
  nand g2010 (n_2132, n_727, n_726);
  nand g2011 (n_2133, n_725, n_727);
  nand g2012 (n_745, n_2131, n_2132, n_2133);
  xor g2013 (n_2134, n_728, n_729);
  xor g2014 (n_734, n_2134, n_730);
  nand g2015 (n_2135, n_728, n_729);
  nand g2016 (n_2136, n_730, n_729);
  nand g2017 (n_2137, n_728, n_730);
  nand g2018 (n_747, n_2135, n_2136, n_2137);
  xor g2019 (n_2138, n_731, n_732);
  xor g2020 (n_735, n_2138, n_733);
  nand g2021 (n_2139, n_731, n_732);
  nand g2022 (n_2140, n_733, n_732);
  nand g2023 (n_2141, n_731, n_733);
  nand g2024 (n_750, n_2139, n_2140, n_2141);
  xor g2025 (n_2142, n_734, n_735);
  xor g2026 (n_178, n_2142, n_736);
  nand g2027 (n_2143, n_734, n_735);
  nand g2028 (n_2144, n_736, n_735);
  nand g2029 (n_2145, n_734, n_736);
  nand g2030 (n_97, n_2143, n_2144, n_2145);
  xor g2031 (n_2146, A[44], A[42]);
  xor g2032 (n_741, n_2146, A[38]);
  nand g2033 (n_2147, A[44], A[42]);
  nand g2034 (n_2148, A[38], A[42]);
  nand g2035 (n_2149, A[44], A[38]);
  nand g2036 (n_751, n_2147, n_2148, n_2149);
  xor g2038 (n_742, n_1698, A[36]);
  nand g2040 (n_2152, A[36], A[28]);
  nand g2042 (n_752, n_1699, n_2152, n_1893);
  xor g2043 (n_2154, A[26], A[40]);
  xor g2044 (n_740, n_2154, A[34]);
  nand g2045 (n_2155, A[26], A[40]);
  nand g2048 (n_753, n_2155, n_2021, n_2088);
  xor g2049 (n_2158, A[32], n_737);
  xor g2050 (n_744, n_2158, n_738);
  nand g2051 (n_2159, A[32], n_737);
  nand g2052 (n_2160, n_738, n_737);
  nand g2053 (n_2161, A[32], n_738);
  nand g2054 (n_757, n_2159, n_2160, n_2161);
  xor g2055 (n_2162, n_739, n_740);
  xor g2056 (n_746, n_2162, n_741);
  nand g2057 (n_2163, n_739, n_740);
  nand g2058 (n_2164, n_741, n_740);
  nand g2059 (n_2165, n_739, n_741);
  nand g2060 (n_759, n_2163, n_2164, n_2165);
  xor g2061 (n_2166, n_742, n_743);
  xor g2062 (n_748, n_2166, n_744);
  nand g2063 (n_2167, n_742, n_743);
  nand g2064 (n_2168, n_744, n_743);
  nand g2065 (n_2169, n_742, n_744);
  nand g2066 (n_761, n_2167, n_2168, n_2169);
  xor g2067 (n_2170, n_745, n_746);
  xor g2068 (n_749, n_2170, n_747);
  nand g2069 (n_2171, n_745, n_746);
  nand g2070 (n_2172, n_747, n_746);
  nand g2071 (n_2173, n_745, n_747);
  nand g2072 (n_764, n_2171, n_2172, n_2173);
  xor g2073 (n_2174, n_748, n_749);
  xor g2074 (n_177, n_2174, n_750);
  nand g2075 (n_2175, n_748, n_749);
  nand g2076 (n_2176, n_750, n_749);
  nand g2077 (n_2177, n_748, n_750);
  nand g2078 (n_96, n_2175, n_2176, n_2177);
  xor g2079 (n_2178, A[45], A[43]);
  xor g2080 (n_755, n_2178, A[39]);
  nand g2081 (n_2179, A[45], A[43]);
  nand g2082 (n_2180, A[39], A[43]);
  nand g2083 (n_2181, A[45], A[39]);
  nand g2084 (n_765, n_2179, n_2180, n_2181);
  xor g2086 (n_756, n_1730, A[37]);
  nand g2088 (n_2184, A[37], A[29]);
  nand g2090 (n_766, n_1731, n_2184, n_1925);
  xor g2091 (n_2186, A[27], A[41]);
  xor g2092 (n_754, n_2186, A[35]);
  nand g2093 (n_2187, A[27], A[41]);
  nand g2096 (n_767, n_2187, n_2053, n_2120);
  xor g2097 (n_2190, A[33], n_751);
  xor g2098 (n_758, n_2190, n_752);
  nand g2099 (n_2191, A[33], n_751);
  nand g2100 (n_2192, n_752, n_751);
  nand g2101 (n_2193, A[33], n_752);
  nand g2102 (n_771, n_2191, n_2192, n_2193);
  xor g2103 (n_2194, n_753, n_754);
  xor g2104 (n_760, n_2194, n_755);
  nand g2105 (n_2195, n_753, n_754);
  nand g2106 (n_2196, n_755, n_754);
  nand g2107 (n_2197, n_753, n_755);
  nand g2108 (n_773, n_2195, n_2196, n_2197);
  xor g2109 (n_2198, n_756, n_757);
  xor g2110 (n_762, n_2198, n_758);
  nand g2111 (n_2199, n_756, n_757);
  nand g2112 (n_2200, n_758, n_757);
  nand g2113 (n_2201, n_756, n_758);
  nand g2114 (n_775, n_2199, n_2200, n_2201);
  xor g2115 (n_2202, n_759, n_760);
  xor g2116 (n_763, n_2202, n_761);
  nand g2117 (n_2203, n_759, n_760);
  nand g2118 (n_2204, n_761, n_760);
  nand g2119 (n_2205, n_759, n_761);
  nand g2120 (n_778, n_2203, n_2204, n_2205);
  xor g2121 (n_2206, n_762, n_763);
  xor g2122 (n_176, n_2206, n_764);
  nand g2123 (n_2207, n_762, n_763);
  nand g2124 (n_2208, n_764, n_763);
  nand g2125 (n_2209, n_762, n_764);
  nand g2126 (n_95, n_2207, n_2208, n_2209);
  xor g2127 (n_2210, A[46], A[44]);
  xor g2128 (n_769, n_2210, A[40]);
  nand g2129 (n_2211, A[46], A[44]);
  nand g2130 (n_2212, A[40], A[44]);
  nand g2131 (n_2213, A[46], A[40]);
  nand g2132 (n_779, n_2211, n_2212, n_2213);
  xor g2134 (n_770, n_1762, A[38]);
  nand g2136 (n_2216, A[38], A[30]);
  nand g2138 (n_780, n_1763, n_2216, n_1957);
  xor g2139 (n_2218, A[28], A[42]);
  xor g2140 (n_768, n_2218, A[36]);
  nand g2141 (n_2219, A[28], A[42]);
  nand g2144 (n_781, n_2219, n_2085, n_2152);
  xor g2145 (n_2222, A[34], n_765);
  xor g2146 (n_772, n_2222, n_766);
  nand g2147 (n_2223, A[34], n_765);
  nand g2148 (n_2224, n_766, n_765);
  nand g2149 (n_2225, A[34], n_766);
  nand g2150 (n_785, n_2223, n_2224, n_2225);
  xor g2151 (n_2226, n_767, n_768);
  xor g2152 (n_774, n_2226, n_769);
  nand g2153 (n_2227, n_767, n_768);
  nand g2154 (n_2228, n_769, n_768);
  nand g2155 (n_2229, n_767, n_769);
  nand g2156 (n_787, n_2227, n_2228, n_2229);
  xor g2157 (n_2230, n_770, n_771);
  xor g2158 (n_776, n_2230, n_772);
  nand g2159 (n_2231, n_770, n_771);
  nand g2160 (n_2232, n_772, n_771);
  nand g2161 (n_2233, n_770, n_772);
  nand g2162 (n_789, n_2231, n_2232, n_2233);
  xor g2163 (n_2234, n_773, n_774);
  xor g2164 (n_777, n_2234, n_775);
  nand g2165 (n_2235, n_773, n_774);
  nand g2166 (n_2236, n_775, n_774);
  nand g2167 (n_2237, n_773, n_775);
  nand g2168 (n_792, n_2235, n_2236, n_2237);
  xor g2169 (n_2238, n_776, n_777);
  xor g2170 (n_175, n_2238, n_778);
  nand g2171 (n_2239, n_776, n_777);
  nand g2172 (n_2240, n_778, n_777);
  nand g2173 (n_2241, n_776, n_778);
  nand g2174 (n_94, n_2239, n_2240, n_2241);
  xor g2175 (n_2242, A[47], A[45]);
  xor g2176 (n_783, n_2242, A[41]);
  nand g2177 (n_2243, A[47], A[45]);
  nand g2178 (n_2244, A[41], A[45]);
  nand g2179 (n_2245, A[47], A[41]);
  nand g2180 (n_793, n_2243, n_2244, n_2245);
  xor g2182 (n_784, n_1794, A[39]);
  nand g2184 (n_2248, A[39], A[31]);
  nand g2186 (n_795, n_1795, n_2248, n_1989);
  xor g2187 (n_2250, A[29], A[43]);
  xor g2188 (n_782, n_2250, A[37]);
  nand g2189 (n_2251, A[29], A[43]);
  nand g2192 (n_794, n_2251, n_2117, n_2184);
  xor g2193 (n_2254, A[35], n_779);
  xor g2194 (n_786, n_2254, n_780);
  nand g2195 (n_2255, A[35], n_779);
  nand g2196 (n_2256, n_780, n_779);
  nand g2197 (n_2257, A[35], n_780);
  nand g2198 (n_799, n_2255, n_2256, n_2257);
  xor g2199 (n_2258, n_781, n_782);
  xor g2200 (n_788, n_2258, n_783);
  nand g2201 (n_2259, n_781, n_782);
  nand g2202 (n_2260, n_783, n_782);
  nand g2203 (n_2261, n_781, n_783);
  nand g2204 (n_801, n_2259, n_2260, n_2261);
  xor g2205 (n_2262, n_784, n_785);
  xor g2206 (n_790, n_2262, n_786);
  nand g2207 (n_2263, n_784, n_785);
  nand g2208 (n_2264, n_786, n_785);
  nand g2209 (n_2265, n_784, n_786);
  nand g2210 (n_804, n_2263, n_2264, n_2265);
  xor g2211 (n_2266, n_787, n_788);
  xor g2212 (n_791, n_2266, n_789);
  nand g2213 (n_2267, n_787, n_788);
  nand g2214 (n_2268, n_789, n_788);
  nand g2215 (n_2269, n_787, n_789);
  nand g2216 (n_806, n_2267, n_2268, n_2269);
  xor g2217 (n_2270, n_790, n_791);
  xor g2218 (n_174, n_2270, n_792);
  nand g2219 (n_2271, n_790, n_791);
  nand g2220 (n_2272, n_792, n_791);
  nand g2221 (n_2273, n_790, n_792);
  nand g2222 (n_93, n_2271, n_2272, n_2273);
  xor g2223 (n_2274, A[46], A[42]);
  xor g2224 (n_797, n_2274, A[34]);
  nand g2225 (n_2275, A[46], A[42]);
  nand g2226 (n_2276, A[34], A[42]);
  nand g2227 (n_2277, A[46], A[34]);
  nand g2228 (n_807, n_2275, n_2276, n_2277);
  xor g2229 (n_2278, A[32], A[40]);
  xor g2230 (n_798, n_2278, A[30]);
  nand g2231 (n_2279, A[32], A[40]);
  nand g2232 (n_2280, A[30], A[40]);
  nand g2234 (n_809, n_2279, n_2280, n_1763);
  xor g2235 (n_2282, A[44], A[38]);
  xor g2236 (n_796, n_2282, A[36]);
  nand g2239 (n_2285, A[44], A[36]);
  nand g2240 (n_808, n_2149, n_1955, n_2285);
  xor g2241 (n_2286, A[48], n_793);
  xor g2242 (n_800, n_2286, n_794);
  nand g2243 (n_2287, A[48], n_793);
  nand g2244 (n_2288, n_794, n_793);
  nand g2245 (n_2289, A[48], n_794);
  nand g2246 (n_813, n_2287, n_2288, n_2289);
  xor g2247 (n_2290, n_795, n_796);
  xor g2248 (n_802, n_2290, n_797);
  nand g2249 (n_2291, n_795, n_796);
  nand g2250 (n_2292, n_797, n_796);
  nand g2251 (n_2293, n_795, n_797);
  nand g2252 (n_815, n_2291, n_2292, n_2293);
  xor g2253 (n_2294, n_798, n_799);
  xor g2254 (n_803, n_2294, n_800);
  nand g2255 (n_2295, n_798, n_799);
  nand g2256 (n_2296, n_800, n_799);
  nand g2257 (n_2297, n_798, n_800);
  nand g2258 (n_818, n_2295, n_2296, n_2297);
  xor g2259 (n_2298, n_801, n_802);
  xor g2260 (n_805, n_2298, n_803);
  nand g2261 (n_2299, n_801, n_802);
  nand g2262 (n_2300, n_803, n_802);
  nand g2263 (n_2301, n_801, n_803);
  nand g2264 (n_820, n_2299, n_2300, n_2301);
  xor g2265 (n_2302, n_804, n_805);
  xor g2266 (n_173, n_2302, n_806);
  nand g2267 (n_2303, n_804, n_805);
  nand g2268 (n_2304, n_806, n_805);
  nand g2269 (n_2305, n_804, n_806);
  nand g2270 (n_92, n_2303, n_2304, n_2305);
  xor g2271 (n_2306, A[47], A[43]);
  xor g2272 (n_811, n_2306, A[35]);
  nand g2273 (n_2307, A[47], A[43]);
  nand g2274 (n_2308, A[35], A[43]);
  nand g2275 (n_2309, A[47], A[35]);
  nand g2276 (n_822, n_2307, n_2308, n_2309);
  xor g2277 (n_2310, A[33], A[41]);
  xor g2278 (n_812, n_2310, A[31]);
  nand g2279 (n_2311, A[33], A[41]);
  nand g2280 (n_2312, A[31], A[41]);
  nand g2282 (n_823, n_2311, n_2312, n_1795);
  xor g2283 (n_2314, A[45], A[39]);
  xor g2284 (n_810, n_2314, A[37]);
  nand g2287 (n_2317, A[45], A[37]);
  nand g2288 (n_821, n_2181, n_1987, n_2317);
  xor g2289 (n_2318, A[49], n_807);
  xor g2290 (n_814, n_2318, n_808);
  nand g2291 (n_2319, A[49], n_807);
  nand g2292 (n_2320, n_808, n_807);
  nand g2293 (n_2321, A[49], n_808);
  nand g2294 (n_827, n_2319, n_2320, n_2321);
  xor g2295 (n_2322, n_809, n_810);
  xor g2296 (n_816, n_2322, n_811);
  nand g2297 (n_2323, n_809, n_810);
  nand g2298 (n_2324, n_811, n_810);
  nand g2299 (n_2325, n_809, n_811);
  nand g2300 (n_828, n_2323, n_2324, n_2325);
  xor g2301 (n_2326, n_812, n_813);
  xor g2302 (n_817, n_2326, n_814);
  nand g2303 (n_2327, n_812, n_813);
  nand g2304 (n_2328, n_814, n_813);
  nand g2305 (n_2329, n_812, n_814);
  nand g2306 (n_832, n_2327, n_2328, n_2329);
  xor g2307 (n_2330, n_815, n_816);
  xor g2308 (n_819, n_2330, n_817);
  nand g2309 (n_2331, n_815, n_816);
  nand g2310 (n_2332, n_817, n_816);
  nand g2311 (n_2333, n_815, n_817);
  nand g2312 (n_834, n_2331, n_2332, n_2333);
  xor g2313 (n_2334, n_818, n_819);
  xor g2314 (n_172, n_2334, n_820);
  nand g2315 (n_2335, n_818, n_819);
  nand g2316 (n_2336, n_820, n_819);
  nand g2317 (n_2337, n_818, n_820);
  nand g2318 (n_91, n_2335, n_2336, n_2337);
  xor g2320 (n_824, n_2210, A[36]);
  nand g2323 (n_2341, A[46], A[36]);
  nand g2324 (n_835, n_2211, n_2285, n_2341);
  xor g2325 (n_2342, A[34], A[42]);
  xor g2326 (n_826, n_2342, A[32]);
  nand g2328 (n_2344, A[32], A[42]);
  nand g2330 (n_836, n_2276, n_2344, n_1827);
  xor g2332 (n_825, n_2018, A[48]);
  nand g2334 (n_2348, A[48], A[38]);
  nand g2335 (n_2349, A[40], A[48]);
  nand g2336 (n_838, n_2019, n_2348, n_2349);
  xor g2337 (n_2350, A[50], n_821);
  xor g2338 (n_829, n_2350, n_822);
  nand g2339 (n_2351, A[50], n_821);
  nand g2340 (n_2352, n_822, n_821);
  nand g2341 (n_2353, A[50], n_822);
  nand g2342 (n_841, n_2351, n_2352, n_2353);
  xor g2343 (n_2354, n_823, n_824);
  xor g2344 (n_830, n_2354, n_825);
  nand g2345 (n_2355, n_823, n_824);
  nand g2346 (n_2356, n_825, n_824);
  nand g2347 (n_2357, n_823, n_825);
  nand g2348 (n_842, n_2355, n_2356, n_2357);
  xor g2349 (n_2358, n_826, n_827);
  xor g2350 (n_831, n_2358, n_828);
  nand g2351 (n_2359, n_826, n_827);
  nand g2352 (n_2360, n_828, n_827);
  nand g2353 (n_2361, n_826, n_828);
  nand g2354 (n_846, n_2359, n_2360, n_2361);
  xor g2355 (n_2362, n_829, n_830);
  xor g2356 (n_833, n_2362, n_831);
  nand g2357 (n_2363, n_829, n_830);
  nand g2358 (n_2364, n_831, n_830);
  nand g2359 (n_2365, n_829, n_831);
  nand g2360 (n_848, n_2363, n_2364, n_2365);
  xor g2361 (n_2366, n_832, n_833);
  xor g2362 (n_171, n_2366, n_834);
  nand g2363 (n_2367, n_832, n_833);
  nand g2364 (n_2368, n_834, n_833);
  nand g2365 (n_2369, n_832, n_834);
  nand g2366 (n_90, n_2367, n_2368, n_2369);
  xor g2368 (n_837, n_2242, A[37]);
  nand g2371 (n_2373, A[47], A[37]);
  nand g2372 (n_849, n_2243, n_2317, n_2373);
  xor g2373 (n_2374, A[35], A[43]);
  xor g2374 (n_840, n_2374, A[33]);
  nand g2376 (n_2376, A[33], A[43]);
  nand g2378 (n_850, n_2308, n_2376, n_1859);
  xor g2380 (n_839, n_2050, A[49]);
  nand g2382 (n_2380, A[49], A[39]);
  nand g2383 (n_2381, A[41], A[49]);
  nand g2384 (n_852, n_2051, n_2380, n_2381);
  xor g2385 (n_2382, A[51], n_835);
  xor g2386 (n_843, n_2382, n_836);
  nand g2387 (n_2383, A[51], n_835);
  nand g2388 (n_2384, n_836, n_835);
  nand g2389 (n_2385, A[51], n_836);
  nand g2390 (n_855, n_2383, n_2384, n_2385);
  xor g2391 (n_2386, n_837, n_838);
  xor g2392 (n_844, n_2386, n_839);
  nand g2393 (n_2387, n_837, n_838);
  nand g2394 (n_2388, n_839, n_838);
  nand g2395 (n_2389, n_837, n_839);
  nand g2396 (n_856, n_2387, n_2388, n_2389);
  xor g2397 (n_2390, n_840, n_841);
  xor g2398 (n_845, n_2390, n_842);
  nand g2399 (n_2391, n_840, n_841);
  nand g2400 (n_2392, n_842, n_841);
  nand g2401 (n_2393, n_840, n_842);
  nand g2402 (n_860, n_2391, n_2392, n_2393);
  xor g2403 (n_2394, n_843, n_844);
  xor g2404 (n_847, n_2394, n_845);
  nand g2405 (n_2395, n_843, n_844);
  nand g2406 (n_2396, n_845, n_844);
  nand g2407 (n_2397, n_843, n_845);
  nand g2408 (n_862, n_2395, n_2396, n_2397);
  xor g2409 (n_2398, n_846, n_847);
  xor g2410 (n_170, n_2398, n_848);
  nand g2411 (n_2399, n_846, n_847);
  nand g2412 (n_2400, n_848, n_847);
  nand g2413 (n_2401, n_846, n_848);
  nand g2414 (n_89, n_2399, n_2400, n_2401);
  xor g2416 (n_851, n_2210, A[38]);
  nand g2419 (n_2405, A[46], A[38]);
  nand g2420 (n_863, n_2211, n_2149, n_2405);
  xor g2422 (n_853, n_1890, A[42]);
  nand g2426 (n_864, n_1891, n_2276, n_2085);
  xor g2427 (n_2410, A[40], A[50]);
  xor g2428 (n_854, n_2410, A[52]);
  nand g2429 (n_2411, A[40], A[50]);
  nand g2430 (n_2412, A[52], A[50]);
  nand g2431 (n_2413, A[40], A[52]);
  nand g2432 (n_866, n_2411, n_2412, n_2413);
  xor g2433 (n_2414, A[48], n_849);
  xor g2434 (n_857, n_2414, n_850);
  nand g2435 (n_2415, A[48], n_849);
  nand g2436 (n_2416, n_850, n_849);
  nand g2437 (n_2417, A[48], n_850);
  nand g2438 (n_869, n_2415, n_2416, n_2417);
  xor g2439 (n_2418, n_851, n_852);
  xor g2440 (n_858, n_2418, n_853);
  nand g2441 (n_2419, n_851, n_852);
  nand g2442 (n_2420, n_853, n_852);
  nand g2443 (n_2421, n_851, n_853);
  nand g2444 (n_870, n_2419, n_2420, n_2421);
  xor g2445 (n_2422, n_854, n_855);
  xor g2446 (n_859, n_2422, n_856);
  nand g2447 (n_2423, n_854, n_855);
  nand g2448 (n_2424, n_856, n_855);
  nand g2449 (n_2425, n_854, n_856);
  nand g2450 (n_874, n_2423, n_2424, n_2425);
  xor g2451 (n_2426, n_857, n_858);
  xor g2452 (n_861, n_2426, n_859);
  nand g2453 (n_2427, n_857, n_858);
  nand g2454 (n_2428, n_859, n_858);
  nand g2455 (n_2429, n_857, n_859);
  nand g2456 (n_876, n_2427, n_2428, n_2429);
  xor g2457 (n_2430, n_860, n_861);
  xor g2458 (n_169, n_2430, n_862);
  nand g2459 (n_2431, n_860, n_861);
  nand g2460 (n_2432, n_862, n_861);
  nand g2461 (n_2433, n_860, n_862);
  nand g2462 (n_88, n_2431, n_2432, n_2433);
  xor g2464 (n_865, n_2242, A[39]);
  nand g2467 (n_2437, A[47], A[39]);
  nand g2468 (n_877, n_2243, n_2181, n_2437);
  xor g2470 (n_867, n_1922, A[43]);
  nand g2474 (n_878, n_1923, n_2308, n_2117);
  xor g2475 (n_2442, A[41], A[51]);
  xor g2476 (n_868, n_2442, A[53]);
  nand g2477 (n_2443, A[41], A[51]);
  nand g2478 (n_2444, A[53], A[51]);
  nand g2479 (n_2445, A[41], A[53]);
  nand g2480 (n_880, n_2443, n_2444, n_2445);
  xor g2481 (n_2446, A[49], n_863);
  xor g2482 (n_871, n_2446, n_864);
  nand g2483 (n_2447, A[49], n_863);
  nand g2484 (n_2448, n_864, n_863);
  nand g2485 (n_2449, A[49], n_864);
  nand g2486 (n_883, n_2447, n_2448, n_2449);
  xor g2487 (n_2450, n_865, n_866);
  xor g2488 (n_872, n_2450, n_867);
  nand g2489 (n_2451, n_865, n_866);
  nand g2490 (n_2452, n_867, n_866);
  nand g2491 (n_2453, n_865, n_867);
  nand g2492 (n_884, n_2451, n_2452, n_2453);
  xor g2493 (n_2454, n_868, n_869);
  xor g2494 (n_873, n_2454, n_870);
  nand g2495 (n_2455, n_868, n_869);
  nand g2496 (n_2456, n_870, n_869);
  nand g2497 (n_2457, n_868, n_870);
  nand g2498 (n_888, n_2455, n_2456, n_2457);
  xor g2499 (n_2458, n_871, n_872);
  xor g2500 (n_875, n_2458, n_873);
  nand g2501 (n_2459, n_871, n_872);
  nand g2502 (n_2460, n_873, n_872);
  nand g2503 (n_2461, n_871, n_873);
  nand g2504 (n_890, n_2459, n_2460, n_2461);
  xor g2505 (n_2462, n_874, n_875);
  xor g2506 (n_168, n_2462, n_876);
  nand g2507 (n_2463, n_874, n_875);
  nand g2508 (n_2464, n_876, n_875);
  nand g2509 (n_2465, n_874, n_876);
  nand g2510 (n_87, n_2463, n_2464, n_2465);
  xor g2511 (n_2466, A[46], A[40]);
  xor g2512 (n_879, n_2466, A[38]);
  nand g2516 (n_891, n_2213, n_2019, n_2405);
  xor g2517 (n_2470, A[36], A[44]);
  xor g2518 (n_881, n_2470, A[42]);
  nand g2522 (n_892, n_2285, n_2147, n_2085);
  xor g2523 (n_2474, A[48], A[54]);
  xor g2524 (n_882, n_2474, A[52]);
  nand g2525 (n_2475, A[48], A[54]);
  nand g2526 (n_2476, A[52], A[54]);
  nand g2527 (n_2477, A[48], A[52]);
  nand g2528 (n_894, n_2475, n_2476, n_2477);
  xor g2529 (n_2478, A[50], n_877);
  xor g2530 (n_885, n_2478, n_878);
  nand g2531 (n_2479, A[50], n_877);
  nand g2532 (n_2480, n_878, n_877);
  nand g2533 (n_2481, A[50], n_878);
  nand g2534 (n_897, n_2479, n_2480, n_2481);
  xor g2535 (n_2482, n_879, n_880);
  xor g2536 (n_886, n_2482, n_881);
  nand g2537 (n_2483, n_879, n_880);
  nand g2538 (n_2484, n_881, n_880);
  nand g2539 (n_2485, n_879, n_881);
  nand g2540 (n_898, n_2483, n_2484, n_2485);
  xor g2541 (n_2486, n_882, n_883);
  xor g2542 (n_887, n_2486, n_884);
  nand g2543 (n_2487, n_882, n_883);
  nand g2544 (n_2488, n_884, n_883);
  nand g2545 (n_2489, n_882, n_884);
  nand g2546 (n_902, n_2487, n_2488, n_2489);
  xor g2547 (n_2490, n_885, n_886);
  xor g2548 (n_889, n_2490, n_887);
  nand g2549 (n_2491, n_885, n_886);
  nand g2550 (n_2492, n_887, n_886);
  nand g2551 (n_2493, n_885, n_887);
  nand g2552 (n_904, n_2491, n_2492, n_2493);
  xor g2553 (n_2494, n_888, n_889);
  xor g2554 (n_167, n_2494, n_890);
  nand g2555 (n_2495, n_888, n_889);
  nand g2556 (n_2496, n_890, n_889);
  nand g2557 (n_2497, n_888, n_890);
  nand g2558 (n_86, n_2495, n_2496, n_2497);
  xor g2559 (n_2498, A[47], A[41]);
  xor g2560 (n_893, n_2498, A[39]);
  nand g2564 (n_905, n_2245, n_2051, n_2437);
  xor g2565 (n_2502, A[37], A[45]);
  xor g2566 (n_895, n_2502, A[43]);
  nand g2570 (n_906, n_2317, n_2179, n_2117);
  xor g2571 (n_2506, A[49], A[55]);
  xor g2572 (n_896, n_2506, A[53]);
  nand g2573 (n_2507, A[49], A[55]);
  nand g2574 (n_2508, A[53], A[55]);
  nand g2575 (n_2509, A[49], A[53]);
  nand g2576 (n_909, n_2507, n_2508, n_2509);
  xor g2577 (n_2510, A[51], n_891);
  xor g2578 (n_899, n_2510, n_892);
  nand g2579 (n_2511, A[51], n_891);
  nand g2580 (n_2512, n_892, n_891);
  nand g2581 (n_2513, A[51], n_892);
  nand g2582 (n_911, n_2511, n_2512, n_2513);
  xor g2583 (n_2514, n_893, n_894);
  xor g2584 (n_900, n_2514, n_895);
  nand g2585 (n_2515, n_893, n_894);
  nand g2586 (n_2516, n_895, n_894);
  nand g2587 (n_2517, n_893, n_895);
  nand g2588 (n_912, n_2515, n_2516, n_2517);
  xor g2589 (n_2518, n_896, n_897);
  xor g2590 (n_901, n_2518, n_898);
  nand g2591 (n_2519, n_896, n_897);
  nand g2592 (n_2520, n_898, n_897);
  nand g2593 (n_2521, n_896, n_898);
  nand g2594 (n_916, n_2519, n_2520, n_2521);
  xor g2595 (n_2522, n_899, n_900);
  xor g2596 (n_903, n_2522, n_901);
  nand g2597 (n_2523, n_899, n_900);
  nand g2598 (n_2524, n_901, n_900);
  nand g2599 (n_2525, n_899, n_901);
  nand g2600 (n_918, n_2523, n_2524, n_2525);
  xor g2601 (n_2526, n_902, n_903);
  xor g2602 (n_166, n_2526, n_904);
  nand g2603 (n_2527, n_902, n_903);
  nand g2604 (n_2528, n_904, n_903);
  nand g2605 (n_2529, n_902, n_904);
  nand g2606 (n_85, n_2527, n_2528, n_2529);
  xor g2608 (n_907, n_2274, A[40]);
  nand g2612 (n_919, n_2275, n_2083, n_2213);
  xor g2614 (n_908, n_2282, A[50]);
  nand g2616 (n_2536, A[50], A[44]);
  nand g2617 (n_2537, A[38], A[50]);
  nand g2618 (n_922, n_2149, n_2536, n_2537);
  xor g2625 (n_2542, A[56], n_905);
  xor g2626 (n_913, n_2542, n_906);
  nand g2627 (n_2543, A[56], n_905);
  nand g2628 (n_2544, n_906, n_905);
  nand g2629 (n_2545, A[56], n_906);
  nand g2630 (n_925, n_2543, n_2544, n_2545);
  xor g2631 (n_2546, n_907, n_908);
  xor g2632 (n_914, n_2546, n_909);
  nand g2633 (n_2547, n_907, n_908);
  nand g2634 (n_2548, n_909, n_908);
  nand g2635 (n_2549, n_907, n_909);
  nand g2636 (n_926, n_2547, n_2548, n_2549);
  xor g2637 (n_2550, n_882, n_911);
  xor g2638 (n_915, n_2550, n_912);
  nand g2639 (n_2551, n_882, n_911);
  nand g2640 (n_2552, n_912, n_911);
  nand g2641 (n_2553, n_882, n_912);
  nand g2642 (n_930, n_2551, n_2552, n_2553);
  xor g2643 (n_2554, n_913, n_914);
  xor g2644 (n_917, n_2554, n_915);
  nand g2645 (n_2555, n_913, n_914);
  nand g2646 (n_2556, n_915, n_914);
  nand g2647 (n_2557, n_913, n_915);
  nand g2648 (n_932, n_2555, n_2556, n_2557);
  xor g2649 (n_2558, n_916, n_917);
  xor g2650 (n_165, n_2558, n_918);
  nand g2651 (n_2559, n_916, n_917);
  nand g2652 (n_2560, n_918, n_917);
  nand g2653 (n_2561, n_916, n_918);
  nand g2654 (n_84, n_2559, n_2560, n_2561);
  xor g2656 (n_920, n_2306, A[41]);
  nand g2660 (n_933, n_2307, n_2115, n_2245);
  xor g2662 (n_921, n_2314, A[51]);
  nand g2664 (n_2568, A[51], A[45]);
  nand g2665 (n_2569, A[39], A[51]);
  nand g2666 (n_935, n_2181, n_2568, n_2569);
  xor g2673 (n_2574, A[57], n_919);
  xor g2674 (n_927, n_2574, n_920);
  nand g2675 (n_2575, A[57], n_919);
  nand g2676 (n_2576, n_920, n_919);
  nand g2677 (n_2577, A[57], n_920);
  nand g2678 (n_940, n_2575, n_2576, n_2577);
  xor g2679 (n_2578, n_921, n_922);
  xor g2680 (n_928, n_2578, n_894);
  nand g2681 (n_2579, n_921, n_922);
  nand g2682 (n_2580, n_894, n_922);
  nand g2683 (n_2581, n_921, n_894);
  nand g2684 (n_939, n_2579, n_2580, n_2581);
  xor g2685 (n_2582, n_896, n_925);
  xor g2686 (n_929, n_2582, n_926);
  nand g2687 (n_2583, n_896, n_925);
  nand g2688 (n_2584, n_926, n_925);
  nand g2689 (n_2585, n_896, n_926);
  nand g2690 (n_943, n_2583, n_2584, n_2585);
  xor g2691 (n_2586, n_927, n_928);
  xor g2692 (n_931, n_2586, n_929);
  nand g2693 (n_2587, n_927, n_928);
  nand g2694 (n_2588, n_929, n_928);
  nand g2695 (n_2589, n_927, n_929);
  nand g2696 (n_946, n_2587, n_2588, n_2589);
  xor g2697 (n_2590, n_930, n_931);
  xor g2698 (n_164, n_2590, n_932);
  nand g2699 (n_2591, n_930, n_931);
  nand g2700 (n_2592, n_932, n_931);
  nand g2701 (n_2593, n_930, n_932);
  nand g2702 (n_83, n_2591, n_2592, n_2593);
  xor g2704 (n_934, n_2210, A[42]);
  nand g2708 (n_947, n_2211, n_2147, n_2275);
  xor g2709 (n_2598, A[40], A[52]);
  xor g2710 (n_938, n_2598, A[56]);
  nand g2712 (n_2600, A[56], A[52]);
  nand g2713 (n_2601, A[40], A[56]);
  nand g2714 (n_949, n_2413, n_2600, n_2601);
  xor g2715 (n_2602, A[50], A[58]);
  xor g2716 (n_937, n_2602, A[48]);
  nand g2717 (n_2603, A[50], A[58]);
  nand g2718 (n_2604, A[48], A[58]);
  nand g2719 (n_2605, A[50], A[48]);
  nand g2720 (n_950, n_2603, n_2604, n_2605);
  xor g2721 (n_2606, A[54], n_933);
  xor g2722 (n_941, n_2606, n_934);
  nand g2723 (n_2607, A[54], n_933);
  nand g2724 (n_2608, n_934, n_933);
  nand g2725 (n_2609, A[54], n_934);
  nand g2726 (n_953, n_2607, n_2608, n_2609);
  xor g2727 (n_2610, n_935, n_909);
  xor g2728 (n_942, n_2610, n_937);
  nand g2729 (n_2611, n_935, n_909);
  nand g2730 (n_2612, n_937, n_909);
  nand g2731 (n_2613, n_935, n_937);
  nand g2732 (n_956, n_2611, n_2612, n_2613);
  xor g2733 (n_2614, n_938, n_939);
  xor g2734 (n_944, n_2614, n_940);
  nand g2735 (n_2615, n_938, n_939);
  nand g2736 (n_2616, n_940, n_939);
  nand g2737 (n_2617, n_938, n_940);
  nand g2738 (n_957, n_2615, n_2616, n_2617);
  xor g2739 (n_2618, n_941, n_942);
  xor g2740 (n_945, n_2618, n_943);
  nand g2741 (n_2619, n_941, n_942);
  nand g2742 (n_2620, n_943, n_942);
  nand g2743 (n_2621, n_941, n_943);
  nand g2744 (n_960, n_2619, n_2620, n_2621);
  xor g2745 (n_2622, n_944, n_945);
  xor g2746 (n_163, n_2622, n_946);
  nand g2747 (n_2623, n_944, n_945);
  nand g2748 (n_2624, n_946, n_945);
  nand g2749 (n_2625, n_944, n_946);
  nand g2750 (n_82, n_2623, n_2624, n_2625);
  xor g2752 (n_948, n_2242, A[43]);
  nand g2756 (n_963, n_2243, n_2179, n_2307);
  xor g2757 (n_2630, A[41], A[53]);
  xor g2758 (n_952, n_2630, A[57]);
  nand g2760 (n_2632, A[57], A[53]);
  nand g2761 (n_2633, A[41], A[57]);
  nand g2762 (n_966, n_2445, n_2632, n_2633);
  xor g2763 (n_2634, A[51], A[59]);
  xor g2764 (n_951, n_2634, A[49]);
  nand g2765 (n_2635, A[51], A[59]);
  nand g2766 (n_2636, A[49], A[59]);
  nand g2767 (n_2637, A[51], A[49]);
  nand g2768 (n_964, n_2635, n_2636, n_2637);
  xor g2769 (n_2638, A[55], n_947);
  xor g2770 (n_954, n_2638, n_948);
  nand g2771 (n_2639, A[55], n_947);
  nand g2772 (n_2640, n_948, n_947);
  nand g2773 (n_2641, A[55], n_948);
  nand g2774 (n_969, n_2639, n_2640, n_2641);
  xor g2775 (n_2642, n_949, n_950);
  xor g2776 (n_955, n_2642, n_951);
  nand g2777 (n_2643, n_949, n_950);
  nand g2778 (n_2644, n_951, n_950);
  nand g2779 (n_2645, n_949, n_951);
  nand g2780 (n_971, n_2643, n_2644, n_2645);
  xor g2781 (n_2646, n_952, n_953);
  xor g2782 (n_958, n_2646, n_954);
  nand g2783 (n_2647, n_952, n_953);
  nand g2784 (n_2648, n_954, n_953);
  nand g2785 (n_2649, n_952, n_954);
  nand g2786 (n_973, n_2647, n_2648, n_2649);
  xor g2787 (n_2650, n_955, n_956);
  xor g2788 (n_959, n_2650, n_957);
  nand g2789 (n_2651, n_955, n_956);
  nand g2790 (n_2652, n_957, n_956);
  nand g2791 (n_2653, n_955, n_957);
  nand g2792 (n_976, n_2651, n_2652, n_2653);
  xor g2793 (n_2654, n_958, n_959);
  xor g2794 (n_162, n_2654, n_960);
  nand g2795 (n_2655, n_958, n_959);
  nand g2796 (n_2656, n_960, n_959);
  nand g2797 (n_2657, n_958, n_960);
  nand g2798 (n_81, n_2655, n_2656, n_2657);
  xor g2801 (n_2658, A[60], A[44]);
  xor g2802 (n_965, n_2658, A[46]);
  nand g2803 (n_2659, A[60], A[44]);
  nand g2805 (n_2661, A[60], A[46]);
  nand g2806 (n_980, n_2659, n_2211, n_2661);
  xor g2807 (n_2662, A[42], A[58]);
  xor g2808 (n_967, n_2662, A[54]);
  nand g2809 (n_2663, A[42], A[58]);
  nand g2810 (n_2664, A[54], A[58]);
  nand g2811 (n_2665, A[42], A[54]);
  nand g2812 (n_983, n_2663, n_2664, n_2665);
  xor g2813 (n_2666, A[52], A[56]);
  xor g2814 (n_968, n_2666, A[50]);
  nand g2816 (n_2668, A[50], A[56]);
  nand g2818 (n_981, n_2600, n_2668, n_2412);
  xor g2819 (n_2670, A[48], n_963);
  xor g2820 (n_970, n_2670, n_964);
  nand g2821 (n_2671, A[48], n_963);
  nand g2822 (n_2672, n_964, n_963);
  nand g2823 (n_2673, A[48], n_964);
  nand g2824 (n_986, n_2671, n_2672, n_2673);
  xor g2825 (n_2674, n_965, n_966);
  xor g2826 (n_972, n_2674, n_967);
  nand g2827 (n_2675, n_965, n_966);
  nand g2828 (n_2676, n_967, n_966);
  nand g2829 (n_2677, n_965, n_967);
  nand g2830 (n_988, n_2675, n_2676, n_2677);
  xor g2831 (n_2678, n_968, n_969);
  xor g2832 (n_974, n_2678, n_970);
  nand g2833 (n_2679, n_968, n_969);
  nand g2834 (n_2680, n_970, n_969);
  nand g2835 (n_2681, n_968, n_970);
  nand g2836 (n_990, n_2679, n_2680, n_2681);
  xor g2837 (n_2682, n_971, n_972);
  xor g2838 (n_975, n_2682, n_973);
  nand g2839 (n_2683, n_971, n_972);
  nand g2840 (n_2684, n_973, n_972);
  nand g2841 (n_2685, n_971, n_973);
  nand g2842 (n_993, n_2683, n_2684, n_2685);
  xor g2843 (n_2686, n_974, n_975);
  xor g2844 (n_161, n_2686, n_976);
  nand g2845 (n_2687, n_974, n_975);
  nand g2846 (n_2688, n_976, n_975);
  nand g2847 (n_2689, n_974, n_976);
  nand g2848 (n_80, n_2687, n_2688, n_2689);
  xor g2852 (n_982, n_2306, A[60]);
  nand g2854 (n_2692, A[60], A[47]);
  nand g2855 (n_2693, A[43], A[60]);
  nand g2856 (n_995, n_2307, n_2692, n_2693);
  xor g2857 (n_2694, A[45], A[57]);
  xor g2858 (n_984, n_2694, A[53]);
  nand g2859 (n_2695, A[45], A[57]);
  nand g2861 (n_2697, A[45], A[53]);
  nand g2862 (n_997, n_2695, n_2632, n_2697);
  xor g2869 (n_2702, A[55], n_980);
  xor g2870 (n_987, n_2702, n_981);
  nand g2871 (n_2703, A[55], n_980);
  nand g2872 (n_2704, n_981, n_980);
  nand g2873 (n_2705, A[55], n_981);
  nand g2874 (n_1001, n_2703, n_2704, n_2705);
  xor g2875 (n_2706, n_982, n_983);
  xor g2876 (n_989, n_2706, n_984);
  nand g2877 (n_2707, n_982, n_983);
  nand g2878 (n_2708, n_984, n_983);
  nand g2879 (n_2709, n_982, n_984);
  nand g2880 (n_1004, n_2707, n_2708, n_2709);
  xor g2881 (n_2710, n_951, n_986);
  xor g2882 (n_991, n_2710, n_987);
  nand g2883 (n_2711, n_951, n_986);
  nand g2884 (n_2712, n_987, n_986);
  nand g2885 (n_2713, n_951, n_987);
  nand g2886 (n_1005, n_2711, n_2712, n_2713);
  xor g2887 (n_2714, n_988, n_989);
  xor g2888 (n_992, n_2714, n_990);
  nand g2889 (n_2715, n_988, n_989);
  nand g2890 (n_2716, n_990, n_989);
  nand g2891 (n_2717, n_988, n_990);
  nand g2892 (n_1008, n_2715, n_2716, n_2717);
  xor g2893 (n_2718, n_991, n_992);
  xor g2894 (n_160, n_2718, n_993);
  nand g2895 (n_2719, n_991, n_992);
  nand g2896 (n_2720, n_993, n_992);
  nand g2897 (n_2721, n_991, n_993);
  nand g2898 (n_79, n_2719, n_2720, n_2721);
  xor g2900 (n_996, n_2722, A[44]);
  nand g2904 (n_1011, n_2723, n_2211, n_2725);
  xor g2906 (n_1000, n_2726, A[58]);
  xor g2917 (n_2734, A[48], n_995);
  xor g2918 (n_1002, n_2734, n_996);
  nand g2919 (n_2735, A[48], n_995);
  nand g2920 (n_2736, n_996, n_995);
  nand g2921 (n_2737, A[48], n_996);
  nand g2922 (n_1017, n_2735, n_2736, n_2737);
  xor g2923 (n_2738, n_997, n_964);
  xor g2924 (n_1003, n_2738, n_968);
  nand g2925 (n_2739, n_997, n_964);
  nand g2926 (n_2740, n_968, n_964);
  nand g2927 (n_2741, n_997, n_968);
  nand g2928 (n_1019, n_2739, n_2740, n_2741);
  xor g2929 (n_2742, n_1000, n_1001);
  xor g2930 (n_1006, n_2742, n_1002);
  nand g2931 (n_2743, n_1000, n_1001);
  nand g2932 (n_2744, n_1002, n_1001);
  nand g2933 (n_2745, n_1000, n_1002);
  nand g2934 (n_1021, n_2743, n_2744, n_2745);
  xor g2935 (n_2746, n_1003, n_1004);
  xor g2936 (n_1007, n_2746, n_1005);
  nand g2937 (n_2747, n_1003, n_1004);
  nand g2938 (n_2748, n_1005, n_1004);
  nand g2939 (n_2749, n_1003, n_1005);
  nand g2940 (n_1023, n_2747, n_2748, n_2749);
  xor g2941 (n_2750, n_1006, n_1007);
  xor g2942 (n_159, n_2750, n_1008);
  nand g2943 (n_2751, n_1006, n_1007);
  nand g2944 (n_2752, n_1008, n_1007);
  nand g2945 (n_2753, n_1006, n_1008);
  nand g2946 (n_78, n_2751, n_2752, n_2753);
  xor g2949 (n_2754, A[45], A[53]);
  xor g2950 (n_1015, n_2754, A[57]);
  xor g2962 (n_1016, n_2762, n_1011);
  nand g2965 (n_2765, A[55], n_1011);
  nand g2966 (n_1030, n_2763, n_2764, n_2765);
  xor g2968 (n_1018, n_2766, n_951);
  nand g2970 (n_2768, n_951, n_981);
  nand g2971 (n_2769, n_1012, n_951);
  nand g2972 (n_1032, n_2767, n_2768, n_2769);
  xor g2973 (n_2770, n_1015, n_1016);
  xor g2974 (n_1020, n_2770, n_1017);
  nand g2975 (n_2771, n_1015, n_1016);
  nand g2976 (n_2772, n_1017, n_1016);
  nand g2977 (n_2773, n_1015, n_1017);
  nand g2978 (n_1034, n_2771, n_2772, n_2773);
  xor g2979 (n_2774, n_1018, n_1019);
  xor g2980 (n_1022, n_2774, n_1020);
  nand g2981 (n_2775, n_1018, n_1019);
  nand g2982 (n_2776, n_1020, n_1019);
  nand g2983 (n_2777, n_1018, n_1020);
  nand g2984 (n_1036, n_2775, n_2776, n_2777);
  xor g2985 (n_2778, n_1021, n_1022);
  xor g2986 (n_158, n_2778, n_1023);
  nand g2987 (n_2779, n_1021, n_1022);
  nand g2988 (n_2780, n_1023, n_1022);
  nand g2989 (n_2781, n_1021, n_1023);
  nand g2990 (n_77, n_2779, n_2780, n_2781);
  xor g2992 (n_1026, n_2722, A[58]);
  nand g2994 (n_2784, A[58], A[46]);
  nand g2996 (n_1039, n_2723, n_2784, n_2729);
  xor g2997 (n_2786, A[54], A[52]);
  xor g2998 (n_1029, n_2786, A[56]);
  nand g3001 (n_2789, A[54], A[56]);
  nand g3002 (n_1040, n_2476, n_2600, n_2789);
  xor g3003 (n_2790, A[50], A[48]);
  xor g3004 (n_1028, n_2790, A[47]);
  nand g3006 (n_2792, A[47], A[48]);
  nand g3007 (n_2793, A[50], A[47]);
  nand g3008 (n_1042, n_2605, n_2792, n_2793);
  xor g3009 (n_2794, n_964, n_1026);
  xor g3010 (n_1031, n_2794, n_997);
  nand g3011 (n_2795, n_964, n_1026);
  nand g3012 (n_2796, n_997, n_1026);
  nand g3014 (n_1044, n_2795, n_2796, n_2739);
  xor g3015 (n_2798, n_1028, n_1029);
  xor g3016 (n_1033, n_2798, n_1030);
  nand g3017 (n_2799, n_1028, n_1029);
  nand g3018 (n_2800, n_1030, n_1029);
  nand g3019 (n_2801, n_1028, n_1030);
  nand g3020 (n_1046, n_2799, n_2800, n_2801);
  xor g3021 (n_2802, n_1031, n_1032);
  xor g3022 (n_1035, n_2802, n_1033);
  nand g3023 (n_2803, n_1031, n_1032);
  nand g3024 (n_2804, n_1033, n_1032);
  nand g3025 (n_2805, n_1031, n_1033);
  nand g3026 (n_1049, n_2803, n_2804, n_2805);
  xor g3027 (n_2806, n_1034, n_1035);
  xor g3028 (n_157, n_2806, n_1036);
  nand g3029 (n_2807, n_1034, n_1035);
  nand g3030 (n_2808, n_1036, n_1035);
  nand g3031 (n_2809, n_1034, n_1036);
  nand g3032 (n_76, n_2807, n_2808, n_2809);
  xor g3035 (n_2810, A[57], A[53]);
  xor g3036 (n_1043, n_2810, A[51]);
  nand g3039 (n_2813, A[57], A[51]);
  nand g3040 (n_1051, n_2632, n_2444, n_2813);
  xor g3041 (n_2814, A[59], A[49]);
  xor g3042 (n_1041, n_2814, A[55]);
  nand g3045 (n_2817, A[59], A[55]);
  nand g3046 (n_1052, n_2636, n_2507, n_2817);
  xor g3048 (n_1045, n_2818, n_1040);
  nand g3050 (n_2820, n_1040, n_1039);
  nand g3052 (n_1056, n_2819, n_2820, n_2821);
  xor g3053 (n_2822, n_1041, n_1042);
  xor g3054 (n_1047, n_2822, n_1043);
  nand g3055 (n_2823, n_1041, n_1042);
  nand g3056 (n_2824, n_1043, n_1042);
  nand g3057 (n_2825, n_1041, n_1043);
  nand g3058 (n_1057, n_2823, n_2824, n_2825);
  xor g3059 (n_2826, n_1044, n_1045);
  xor g3060 (n_1048, n_2826, n_1046);
  nand g3061 (n_2827, n_1044, n_1045);
  nand g3062 (n_2828, n_1046, n_1045);
  nand g3063 (n_2829, n_1044, n_1046);
  nand g3064 (n_1060, n_2827, n_2828, n_2829);
  xor g3065 (n_2830, n_1047, n_1048);
  xor g3066 (n_156, n_2830, n_1049);
  nand g3067 (n_2831, n_1047, n_1048);
  nand g3068 (n_2832, n_1049, n_1048);
  nand g3069 (n_2833, n_1047, n_1049);
  nand g3070 (n_75, n_2831, n_2832, n_2833);
  xor g3072 (n_1054, n_2834, A[54]);
  nand g3076 (n_1012, n_2729, n_2664, n_2727);
  xor g3083 (n_2842, A[48], A[47]);
  xor g3084 (n_1055, n_2842, n_1051);
  nand g3086 (n_2844, n_1051, A[47]);
  nand g3087 (n_2845, A[48], n_1051);
  nand g3088 (n_1067, n_2792, n_2844, n_2845);
  xor g3089 (n_2846, n_1052, n_968);
  xor g3090 (n_1058, n_2846, n_1054);
  nand g3091 (n_2847, n_1052, n_968);
  nand g3092 (n_2848, n_1054, n_968);
  nand g3093 (n_2849, n_1052, n_1054);
  nand g3094 (n_1068, n_2847, n_2848, n_2849);
  xor g3095 (n_2850, n_1055, n_1056);
  xor g3096 (n_1059, n_2850, n_1057);
  nand g3097 (n_2851, n_1055, n_1056);
  nand g3098 (n_2852, n_1057, n_1056);
  nand g3099 (n_2853, n_1055, n_1057);
  nand g3100 (n_1071, n_2851, n_2852, n_2853);
  xor g3101 (n_2854, n_1058, n_1059);
  xor g3102 (n_155, n_2854, n_1060);
  nand g3103 (n_2855, n_1058, n_1059);
  nand g3104 (n_2856, n_1060, n_1059);
  nand g3105 (n_2857, n_1058, n_1060);
  nand g3106 (n_74, n_2855, n_2856, n_2857);
  xor g3109 (n_2858, A[53], A[51]);
  xor g3110 (n_1065, n_2858, A[59]);
  nand g3113 (n_2861, A[53], A[59]);
  nand g3114 (n_1073, n_2444, n_2635, n_2861);
  nand g3120 (n_1076, n_2507, n_2864, n_2865);
  xor g3121 (n_2766, n_981, n_1012);
  xor g3122 (n_1069, n_2766, n_1065);
  nand g3123 (n_2767, n_981, n_1012);
  nand g3124 (n_2868, n_1065, n_1012);
  nand g3125 (n_2869, n_981, n_1065);
  nand g3126 (n_1078, n_2767, n_2868, n_2869);
  xor g3127 (n_2870, n_1066, n_1067);
  xor g3128 (n_1070, n_2870, n_1068);
  nand g3129 (n_2871, n_1066, n_1067);
  nand g3130 (n_2872, n_1068, n_1067);
  nand g3131 (n_2873, n_1066, n_1068);
  nand g3132 (n_1080, n_2871, n_2872, n_2873);
  xor g3133 (n_2874, n_1069, n_1070);
  xor g3134 (n_154, n_2874, n_1071);
  nand g3135 (n_2875, n_1069, n_1070);
  nand g3136 (n_2876, n_1071, n_1070);
  nand g3137 (n_2877, n_1069, n_1071);
  nand g3138 (n_73, n_2875, n_2876, n_2877);
  xor g3151 (n_2886, A[57], n_1073);
  xor g3152 (n_1077, n_2886, n_968);
  nand g3153 (n_2887, A[57], n_1073);
  nand g3154 (n_2888, n_968, n_1073);
  nand g3155 (n_2889, A[57], n_968);
  nand g3156 (n_1087, n_2887, n_2888, n_2889);
  xor g3157 (n_2890, n_1054, n_1076);
  xor g3158 (n_1079, n_2890, n_1077);
  nand g3159 (n_2891, n_1054, n_1076);
  nand g3160 (n_2892, n_1077, n_1076);
  nand g3161 (n_2893, n_1054, n_1077);
  nand g3162 (n_1089, n_2891, n_2892, n_2893);
  xor g3163 (n_2894, n_1078, n_1079);
  xor g3164 (n_153, n_2894, n_1080);
  nand g3165 (n_2895, n_1078, n_1079);
  nand g3166 (n_2896, n_1080, n_1079);
  nand g3167 (n_2897, n_1078, n_1080);
  nand g3168 (n_72, n_2895, n_2896, n_2897);
  nand g3182 (n_1094, n_2864, n_2904, n_2705);
  xor g3183 (n_2906, n_1012, n_1065);
  xor g3184 (n_1088, n_2906, n_1086);
  nand g3186 (n_2908, n_1086, n_1065);
  nand g3187 (n_2909, n_1012, n_1086);
  nand g3188 (n_1096, n_2868, n_2908, n_2909);
  xor g3189 (n_2910, n_1087, n_1088);
  xor g3190 (n_152, n_2910, n_1089);
  nand g3191 (n_2911, n_1087, n_1088);
  nand g3192 (n_2912, n_1089, n_1088);
  nand g3193 (n_2913, n_1087, n_1089);
  nand g3194 (n_151, n_2911, n_2912, n_2913);
  xor g3202 (n_1093, n_2666, A[57]);
  nand g3204 (n_2920, A[57], A[56]);
  nand g3205 (n_2921, A[52], A[57]);
  nand g3206 (n_1101, n_2600, n_2920, n_2921);
  xor g3207 (n_2922, n_1073, n_1054);
  xor g3208 (n_1095, n_2922, n_1093);
  nand g3209 (n_2923, n_1073, n_1054);
  nand g3210 (n_2924, n_1093, n_1054);
  nand g3211 (n_2925, n_1073, n_1093);
  nand g3212 (n_1103, n_2923, n_2924, n_2925);
  xor g3213 (n_2926, n_1094, n_1095);
  xor g3214 (n_71, n_2926, n_1096);
  nand g3215 (n_2927, n_1094, n_1095);
  nand g3216 (n_2928, n_1096, n_1095);
  nand g3217 (n_2929, n_1094, n_1096);
  nand g3218 (n_150, n_2927, n_2928, n_2929);
  xor g3222 (n_1100, n_2810, A[55]);
  nand g3224 (n_2932, A[55], A[57]);
  nand g3226 (n_1105, n_2632, n_2932, n_2508);
  xor g3228 (n_1102, n_2934, n_1100);
  nand g3230 (n_2936, n_1100, n_1012);
  nand g3232 (n_1108, n_2935, n_2936, n_2937);
  xor g3233 (n_2938, n_1101, n_1102);
  xor g3234 (n_70, n_2938, n_1103);
  nand g3235 (n_2939, n_1101, n_1102);
  nand g3236 (n_2940, n_1103, n_1102);
  nand g3237 (n_2941, n_1101, n_1103);
  nand g3238 (n_149, n_2939, n_2940, n_2941);
  xor g3245 (n_2946, A[56], A[59]);
  xor g3246 (n_1107, n_2946, n_1105);
  nand g3247 (n_2947, A[56], A[59]);
  nand g3248 (n_2948, n_1105, A[59]);
  nand g3249 (n_2949, A[56], n_1105);
  nand g3250 (n_1113, n_2947, n_2948, n_2949);
  xor g3251 (n_2950, n_1054, n_1107);
  xor g3252 (n_69, n_2950, n_1108);
  nand g3253 (n_2951, n_1054, n_1107);
  nand g3254 (n_2952, n_1108, n_1107);
  nand g3255 (n_2953, n_1054, n_1108);
  nand g3256 (n_148, n_2951, n_2952, n_2953);
  xor g3259 (n_2954, A[57], A[55]);
  nand g3264 (n_1116, n_2932, n_2956, n_2957);
  xor g3265 (n_2958, n_1012, n_1112);
  xor g3266 (n_68, n_2958, n_1113);
  nand g3267 (n_2959, n_1012, n_1112);
  nand g3268 (n_2960, n_1113, n_1112);
  nand g3269 (n_2961, n_1012, n_1113);
  nand g3270 (n_147, n_2959, n_2960, n_2961);
  xor g3272 (n_1115, n_2834, A[56]);
  nand g3274 (n_2964, A[56], A[58]);
  nand g3276 (n_1119, n_2729, n_2964, n_2965);
  xor g3277 (n_2966, A[59], n_1115);
  xor g3278 (n_67, n_2966, n_1116);
  nand g3279 (n_2967, A[59], n_1115);
  nand g3280 (n_2968, n_1116, n_1115);
  nand g3281 (n_2969, A[59], n_1116);
  nand g3282 (n_146, n_2967, n_2968, n_2969);
  xor g3286 (n_66, n_2970, n_1119);
  nand g3289 (n_2973, A[59], n_1119);
  nand g3290 (n_145, n_2971, n_2972, n_2973);
  xor g3292 (n_65, n_2834, A[57]);
  nand g3294 (n_2976, A[57], A[58]);
  nand g3296 (n_144, n_2729, n_2976, n_2977);
  nor g11 (n_2993, A[2], A[0]);
  nor g13 (n_2989, A[1], A[3]);
  nor g15 (n_2999, A[2], n_217);
  nand g16 (n_2994, A[2], n_217);
  nor g17 (n_2995, n_136, n_216);
  nand g18 (n_2996, n_136, n_216);
  nor g19 (n_3005, n_135, n_215);
  nand g20 (n_3000, n_135, n_215);
  nor g21 (n_3001, n_134, n_214);
  nand g22 (n_3002, n_134, n_214);
  nor g23 (n_3011, n_133, n_213);
  nand g24 (n_3006, n_133, n_213);
  nor g25 (n_3007, n_132, n_212);
  nand g26 (n_3008, n_132, n_212);
  nor g27 (n_3017, n_131, n_211);
  nand g28 (n_3012, n_131, n_211);
  nor g29 (n_3013, n_130, n_210);
  nand g30 (n_3014, n_130, n_210);
  nor g31 (n_3023, n_129, n_209);
  nand g32 (n_3018, n_129, n_209);
  nor g33 (n_3019, n_128, n_208);
  nand g34 (n_3020, n_128, n_208);
  nor g35 (n_3029, n_127, n_207);
  nand g36 (n_3024, n_127, n_207);
  nor g37 (n_3025, n_126, n_206);
  nand g38 (n_3026, n_126, n_206);
  nor g39 (n_3035, n_125, n_205);
  nand g40 (n_3030, n_125, n_205);
  nor g41 (n_3031, n_124, n_204);
  nand g42 (n_3032, n_124, n_204);
  nor g43 (n_3041, n_123, n_203);
  nand g44 (n_3036, n_123, n_203);
  nor g45 (n_3037, n_122, n_202);
  nand g46 (n_3038, n_122, n_202);
  nor g47 (n_3047, n_121, n_201);
  nand g48 (n_3042, n_121, n_201);
  nor g49 (n_3043, n_120, n_200);
  nand g50 (n_3044, n_120, n_200);
  nor g51 (n_3053, n_119, n_199);
  nand g52 (n_3048, n_119, n_199);
  nor g53 (n_3049, n_118, n_198);
  nand g54 (n_3050, n_118, n_198);
  nor g55 (n_3059, n_117, n_197);
  nand g56 (n_3054, n_117, n_197);
  nor g57 (n_3055, n_116, n_196);
  nand g58 (n_3056, n_116, n_196);
  nor g59 (n_3065, n_115, n_195);
  nand g60 (n_3060, n_115, n_195);
  nor g61 (n_3061, n_114, n_194);
  nand g62 (n_3062, n_114, n_194);
  nor g63 (n_3071, n_113, n_193);
  nand g64 (n_3066, n_113, n_193);
  nor g65 (n_3067, n_112, n_192);
  nand g66 (n_3068, n_112, n_192);
  nor g67 (n_3077, n_111, n_191);
  nand g68 (n_3072, n_111, n_191);
  nor g69 (n_3073, n_110, n_190);
  nand g70 (n_3074, n_110, n_190);
  nor g71 (n_3083, n_109, n_189);
  nand g72 (n_3078, n_109, n_189);
  nor g73 (n_3079, n_108, n_188);
  nand g74 (n_3080, n_108, n_188);
  nor g75 (n_3089, n_107, n_187);
  nand g76 (n_3084, n_107, n_187);
  nor g77 (n_3085, n_106, n_186);
  nand g78 (n_3086, n_106, n_186);
  nor g79 (n_3095, n_105, n_185);
  nand g80 (n_3090, n_105, n_185);
  nor g81 (n_3091, n_104, n_184);
  nand g82 (n_3092, n_104, n_184);
  nor g83 (n_3101, n_103, n_183);
  nand g84 (n_3096, n_103, n_183);
  nor g85 (n_3097, n_102, n_182);
  nand g86 (n_3098, n_102, n_182);
  nor g87 (n_3107, n_101, n_181);
  nand g88 (n_3102, n_101, n_181);
  nor g89 (n_3103, n_100, n_180);
  nand g90 (n_3104, n_100, n_180);
  nor g91 (n_3113, n_99, n_179);
  nand g92 (n_3108, n_99, n_179);
  nor g93 (n_3109, n_98, n_178);
  nand g94 (n_3110, n_98, n_178);
  nor g95 (n_3119, n_97, n_177);
  nand g96 (n_3114, n_97, n_177);
  nor g97 (n_3115, n_96, n_176);
  nand g98 (n_3116, n_96, n_176);
  nor g99 (n_3125, n_95, n_175);
  nand g100 (n_3120, n_95, n_175);
  nor g101 (n_3121, n_94, n_174);
  nand g102 (n_3122, n_94, n_174);
  nor g103 (n_3131, n_93, n_173);
  nand g104 (n_3126, n_93, n_173);
  nor g105 (n_3127, n_92, n_172);
  nand g106 (n_3128, n_92, n_172);
  nor g107 (n_3137, n_91, n_171);
  nand g108 (n_3132, n_91, n_171);
  nor g109 (n_3133, n_90, n_170);
  nand g110 (n_3134, n_90, n_170);
  nor g111 (n_3143, n_89, n_169);
  nand g112 (n_3138, n_89, n_169);
  nor g113 (n_3139, n_88, n_168);
  nand g114 (n_3140, n_88, n_168);
  nor g115 (n_3149, n_87, n_167);
  nand g116 (n_3144, n_87, n_167);
  nor g117 (n_3145, n_86, n_166);
  nand g118 (n_3146, n_86, n_166);
  nor g119 (n_3155, n_85, n_165);
  nand g120 (n_3150, n_85, n_165);
  nor g121 (n_3151, n_84, n_164);
  nand g122 (n_3152, n_84, n_164);
  nor g123 (n_3161, n_83, n_163);
  nand g124 (n_3156, n_83, n_163);
  nor g125 (n_3157, n_82, n_162);
  nand g126 (n_3158, n_82, n_162);
  nor g127 (n_3167, n_81, n_161);
  nand g128 (n_3162, n_81, n_161);
  nor g129 (n_3163, n_80, n_160);
  nand g130 (n_3164, n_80, n_160);
  nor g131 (n_3173, n_79, n_159);
  nand g132 (n_3168, n_79, n_159);
  nor g133 (n_3169, n_78, n_158);
  nand g134 (n_3170, n_78, n_158);
  nor g135 (n_3179, n_77, n_157);
  nand g136 (n_3174, n_77, n_157);
  nor g137 (n_3175, n_76, n_156);
  nand g138 (n_3176, n_76, n_156);
  nor g139 (n_3185, n_75, n_155);
  nand g140 (n_3180, n_75, n_155);
  nor g141 (n_3181, n_74, n_154);
  nand g142 (n_3182, n_74, n_154);
  nor g143 (n_3191, n_73, n_153);
  nand g144 (n_3186, n_73, n_153);
  nor g145 (n_3187, n_72, n_152);
  nand g146 (n_3188, n_72, n_152);
  nor g147 (n_3197, n_71, n_151);
  nand g148 (n_3192, n_71, n_151);
  nor g149 (n_3193, n_70, n_150);
  nand g150 (n_3194, n_70, n_150);
  nor g151 (n_3203, n_69, n_149);
  nand g152 (n_3198, n_69, n_149);
  nor g153 (n_3199, n_68, n_148);
  nand g154 (n_3200, n_68, n_148);
  nor g155 (n_3209, n_67, n_147);
  nand g156 (n_3204, n_67, n_147);
  nor g157 (n_3205, n_66, n_146);
  nand g158 (n_3206, n_66, n_146);
  nor g159 (n_3215, n_65, n_145);
  nand g160 (n_3210, n_65, n_145);
  nor g170 (n_2991, n_1127, n_2989);
  nor g174 (n_2997, n_2994, n_2995);
  nor g177 (n_3230, n_2999, n_2995);
  nor g178 (n_3003, n_3000, n_3001);
  nor g181 (n_3224, n_3005, n_3001);
  nor g182 (n_3009, n_3006, n_3007);
  nor g185 (n_3237, n_3011, n_3007);
  nor g186 (n_3015, n_3012, n_3013);
  nor g189 (n_3231, n_3017, n_3013);
  nor g190 (n_3021, n_3018, n_3019);
  nor g193 (n_3244, n_3023, n_3019);
  nor g194 (n_3027, n_3024, n_3025);
  nor g197 (n_3238, n_3029, n_3025);
  nor g198 (n_3033, n_3030, n_3031);
  nor g201 (n_3251, n_3035, n_3031);
  nor g202 (n_3039, n_3036, n_3037);
  nor g205 (n_3245, n_3041, n_3037);
  nor g206 (n_3045, n_3042, n_3043);
  nor g209 (n_3258, n_3047, n_3043);
  nor g210 (n_3051, n_3048, n_3049);
  nor g213 (n_3252, n_3053, n_3049);
  nor g214 (n_3057, n_3054, n_3055);
  nor g217 (n_3265, n_3059, n_3055);
  nor g218 (n_3063, n_3060, n_3061);
  nor g221 (n_3259, n_3065, n_3061);
  nor g222 (n_3069, n_3066, n_3067);
  nor g225 (n_3272, n_3071, n_3067);
  nor g226 (n_3075, n_3072, n_3073);
  nor g229 (n_3266, n_3077, n_3073);
  nor g230 (n_3081, n_3078, n_3079);
  nor g233 (n_3279, n_3083, n_3079);
  nor g234 (n_3087, n_3084, n_3085);
  nor g237 (n_3273, n_3089, n_3085);
  nor g238 (n_3093, n_3090, n_3091);
  nor g241 (n_3286, n_3095, n_3091);
  nor g242 (n_3099, n_3096, n_3097);
  nor g245 (n_3280, n_3101, n_3097);
  nor g246 (n_3105, n_3102, n_3103);
  nor g249 (n_3293, n_3107, n_3103);
  nor g250 (n_3111, n_3108, n_3109);
  nor g253 (n_3287, n_3113, n_3109);
  nor g254 (n_3117, n_3114, n_3115);
  nor g257 (n_3300, n_3119, n_3115);
  nor g258 (n_3123, n_3120, n_3121);
  nor g261 (n_3294, n_3125, n_3121);
  nor g262 (n_3129, n_3126, n_3127);
  nor g265 (n_3307, n_3131, n_3127);
  nor g266 (n_3135, n_3132, n_3133);
  nor g269 (n_3301, n_3137, n_3133);
  nor g270 (n_3141, n_3138, n_3139);
  nor g273 (n_3314, n_3143, n_3139);
  nor g274 (n_3147, n_3144, n_3145);
  nor g277 (n_3308, n_3149, n_3145);
  nor g278 (n_3153, n_3150, n_3151);
  nor g281 (n_3321, n_3155, n_3151);
  nor g282 (n_3159, n_3156, n_3157);
  nor g285 (n_3315, n_3161, n_3157);
  nor g286 (n_3165, n_3162, n_3163);
  nor g289 (n_3328, n_3167, n_3163);
  nor g290 (n_3171, n_3168, n_3169);
  nor g293 (n_3322, n_3173, n_3169);
  nor g294 (n_3177, n_3174, n_3175);
  nor g297 (n_3335, n_3179, n_3175);
  nor g298 (n_3183, n_3180, n_3181);
  nor g301 (n_3329, n_3185, n_3181);
  nor g302 (n_3189, n_3186, n_3187);
  nor g305 (n_3342, n_3191, n_3187);
  nor g306 (n_3195, n_3192, n_3193);
  nor g309 (n_3336, n_3197, n_3193);
  nor g310 (n_3201, n_3198, n_3199);
  nor g313 (n_3349, n_3203, n_3199);
  nor g314 (n_3207, n_3204, n_3205);
  nor g317 (n_3343, n_3209, n_3205);
  nor g318 (n_3213, n_3210, n_3211);
  nor g321 (n_3351, n_3215, n_3211);
  nand g332 (n_3352, n_3230, n_3224);
  nand g337 (n_3362, n_3237, n_3231);
  nand g342 (n_3357, n_3244, n_3238);
  nand g347 (n_3368, n_3251, n_3245);
  nand g352 (n_3363, n_3258, n_3252);
  nand g357 (n_3374, n_3265, n_3259);
  nand g362 (n_3369, n_3272, n_3266);
  nand g367 (n_3380, n_3279, n_3273);
  nand g372 (n_3375, n_3286, n_3280);
  nand g377 (n_3386, n_3293, n_3287);
  nand g382 (n_3381, n_3300, n_3294);
  nand g387 (n_3392, n_3307, n_3301);
  nand g392 (n_3387, n_3314, n_3308);
  nand g397 (n_3398, n_3321, n_3315);
  nand g402 (n_3393, n_3328, n_3322);
  nand g407 (n_3404, n_3335, n_3329);
  nand g412 (n_3399, n_3342, n_3336);
  nand g417 (n_3406, n_3349, n_3343);
  nand g425 (n_3408, n_3355, n_3356);
  nor g426 (n_3360, n_3357, n_3358);
  nor g429 (n_3407, n_3362, n_3357);
  nor g430 (n_3366, n_3363, n_3364);
  nor g433 (n_3417, n_3368, n_3363);
  nor g434 (n_3372, n_3369, n_3370);
  nor g437 (n_3411, n_3374, n_3369);
  nor g438 (n_3378, n_3375, n_3376);
  nor g441 (n_3424, n_3380, n_3375);
  nor g442 (n_3384, n_3381, n_3382);
  nor g445 (n_3418, n_3386, n_3381);
  nor g446 (n_3390, n_3387, n_3388);
  nor g449 (n_3431, n_3392, n_3387);
  nor g450 (n_3396, n_3393, n_3394);
  nor g453 (n_3425, n_3398, n_3393);
  nor g454 (n_3402, n_3399, n_3400);
  nor g457 (n_3433, n_3404, n_3399);
  nand g462 (n_3410, n_3407, n_3408);
  nand g463 (n_3435, n_3409, n_3410);
  nand g468 (n_3434, n_3417, n_3411);
  nand g473 (n_3444, n_3424, n_3418);
  nand g478 (n_3439, n_3431, n_3425);
  nand g3306 (n_3446, n_3437, n_3438);
  nor g3307 (n_3442, n_3439, n_3440);
  nor g3310 (n_3445, n_3444, n_3439);
  nand g3311 (n_3448, n_3445, n_3446);
  nand g3312 (n_3451, n_3447, n_3448);
  nand g3315 (n_3454, n_3440, n_3450);
  nand g3316 (n_3452, n_3417, n_3435);
  nand g3317 (n_3461, n_3412, n_3452);
  nand g3318 (n_3453, n_3424, n_3446);
  nand g3319 (n_3466, n_3419, n_3453);
  nand g3320 (n_3455, n_3431, n_3454);
  nand g3321 (n_3471, n_3426, n_3455);
  nand g3322 (n_3456, n_3433, n_3451);
  nand g3323 (n_3476, n_3432, n_3456);
  nand g3326 (n_3481, n_3358, n_3458);
  nand g3329 (n_3484, n_3364, n_3460);
  nand g3332 (n_3487, n_3370, n_3463);
  nand g3335 (n_3490, n_3376, n_3465);
  nand g3338 (n_3493, n_3382, n_3468);
  nand g3341 (n_3496, n_3388, n_3470);
  nand g3344 (n_3499, n_3394, n_3473);
  nand g3347 (n_3502, n_3400, n_3475);
  nand g3350 (n_3505, n_3405, n_3478);
  nand g3352 (n_3511, n_3225, n_3479);
  nand g3353 (n_3480, n_3237, n_3408);
  nand g3354 (n_3516, n_3232, n_3480);
  nand g3355 (n_3482, n_3244, n_3481);
  nand g3356 (n_3521, n_3239, n_3482);
  nand g3357 (n_3483, n_3251, n_3435);
  nand g3358 (n_3526, n_3246, n_3483);
  nand g3359 (n_3485, n_3258, n_3484);
  nand g3360 (n_3531, n_3253, n_3485);
  nand g3361 (n_3486, n_3265, n_3461);
  nand g3362 (n_3536, n_3260, n_3486);
  nand g3363 (n_3488, n_3272, n_3487);
  nand g3364 (n_3541, n_3267, n_3488);
  nand g3365 (n_3489, n_3279, n_3446);
  nand g3366 (n_3546, n_3274, n_3489);
  nand g3367 (n_3491, n_3286, n_3490);
  nand g3368 (n_3551, n_3281, n_3491);
  nand g3369 (n_3492, n_3293, n_3466);
  nand g3370 (n_3556, n_3288, n_3492);
  nand g3371 (n_3494, n_3300, n_3493);
  nand g3372 (n_3561, n_3295, n_3494);
  nand g3373 (n_3495, n_3307, n_3454);
  nand g3374 (n_3566, n_3302, n_3495);
  nand g3375 (n_3497, n_3314, n_3496);
  nand g3376 (n_3571, n_3309, n_3497);
  nand g3377 (n_3498, n_3321, n_3471);
  nand g3378 (n_3576, n_3316, n_3498);
  nand g3379 (n_3500, n_3328, n_3499);
  nand g3380 (n_3581, n_3323, n_3500);
  nand g3381 (n_3501, n_3335, n_3451);
  nand g3382 (n_3586, n_3330, n_3501);
  nand g3383 (n_3503, n_3342, n_3502);
  nand g3384 (n_3591, n_3337, n_3503);
  nand g3385 (n_3504, n_3349, n_3476);
  nand g3386 (n_3596, n_3344, n_3504);
  nand g3387 (n_3506, n_3351, n_3505);
  nand g3388 (n_3601, n_3350, n_3506);
  nand g3394 (n_3611, n_2994, n_3510);
  nand g3397 (n_3615, n_3000, n_3513);
  nand g3400 (n_3619, n_3006, n_3515);
  nand g3403 (n_3623, n_3012, n_3518);
  nand g3406 (n_3627, n_3018, n_3520);
  nand g3409 (n_3631, n_3024, n_3523);
  nand g3412 (n_3635, n_3030, n_3525);
  nand g3415 (n_3639, n_3036, n_3528);
  nand g3418 (n_3643, n_3042, n_3530);
  nand g3421 (n_3647, n_3048, n_3533);
  nand g3424 (n_3651, n_3054, n_3535);
  nand g3427 (n_3655, n_3060, n_3538);
  nand g3430 (n_3659, n_3066, n_3540);
  nand g3433 (n_3663, n_3072, n_3543);
  nand g3436 (n_3667, n_3078, n_3545);
  nand g3439 (n_3671, n_3084, n_3548);
  nand g3442 (n_3675, n_3090, n_3550);
  nand g3445 (n_3679, n_3096, n_3553);
  nand g3448 (n_3683, n_3102, n_3555);
  nand g3451 (n_3687, n_3108, n_3558);
  nand g3454 (n_3691, n_3114, n_3560);
  nand g3457 (n_3695, n_3120, n_3563);
  nand g3460 (n_3699, n_3126, n_3565);
  nand g3463 (n_3703, n_3132, n_3568);
  nand g3466 (n_3707, n_3138, n_3570);
  nand g3469 (n_3711, n_3144, n_3573);
  nand g3472 (n_3715, n_3150, n_3575);
  nand g3475 (n_3719, n_3156, n_3578);
  nand g3478 (n_3723, n_3162, n_3580);
  nand g3481 (n_3727, n_3168, n_3583);
  nand g3484 (n_3731, n_3174, n_3585);
  nand g3487 (n_3735, n_3180, n_3588);
  nand g3490 (n_3739, n_3186, n_3590);
  nand g3493 (n_3743, n_3192, n_3593);
  nand g3496 (n_3747, n_3198, n_3595);
  nand g3499 (n_3751, n_3204, n_3598);
  nand g3502 (n_3755, n_3210, n_3600);
  nand g3505 (n_3759, n_3216, n_3603);
  xnor g3517 (Z[5], n_3611, n_3612);
  xnor g3519 (Z[6], n_3511, n_3613);
  xnor g3522 (Z[7], n_3615, n_3616);
  xnor g3524 (Z[8], n_3408, n_3617);
  xnor g3527 (Z[9], n_3619, n_3620);
  xnor g3529 (Z[10], n_3516, n_3621);
  xnor g3532 (Z[11], n_3623, n_3624);
  xnor g3534 (Z[12], n_3481, n_3625);
  xnor g3537 (Z[13], n_3627, n_3628);
  xnor g3539 (Z[14], n_3521, n_3629);
  xnor g3542 (Z[15], n_3631, n_3632);
  xnor g3544 (Z[16], n_3435, n_3633);
  xnor g3547 (Z[17], n_3635, n_3636);
  xnor g3549 (Z[18], n_3526, n_3637);
  xnor g3552 (Z[19], n_3639, n_3640);
  xnor g3554 (Z[20], n_3484, n_3641);
  xnor g3557 (Z[21], n_3643, n_3644);
  xnor g3559 (Z[22], n_3531, n_3645);
  xnor g3562 (Z[23], n_3647, n_3648);
  xnor g3564 (Z[24], n_3461, n_3649);
  xnor g3567 (Z[25], n_3651, n_3652);
  xnor g3569 (Z[26], n_3536, n_3653);
  xnor g3572 (Z[27], n_3655, n_3656);
  xnor g3574 (Z[28], n_3487, n_3657);
  xnor g3577 (Z[29], n_3659, n_3660);
  xnor g3579 (Z[30], n_3541, n_3661);
  xnor g3582 (Z[31], n_3663, n_3664);
  xnor g3584 (Z[32], n_3446, n_3665);
  xnor g3587 (Z[33], n_3667, n_3668);
  xnor g3589 (Z[34], n_3546, n_3669);
  xnor g3592 (Z[35], n_3671, n_3672);
  xnor g3594 (Z[36], n_3490, n_3673);
  xnor g3597 (Z[37], n_3675, n_3676);
  xnor g3599 (Z[38], n_3551, n_3677);
  xnor g3602 (Z[39], n_3679, n_3680);
  xnor g3604 (Z[40], n_3466, n_3681);
  xnor g3607 (Z[41], n_3683, n_3684);
  xnor g3609 (Z[42], n_3556, n_3685);
  xnor g3612 (Z[43], n_3687, n_3688);
  xnor g3614 (Z[44], n_3493, n_3689);
  xnor g3617 (Z[45], n_3691, n_3692);
  xnor g3619 (Z[46], n_3561, n_3693);
  xnor g3622 (Z[47], n_3695, n_3696);
  xnor g3624 (Z[48], n_3454, n_3697);
  xnor g3627 (Z[49], n_3699, n_3700);
  xnor g3629 (Z[50], n_3566, n_3701);
  xnor g3632 (Z[51], n_3703, n_3704);
  xnor g3634 (Z[52], n_3496, n_3705);
  xnor g3637 (Z[53], n_3707, n_3708);
  xnor g3639 (Z[54], n_3571, n_3709);
  xnor g3642 (Z[55], n_3711, n_3712);
  xnor g3644 (Z[56], n_3471, n_3713);
  xnor g3647 (Z[57], n_3715, n_3716);
  xnor g3649 (Z[58], n_3576, n_3717);
  xnor g3652 (Z[59], n_3719, n_3720);
  xnor g3654 (Z[60], n_3499, n_3721);
  xnor g3657 (Z[61], n_3723, n_3724);
  xnor g3659 (Z[62], n_3581, n_3725);
  xnor g3662 (Z[63], n_3727, n_3728);
  xnor g3664 (Z[64], n_3451, n_3729);
  xnor g3667 (Z[65], n_3731, n_3732);
  xnor g3669 (Z[66], n_3586, n_3733);
  xnor g3672 (Z[67], n_3735, n_3736);
  xnor g3674 (Z[68], n_3502, n_3737);
  xnor g3677 (Z[69], n_3739, n_3740);
  xnor g3679 (Z[70], n_3591, n_3741);
  xnor g3682 (Z[71], n_3743, n_3744);
  xnor g3684 (Z[72], n_3476, n_3745);
  xnor g3687 (Z[73], n_3747, n_3748);
  xnor g3689 (Z[74], n_3596, n_3749);
  xnor g3692 (Z[75], n_3751, n_3752);
  xnor g3694 (Z[76], n_3505, n_3753);
  xnor g3697 (Z[77], n_3755, n_3756);
  xnor g3699 (Z[78], n_3601, n_3757);
  or g3716 (n_310, wc, wc0, n_136);
  not gc0 (wc0, n_1127);
  not gc (wc, n_1141);
  or g3717 (n_319, wc1, wc2, n_304);
  not gc2 (wc2, n_1141);
  not gc1 (wc1, n_1160);
  or g3718 (n_332, wc3, n_309, n_304);
  not gc3 (wc3, n_1188);
  or g3719 (n_349, wc4, wc5, n_309);
  not gc5 (wc5, n_1223);
  not gc4 (wc4, n_1224);
  or g3720 (n_371, wc6, wc7, n_309);
  not gc7 (wc7, n_1271);
  not gc6 (wc6, n_1272);
  or g3721 (n_418, wc8, wc9, n_304);
  not gc9 (wc9, n_1272);
  not gc8 (wc8, n_1319);
  or g3722 (n_446, wc10, wc11, n_309);
  not gc11 (wc11, n_1448);
  not gc10 (wc10, n_1449);
  or g3723 (n_474, wc12, wc13, n_318);
  not gc13 (wc13, n_1388);
  not gc12 (wc12, n_1512);
  or g3724 (n_500, wc14, wc15, n_331);
  not gc15 (wc15, n_1452);
  not gc14 (wc14, n_1576);
  or g3725 (n_528, wc16, wc17, n_348);
  not gc17 (wc17, n_1381);
  not gc16 (wc16, n_1640);
  or g3726 (n_556, wc18, wc19, n_369);
  not gc19 (wc19, n_1445);
  not gc18 (wc18, n_1704);
  or g3727 (n_584, wc20, wc21, n_394);
  not gc21 (wc21, n_1509);
  not gc20 (wc20, n_1768);
  xnor g3728 (n_2722, A[60], A[46]);
  or g3729 (n_2723, wc22, A[60]);
  not gc22 (wc22, A[46]);
  or g3730 (n_2725, wc23, A[60]);
  not gc23 (wc23, A[44]);
  xnor g3731 (n_2762, A[55], A[47]);
  or g3732 (n_2763, A[47], wc24);
  not gc24 (wc24, A[55]);
  or g3733 (n_2729, wc25, A[60]);
  not gc25 (wc25, A[58]);
  xnor g3734 (n_2834, A[60], A[58]);
  or g3735 (n_2727, wc26, A[60]);
  not gc26 (wc26, A[54]);
  xnor g3736 (n_1066, n_2506, A[57]);
  or g3737 (n_2864, wc27, A[57]);
  not gc27 (wc27, A[55]);
  or g3738 (n_2865, wc28, A[57]);
  not gc28 (wc28, A[49]);
  xnor g3740 (n_1112, n_2954, A[59]);
  or g3741 (n_2956, wc29, A[59]);
  not gc29 (wc29, A[55]);
  or g3742 (n_2957, wc30, A[59]);
  not gc30 (wc30, A[57]);
  or g3743 (n_2965, wc31, A[60]);
  not gc31 (wc31, A[56]);
  xnor g3744 (n_2970, A[59], A[57]);
  or g3745 (n_2971, A[57], wc32);
  not gc32 (wc32, A[59]);
  or g3746 (n_2977, wc33, A[60]);
  not gc33 (wc33, A[57]);
  and g3747 (n_3219, wc34, A[60]);
  not gc34 (wc34, A[59]);
  or g3748 (n_3216, wc35, A[60]);
  not gc35 (wc35, A[59]);
  or g3749 (n_400, wc36, wc37, n_309);
  not gc37 (wc37, n_1328);
  not gc36 (wc36, n_1329);
  or g3750 (n_2821, A[47], wc38);
  not gc38 (wc38, n_1040);
  xnor g3751 (n_1086, n_981, n_2954);
  or g3752 (n_2904, A[57], wc39);
  not gc39 (wc39, n_981);
  or g3753 (n_2937, A[59], wc40);
  not gc40 (wc40, n_1100);
  and g3754 (n_3222, wc41, n_1123);
  not gc41 (wc41, n_2991);
  or g3756 (n_3605, n_2993, wc42);
  not gc42 (wc42, n_1127);
  or g3757 (n_3608, n_2989, wc43);
  not gc43 (wc43, n_1123);
  xnor g3758 (n_2726, A[60], A[54]);
  or g3759 (n_2764, A[47], wc44);
  not gc44 (wc44, n_1011);
  xnor g3760 (n_2818, n_1039, A[47]);
  or g3761 (n_2819, A[47], wc45);
  not gc45 (wc45, n_1039);
  xnor g3762 (n_2934, n_1012, A[59]);
  or g3763 (n_2935, A[59], wc46);
  not gc46 (wc46, n_1012);
  or g3764 (n_2972, A[57], wc47);
  not gc47 (wc47, n_1119);
  and g3765 (n_3211, A[59], wc48);
  not gc48 (wc48, n_144);
  or g3766 (n_3212, A[59], wc49);
  not gc49 (wc49, n_144);
  or g3767 (n_3609, wc50, n_2999);
  not gc50 (wc50, n_2994);
  or g3768 (n_3757, wc51, n_3219);
  not gc51 (wc51, n_3216);
  and g3769 (n_3225, wc52, n_2996);
  not gc52 (wc52, n_2997);
  not g3770 (Z[2], n_3605);
  or g3771 (n_3612, wc53, n_2995);
  not gc53 (wc53, n_2996);
  or g3772 (n_3613, wc54, n_3005);
  not gc54 (wc54, n_3000);
  and g3773 (n_3227, wc55, n_3002);
  not gc55 (wc55, n_3003);
  or g3776 (n_3616, wc56, n_3001);
  not gc56 (wc56, n_3002);
  or g3777 (n_3756, wc57, n_3211);
  not gc57 (wc57, n_3212);
  and g3778 (n_3232, wc58, n_3008);
  not gc58 (wc58, n_3009);
  and g3779 (n_3228, wc59, n_3224);
  not gc59 (wc59, n_3225);
  or g3780 (n_3479, n_3222, wc60);
  not gc60 (wc60, n_3230);
  or g3781 (n_3510, n_2999, n_3222);
  xor g3782 (Z[3], n_1127, n_3608);
  xor g3783 (Z[4], n_3222, n_3609);
  or g3784 (n_3617, wc61, n_3011);
  not gc61 (wc61, n_3006);
  or g3785 (n_3620, wc62, n_3007);
  not gc62 (wc62, n_3008);
  and g3786 (n_3350, n_3212, wc63);
  not gc63 (wc63, n_3213);
  and g3787 (n_3355, wc64, n_3227);
  not gc64 (wc64, n_3228);
  or g3788 (n_3356, n_3352, n_3222);
  or g3789 (n_3621, wc65, n_3017);
  not gc65 (wc65, n_3012);
  or g3790 (n_3752, wc66, n_3205);
  not gc66 (wc66, n_3206);
  or g3791 (n_3753, wc67, n_3215);
  not gc67 (wc67, n_3210);
  and g3792 (n_3234, wc68, n_3014);
  not gc68 (wc68, n_3015);
  and g3793 (n_3239, wc69, n_3020);
  not gc69 (wc69, n_3021);
  and g3794 (n_3346, wc70, n_3206);
  not gc70 (wc70, n_3207);
  or g3795 (n_3513, wc71, n_3005);
  not gc71 (wc71, n_3511);
  or g3796 (n_3624, wc72, n_3013);
  not gc72 (wc72, n_3014);
  or g3797 (n_3625, wc73, n_3023);
  not gc73 (wc73, n_3018);
  or g3798 (n_3628, wc74, n_3019);
  not gc74 (wc74, n_3020);
  or g3799 (n_3749, wc75, n_3209);
  not gc75 (wc75, n_3204);
  and g3800 (n_3241, wc76, n_3026);
  not gc76 (wc76, n_3027);
  and g3801 (n_3344, wc77, n_3200);
  not gc77 (wc77, n_3201);
  and g3802 (n_3235, wc78, n_3231);
  not gc78 (wc78, n_3232);
  or g3803 (n_3515, wc79, n_3011);
  not gc79 (wc79, n_3408);
  or g3804 (n_3629, wc80, n_3029);
  not gc80 (wc80, n_3024);
  or g3805 (n_3632, wc81, n_3025);
  not gc81 (wc81, n_3026);
  or g3806 (n_3744, wc82, n_3193);
  not gc82 (wc82, n_3194);
  or g3807 (n_3745, wc83, n_3203);
  not gc83 (wc83, n_3198);
  or g3808 (n_3748, wc84, n_3199);
  not gc84 (wc84, n_3200);
  and g3809 (n_3246, wc85, n_3032);
  not gc85 (wc85, n_3033);
  and g3810 (n_3248, wc86, n_3038);
  not gc86 (wc86, n_3039);
  and g3811 (n_3339, wc87, n_3194);
  not gc87 (wc87, n_3195);
  and g3812 (n_3358, wc88, n_3234);
  not gc88 (wc88, n_3235);
  and g3813 (n_3242, wc89, n_3238);
  not gc89 (wc89, n_3239);
  and g3814 (n_3347, wc90, n_3343);
  not gc90 (wc90, n_3344);
  or g3815 (n_3458, wc91, n_3362);
  not gc91 (wc91, n_3408);
  or g3816 (n_3633, wc92, n_3035);
  not gc92 (wc92, n_3030);
  or g3817 (n_3636, wc93, n_3031);
  not gc93 (wc93, n_3032);
  or g3818 (n_3637, wc94, n_3041);
  not gc94 (wc94, n_3036);
  or g3819 (n_3640, wc95, n_3037);
  not gc95 (wc95, n_3038);
  or g3820 (n_3641, wc96, n_3047);
  not gc96 (wc96, n_3042);
  or g3821 (n_3741, wc97, n_3197);
  not gc97 (wc97, n_3192);
  and g3822 (n_3253, wc98, n_3044);
  not gc98 (wc98, n_3045);
  and g3823 (n_3337, wc99, n_3188);
  not gc99 (wc99, n_3189);
  and g3824 (n_3359, wc100, n_3241);
  not gc100 (wc100, n_3242);
  and g3825 (n_3249, wc101, n_3245);
  not gc101 (wc101, n_3246);
  and g3826 (n_3405, wc102, n_3346);
  not gc102 (wc102, n_3347);
  or g3827 (n_3518, wc103, n_3017);
  not gc103 (wc103, n_3516);
  or g3828 (n_3644, wc104, n_3043);
  not gc104 (wc104, n_3044);
  or g3829 (n_3645, wc105, n_3053);
  not gc105 (wc105, n_3048);
  or g3830 (n_3737, wc106, n_3191);
  not gc106 (wc106, n_3186);
  or g3831 (n_3740, wc107, n_3187);
  not gc107 (wc107, n_3188);
  and g3832 (n_3255, wc108, n_3050);
  not gc108 (wc108, n_3051);
  and g3833 (n_3260, wc109, n_3056);
  not gc109 (wc109, n_3057);
  and g3834 (n_3262, wc110, n_3062);
  not gc110 (wc110, n_3063);
  and g3835 (n_3267, wc111, n_3068);
  not gc111 (wc111, n_3069);
  and g3836 (n_3269, wc112, n_3074);
  not gc112 (wc112, n_3075);
  and g3837 (n_3274, wc113, n_3080);
  not gc113 (wc113, n_3081);
  and g3838 (n_3276, wc114, n_3086);
  not gc114 (wc114, n_3087);
  and g3839 (n_3281, wc115, n_3092);
  not gc115 (wc115, n_3093);
  and g3840 (n_3283, wc116, n_3098);
  not gc116 (wc116, n_3099);
  and g3841 (n_3288, wc117, n_3104);
  not gc117 (wc117, n_3105);
  and g3842 (n_3290, wc118, n_3110);
  not gc118 (wc118, n_3111);
  and g3843 (n_3295, wc119, n_3116);
  not gc119 (wc119, n_3117);
  and g3844 (n_3297, wc120, n_3122);
  not gc120 (wc120, n_3123);
  and g3845 (n_3302, wc121, n_3128);
  not gc121 (wc121, n_3129);
  and g3846 (n_3304, wc122, n_3134);
  not gc122 (wc122, n_3135);
  and g3847 (n_3309, wc123, n_3140);
  not gc123 (wc123, n_3141);
  and g3848 (n_3311, wc124, n_3146);
  not gc124 (wc124, n_3147);
  and g3849 (n_3316, wc125, n_3152);
  not gc125 (wc125, n_3153);
  and g3850 (n_3318, wc126, n_3158);
  not gc126 (wc126, n_3159);
  and g3851 (n_3323, wc127, n_3164);
  not gc127 (wc127, n_3165);
  and g3852 (n_3364, wc128, n_3248);
  not gc128 (wc128, n_3249);
  and g3853 (n_3340, wc129, n_3336);
  not gc129 (wc129, n_3337);
  or g3854 (n_3520, wc130, n_3023);
  not gc130 (wc130, n_3481);
  or g3855 (n_3648, wc131, n_3049);
  not gc131 (wc131, n_3050);
  or g3856 (n_3649, wc132, n_3059);
  not gc132 (wc132, n_3054);
  or g3857 (n_3652, wc133, n_3055);
  not gc133 (wc133, n_3056);
  or g3858 (n_3653, wc134, n_3065);
  not gc134 (wc134, n_3060);
  or g3859 (n_3656, wc135, n_3061);
  not gc135 (wc135, n_3062);
  or g3860 (n_3657, wc136, n_3071);
  not gc136 (wc136, n_3066);
  or g3861 (n_3660, wc137, n_3067);
  not gc137 (wc137, n_3068);
  or g3862 (n_3661, wc138, n_3077);
  not gc138 (wc138, n_3072);
  or g3863 (n_3664, wc139, n_3073);
  not gc139 (wc139, n_3074);
  or g3864 (n_3665, wc140, n_3083);
  not gc140 (wc140, n_3078);
  or g3865 (n_3668, wc141, n_3079);
  not gc141 (wc141, n_3080);
  or g3866 (n_3669, wc142, n_3089);
  not gc142 (wc142, n_3084);
  or g3867 (n_3672, wc143, n_3085);
  not gc143 (wc143, n_3086);
  or g3868 (n_3673, wc144, n_3095);
  not gc144 (wc144, n_3090);
  or g3869 (n_3676, wc145, n_3091);
  not gc145 (wc145, n_3092);
  or g3870 (n_3677, wc146, n_3101);
  not gc146 (wc146, n_3096);
  or g3871 (n_3680, wc147, n_3097);
  not gc147 (wc147, n_3098);
  or g3872 (n_3681, wc148, n_3107);
  not gc148 (wc148, n_3102);
  or g3873 (n_3684, wc149, n_3103);
  not gc149 (wc149, n_3104);
  or g3874 (n_3685, wc150, n_3113);
  not gc150 (wc150, n_3108);
  or g3875 (n_3688, wc151, n_3109);
  not gc151 (wc151, n_3110);
  or g3876 (n_3689, wc152, n_3119);
  not gc152 (wc152, n_3114);
  or g3877 (n_3692, wc153, n_3115);
  not gc153 (wc153, n_3116);
  or g3878 (n_3693, wc154, n_3125);
  not gc154 (wc154, n_3120);
  or g3879 (n_3696, wc155, n_3121);
  not gc155 (wc155, n_3122);
  or g3880 (n_3697, wc156, n_3131);
  not gc156 (wc156, n_3126);
  or g3881 (n_3700, wc157, n_3127);
  not gc157 (wc157, n_3128);
  or g3882 (n_3701, wc158, n_3137);
  not gc158 (wc158, n_3132);
  or g3883 (n_3704, wc159, n_3133);
  not gc159 (wc159, n_3134);
  or g3884 (n_3705, wc160, n_3143);
  not gc160 (wc160, n_3138);
  or g3885 (n_3708, wc161, n_3139);
  not gc161 (wc161, n_3140);
  or g3886 (n_3709, wc162, n_3149);
  not gc162 (wc162, n_3144);
  or g3887 (n_3712, wc163, n_3145);
  not gc163 (wc163, n_3146);
  or g3888 (n_3713, wc164, n_3155);
  not gc164 (wc164, n_3150);
  or g3889 (n_3716, wc165, n_3151);
  not gc165 (wc165, n_3152);
  or g3890 (n_3717, wc166, n_3161);
  not gc166 (wc166, n_3156);
  or g3891 (n_3720, wc167, n_3157);
  not gc167 (wc167, n_3158);
  or g3892 (n_3721, wc168, n_3167);
  not gc168 (wc168, n_3162);
  or g3893 (n_3724, wc169, n_3163);
  not gc169 (wc169, n_3164);
  and g3894 (n_3325, wc170, n_3170);
  not gc170 (wc170, n_3171);
  and g3895 (n_3332, wc171, n_3182);
  not gc171 (wc171, n_3183);
  and g3896 (n_3256, wc172, n_3252);
  not gc172 (wc172, n_3253);
  and g3897 (n_3263, wc173, n_3259);
  not gc173 (wc173, n_3260);
  and g3898 (n_3270, wc174, n_3266);
  not gc174 (wc174, n_3267);
  and g3899 (n_3277, wc175, n_3273);
  not gc175 (wc175, n_3274);
  and g3900 (n_3284, wc176, n_3280);
  not gc176 (wc176, n_3281);
  and g3901 (n_3291, wc177, n_3287);
  not gc177 (wc177, n_3288);
  and g3902 (n_3298, wc178, n_3294);
  not gc178 (wc178, n_3295);
  and g3903 (n_3305, wc179, n_3301);
  not gc179 (wc179, n_3302);
  and g3904 (n_3312, wc180, n_3308);
  not gc180 (wc180, n_3309);
  and g3905 (n_3319, wc181, n_3315);
  not gc181 (wc181, n_3316);
  and g3906 (n_3401, wc182, n_3339);
  not gc182 (wc182, n_3340);
  and g3907 (n_3409, n_3359, wc183);
  not gc183 (wc183, n_3360);
  or g3908 (n_3725, wc184, n_3173);
  not gc184 (wc184, n_3168);
  or g3909 (n_3728, wc185, n_3169);
  not gc185 (wc185, n_3170);
  or g3910 (n_3733, wc186, n_3185);
  not gc186 (wc186, n_3180);
  or g3911 (n_3736, wc187, n_3181);
  not gc187 (wc187, n_3182);
  and g3912 (n_3330, wc188, n_3176);
  not gc188 (wc188, n_3177);
  and g3913 (n_3365, wc189, n_3255);
  not gc189 (wc189, n_3256);
  and g3914 (n_3370, wc190, n_3262);
  not gc190 (wc190, n_3263);
  and g3915 (n_3371, wc191, n_3269);
  not gc191 (wc191, n_3270);
  and g3916 (n_3376, wc192, n_3276);
  not gc192 (wc192, n_3277);
  and g3917 (n_3377, wc193, n_3283);
  not gc193 (wc193, n_3284);
  and g3918 (n_3382, wc194, n_3290);
  not gc194 (wc194, n_3291);
  and g3919 (n_3383, wc195, n_3297);
  not gc195 (wc195, n_3298);
  and g3920 (n_3388, wc196, n_3304);
  not gc196 (wc196, n_3305);
  and g3921 (n_3389, wc197, n_3311);
  not gc197 (wc197, n_3312);
  and g3922 (n_3394, wc198, n_3318);
  not gc198 (wc198, n_3319);
  and g3923 (n_3326, wc199, n_3322);
  not gc199 (wc199, n_3323);
  or g3924 (n_3523, wc200, n_3029);
  not gc200 (wc200, n_3521);
  or g3925 (n_3729, wc201, n_3179);
  not gc201 (wc201, n_3174);
  or g3926 (n_3732, wc202, n_3175);
  not gc202 (wc202, n_3176);
  and g3927 (n_3395, wc203, n_3325);
  not gc203 (wc203, n_3326);
  and g3928 (n_3333, wc204, n_3329);
  not gc204 (wc204, n_3330);
  or g3929 (n_3460, wc205, n_3368);
  not gc205 (wc205, n_3435);
  or g3930 (n_3525, wc206, n_3035);
  not gc206 (wc206, n_3435);
  and g3931 (n_3400, wc207, n_3332);
  not gc207 (wc207, n_3333);
  and g3932 (n_3412, n_3365, wc208);
  not gc208 (wc208, n_3366);
  and g3933 (n_3414, n_3371, wc209);
  not gc209 (wc209, n_3372);
  and g3934 (n_3419, n_3377, wc210);
  not gc210 (wc210, n_3378);
  and g3935 (n_3421, n_3383, wc211);
  not gc211 (wc211, n_3384);
  and g3936 (n_3426, n_3389, wc212);
  not gc212 (wc212, n_3390);
  or g3937 (n_3438, n_3434, wc213);
  not gc213 (wc213, n_3435);
  and g3938 (n_3428, n_3395, wc214);
  not gc214 (wc214, n_3396);
  and g3939 (n_3415, wc215, n_3411);
  not gc215 (wc215, n_3412);
  and g3940 (n_3422, wc216, n_3418);
  not gc216 (wc216, n_3419);
  and g3941 (n_3429, wc217, n_3425);
  not gc217 (wc217, n_3426);
  or g3942 (n_3528, wc218, n_3041);
  not gc218 (wc218, n_3526);
  or g3943 (n_3530, wc219, n_3047);
  not gc219 (wc219, n_3484);
  and g3944 (n_3432, n_3401, wc220);
  not gc220 (wc220, n_3402);
  and g3945 (n_3437, wc221, n_3414);
  not gc221 (wc221, n_3415);
  and g3946 (n_3440, wc222, n_3421);
  not gc222 (wc222, n_3422);
  or g3947 (n_3463, wc223, n_3374);
  not gc223 (wc223, n_3461);
  or g3948 (n_3535, wc224, n_3059);
  not gc224 (wc224, n_3461);
  and g3949 (n_3441, wc225, n_3428);
  not gc225 (wc225, n_3429);
  or g3950 (n_3533, wc226, n_3053);
  not gc226 (wc226, n_3531);
  or g3951 (n_3450, wc227, n_3444);
  not gc227 (wc227, n_3446);
  or g3952 (n_3465, wc228, n_3380);
  not gc228 (wc228, n_3446);
  or g3953 (n_3538, wc229, n_3065);
  not gc229 (wc229, n_3536);
  or g3954 (n_3540, wc230, n_3071);
  not gc230 (wc230, n_3487);
  or g3955 (n_3545, wc231, n_3083);
  not gc231 (wc231, n_3446);
  and g3956 (n_3447, n_3441, wc232);
  not gc232 (wc232, n_3442);
  or g3957 (n_3468, wc233, n_3386);
  not gc233 (wc233, n_3466);
  or g3958 (n_3470, wc234, n_3392);
  not gc234 (wc234, n_3454);
  or g3959 (n_3543, wc235, n_3077);
  not gc235 (wc235, n_3541);
  or g3960 (n_3548, wc236, n_3089);
  not gc236 (wc236, n_3546);
  or g3961 (n_3550, wc237, n_3095);
  not gc237 (wc237, n_3490);
  or g3962 (n_3555, wc238, n_3107);
  not gc238 (wc238, n_3466);
  or g3963 (n_3565, wc239, n_3131);
  not gc239 (wc239, n_3454);
  or g3964 (n_3475, wc240, n_3404);
  not gc240 (wc240, n_3451);
  or g3965 (n_3585, wc241, n_3179);
  not gc241 (wc241, n_3451);
  or g3966 (n_3473, wc242, n_3398);
  not gc242 (wc242, n_3471);
  or g3967 (n_3553, wc243, n_3101);
  not gc243 (wc243, n_3551);
  or g3968 (n_3558, wc244, n_3113);
  not gc244 (wc244, n_3556);
  or g3969 (n_3560, wc245, n_3119);
  not gc245 (wc245, n_3493);
  or g3970 (n_3568, wc246, n_3137);
  not gc246 (wc246, n_3566);
  or g3971 (n_3570, wc247, n_3143);
  not gc247 (wc247, n_3496);
  or g3972 (n_3575, wc248, n_3155);
  not gc248 (wc248, n_3471);
  or g3973 (n_3478, wc249, n_3406);
  not gc249 (wc249, n_3476);
  or g3974 (n_3588, wc250, n_3185);
  not gc250 (wc250, n_3586);
  or g3975 (n_3590, wc251, n_3191);
  not gc251 (wc251, n_3502);
  or g3976 (n_3595, wc252, n_3203);
  not gc252 (wc252, n_3476);
  or g3977 (n_3563, wc253, n_3125);
  not gc253 (wc253, n_3561);
  or g3978 (n_3573, wc254, n_3149);
  not gc254 (wc254, n_3571);
  or g3979 (n_3578, wc255, n_3161);
  not gc255 (wc255, n_3576);
  or g3980 (n_3580, wc256, n_3167);
  not gc256 (wc256, n_3499);
  or g3981 (n_3593, wc257, n_3197);
  not gc257 (wc257, n_3591);
  or g3982 (n_3598, wc258, n_3209);
  not gc258 (wc258, n_3596);
  or g3983 (n_3600, wc259, n_3215);
  not gc259 (wc259, n_3505);
  or g3984 (n_3583, wc260, n_3173);
  not gc260 (wc260, n_3581);
  or g3985 (n_3603, n_3219, wc261);
  not gc261 (wc261, n_3601);
  not g3986 (Z[79], n_3759);
endmodule

module mult_signed_const_14241_GENERIC(A, Z);
  input [60:0] A;
  output [79:0] Z;
  wire [60:0] A;
  wire [79:0] Z;
  mult_signed_const_14241_GENERIC_REAL g1(.A ({A[60:2], A[0], A[0]}),
       .Z (Z));
endmodule

module mult_signed_const_14732_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [61:0] A;
  output [80:0] Z;
  wire [61:0] A;
  wire [80:0] Z;
  wire n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_143, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212;
  wire n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220;
  wire n_221, n_222, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593;
  wire n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601;
  wire n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609;
  wire n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617;
  wire n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681;
  wire n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697;
  wire n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705;
  wire n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721;
  wire n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729;
  wire n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737;
  wire n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745;
  wire n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753;
  wire n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761;
  wire n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769;
  wire n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777;
  wire n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785;
  wire n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793;
  wire n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801;
  wire n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809;
  wire n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817;
  wire n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825;
  wire n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833;
  wire n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841;
  wire n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865;
  wire n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873;
  wire n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897;
  wire n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905;
  wire n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913;
  wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
  wire n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929;
  wire n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937;
  wire n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945;
  wire n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953;
  wire n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961;
  wire n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969;
  wire n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977;
  wire n_978, n_979, n_982, n_983, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006;
  wire n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1014, n_1015;
  wire n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023;
  wire n_1024, n_1025, n_1026, n_1027, n_1030, n_1031, n_1032, n_1033;
  wire n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041;
  wire n_1042, n_1044, n_1045, n_1047, n_1048, n_1049, n_1050, n_1051;
  wire n_1052, n_1053, n_1054, n_1055, n_1059, n_1060, n_1061, n_1062;
  wire n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1070, n_1071;
  wire n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1084, n_1085;
  wire n_1086, n_1087, n_1088, n_1089, n_1090, n_1092, n_1095, n_1096;
  wire n_1097, n_1098, n_1099, n_1105, n_1106, n_1107, n_1108, n_1112;
  wire n_1113, n_1114, n_1115, n_1119, n_1120, n_1121, n_1122, n_1124;
  wire n_1126, n_1127, n_1131, n_1132, n_1134, n_1135, n_1138, n_1141;
  wire n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149;
  wire n_1150, n_1152, n_1153, n_1154, n_1155, n_1156, n_1160, n_1161;
  wire n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169;
  wire n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1179;
  wire n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188;
  wire n_1189, n_1190, n_1191, n_1192, n_1193, n_1197, n_1198, n_1199;
  wire n_1200, n_1201, n_1202, n_1203, n_1204, n_1207, n_1211, n_1212;
  wire n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220;
  wire n_1221, n_1222, n_1223, n_1224, n_1225, n_1229, n_1230, n_1231;
  wire n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239;
  wire n_1240, n_1241, n_1242, n_1243, n_1245, n_1246, n_1248, n_1249;
  wire n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257;
  wire n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265;
  wire n_1268, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
  wire n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285;
  wire n_1288, n_1289, n_1290, n_1291, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304;
  wire n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312;
  wire n_1313, n_1315, n_1317, n_1320, n_1321, n_1322, n_1323, n_1324;
  wire n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332;
  wire n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1340, n_1341;
  wire n_1343, n_1344, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352;
  wire n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360;
  wire n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368;
  wire n_1371, n_1373, n_1374, n_1377, n_1378, n_1379, n_1380, n_1381;
  wire n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
  wire n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397;
  wire n_1398, n_1399, n_1400, n_1405, n_1406, n_1407, n_1409, n_1410;
  wire n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418;
  wire n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426;
  wire n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1437, n_1438;
  wire n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448;
  wire n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456;
  wire n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464;
  wire n_1467, n_1468, n_1469, n_1470, n_1471, n_1473, n_1474, n_1475;
  wire n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483;
  wire n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491;
  wire n_1492, n_1493, n_1494, n_1495, n_1496, n_1499, n_1501, n_1502;
  wire n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512;
  wire n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520;
  wire n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528;
  wire n_1531, n_1533, n_1534, n_1537, n_1538, n_1539, n_1540, n_1541;
  wire n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557;
  wire n_1558, n_1559, n_1560, n_1563, n_1565, n_1566, n_1569, n_1570;
  wire n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578;
  wire n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586;
  wire n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1595, n_1597;
  wire n_1598, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607;
  wire n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615;
  wire n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623;
  wire n_1624, n_1627, n_1629, n_1630, n_1633, n_1634, n_1635, n_1636;
  wire n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644;
  wire n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652;
  wire n_1653, n_1654, n_1655, n_1656, n_1659, n_1661, n_1662, n_1665;
  wire n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673;
  wire n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681;
  wire n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1691;
  wire n_1693, n_1694, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702;
  wire n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710;
  wire n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718;
  wire n_1719, n_1720, n_1723, n_1725, n_1726, n_1729, n_1730, n_1731;
  wire n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739;
  wire n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747;
  wire n_1748, n_1749, n_1750, n_1751, n_1752, n_1755, n_1757, n_1758;
  wire n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768;
  wire n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776;
  wire n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784;
  wire n_1787, n_1789, n_1790, n_1793, n_1794, n_1795, n_1796, n_1797;
  wire n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805;
  wire n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813;
  wire n_1814, n_1815, n_1816, n_1819, n_1821, n_1822, n_1825, n_1826;
  wire n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834;
  wire n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842;
  wire n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1851, n_1853;
  wire n_1854, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863;
  wire n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871;
  wire n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879;
  wire n_1880, n_1883, n_1885, n_1886, n_1889, n_1890, n_1891, n_1892;
  wire n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900;
  wire n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908;
  wire n_1909, n_1910, n_1911, n_1912, n_1915, n_1917, n_1918, n_1921;
  wire n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929;
  wire n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937;
  wire n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1947;
  wire n_1949, n_1950, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958;
  wire n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966;
  wire n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974;
  wire n_1975, n_1976, n_1979, n_1981, n_1982, n_1985, n_1986, n_1987;
  wire n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995;
  wire n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003;
  wire n_2004, n_2005, n_2006, n_2007, n_2008, n_2011, n_2013, n_2014;
  wire n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024;
  wire n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032;
  wire n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040;
  wire n_2043, n_2045, n_2046, n_2049, n_2050, n_2051, n_2052, n_2053;
  wire n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061;
  wire n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069;
  wire n_2070, n_2071, n_2072, n_2075, n_2077, n_2078, n_2081, n_2082;
  wire n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090;
  wire n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098;
  wire n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2107, n_2109;
  wire n_2110, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119;
  wire n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127;
  wire n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135;
  wire n_2136, n_2139, n_2141, n_2142, n_2145, n_2146, n_2147, n_2148;
  wire n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156;
  wire n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164;
  wire n_2165, n_2166, n_2167, n_2168, n_2171, n_2173, n_2174, n_2177;
  wire n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185;
  wire n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193;
  wire n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2203;
  wire n_2205, n_2206, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214;
  wire n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222;
  wire n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230;
  wire n_2231, n_2232, n_2235, n_2237, n_2238, n_2241, n_2242, n_2243;
  wire n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251;
  wire n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259;
  wire n_2260, n_2261, n_2262, n_2263, n_2264, n_2267, n_2269, n_2270;
  wire n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280;
  wire n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288;
  wire n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296;
  wire n_2299, n_2301, n_2302, n_2305, n_2306, n_2307, n_2308, n_2309;
  wire n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317;
  wire n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325;
  wire n_2326, n_2327, n_2328, n_2331, n_2333, n_2334, n_2337, n_2338;
  wire n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346;
  wire n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354;
  wire n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2363, n_2365;
  wire n_2366, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375;
  wire n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383;
  wire n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391;
  wire n_2392, n_2395, n_2397, n_2398, n_2401, n_2402, n_2403, n_2404;
  wire n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412;
  wire n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420;
  wire n_2421, n_2422, n_2423, n_2424, n_2427, n_2429, n_2430, n_2433;
  wire n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441;
  wire n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449;
  wire n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2459;
  wire n_2461, n_2462, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470;
  wire n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478;
  wire n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486;
  wire n_2487, n_2488, n_2491, n_2493, n_2494, n_2497, n_2498, n_2499;
  wire n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507;
  wire n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515;
  wire n_2516, n_2517, n_2518, n_2519, n_2520, n_2523, n_2525, n_2526;
  wire n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536;
  wire n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544;
  wire n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552;
  wire n_2555, n_2557, n_2558, n_2561, n_2562, n_2563, n_2564, n_2565;
  wire n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573;
  wire n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581;
  wire n_2582, n_2583, n_2584, n_2587, n_2589, n_2590, n_2593, n_2594;
  wire n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602;
  wire n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610;
  wire n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2619, n_2621;
  wire n_2622, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631;
  wire n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639;
  wire n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647;
  wire n_2648, n_2651, n_2653, n_2654, n_2657, n_2658, n_2659, n_2660;
  wire n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668;
  wire n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676;
  wire n_2677, n_2678, n_2679, n_2680, n_2683, n_2685, n_2686, n_2689;
  wire n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697;
  wire n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, n_2705;
  wire n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713;
  wire n_2714, n_2715, n_2717, n_2721, n_2722, n_2723, n_2724, n_2725;
  wire n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733;
  wire n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, n_2741;
  wire n_2742, n_2744, n_2745, n_2746, n_2747, n_2748, n_2752, n_2753;
  wire n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761;
  wire n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769;
  wire n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, n_2779;
  wire n_2781, n_2782, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789;
  wire n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797;
  wire n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805;
  wire n_2806, n_2809, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818;
  wire n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826;
  wire n_2827, n_2828, n_2829, n_2830, n_2831, n_2832, n_2837, n_2840;
  wire n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850;
  wire n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, n_2858;
  wire n_2859, n_2860, n_2861, n_2865, n_2868, n_2869, n_2871, n_2872;
  wire n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880;
  wire n_2881, n_2882, n_2883, n_2884, n_2893, n_2895, n_2896, n_2897;
  wire n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905;
  wire n_2906, n_2907, n_2908, n_2915, n_2916, n_2917, n_2918, n_2919;
  wire n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927;
  wire n_2928, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943;
  wire n_2944, n_2945, n_2946, n_2947, n_2948, n_2955, n_2956, n_2957;
  wire n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2971, n_2972;
  wire n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980;
  wire n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, n_2997, n_2998;
  wire n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3007, n_3008;
  wire n_3009, n_3010, n_3011, n_3012, n_3017, n_3018, n_3019, n_3020;
  wire n_3022, n_3023, n_3024, n_3027, n_3028, n_3040, n_3042, n_3044;
  wire n_3045, n_3046, n_3047, n_3048, n_3050, n_3051, n_3052, n_3053;
  wire n_3054, n_3056, n_3057, n_3058, n_3059, n_3060, n_3062, n_3063;
  wire n_3064, n_3065, n_3066, n_3068, n_3069, n_3070, n_3071, n_3072;
  wire n_3074, n_3075, n_3076, n_3077, n_3078, n_3080, n_3081, n_3082;
  wire n_3083, n_3084, n_3086, n_3087, n_3088, n_3089, n_3090, n_3092;
  wire n_3093, n_3094, n_3095, n_3096, n_3098, n_3099, n_3100, n_3101;
  wire n_3102, n_3104, n_3105, n_3106, n_3107, n_3108, n_3110, n_3111;
  wire n_3112, n_3113, n_3114, n_3116, n_3117, n_3118, n_3119, n_3120;
  wire n_3122, n_3123, n_3124, n_3125, n_3126, n_3128, n_3129, n_3130;
  wire n_3131, n_3132, n_3134, n_3135, n_3136, n_3137, n_3138, n_3140;
  wire n_3141, n_3142, n_3143, n_3144, n_3146, n_3147, n_3148, n_3149;
  wire n_3150, n_3152, n_3153, n_3154, n_3155, n_3156, n_3158, n_3159;
  wire n_3160, n_3161, n_3162, n_3164, n_3165, n_3166, n_3167, n_3168;
  wire n_3170, n_3171, n_3172, n_3173, n_3174, n_3176, n_3177, n_3178;
  wire n_3179, n_3180, n_3182, n_3183, n_3184, n_3185, n_3186, n_3188;
  wire n_3189, n_3190, n_3191, n_3192, n_3194, n_3195, n_3196, n_3197;
  wire n_3198, n_3200, n_3201, n_3202, n_3203, n_3204, n_3206, n_3207;
  wire n_3208, n_3209, n_3210, n_3212, n_3213, n_3214, n_3215, n_3216;
  wire n_3218, n_3219, n_3220, n_3221, n_3222, n_3224, n_3225, n_3226;
  wire n_3227, n_3228, n_3230, n_3231, n_3232, n_3233, n_3234, n_3236;
  wire n_3237, n_3238, n_3239, n_3240, n_3242, n_3243, n_3244, n_3245;
  wire n_3246, n_3248, n_3249, n_3250, n_3251, n_3252, n_3254, n_3255;
  wire n_3256, n_3257, n_3258, n_3260, n_3261, n_3262, n_3263, n_3264;
  wire n_3266, n_3267, n_3268, n_3269, n_3270, n_3272, n_3275, n_3277;
  wire n_3278, n_3280, n_3281, n_3283, n_3284, n_3285, n_3287, n_3288;
  wire n_3290, n_3291, n_3292, n_3294, n_3295, n_3297, n_3298, n_3299;
  wire n_3301, n_3302, n_3304, n_3305, n_3306, n_3308, n_3309, n_3311;
  wire n_3312, n_3313, n_3315, n_3316, n_3318, n_3319, n_3320, n_3322;
  wire n_3323, n_3325, n_3326, n_3327, n_3329, n_3330, n_3332, n_3333;
  wire n_3334, n_3336, n_3337, n_3339, n_3340, n_3341, n_3343, n_3344;
  wire n_3346, n_3347, n_3348, n_3350, n_3351, n_3353, n_3354, n_3355;
  wire n_3357, n_3358, n_3360, n_3361, n_3362, n_3364, n_3365, n_3367;
  wire n_3368, n_3369, n_3371, n_3372, n_3374, n_3375, n_3376, n_3378;
  wire n_3379, n_3381, n_3382, n_3383, n_3385, n_3386, n_3388, n_3389;
  wire n_3390, n_3392, n_3393, n_3395, n_3396, n_3397, n_3399, n_3400;
  wire n_3402, n_3403, n_3404, n_3406, n_3407, n_3409, n_3410, n_3413;
  wire n_3414, n_3415, n_3416, n_3417, n_3418, n_3420, n_3421, n_3422;
  wire n_3423, n_3424, n_3426, n_3427, n_3428, n_3429, n_3430, n_3432;
  wire n_3433, n_3434, n_3435, n_3436, n_3438, n_3439, n_3440, n_3441;
  wire n_3442, n_3444, n_3445, n_3446, n_3447, n_3448, n_3450, n_3451;
  wire n_3452, n_3453, n_3454, n_3456, n_3457, n_3458, n_3459, n_3460;
  wire n_3462, n_3463, n_3464, n_3465, n_3466, n_3468, n_3469, n_3470;
  wire n_3471, n_3472, n_3473, n_3474, n_3476, n_3477, n_3479, n_3480;
  wire n_3481, n_3483, n_3484, n_3486, n_3487, n_3488, n_3490, n_3491;
  wire n_3493, n_3494, n_3495, n_3497, n_3498, n_3500, n_3501, n_3502;
  wire n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, n_3511, n_3512;
  wire n_3513, n_3514, n_3515, n_3517, n_3518, n_3519, n_3521, n_3522;
  wire n_3523, n_3524, n_3525, n_3526, n_3527, n_3529, n_3531, n_3532;
  wire n_3534, n_3536, n_3537, n_3539, n_3541, n_3542, n_3544, n_3546;
  wire n_3547, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, n_3555;
  wire n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563;
  wire n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571;
  wire n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3581, n_3582;
  wire n_3584, n_3586, n_3587, n_3589, n_3591, n_3592, n_3594, n_3596;
  wire n_3597, n_3599, n_3601, n_3602, n_3604, n_3606, n_3607, n_3609;
  wire n_3611, n_3612, n_3614, n_3616, n_3617, n_3619, n_3621, n_3622;
  wire n_3624, n_3626, n_3627, n_3629, n_3631, n_3632, n_3634, n_3636;
  wire n_3637, n_3639, n_3641, n_3642, n_3644, n_3646, n_3647, n_3649;
  wire n_3651, n_3652, n_3654, n_3656, n_3657, n_3659, n_3661, n_3662;
  wire n_3664, n_3666, n_3667, n_3669, n_3671, n_3672, n_3674, n_3676;
  wire n_3680, n_3683, n_3684, n_3686, n_3687, n_3688, n_3690, n_3691;
  wire n_3692, n_3694, n_3695, n_3696, n_3698, n_3699, n_3700, n_3702;
  wire n_3703, n_3704, n_3706, n_3707, n_3708, n_3710, n_3711, n_3712;
  wire n_3714, n_3715, n_3716, n_3718, n_3719, n_3720, n_3722, n_3723;
  wire n_3724, n_3726, n_3727, n_3728, n_3730, n_3731, n_3732, n_3734;
  wire n_3735, n_3736, n_3738, n_3739, n_3740, n_3742, n_3743, n_3744;
  wire n_3746, n_3747, n_3748, n_3750, n_3751, n_3752, n_3754, n_3755;
  wire n_3756, n_3758, n_3759, n_3760, n_3762, n_3763, n_3764, n_3766;
  wire n_3767, n_3768, n_3770, n_3771, n_3772, n_3774, n_3775, n_3776;
  wire n_3778, n_3779, n_3780, n_3782, n_3783, n_3784, n_3786, n_3787;
  wire n_3788, n_3790, n_3791, n_3792, n_3794, n_3795, n_3796, n_3798;
  wire n_3799, n_3800, n_3802, n_3803, n_3804, n_3806, n_3807, n_3808;
  wire n_3810, n_3811, n_3812, n_3814, n_3815, n_3816, n_3818, n_3819;
  wire n_3820, n_3822, n_3823, n_3824, n_3826, n_3827, n_3828, n_3830;
  wire n_3831, n_3832, n_3834, n_3835;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g492 (n_220, A[4], A[0]);
  and g2 (n_138, A[4], A[0]);
  xor g493 (n_1141, A[5], A[3]);
  xor g494 (n_219, n_1141, A[1]);
  nand g3 (n_1142, A[5], A[3]);
  nand g495 (n_1143, A[1], A[3]);
  nand g496 (n_1144, A[5], A[1]);
  nand g497 (n_137, n_1142, n_1143, n_1144);
  xor g498 (n_307, A[6], A[4]);
  and g499 (n_308, A[6], A[4]);
  xor g500 (n_1145, A[0], A[2]);
  xor g501 (n_218, n_1145, n_307);
  nand g502 (n_1146, A[0], A[2]);
  nand g4 (n_1147, n_307, A[2]);
  nand g5 (n_1148, A[0], n_307);
  nand g503 (n_136, n_1146, n_1147, n_1148);
  xor g504 (n_1149, A[7], A[5]);
  xor g505 (n_309, n_1149, A[1]);
  nand g506 (n_1150, A[7], A[5]);
  nand g508 (n_1152, A[7], A[1]);
  nand g6 (n_311, n_1150, n_1144, n_1152);
  xor g509 (n_1153, A[3], n_308);
  xor g510 (n_217, n_1153, n_309);
  nand g511 (n_1154, A[3], n_308);
  nand g512 (n_1155, n_309, n_308);
  nand g513 (n_1156, A[3], n_309);
  nand g514 (n_135, n_1154, n_1155, n_1156);
  xor g515 (n_310, A[8], A[6]);
  and g516 (n_313, A[8], A[6]);
  xor g518 (n_312, n_1145, A[4]);
  nand g521 (n_1160, A[2], A[4]);
  xor g523 (n_1161, n_310, n_311);
  xor g524 (n_216, n_1161, n_312);
  nand g525 (n_1162, n_310, n_311);
  nand g526 (n_1163, n_312, n_311);
  nand g527 (n_1164, n_310, n_312);
  nand g528 (n_134, n_1162, n_1163, n_1164);
  xor g529 (n_1165, A[9], A[7]);
  xor g530 (n_315, n_1165, A[3]);
  nand g531 (n_1166, A[9], A[7]);
  nand g532 (n_1167, A[3], A[7]);
  nand g533 (n_1168, A[9], A[3]);
  nand g534 (n_318, n_1166, n_1167, n_1168);
  xor g535 (n_1169, A[1], A[5]);
  xor g536 (n_316, n_1169, n_313);
  nand g538 (n_1171, n_313, A[5]);
  nand g539 (n_1172, A[1], n_313);
  nand g540 (n_320, n_1144, n_1171, n_1172);
  xor g541 (n_1173, n_314, n_315);
  xor g542 (n_215, n_1173, n_316);
  nand g543 (n_1174, n_314, n_315);
  nand g544 (n_1175, n_316, n_315);
  nand g545 (n_1176, n_314, n_316);
  nand g546 (n_133, n_1174, n_1175, n_1176);
  xor g547 (n_317, A[10], A[8]);
  and g548 (n_322, A[10], A[8]);
  xor g549 (n_1177, A[4], A[2]);
  xor g550 (n_319, n_1177, A[6]);
  nand g552 (n_1179, A[6], A[2]);
  xor g555 (n_1181, A[0], n_317);
  xor g556 (n_321, n_1181, n_318);
  nand g557 (n_1182, A[0], n_317);
  nand g558 (n_1183, n_318, n_317);
  nand g559 (n_1184, A[0], n_318);
  nand g560 (n_326, n_1182, n_1183, n_1184);
  xor g561 (n_1185, n_319, n_320);
  xor g562 (n_214, n_1185, n_321);
  nand g563 (n_1186, n_319, n_320);
  nand g564 (n_1187, n_321, n_320);
  nand g565 (n_1188, n_319, n_321);
  nand g566 (n_132, n_1186, n_1187, n_1188);
  xor g567 (n_1189, A[11], A[9]);
  xor g568 (n_324, n_1189, A[5]);
  nand g569 (n_1190, A[11], A[9]);
  nand g570 (n_1191, A[5], A[9]);
  nand g571 (n_1192, A[11], A[5]);
  nand g572 (n_329, n_1190, n_1191, n_1192);
  xor g573 (n_1193, A[3], A[7]);
  xor g574 (n_325, n_1193, A[1]);
  nand g578 (n_330, n_1167, n_1152, n_1143);
  xor g579 (n_1197, n_322, n_323);
  xor g580 (n_327, n_1197, n_324);
  nand g581 (n_1198, n_322, n_323);
  nand g582 (n_1199, n_324, n_323);
  nand g583 (n_1200, n_322, n_324);
  nand g584 (n_334, n_1198, n_1199, n_1200);
  xor g585 (n_1201, n_325, n_326);
  xor g586 (n_213, n_1201, n_327);
  nand g587 (n_1202, n_325, n_326);
  nand g588 (n_1203, n_327, n_326);
  nand g589 (n_1204, n_325, n_327);
  nand g590 (n_131, n_1202, n_1203, n_1204);
  xor g591 (n_328, A[12], A[10]);
  and g592 (n_335, A[12], A[10]);
  xor g594 (n_331, n_307, A[8]);
  nand g596 (n_1207, A[8], A[4]);
  xor g600 (n_332, n_1145, n_328);
  nand g602 (n_1211, n_328, A[0]);
  nand g603 (n_1212, A[2], n_328);
  nand g604 (n_339, n_1146, n_1211, n_1212);
  xor g605 (n_1213, n_329, n_330);
  xor g606 (n_333, n_1213, n_331);
  nand g607 (n_1214, n_329, n_330);
  nand g608 (n_1215, n_331, n_330);
  nand g609 (n_1216, n_329, n_331);
  nand g610 (n_341, n_1214, n_1215, n_1216);
  xor g611 (n_1217, n_332, n_333);
  xor g612 (n_212, n_1217, n_334);
  nand g613 (n_1218, n_332, n_333);
  nand g614 (n_1219, n_334, n_333);
  nand g615 (n_1220, n_332, n_334);
  nand g616 (n_130, n_1218, n_1219, n_1220);
  xor g617 (n_1221, A[13], A[11]);
  xor g618 (n_338, n_1221, A[7]);
  nand g619 (n_1222, A[13], A[11]);
  nand g620 (n_1223, A[7], A[11]);
  nand g621 (n_1224, A[13], A[7]);
  nand g622 (n_344, n_1222, n_1223, n_1224);
  xor g623 (n_1225, A[5], A[9]);
  xor g624 (n_337, n_1225, A[3]);
  nand g628 (n_345, n_1191, n_1168, n_1142);
  xor g629 (n_1229, A[1], n_335);
  xor g630 (n_340, n_1229, n_336);
  nand g631 (n_1230, A[1], n_335);
  nand g632 (n_1231, n_336, n_335);
  nand g633 (n_1232, A[1], n_336);
  nand g634 (n_348, n_1230, n_1231, n_1232);
  xor g635 (n_1233, n_337, n_338);
  xor g636 (n_342, n_1233, n_339);
  nand g637 (n_1234, n_337, n_338);
  nand g638 (n_1235, n_339, n_338);
  nand g639 (n_1236, n_337, n_339);
  nand g640 (n_350, n_1234, n_1235, n_1236);
  xor g641 (n_1237, n_340, n_341);
  xor g642 (n_211, n_1237, n_342);
  nand g643 (n_1238, n_340, n_341);
  nand g644 (n_1239, n_342, n_341);
  nand g645 (n_1240, n_340, n_342);
  nand g646 (n_129, n_1238, n_1239, n_1240);
  xor g647 (n_343, A[14], A[12]);
  and g648 (n_352, A[14], A[12]);
  xor g649 (n_1241, A[8], A[0]);
  xor g650 (n_347, n_1241, A[6]);
  nand g651 (n_1242, A[8], A[0]);
  nand g652 (n_1243, A[6], A[0]);
  xor g655 (n_1245, A[10], A[4]);
  xor g656 (n_346, n_1245, A[2]);
  nand g657 (n_1246, A[10], A[4]);
  nand g659 (n_1248, A[10], A[2]);
  nand g660 (n_354, n_1246, n_1160, n_1248);
  xor g661 (n_1249, n_343, n_344);
  xor g662 (n_349, n_1249, n_345);
  nand g663 (n_1250, n_343, n_344);
  nand g664 (n_1251, n_345, n_344);
  nand g665 (n_1252, n_343, n_345);
  nand g666 (n_358, n_1250, n_1251, n_1252);
  xor g667 (n_1253, n_346, n_347);
  xor g668 (n_351, n_1253, n_348);
  nand g669 (n_1254, n_346, n_347);
  nand g670 (n_1255, n_348, n_347);
  nand g671 (n_1256, n_346, n_348);
  nand g672 (n_361, n_1254, n_1255, n_1256);
  xor g673 (n_1257, n_349, n_350);
  xor g674 (n_210, n_1257, n_351);
  nand g675 (n_1258, n_349, n_350);
  nand g676 (n_1259, n_351, n_350);
  nand g677 (n_1260, n_349, n_351);
  nand g678 (n_128, n_1258, n_1259, n_1260);
  xor g679 (n_1261, A[15], A[13]);
  xor g680 (n_355, n_1261, A[9]);
  nand g681 (n_1262, A[15], A[13]);
  nand g682 (n_1263, A[9], A[13]);
  nand g683 (n_1264, A[15], A[9]);
  nand g684 (n_363, n_1262, n_1263, n_1264);
  xor g685 (n_1265, A[1], A[7]);
  xor g686 (n_356, n_1265, A[11]);
  nand g689 (n_1268, A[1], A[11]);
  nand g690 (n_364, n_1152, n_1223, n_1268);
  xor g692 (n_357, n_1141, n_352);
  nand g694 (n_1271, n_352, A[3]);
  nand g695 (n_1272, A[5], n_352);
  nand g696 (n_367, n_1142, n_1271, n_1272);
  xor g697 (n_1273, n_353, n_354);
  xor g698 (n_359, n_1273, n_355);
  nand g699 (n_1274, n_353, n_354);
  nand g700 (n_1275, n_355, n_354);
  nand g701 (n_1276, n_353, n_355);
  nand g702 (n_369, n_1274, n_1275, n_1276);
  xor g703 (n_1277, n_356, n_357);
  xor g704 (n_360, n_1277, n_358);
  nand g705 (n_1278, n_356, n_357);
  nand g706 (n_1279, n_358, n_357);
  nand g707 (n_1280, n_356, n_358);
  nand g708 (n_371, n_1278, n_1279, n_1280);
  xor g709 (n_1281, n_359, n_360);
  xor g710 (n_209, n_1281, n_361);
  nand g711 (n_1282, n_359, n_360);
  nand g712 (n_1283, n_361, n_360);
  nand g713 (n_1284, n_359, n_361);
  nand g714 (n_127, n_1282, n_1283, n_1284);
  xor g715 (n_362, A[16], A[14]);
  and g716 (n_373, A[16], A[14]);
  xor g717 (n_1285, A[10], A[2]);
  xor g718 (n_366, n_1285, A[0]);
  nand g721 (n_1288, A[10], A[0]);
  nand g722 (n_374, n_1248, n_1146, n_1288);
  xor g723 (n_1289, A[8], A[12]);
  xor g724 (n_365, n_1289, A[6]);
  nand g725 (n_1290, A[8], A[12]);
  nand g726 (n_1291, A[6], A[12]);
  xor g729 (n_1293, A[4], n_362);
  xor g730 (n_368, n_1293, n_363);
  nand g731 (n_1294, A[4], n_362);
  nand g732 (n_1295, n_363, n_362);
  nand g733 (n_1296, A[4], n_363);
  nand g734 (n_379, n_1294, n_1295, n_1296);
  xor g735 (n_1297, n_364, n_365);
  xor g736 (n_370, n_1297, n_366);
  nand g737 (n_1298, n_364, n_365);
  nand g738 (n_1299, n_366, n_365);
  nand g739 (n_1300, n_364, n_366);
  nand g740 (n_381, n_1298, n_1299, n_1300);
  xor g741 (n_1301, n_367, n_368);
  xor g742 (n_372, n_1301, n_369);
  nand g743 (n_1302, n_367, n_368);
  nand g744 (n_1303, n_369, n_368);
  nand g745 (n_1304, n_367, n_369);
  nand g746 (n_383, n_1302, n_1303, n_1304);
  xor g747 (n_1305, n_370, n_371);
  xor g748 (n_208, n_1305, n_372);
  nand g749 (n_1306, n_370, n_371);
  nand g750 (n_1307, n_372, n_371);
  nand g751 (n_1308, n_370, n_372);
  nand g752 (n_126, n_1306, n_1307, n_1308);
  xor g753 (n_1309, A[17], A[15]);
  xor g754 (n_377, n_1309, A[11]);
  nand g755 (n_1310, A[17], A[15]);
  nand g756 (n_1311, A[11], A[15]);
  nand g757 (n_1312, A[17], A[11]);
  nand g758 (n_386, n_1310, n_1311, n_1312);
  xor g759 (n_1313, A[3], A[1]);
  xor g760 (n_378, n_1313, A[9]);
  nand g762 (n_1315, A[9], A[1]);
  nand g764 (n_388, n_1143, n_1315, n_1168);
  xor g765 (n_1317, A[13], A[7]);
  xor g766 (n_376, n_1317, A[5]);
  nand g769 (n_1320, A[13], A[5]);
  nand g770 (n_387, n_1224, n_1150, n_1320);
  xor g771 (n_1321, n_373, n_374);
  xor g772 (n_380, n_1321, n_375);
  nand g773 (n_1322, n_373, n_374);
  nand g774 (n_1323, n_375, n_374);
  nand g775 (n_1324, n_373, n_375);
  nand g776 (n_392, n_1322, n_1323, n_1324);
  xor g777 (n_1325, n_376, n_377);
  xor g778 (n_382, n_1325, n_378);
  nand g779 (n_1326, n_376, n_377);
  nand g780 (n_1327, n_378, n_377);
  nand g781 (n_1328, n_376, n_378);
  nand g782 (n_394, n_1326, n_1327, n_1328);
  xor g783 (n_1329, n_379, n_380);
  xor g784 (n_384, n_1329, n_381);
  nand g785 (n_1330, n_379, n_380);
  nand g786 (n_1331, n_381, n_380);
  nand g787 (n_1332, n_379, n_381);
  nand g788 (n_396, n_1330, n_1331, n_1332);
  xor g789 (n_1333, n_382, n_383);
  xor g790 (n_207, n_1333, n_384);
  nand g791 (n_1334, n_382, n_383);
  nand g792 (n_1335, n_384, n_383);
  nand g793 (n_1336, n_382, n_384);
  nand g794 (n_125, n_1334, n_1335, n_1336);
  xor g795 (n_385, A[18], A[16]);
  and g796 (n_398, A[18], A[16]);
  xor g797 (n_1337, A[12], A[4]);
  xor g798 (n_389, n_1337, A[2]);
  nand g799 (n_1338, A[12], A[4]);
  nand g801 (n_1340, A[12], A[2]);
  nand g802 (n_399, n_1338, n_1160, n_1340);
  xor g803 (n_1341, A[10], A[0]);
  xor g804 (n_390, n_1341, A[14]);
  nand g806 (n_1343, A[14], A[0]);
  nand g807 (n_1344, A[10], A[14]);
  nand g808 (n_400, n_1288, n_1343, n_1344);
  xor g810 (n_391, n_310, n_385);
  nand g812 (n_1347, n_385, A[6]);
  nand g813 (n_1348, A[8], n_385);
  xor g815 (n_1349, n_386, n_387);
  xor g816 (n_393, n_1349, n_388);
  nand g817 (n_1350, n_386, n_387);
  nand g818 (n_1351, n_388, n_387);
  nand g819 (n_1352, n_386, n_388);
  nand g820 (n_406, n_1350, n_1351, n_1352);
  xor g821 (n_1353, n_389, n_390);
  xor g822 (n_395, n_1353, n_391);
  nand g823 (n_1354, n_389, n_390);
  nand g824 (n_1355, n_391, n_390);
  nand g825 (n_1356, n_389, n_391);
  nand g826 (n_407, n_1354, n_1355, n_1356);
  xor g827 (n_1357, n_392, n_393);
  xor g828 (n_397, n_1357, n_394);
  nand g829 (n_1358, n_392, n_393);
  nand g830 (n_1359, n_394, n_393);
  nand g831 (n_1360, n_392, n_394);
  nand g832 (n_410, n_1358, n_1359, n_1360);
  xor g833 (n_1361, n_395, n_396);
  xor g834 (n_206, n_1361, n_397);
  nand g835 (n_1362, n_395, n_396);
  nand g836 (n_1363, n_397, n_396);
  nand g837 (n_1364, n_395, n_397);
  nand g838 (n_124, n_1362, n_1363, n_1364);
  xor g839 (n_1365, A[19], A[17]);
  xor g840 (n_402, n_1365, A[13]);
  nand g841 (n_1366, A[19], A[17]);
  nand g842 (n_1367, A[13], A[17]);
  nand g843 (n_1368, A[19], A[13]);
  nand g844 (n_412, n_1366, n_1367, n_1368);
  xor g846 (n_403, n_1141, A[11]);
  nand g848 (n_1371, A[11], A[3]);
  nand g850 (n_413, n_1142, n_1371, n_1192);
  xor g851 (n_1373, A[1], A[15]);
  xor g852 (n_401, n_1373, A[9]);
  nand g853 (n_1374, A[1], A[15]);
  nand g856 (n_414, n_1374, n_1264, n_1315);
  xor g857 (n_1377, A[7], n_398);
  xor g858 (n_405, n_1377, n_399);
  nand g859 (n_1378, A[7], n_398);
  nand g860 (n_1379, n_399, n_398);
  nand g861 (n_1380, A[7], n_399);
  nand g862 (n_418, n_1378, n_1379, n_1380);
  xor g863 (n_1381, n_400, n_401);
  xor g864 (n_408, n_1381, n_402);
  nand g865 (n_1382, n_400, n_401);
  nand g866 (n_1383, n_402, n_401);
  nand g867 (n_1384, n_400, n_402);
  nand g868 (n_420, n_1382, n_1383, n_1384);
  xor g869 (n_1385, n_403, n_404);
  xor g870 (n_409, n_1385, n_405);
  nand g871 (n_1386, n_403, n_404);
  nand g872 (n_1387, n_405, n_404);
  nand g873 (n_1388, n_403, n_405);
  nand g874 (n_422, n_1386, n_1387, n_1388);
  xor g875 (n_1389, n_406, n_407);
  xor g876 (n_411, n_1389, n_408);
  nand g877 (n_1390, n_406, n_407);
  nand g878 (n_1391, n_408, n_407);
  nand g879 (n_1392, n_406, n_408);
  nand g880 (n_140, n_1390, n_1391, n_1392);
  xor g881 (n_1393, n_409, n_410);
  xor g882 (n_205, n_1393, n_411);
  nand g883 (n_1394, n_409, n_410);
  nand g884 (n_1395, n_411, n_410);
  nand g885 (n_1396, n_409, n_411);
  nand g886 (n_123, n_1394, n_1395, n_1396);
  xor g887 (n_1397, A[20], A[18]);
  xor g888 (n_416, n_1397, A[14]);
  nand g889 (n_1398, A[20], A[18]);
  nand g890 (n_1399, A[14], A[18]);
  nand g891 (n_1400, A[20], A[14]);
  nand g892 (n_143, n_1398, n_1399, n_1400);
  xor g894 (n_417, n_307, A[12]);
  xor g899 (n_1405, A[2], A[16]);
  xor g900 (n_415, n_1405, A[10]);
  nand g901 (n_1406, A[2], A[16]);
  nand g902 (n_1407, A[10], A[16]);
  nand g904 (n_424, n_1406, n_1407, n_1248);
  xor g905 (n_1409, A[8], n_412);
  xor g906 (n_419, n_1409, n_413);
  nand g907 (n_1410, A[8], n_412);
  nand g908 (n_1411, n_413, n_412);
  nand g909 (n_1412, A[8], n_413);
  nand g910 (n_428, n_1410, n_1411, n_1412);
  xor g911 (n_1413, n_414, n_415);
  xor g912 (n_421, n_1413, n_416);
  nand g913 (n_1414, n_414, n_415);
  nand g914 (n_1415, n_416, n_415);
  nand g915 (n_1416, n_414, n_416);
  nand g916 (n_430, n_1414, n_1415, n_1416);
  xor g917 (n_1417, n_417, n_418);
  xor g918 (n_139, n_1417, n_419);
  nand g919 (n_1418, n_417, n_418);
  nand g920 (n_1419, n_419, n_418);
  nand g921 (n_1420, n_417, n_419);
  nand g922 (n_432, n_1418, n_1419, n_1420);
  xor g923 (n_1421, n_420, n_421);
  xor g924 (n_141, n_1421, n_422);
  nand g925 (n_1422, n_420, n_421);
  nand g926 (n_1423, n_422, n_421);
  nand g927 (n_1424, n_420, n_422);
  nand g928 (n_434, n_1422, n_1423, n_1424);
  xor g929 (n_1425, n_139, n_140);
  xor g930 (n_204, n_1425, n_141);
  nand g931 (n_1426, n_139, n_140);
  nand g932 (n_1427, n_141, n_140);
  nand g933 (n_1428, n_139, n_141);
  nand g934 (n_122, n_1426, n_1427, n_1428);
  xor g935 (n_1429, A[21], A[19]);
  xor g936 (n_426, n_1429, A[15]);
  nand g937 (n_1430, A[21], A[19]);
  nand g938 (n_1431, A[15], A[19]);
  nand g939 (n_1432, A[21], A[15]);
  nand g940 (n_436, n_1430, n_1431, n_1432);
  xor g942 (n_427, n_1149, A[13]);
  xor g947 (n_1437, A[3], A[17]);
  xor g948 (n_425, n_1437, A[11]);
  nand g949 (n_1438, A[3], A[17]);
  nand g952 (n_438, n_1438, n_1312, n_1371);
  xor g953 (n_1441, A[9], n_143);
  xor g954 (n_429, n_1441, n_423);
  nand g955 (n_1442, A[9], n_143);
  nand g956 (n_1443, n_423, n_143);
  nand g957 (n_1444, A[9], n_423);
  nand g958 (n_442, n_1442, n_1443, n_1444);
  xor g959 (n_1445, n_424, n_425);
  xor g960 (n_431, n_1445, n_426);
  nand g961 (n_1446, n_424, n_425);
  nand g962 (n_1447, n_426, n_425);
  nand g963 (n_1448, n_424, n_426);
  nand g964 (n_444, n_1446, n_1447, n_1448);
  xor g965 (n_1449, n_427, n_428);
  xor g966 (n_433, n_1449, n_429);
  nand g967 (n_1450, n_427, n_428);
  nand g968 (n_1451, n_429, n_428);
  nand g969 (n_1452, n_427, n_429);
  nand g970 (n_446, n_1450, n_1451, n_1452);
  xor g971 (n_1453, n_430, n_431);
  xor g972 (n_435, n_1453, n_432);
  nand g973 (n_1454, n_430, n_431);
  nand g974 (n_1455, n_432, n_431);
  nand g975 (n_1456, n_430, n_432);
  nand g976 (n_449, n_1454, n_1455, n_1456);
  xor g977 (n_1457, n_433, n_434);
  xor g978 (n_203, n_1457, n_435);
  nand g979 (n_1458, n_433, n_434);
  nand g980 (n_1459, n_435, n_434);
  nand g981 (n_1460, n_433, n_435);
  nand g982 (n_121, n_1458, n_1459, n_1460);
  xor g983 (n_1461, A[22], A[20]);
  xor g984 (n_440, n_1461, A[16]);
  nand g985 (n_1462, A[22], A[20]);
  nand g986 (n_1463, A[16], A[20]);
  nand g987 (n_1464, A[22], A[16]);
  nand g988 (n_450, n_1462, n_1463, n_1464);
  xor g990 (n_441, n_310, A[14]);
  nand g992 (n_1467, A[14], A[6]);
  nand g993 (n_1468, A[8], A[14]);
  xor g995 (n_1469, A[4], A[18]);
  xor g996 (n_439, n_1469, A[12]);
  nand g997 (n_1470, A[4], A[18]);
  nand g998 (n_1471, A[12], A[18]);
  nand g1000 (n_452, n_1470, n_1471, n_1338);
  xor g1001 (n_1473, A[10], n_436);
  xor g1002 (n_443, n_1473, n_387);
  nand g1003 (n_1474, A[10], n_436);
  nand g1004 (n_1475, n_387, n_436);
  nand g1005 (n_1476, A[10], n_387);
  nand g1006 (n_456, n_1474, n_1475, n_1476);
  xor g1007 (n_1477, n_438, n_439);
  xor g1008 (n_445, n_1477, n_440);
  nand g1009 (n_1478, n_438, n_439);
  nand g1010 (n_1479, n_440, n_439);
  nand g1011 (n_1480, n_438, n_440);
  nand g1012 (n_458, n_1478, n_1479, n_1480);
  xor g1013 (n_1481, n_441, n_442);
  xor g1014 (n_447, n_1481, n_443);
  nand g1015 (n_1482, n_441, n_442);
  nand g1016 (n_1483, n_443, n_442);
  nand g1017 (n_1484, n_441, n_443);
  nand g1018 (n_460, n_1482, n_1483, n_1484);
  xor g1019 (n_1485, n_444, n_445);
  xor g1020 (n_448, n_1485, n_446);
  nand g1021 (n_1486, n_444, n_445);
  nand g1022 (n_1487, n_446, n_445);
  nand g1023 (n_1488, n_444, n_446);
  nand g1024 (n_463, n_1486, n_1487, n_1488);
  xor g1025 (n_1489, n_447, n_448);
  xor g1026 (n_202, n_1489, n_449);
  nand g1027 (n_1490, n_447, n_448);
  nand g1028 (n_1491, n_449, n_448);
  nand g1029 (n_1492, n_447, n_449);
  nand g1030 (n_120, n_1490, n_1491, n_1492);
  xor g1031 (n_1493, A[23], A[21]);
  xor g1032 (n_454, n_1493, A[17]);
  nand g1033 (n_1494, A[23], A[21]);
  nand g1034 (n_1495, A[17], A[21]);
  nand g1035 (n_1496, A[23], A[17]);
  nand g1036 (n_464, n_1494, n_1495, n_1496);
  xor g1038 (n_455, n_1165, A[15]);
  nand g1040 (n_1499, A[15], A[7]);
  nand g1042 (n_465, n_1166, n_1499, n_1264);
  xor g1043 (n_1501, A[5], A[19]);
  xor g1044 (n_453, n_1501, A[13]);
  nand g1045 (n_1502, A[5], A[19]);
  nand g1048 (n_466, n_1502, n_1368, n_1320);
  xor g1049 (n_1505, A[11], n_450);
  xor g1050 (n_457, n_1505, n_451);
  nand g1051 (n_1506, A[11], n_450);
  nand g1052 (n_1507, n_451, n_450);
  nand g1053 (n_1508, A[11], n_451);
  nand g1054 (n_470, n_1506, n_1507, n_1508);
  xor g1055 (n_1509, n_452, n_453);
  xor g1056 (n_459, n_1509, n_454);
  nand g1057 (n_1510, n_452, n_453);
  nand g1058 (n_1511, n_454, n_453);
  nand g1059 (n_1512, n_452, n_454);
  nand g1060 (n_472, n_1510, n_1511, n_1512);
  xor g1061 (n_1513, n_455, n_456);
  xor g1062 (n_461, n_1513, n_457);
  nand g1063 (n_1514, n_455, n_456);
  nand g1064 (n_1515, n_457, n_456);
  nand g1065 (n_1516, n_455, n_457);
  nand g1066 (n_474, n_1514, n_1515, n_1516);
  xor g1067 (n_1517, n_458, n_459);
  xor g1068 (n_462, n_1517, n_460);
  nand g1069 (n_1518, n_458, n_459);
  nand g1070 (n_1519, n_460, n_459);
  nand g1071 (n_1520, n_458, n_460);
  nand g1072 (n_477, n_1518, n_1519, n_1520);
  xor g1073 (n_1521, n_461, n_462);
  xor g1074 (n_201, n_1521, n_463);
  nand g1075 (n_1522, n_461, n_462);
  nand g1076 (n_1523, n_463, n_462);
  nand g1077 (n_1524, n_461, n_463);
  nand g1078 (n_119, n_1522, n_1523, n_1524);
  xor g1079 (n_1525, A[24], A[22]);
  xor g1080 (n_468, n_1525, A[18]);
  nand g1081 (n_1526, A[24], A[22]);
  nand g1082 (n_1527, A[18], A[22]);
  nand g1083 (n_1528, A[24], A[18]);
  nand g1084 (n_478, n_1526, n_1527, n_1528);
  xor g1086 (n_469, n_317, A[16]);
  nand g1088 (n_1531, A[16], A[8]);
  xor g1091 (n_1533, A[6], A[20]);
  xor g1092 (n_467, n_1533, A[14]);
  nand g1093 (n_1534, A[6], A[20]);
  nand g1096 (n_480, n_1534, n_1400, n_1467);
  xor g1097 (n_1537, A[12], n_464);
  xor g1098 (n_471, n_1537, n_465);
  nand g1099 (n_1538, A[12], n_464);
  nand g1100 (n_1539, n_465, n_464);
  nand g1101 (n_1540, A[12], n_465);
  nand g1102 (n_484, n_1538, n_1539, n_1540);
  xor g1103 (n_1541, n_466, n_467);
  xor g1104 (n_473, n_1541, n_468);
  nand g1105 (n_1542, n_466, n_467);
  nand g1106 (n_1543, n_468, n_467);
  nand g1107 (n_1544, n_466, n_468);
  nand g1108 (n_486, n_1542, n_1543, n_1544);
  xor g1109 (n_1545, n_469, n_470);
  xor g1110 (n_475, n_1545, n_471);
  nand g1111 (n_1546, n_469, n_470);
  nand g1112 (n_1547, n_471, n_470);
  nand g1113 (n_1548, n_469, n_471);
  nand g1114 (n_488, n_1546, n_1547, n_1548);
  xor g1115 (n_1549, n_472, n_473);
  xor g1116 (n_476, n_1549, n_474);
  nand g1117 (n_1550, n_472, n_473);
  nand g1118 (n_1551, n_474, n_473);
  nand g1119 (n_1552, n_472, n_474);
  nand g1120 (n_491, n_1550, n_1551, n_1552);
  xor g1121 (n_1553, n_475, n_476);
  xor g1122 (n_200, n_1553, n_477);
  nand g1123 (n_1554, n_475, n_476);
  nand g1124 (n_1555, n_477, n_476);
  nand g1125 (n_1556, n_475, n_477);
  nand g1126 (n_118, n_1554, n_1555, n_1556);
  xor g1127 (n_1557, A[25], A[23]);
  xor g1128 (n_482, n_1557, A[19]);
  nand g1129 (n_1558, A[25], A[23]);
  nand g1130 (n_1559, A[19], A[23]);
  nand g1131 (n_1560, A[25], A[19]);
  nand g1132 (n_492, n_1558, n_1559, n_1560);
  xor g1134 (n_483, n_1189, A[17]);
  nand g1136 (n_1563, A[17], A[9]);
  nand g1138 (n_493, n_1190, n_1563, n_1312);
  xor g1139 (n_1565, A[7], A[21]);
  xor g1140 (n_481, n_1565, A[15]);
  nand g1141 (n_1566, A[7], A[21]);
  nand g1144 (n_494, n_1566, n_1432, n_1499);
  xor g1145 (n_1569, A[13], n_478);
  xor g1146 (n_485, n_1569, n_479);
  nand g1147 (n_1570, A[13], n_478);
  nand g1148 (n_1571, n_479, n_478);
  nand g1149 (n_1572, A[13], n_479);
  nand g1150 (n_496, n_1570, n_1571, n_1572);
  xor g1151 (n_1573, n_480, n_481);
  xor g1152 (n_487, n_1573, n_482);
  nand g1153 (n_1574, n_480, n_481);
  nand g1154 (n_1575, n_482, n_481);
  nand g1155 (n_1576, n_480, n_482);
  nand g1156 (n_498, n_1574, n_1575, n_1576);
  xor g1157 (n_1577, n_483, n_484);
  xor g1158 (n_489, n_1577, n_485);
  nand g1159 (n_1578, n_483, n_484);
  nand g1160 (n_1579, n_485, n_484);
  nand g1161 (n_1580, n_483, n_485);
  nand g1162 (n_500, n_1578, n_1579, n_1580);
  xor g1163 (n_1581, n_486, n_487);
  xor g1164 (n_490, n_1581, n_488);
  nand g1165 (n_1582, n_486, n_487);
  nand g1166 (n_1583, n_488, n_487);
  nand g1167 (n_1584, n_486, n_488);
  nand g1168 (n_503, n_1582, n_1583, n_1584);
  xor g1169 (n_1585, n_489, n_490);
  xor g1170 (n_199, n_1585, n_491);
  nand g1171 (n_1586, n_489, n_490);
  nand g1172 (n_1587, n_491, n_490);
  nand g1173 (n_1588, n_489, n_491);
  nand g1174 (n_117, n_1586, n_1587, n_1588);
  xor g1175 (n_1589, A[26], A[24]);
  xor g1176 (n_222, n_1589, A[20]);
  nand g1177 (n_1590, A[26], A[24]);
  nand g1178 (n_1591, A[20], A[24]);
  nand g1179 (n_1592, A[26], A[20]);
  nand g1180 (n_504, n_1590, n_1591, n_1592);
  xor g1182 (n_495, n_328, A[18]);
  nand g1184 (n_1595, A[18], A[10]);
  xor g1187 (n_1597, A[8], A[22]);
  xor g1188 (n_221, n_1597, A[16]);
  nand g1189 (n_1598, A[8], A[22]);
  nand g1192 (n_506, n_1598, n_1464, n_1531);
  xor g1193 (n_1601, A[14], n_492);
  xor g1194 (n_497, n_1601, n_493);
  nand g1195 (n_1602, A[14], n_492);
  nand g1196 (n_1603, n_493, n_492);
  nand g1197 (n_1604, A[14], n_493);
  nand g1198 (n_510, n_1602, n_1603, n_1604);
  xor g1199 (n_1605, n_494, n_221);
  xor g1200 (n_499, n_1605, n_222);
  nand g1201 (n_1606, n_494, n_221);
  nand g1202 (n_1607, n_222, n_221);
  nand g1203 (n_1608, n_494, n_222);
  nand g1204 (n_512, n_1606, n_1607, n_1608);
  xor g1205 (n_1609, n_495, n_496);
  xor g1206 (n_501, n_1609, n_497);
  nand g1207 (n_1610, n_495, n_496);
  nand g1208 (n_1611, n_497, n_496);
  nand g1209 (n_1612, n_495, n_497);
  nand g1210 (n_514, n_1610, n_1611, n_1612);
  xor g1211 (n_1613, n_498, n_499);
  xor g1212 (n_502, n_1613, n_500);
  nand g1213 (n_1614, n_498, n_499);
  nand g1214 (n_1615, n_500, n_499);
  nand g1215 (n_1616, n_498, n_500);
  nand g1216 (n_517, n_1614, n_1615, n_1616);
  xor g1217 (n_1617, n_501, n_502);
  xor g1218 (n_198, n_1617, n_503);
  nand g1219 (n_1618, n_501, n_502);
  nand g1220 (n_1619, n_503, n_502);
  nand g1221 (n_1620, n_501, n_503);
  nand g1222 (n_116, n_1618, n_1619, n_1620);
  xor g1223 (n_1621, A[27], A[25]);
  xor g1224 (n_508, n_1621, A[21]);
  nand g1225 (n_1622, A[27], A[25]);
  nand g1226 (n_1623, A[21], A[25]);
  nand g1227 (n_1624, A[27], A[21]);
  nand g1228 (n_518, n_1622, n_1623, n_1624);
  xor g1230 (n_509, n_1221, A[19]);
  nand g1232 (n_1627, A[19], A[11]);
  nand g1234 (n_519, n_1222, n_1627, n_1368);
  xor g1235 (n_1629, A[9], A[23]);
  xor g1236 (n_507, n_1629, A[17]);
  nand g1237 (n_1630, A[9], A[23]);
  nand g1240 (n_520, n_1630, n_1496, n_1563);
  xor g1241 (n_1633, A[15], n_504);
  xor g1242 (n_511, n_1633, n_505);
  nand g1243 (n_1634, A[15], n_504);
  nand g1244 (n_1635, n_505, n_504);
  nand g1245 (n_1636, A[15], n_505);
  nand g1246 (n_524, n_1634, n_1635, n_1636);
  xor g1247 (n_1637, n_506, n_507);
  xor g1248 (n_513, n_1637, n_508);
  nand g1249 (n_1638, n_506, n_507);
  nand g1250 (n_1639, n_508, n_507);
  nand g1251 (n_1640, n_506, n_508);
  nand g1252 (n_526, n_1638, n_1639, n_1640);
  xor g1253 (n_1641, n_509, n_510);
  xor g1254 (n_515, n_1641, n_511);
  nand g1255 (n_1642, n_509, n_510);
  nand g1256 (n_1643, n_511, n_510);
  nand g1257 (n_1644, n_509, n_511);
  nand g1258 (n_528, n_1642, n_1643, n_1644);
  xor g1259 (n_1645, n_512, n_513);
  xor g1260 (n_516, n_1645, n_514);
  nand g1261 (n_1646, n_512, n_513);
  nand g1262 (n_1647, n_514, n_513);
  nand g1263 (n_1648, n_512, n_514);
  nand g1264 (n_531, n_1646, n_1647, n_1648);
  xor g1265 (n_1649, n_515, n_516);
  xor g1266 (n_197, n_1649, n_517);
  nand g1267 (n_1650, n_515, n_516);
  nand g1268 (n_1651, n_517, n_516);
  nand g1269 (n_1652, n_515, n_517);
  nand g1270 (n_115, n_1650, n_1651, n_1652);
  xor g1271 (n_1653, A[28], A[26]);
  xor g1272 (n_522, n_1653, A[22]);
  nand g1273 (n_1654, A[28], A[26]);
  nand g1274 (n_1655, A[22], A[26]);
  nand g1275 (n_1656, A[28], A[22]);
  nand g1276 (n_532, n_1654, n_1655, n_1656);
  xor g1278 (n_523, n_343, A[20]);
  nand g1280 (n_1659, A[20], A[12]);
  xor g1283 (n_1661, A[10], A[24]);
  xor g1284 (n_521, n_1661, A[18]);
  nand g1285 (n_1662, A[10], A[24]);
  nand g1288 (n_534, n_1662, n_1528, n_1595);
  xor g1289 (n_1665, A[16], n_518);
  xor g1290 (n_525, n_1665, n_519);
  nand g1291 (n_1666, A[16], n_518);
  nand g1292 (n_1667, n_519, n_518);
  nand g1293 (n_1668, A[16], n_519);
  nand g1294 (n_538, n_1666, n_1667, n_1668);
  xor g1295 (n_1669, n_520, n_521);
  xor g1296 (n_527, n_1669, n_522);
  nand g1297 (n_1670, n_520, n_521);
  nand g1298 (n_1671, n_522, n_521);
  nand g1299 (n_1672, n_520, n_522);
  nand g1300 (n_540, n_1670, n_1671, n_1672);
  xor g1301 (n_1673, n_523, n_524);
  xor g1302 (n_529, n_1673, n_525);
  nand g1303 (n_1674, n_523, n_524);
  nand g1304 (n_1675, n_525, n_524);
  nand g1305 (n_1676, n_523, n_525);
  nand g1306 (n_542, n_1674, n_1675, n_1676);
  xor g1307 (n_1677, n_526, n_527);
  xor g1308 (n_530, n_1677, n_528);
  nand g1309 (n_1678, n_526, n_527);
  nand g1310 (n_1679, n_528, n_527);
  nand g1311 (n_1680, n_526, n_528);
  nand g1312 (n_545, n_1678, n_1679, n_1680);
  xor g1313 (n_1681, n_529, n_530);
  xor g1314 (n_196, n_1681, n_531);
  nand g1315 (n_1682, n_529, n_530);
  nand g1316 (n_1683, n_531, n_530);
  nand g1317 (n_1684, n_529, n_531);
  nand g1318 (n_114, n_1682, n_1683, n_1684);
  xor g1319 (n_1685, A[29], A[27]);
  xor g1320 (n_536, n_1685, A[23]);
  nand g1321 (n_1686, A[29], A[27]);
  nand g1322 (n_1687, A[23], A[27]);
  nand g1323 (n_1688, A[29], A[23]);
  nand g1324 (n_546, n_1686, n_1687, n_1688);
  xor g1326 (n_537, n_1261, A[21]);
  nand g1328 (n_1691, A[21], A[13]);
  nand g1330 (n_547, n_1262, n_1691, n_1432);
  xor g1331 (n_1693, A[11], A[25]);
  xor g1332 (n_535, n_1693, A[19]);
  nand g1333 (n_1694, A[11], A[25]);
  nand g1336 (n_548, n_1694, n_1560, n_1627);
  xor g1337 (n_1697, A[17], n_532);
  xor g1338 (n_539, n_1697, n_533);
  nand g1339 (n_1698, A[17], n_532);
  nand g1340 (n_1699, n_533, n_532);
  nand g1341 (n_1700, A[17], n_533);
  nand g1342 (n_552, n_1698, n_1699, n_1700);
  xor g1343 (n_1701, n_534, n_535);
  xor g1344 (n_541, n_1701, n_536);
  nand g1345 (n_1702, n_534, n_535);
  nand g1346 (n_1703, n_536, n_535);
  nand g1347 (n_1704, n_534, n_536);
  nand g1348 (n_554, n_1702, n_1703, n_1704);
  xor g1349 (n_1705, n_537, n_538);
  xor g1350 (n_543, n_1705, n_539);
  nand g1351 (n_1706, n_537, n_538);
  nand g1352 (n_1707, n_539, n_538);
  nand g1353 (n_1708, n_537, n_539);
  nand g1354 (n_556, n_1706, n_1707, n_1708);
  xor g1355 (n_1709, n_540, n_541);
  xor g1356 (n_544, n_1709, n_542);
  nand g1357 (n_1710, n_540, n_541);
  nand g1358 (n_1711, n_542, n_541);
  nand g1359 (n_1712, n_540, n_542);
  nand g1360 (n_559, n_1710, n_1711, n_1712);
  xor g1361 (n_1713, n_543, n_544);
  xor g1362 (n_195, n_1713, n_545);
  nand g1363 (n_1714, n_543, n_544);
  nand g1364 (n_1715, n_545, n_544);
  nand g1365 (n_1716, n_543, n_545);
  nand g1366 (n_113, n_1714, n_1715, n_1716);
  xor g1367 (n_1717, A[30], A[28]);
  xor g1368 (n_550, n_1717, A[24]);
  nand g1369 (n_1718, A[30], A[28]);
  nand g1370 (n_1719, A[24], A[28]);
  nand g1371 (n_1720, A[30], A[24]);
  nand g1372 (n_560, n_1718, n_1719, n_1720);
  xor g1374 (n_551, n_362, A[22]);
  nand g1376 (n_1723, A[22], A[14]);
  xor g1379 (n_1725, A[12], A[26]);
  xor g1380 (n_549, n_1725, A[20]);
  nand g1381 (n_1726, A[12], A[26]);
  nand g1384 (n_562, n_1726, n_1592, n_1659);
  xor g1385 (n_1729, A[18], n_546);
  xor g1386 (n_553, n_1729, n_547);
  nand g1387 (n_1730, A[18], n_546);
  nand g1388 (n_1731, n_547, n_546);
  nand g1389 (n_1732, A[18], n_547);
  nand g1390 (n_566, n_1730, n_1731, n_1732);
  xor g1391 (n_1733, n_548, n_549);
  xor g1392 (n_555, n_1733, n_550);
  nand g1393 (n_1734, n_548, n_549);
  nand g1394 (n_1735, n_550, n_549);
  nand g1395 (n_1736, n_548, n_550);
  nand g1396 (n_568, n_1734, n_1735, n_1736);
  xor g1397 (n_1737, n_551, n_552);
  xor g1398 (n_557, n_1737, n_553);
  nand g1399 (n_1738, n_551, n_552);
  nand g1400 (n_1739, n_553, n_552);
  nand g1401 (n_1740, n_551, n_553);
  nand g1402 (n_570, n_1738, n_1739, n_1740);
  xor g1403 (n_1741, n_554, n_555);
  xor g1404 (n_558, n_1741, n_556);
  nand g1405 (n_1742, n_554, n_555);
  nand g1406 (n_1743, n_556, n_555);
  nand g1407 (n_1744, n_554, n_556);
  nand g1408 (n_573, n_1742, n_1743, n_1744);
  xor g1409 (n_1745, n_557, n_558);
  xor g1410 (n_194, n_1745, n_559);
  nand g1411 (n_1746, n_557, n_558);
  nand g1412 (n_1747, n_559, n_558);
  nand g1413 (n_1748, n_557, n_559);
  nand g1414 (n_112, n_1746, n_1747, n_1748);
  xor g1415 (n_1749, A[31], A[29]);
  xor g1416 (n_564, n_1749, A[25]);
  nand g1417 (n_1750, A[31], A[29]);
  nand g1418 (n_1751, A[25], A[29]);
  nand g1419 (n_1752, A[31], A[25]);
  nand g1420 (n_574, n_1750, n_1751, n_1752);
  xor g1422 (n_565, n_1309, A[23]);
  nand g1424 (n_1755, A[23], A[15]);
  nand g1426 (n_575, n_1310, n_1755, n_1496);
  xor g1427 (n_1757, A[13], A[27]);
  xor g1428 (n_563, n_1757, A[21]);
  nand g1429 (n_1758, A[13], A[27]);
  nand g1432 (n_576, n_1758, n_1624, n_1691);
  xor g1433 (n_1761, A[19], n_560);
  xor g1434 (n_567, n_1761, n_561);
  nand g1435 (n_1762, A[19], n_560);
  nand g1436 (n_1763, n_561, n_560);
  nand g1437 (n_1764, A[19], n_561);
  nand g1438 (n_580, n_1762, n_1763, n_1764);
  xor g1439 (n_1765, n_562, n_563);
  xor g1440 (n_569, n_1765, n_564);
  nand g1441 (n_1766, n_562, n_563);
  nand g1442 (n_1767, n_564, n_563);
  nand g1443 (n_1768, n_562, n_564);
  nand g1444 (n_582, n_1766, n_1767, n_1768);
  xor g1445 (n_1769, n_565, n_566);
  xor g1446 (n_571, n_1769, n_567);
  nand g1447 (n_1770, n_565, n_566);
  nand g1448 (n_1771, n_567, n_566);
  nand g1449 (n_1772, n_565, n_567);
  nand g1450 (n_584, n_1770, n_1771, n_1772);
  xor g1451 (n_1773, n_568, n_569);
  xor g1452 (n_572, n_1773, n_570);
  nand g1453 (n_1774, n_568, n_569);
  nand g1454 (n_1775, n_570, n_569);
  nand g1455 (n_1776, n_568, n_570);
  nand g1456 (n_587, n_1774, n_1775, n_1776);
  xor g1457 (n_1777, n_571, n_572);
  xor g1458 (n_193, n_1777, n_573);
  nand g1459 (n_1778, n_571, n_572);
  nand g1460 (n_1779, n_573, n_572);
  nand g1461 (n_1780, n_571, n_573);
  nand g1462 (n_111, n_1778, n_1779, n_1780);
  xor g1463 (n_1781, A[32], A[30]);
  xor g1464 (n_578, n_1781, A[26]);
  nand g1465 (n_1782, A[32], A[30]);
  nand g1466 (n_1783, A[26], A[30]);
  nand g1467 (n_1784, A[32], A[26]);
  nand g1468 (n_588, n_1782, n_1783, n_1784);
  xor g1470 (n_579, n_385, A[24]);
  nand g1472 (n_1787, A[24], A[16]);
  xor g1475 (n_1789, A[14], A[28]);
  xor g1476 (n_577, n_1789, A[22]);
  nand g1477 (n_1790, A[14], A[28]);
  nand g1480 (n_590, n_1790, n_1656, n_1723);
  xor g1481 (n_1793, A[20], n_574);
  xor g1482 (n_581, n_1793, n_575);
  nand g1483 (n_1794, A[20], n_574);
  nand g1484 (n_1795, n_575, n_574);
  nand g1485 (n_1796, A[20], n_575);
  nand g1486 (n_594, n_1794, n_1795, n_1796);
  xor g1487 (n_1797, n_576, n_577);
  xor g1488 (n_583, n_1797, n_578);
  nand g1489 (n_1798, n_576, n_577);
  nand g1490 (n_1799, n_578, n_577);
  nand g1491 (n_1800, n_576, n_578);
  nand g1492 (n_596, n_1798, n_1799, n_1800);
  xor g1493 (n_1801, n_579, n_580);
  xor g1494 (n_585, n_1801, n_581);
  nand g1495 (n_1802, n_579, n_580);
  nand g1496 (n_1803, n_581, n_580);
  nand g1497 (n_1804, n_579, n_581);
  nand g1498 (n_598, n_1802, n_1803, n_1804);
  xor g1499 (n_1805, n_582, n_583);
  xor g1500 (n_586, n_1805, n_584);
  nand g1501 (n_1806, n_582, n_583);
  nand g1502 (n_1807, n_584, n_583);
  nand g1503 (n_1808, n_582, n_584);
  nand g1504 (n_601, n_1806, n_1807, n_1808);
  xor g1505 (n_1809, n_585, n_586);
  xor g1506 (n_192, n_1809, n_587);
  nand g1507 (n_1810, n_585, n_586);
  nand g1508 (n_1811, n_587, n_586);
  nand g1509 (n_1812, n_585, n_587);
  nand g1510 (n_110, n_1810, n_1811, n_1812);
  xor g1511 (n_1813, A[33], A[31]);
  xor g1512 (n_592, n_1813, A[27]);
  nand g1513 (n_1814, A[33], A[31]);
  nand g1514 (n_1815, A[27], A[31]);
  nand g1515 (n_1816, A[33], A[27]);
  nand g1516 (n_602, n_1814, n_1815, n_1816);
  xor g1518 (n_593, n_1365, A[25]);
  nand g1520 (n_1819, A[25], A[17]);
  nand g1522 (n_603, n_1366, n_1819, n_1560);
  xor g1523 (n_1821, A[15], A[29]);
  xor g1524 (n_591, n_1821, A[23]);
  nand g1525 (n_1822, A[15], A[29]);
  nand g1528 (n_604, n_1822, n_1688, n_1755);
  xor g1529 (n_1825, A[21], n_588);
  xor g1530 (n_595, n_1825, n_589);
  nand g1531 (n_1826, A[21], n_588);
  nand g1532 (n_1827, n_589, n_588);
  nand g1533 (n_1828, A[21], n_589);
  nand g1534 (n_608, n_1826, n_1827, n_1828);
  xor g1535 (n_1829, n_590, n_591);
  xor g1536 (n_597, n_1829, n_592);
  nand g1537 (n_1830, n_590, n_591);
  nand g1538 (n_1831, n_592, n_591);
  nand g1539 (n_1832, n_590, n_592);
  nand g1540 (n_610, n_1830, n_1831, n_1832);
  xor g1541 (n_1833, n_593, n_594);
  xor g1542 (n_599, n_1833, n_595);
  nand g1543 (n_1834, n_593, n_594);
  nand g1544 (n_1835, n_595, n_594);
  nand g1545 (n_1836, n_593, n_595);
  nand g1546 (n_612, n_1834, n_1835, n_1836);
  xor g1547 (n_1837, n_596, n_597);
  xor g1548 (n_600, n_1837, n_598);
  nand g1549 (n_1838, n_596, n_597);
  nand g1550 (n_1839, n_598, n_597);
  nand g1551 (n_1840, n_596, n_598);
  nand g1552 (n_615, n_1838, n_1839, n_1840);
  xor g1553 (n_1841, n_599, n_600);
  xor g1554 (n_191, n_1841, n_601);
  nand g1555 (n_1842, n_599, n_600);
  nand g1556 (n_1843, n_601, n_600);
  nand g1557 (n_1844, n_599, n_601);
  nand g1558 (n_109, n_1842, n_1843, n_1844);
  xor g1559 (n_1845, A[34], A[32]);
  xor g1560 (n_606, n_1845, A[28]);
  nand g1561 (n_1846, A[34], A[32]);
  nand g1562 (n_1847, A[28], A[32]);
  nand g1563 (n_1848, A[34], A[28]);
  nand g1564 (n_616, n_1846, n_1847, n_1848);
  xor g1566 (n_607, n_1397, A[26]);
  nand g1568 (n_1851, A[26], A[18]);
  nand g1570 (n_617, n_1398, n_1851, n_1592);
  xor g1571 (n_1853, A[16], A[30]);
  xor g1572 (n_605, n_1853, A[24]);
  nand g1573 (n_1854, A[16], A[30]);
  nand g1576 (n_618, n_1854, n_1720, n_1787);
  xor g1577 (n_1857, A[22], n_602);
  xor g1578 (n_609, n_1857, n_603);
  nand g1579 (n_1858, A[22], n_602);
  nand g1580 (n_1859, n_603, n_602);
  nand g1581 (n_1860, A[22], n_603);
  nand g1582 (n_622, n_1858, n_1859, n_1860);
  xor g1583 (n_1861, n_604, n_605);
  xor g1584 (n_611, n_1861, n_606);
  nand g1585 (n_1862, n_604, n_605);
  nand g1586 (n_1863, n_606, n_605);
  nand g1587 (n_1864, n_604, n_606);
  nand g1588 (n_624, n_1862, n_1863, n_1864);
  xor g1589 (n_1865, n_607, n_608);
  xor g1590 (n_613, n_1865, n_609);
  nand g1591 (n_1866, n_607, n_608);
  nand g1592 (n_1867, n_609, n_608);
  nand g1593 (n_1868, n_607, n_609);
  nand g1594 (n_626, n_1866, n_1867, n_1868);
  xor g1595 (n_1869, n_610, n_611);
  xor g1596 (n_614, n_1869, n_612);
  nand g1597 (n_1870, n_610, n_611);
  nand g1598 (n_1871, n_612, n_611);
  nand g1599 (n_1872, n_610, n_612);
  nand g1600 (n_629, n_1870, n_1871, n_1872);
  xor g1601 (n_1873, n_613, n_614);
  xor g1602 (n_190, n_1873, n_615);
  nand g1603 (n_1874, n_613, n_614);
  nand g1604 (n_1875, n_615, n_614);
  nand g1605 (n_1876, n_613, n_615);
  nand g1606 (n_108, n_1874, n_1875, n_1876);
  xor g1607 (n_1877, A[35], A[33]);
  xor g1608 (n_620, n_1877, A[29]);
  nand g1609 (n_1878, A[35], A[33]);
  nand g1610 (n_1879, A[29], A[33]);
  nand g1611 (n_1880, A[35], A[29]);
  nand g1612 (n_630, n_1878, n_1879, n_1880);
  xor g1614 (n_621, n_1429, A[27]);
  nand g1616 (n_1883, A[27], A[19]);
  nand g1618 (n_631, n_1430, n_1883, n_1624);
  xor g1619 (n_1885, A[17], A[31]);
  xor g1620 (n_619, n_1885, A[25]);
  nand g1621 (n_1886, A[17], A[31]);
  nand g1624 (n_632, n_1886, n_1752, n_1819);
  xor g1625 (n_1889, A[23], n_616);
  xor g1626 (n_623, n_1889, n_617);
  nand g1627 (n_1890, A[23], n_616);
  nand g1628 (n_1891, n_617, n_616);
  nand g1629 (n_1892, A[23], n_617);
  nand g1630 (n_636, n_1890, n_1891, n_1892);
  xor g1631 (n_1893, n_618, n_619);
  xor g1632 (n_625, n_1893, n_620);
  nand g1633 (n_1894, n_618, n_619);
  nand g1634 (n_1895, n_620, n_619);
  nand g1635 (n_1896, n_618, n_620);
  nand g1636 (n_638, n_1894, n_1895, n_1896);
  xor g1637 (n_1897, n_621, n_622);
  xor g1638 (n_627, n_1897, n_623);
  nand g1639 (n_1898, n_621, n_622);
  nand g1640 (n_1899, n_623, n_622);
  nand g1641 (n_1900, n_621, n_623);
  nand g1642 (n_640, n_1898, n_1899, n_1900);
  xor g1643 (n_1901, n_624, n_625);
  xor g1644 (n_628, n_1901, n_626);
  nand g1645 (n_1902, n_624, n_625);
  nand g1646 (n_1903, n_626, n_625);
  nand g1647 (n_1904, n_624, n_626);
  nand g1648 (n_643, n_1902, n_1903, n_1904);
  xor g1649 (n_1905, n_627, n_628);
  xor g1650 (n_189, n_1905, n_629);
  nand g1651 (n_1906, n_627, n_628);
  nand g1652 (n_1907, n_629, n_628);
  nand g1653 (n_1908, n_627, n_629);
  nand g1654 (n_107, n_1906, n_1907, n_1908);
  xor g1655 (n_1909, A[36], A[34]);
  xor g1656 (n_634, n_1909, A[30]);
  nand g1657 (n_1910, A[36], A[34]);
  nand g1658 (n_1911, A[30], A[34]);
  nand g1659 (n_1912, A[36], A[30]);
  nand g1660 (n_644, n_1910, n_1911, n_1912);
  xor g1662 (n_635, n_1461, A[28]);
  nand g1664 (n_1915, A[28], A[20]);
  nand g1666 (n_645, n_1462, n_1915, n_1656);
  xor g1667 (n_1917, A[18], A[32]);
  xor g1668 (n_633, n_1917, A[26]);
  nand g1669 (n_1918, A[18], A[32]);
  nand g1672 (n_646, n_1918, n_1784, n_1851);
  xor g1673 (n_1921, A[24], n_630);
  xor g1674 (n_637, n_1921, n_631);
  nand g1675 (n_1922, A[24], n_630);
  nand g1676 (n_1923, n_631, n_630);
  nand g1677 (n_1924, A[24], n_631);
  nand g1678 (n_650, n_1922, n_1923, n_1924);
  xor g1679 (n_1925, n_632, n_633);
  xor g1680 (n_639, n_1925, n_634);
  nand g1681 (n_1926, n_632, n_633);
  nand g1682 (n_1927, n_634, n_633);
  nand g1683 (n_1928, n_632, n_634);
  nand g1684 (n_652, n_1926, n_1927, n_1928);
  xor g1685 (n_1929, n_635, n_636);
  xor g1686 (n_641, n_1929, n_637);
  nand g1687 (n_1930, n_635, n_636);
  nand g1688 (n_1931, n_637, n_636);
  nand g1689 (n_1932, n_635, n_637);
  nand g1690 (n_654, n_1930, n_1931, n_1932);
  xor g1691 (n_1933, n_638, n_639);
  xor g1692 (n_642, n_1933, n_640);
  nand g1693 (n_1934, n_638, n_639);
  nand g1694 (n_1935, n_640, n_639);
  nand g1695 (n_1936, n_638, n_640);
  nand g1696 (n_657, n_1934, n_1935, n_1936);
  xor g1697 (n_1937, n_641, n_642);
  xor g1698 (n_188, n_1937, n_643);
  nand g1699 (n_1938, n_641, n_642);
  nand g1700 (n_1939, n_643, n_642);
  nand g1701 (n_1940, n_641, n_643);
  nand g1702 (n_106, n_1938, n_1939, n_1940);
  xor g1703 (n_1941, A[37], A[35]);
  xor g1704 (n_648, n_1941, A[31]);
  nand g1705 (n_1942, A[37], A[35]);
  nand g1706 (n_1943, A[31], A[35]);
  nand g1707 (n_1944, A[37], A[31]);
  nand g1708 (n_658, n_1942, n_1943, n_1944);
  xor g1710 (n_649, n_1493, A[29]);
  nand g1712 (n_1947, A[29], A[21]);
  nand g1714 (n_659, n_1494, n_1947, n_1688);
  xor g1715 (n_1949, A[19], A[33]);
  xor g1716 (n_647, n_1949, A[27]);
  nand g1717 (n_1950, A[19], A[33]);
  nand g1720 (n_660, n_1950, n_1816, n_1883);
  xor g1721 (n_1953, A[25], n_644);
  xor g1722 (n_651, n_1953, n_645);
  nand g1723 (n_1954, A[25], n_644);
  nand g1724 (n_1955, n_645, n_644);
  nand g1725 (n_1956, A[25], n_645);
  nand g1726 (n_664, n_1954, n_1955, n_1956);
  xor g1727 (n_1957, n_646, n_647);
  xor g1728 (n_653, n_1957, n_648);
  nand g1729 (n_1958, n_646, n_647);
  nand g1730 (n_1959, n_648, n_647);
  nand g1731 (n_1960, n_646, n_648);
  nand g1732 (n_666, n_1958, n_1959, n_1960);
  xor g1733 (n_1961, n_649, n_650);
  xor g1734 (n_655, n_1961, n_651);
  nand g1735 (n_1962, n_649, n_650);
  nand g1736 (n_1963, n_651, n_650);
  nand g1737 (n_1964, n_649, n_651);
  nand g1738 (n_668, n_1962, n_1963, n_1964);
  xor g1739 (n_1965, n_652, n_653);
  xor g1740 (n_656, n_1965, n_654);
  nand g1741 (n_1966, n_652, n_653);
  nand g1742 (n_1967, n_654, n_653);
  nand g1743 (n_1968, n_652, n_654);
  nand g1744 (n_671, n_1966, n_1967, n_1968);
  xor g1745 (n_1969, n_655, n_656);
  xor g1746 (n_187, n_1969, n_657);
  nand g1747 (n_1970, n_655, n_656);
  nand g1748 (n_1971, n_657, n_656);
  nand g1749 (n_1972, n_655, n_657);
  nand g1750 (n_105, n_1970, n_1971, n_1972);
  xor g1751 (n_1973, A[38], A[36]);
  xor g1752 (n_662, n_1973, A[32]);
  nand g1753 (n_1974, A[38], A[36]);
  nand g1754 (n_1975, A[32], A[36]);
  nand g1755 (n_1976, A[38], A[32]);
  nand g1756 (n_672, n_1974, n_1975, n_1976);
  xor g1758 (n_663, n_1525, A[30]);
  nand g1760 (n_1979, A[30], A[22]);
  nand g1762 (n_673, n_1526, n_1979, n_1720);
  xor g1763 (n_1981, A[20], A[34]);
  xor g1764 (n_661, n_1981, A[28]);
  nand g1765 (n_1982, A[20], A[34]);
  nand g1768 (n_674, n_1982, n_1848, n_1915);
  xor g1769 (n_1985, A[26], n_658);
  xor g1770 (n_665, n_1985, n_659);
  nand g1771 (n_1986, A[26], n_658);
  nand g1772 (n_1987, n_659, n_658);
  nand g1773 (n_1988, A[26], n_659);
  nand g1774 (n_678, n_1986, n_1987, n_1988);
  xor g1775 (n_1989, n_660, n_661);
  xor g1776 (n_667, n_1989, n_662);
  nand g1777 (n_1990, n_660, n_661);
  nand g1778 (n_1991, n_662, n_661);
  nand g1779 (n_1992, n_660, n_662);
  nand g1780 (n_680, n_1990, n_1991, n_1992);
  xor g1781 (n_1993, n_663, n_664);
  xor g1782 (n_669, n_1993, n_665);
  nand g1783 (n_1994, n_663, n_664);
  nand g1784 (n_1995, n_665, n_664);
  nand g1785 (n_1996, n_663, n_665);
  nand g1786 (n_682, n_1994, n_1995, n_1996);
  xor g1787 (n_1997, n_666, n_667);
  xor g1788 (n_670, n_1997, n_668);
  nand g1789 (n_1998, n_666, n_667);
  nand g1790 (n_1999, n_668, n_667);
  nand g1791 (n_2000, n_666, n_668);
  nand g1792 (n_685, n_1998, n_1999, n_2000);
  xor g1793 (n_2001, n_669, n_670);
  xor g1794 (n_186, n_2001, n_671);
  nand g1795 (n_2002, n_669, n_670);
  nand g1796 (n_2003, n_671, n_670);
  nand g1797 (n_2004, n_669, n_671);
  nand g1798 (n_104, n_2002, n_2003, n_2004);
  xor g1799 (n_2005, A[39], A[37]);
  xor g1800 (n_676, n_2005, A[33]);
  nand g1801 (n_2006, A[39], A[37]);
  nand g1802 (n_2007, A[33], A[37]);
  nand g1803 (n_2008, A[39], A[33]);
  nand g1804 (n_686, n_2006, n_2007, n_2008);
  xor g1806 (n_677, n_1557, A[31]);
  nand g1808 (n_2011, A[31], A[23]);
  nand g1810 (n_687, n_1558, n_2011, n_1752);
  xor g1811 (n_2013, A[21], A[35]);
  xor g1812 (n_675, n_2013, A[29]);
  nand g1813 (n_2014, A[21], A[35]);
  nand g1816 (n_688, n_2014, n_1880, n_1947);
  xor g1817 (n_2017, A[27], n_672);
  xor g1818 (n_679, n_2017, n_673);
  nand g1819 (n_2018, A[27], n_672);
  nand g1820 (n_2019, n_673, n_672);
  nand g1821 (n_2020, A[27], n_673);
  nand g1822 (n_692, n_2018, n_2019, n_2020);
  xor g1823 (n_2021, n_674, n_675);
  xor g1824 (n_681, n_2021, n_676);
  nand g1825 (n_2022, n_674, n_675);
  nand g1826 (n_2023, n_676, n_675);
  nand g1827 (n_2024, n_674, n_676);
  nand g1828 (n_694, n_2022, n_2023, n_2024);
  xor g1829 (n_2025, n_677, n_678);
  xor g1830 (n_683, n_2025, n_679);
  nand g1831 (n_2026, n_677, n_678);
  nand g1832 (n_2027, n_679, n_678);
  nand g1833 (n_2028, n_677, n_679);
  nand g1834 (n_696, n_2026, n_2027, n_2028);
  xor g1835 (n_2029, n_680, n_681);
  xor g1836 (n_684, n_2029, n_682);
  nand g1837 (n_2030, n_680, n_681);
  nand g1838 (n_2031, n_682, n_681);
  nand g1839 (n_2032, n_680, n_682);
  nand g1840 (n_699, n_2030, n_2031, n_2032);
  xor g1841 (n_2033, n_683, n_684);
  xor g1842 (n_185, n_2033, n_685);
  nand g1843 (n_2034, n_683, n_684);
  nand g1844 (n_2035, n_685, n_684);
  nand g1845 (n_2036, n_683, n_685);
  nand g1846 (n_103, n_2034, n_2035, n_2036);
  xor g1847 (n_2037, A[40], A[38]);
  xor g1848 (n_690, n_2037, A[34]);
  nand g1849 (n_2038, A[40], A[38]);
  nand g1850 (n_2039, A[34], A[38]);
  nand g1851 (n_2040, A[40], A[34]);
  nand g1852 (n_700, n_2038, n_2039, n_2040);
  xor g1854 (n_691, n_1589, A[32]);
  nand g1856 (n_2043, A[32], A[24]);
  nand g1858 (n_701, n_1590, n_2043, n_1784);
  xor g1859 (n_2045, A[22], A[36]);
  xor g1860 (n_689, n_2045, A[30]);
  nand g1861 (n_2046, A[22], A[36]);
  nand g1864 (n_702, n_2046, n_1912, n_1979);
  xor g1865 (n_2049, A[28], n_686);
  xor g1866 (n_693, n_2049, n_687);
  nand g1867 (n_2050, A[28], n_686);
  nand g1868 (n_2051, n_687, n_686);
  nand g1869 (n_2052, A[28], n_687);
  nand g1870 (n_706, n_2050, n_2051, n_2052);
  xor g1871 (n_2053, n_688, n_689);
  xor g1872 (n_695, n_2053, n_690);
  nand g1873 (n_2054, n_688, n_689);
  nand g1874 (n_2055, n_690, n_689);
  nand g1875 (n_2056, n_688, n_690);
  nand g1876 (n_708, n_2054, n_2055, n_2056);
  xor g1877 (n_2057, n_691, n_692);
  xor g1878 (n_697, n_2057, n_693);
  nand g1879 (n_2058, n_691, n_692);
  nand g1880 (n_2059, n_693, n_692);
  nand g1881 (n_2060, n_691, n_693);
  nand g1882 (n_710, n_2058, n_2059, n_2060);
  xor g1883 (n_2061, n_694, n_695);
  xor g1884 (n_698, n_2061, n_696);
  nand g1885 (n_2062, n_694, n_695);
  nand g1886 (n_2063, n_696, n_695);
  nand g1887 (n_2064, n_694, n_696);
  nand g1888 (n_713, n_2062, n_2063, n_2064);
  xor g1889 (n_2065, n_697, n_698);
  xor g1890 (n_184, n_2065, n_699);
  nand g1891 (n_2066, n_697, n_698);
  nand g1892 (n_2067, n_699, n_698);
  nand g1893 (n_2068, n_697, n_699);
  nand g1894 (n_102, n_2066, n_2067, n_2068);
  xor g1895 (n_2069, A[41], A[39]);
  xor g1896 (n_704, n_2069, A[35]);
  nand g1897 (n_2070, A[41], A[39]);
  nand g1898 (n_2071, A[35], A[39]);
  nand g1899 (n_2072, A[41], A[35]);
  nand g1900 (n_714, n_2070, n_2071, n_2072);
  xor g1902 (n_705, n_1621, A[33]);
  nand g1904 (n_2075, A[33], A[25]);
  nand g1906 (n_715, n_1622, n_2075, n_1816);
  xor g1907 (n_2077, A[23], A[37]);
  xor g1908 (n_703, n_2077, A[31]);
  nand g1909 (n_2078, A[23], A[37]);
  nand g1912 (n_716, n_2078, n_1944, n_2011);
  xor g1913 (n_2081, A[29], n_700);
  xor g1914 (n_707, n_2081, n_701);
  nand g1915 (n_2082, A[29], n_700);
  nand g1916 (n_2083, n_701, n_700);
  nand g1917 (n_2084, A[29], n_701);
  nand g1918 (n_720, n_2082, n_2083, n_2084);
  xor g1919 (n_2085, n_702, n_703);
  xor g1920 (n_709, n_2085, n_704);
  nand g1921 (n_2086, n_702, n_703);
  nand g1922 (n_2087, n_704, n_703);
  nand g1923 (n_2088, n_702, n_704);
  nand g1924 (n_722, n_2086, n_2087, n_2088);
  xor g1925 (n_2089, n_705, n_706);
  xor g1926 (n_711, n_2089, n_707);
  nand g1927 (n_2090, n_705, n_706);
  nand g1928 (n_2091, n_707, n_706);
  nand g1929 (n_2092, n_705, n_707);
  nand g1930 (n_724, n_2090, n_2091, n_2092);
  xor g1931 (n_2093, n_708, n_709);
  xor g1932 (n_712, n_2093, n_710);
  nand g1933 (n_2094, n_708, n_709);
  nand g1934 (n_2095, n_710, n_709);
  nand g1935 (n_2096, n_708, n_710);
  nand g1936 (n_727, n_2094, n_2095, n_2096);
  xor g1937 (n_2097, n_711, n_712);
  xor g1938 (n_183, n_2097, n_713);
  nand g1939 (n_2098, n_711, n_712);
  nand g1940 (n_2099, n_713, n_712);
  nand g1941 (n_2100, n_711, n_713);
  nand g1942 (n_101, n_2098, n_2099, n_2100);
  xor g1943 (n_2101, A[42], A[40]);
  xor g1944 (n_718, n_2101, A[36]);
  nand g1945 (n_2102, A[42], A[40]);
  nand g1946 (n_2103, A[36], A[40]);
  nand g1947 (n_2104, A[42], A[36]);
  nand g1948 (n_728, n_2102, n_2103, n_2104);
  xor g1950 (n_719, n_1653, A[34]);
  nand g1952 (n_2107, A[34], A[26]);
  nand g1954 (n_729, n_1654, n_2107, n_1848);
  xor g1955 (n_2109, A[24], A[38]);
  xor g1956 (n_717, n_2109, A[32]);
  nand g1957 (n_2110, A[24], A[38]);
  nand g1960 (n_730, n_2110, n_1976, n_2043);
  xor g1961 (n_2113, A[30], n_714);
  xor g1962 (n_721, n_2113, n_715);
  nand g1963 (n_2114, A[30], n_714);
  nand g1964 (n_2115, n_715, n_714);
  nand g1965 (n_2116, A[30], n_715);
  nand g1966 (n_734, n_2114, n_2115, n_2116);
  xor g1967 (n_2117, n_716, n_717);
  xor g1968 (n_723, n_2117, n_718);
  nand g1969 (n_2118, n_716, n_717);
  nand g1970 (n_2119, n_718, n_717);
  nand g1971 (n_2120, n_716, n_718);
  nand g1972 (n_736, n_2118, n_2119, n_2120);
  xor g1973 (n_2121, n_719, n_720);
  xor g1974 (n_725, n_2121, n_721);
  nand g1975 (n_2122, n_719, n_720);
  nand g1976 (n_2123, n_721, n_720);
  nand g1977 (n_2124, n_719, n_721);
  nand g1978 (n_738, n_2122, n_2123, n_2124);
  xor g1979 (n_2125, n_722, n_723);
  xor g1980 (n_726, n_2125, n_724);
  nand g1981 (n_2126, n_722, n_723);
  nand g1982 (n_2127, n_724, n_723);
  nand g1983 (n_2128, n_722, n_724);
  nand g1984 (n_741, n_2126, n_2127, n_2128);
  xor g1985 (n_2129, n_725, n_726);
  xor g1986 (n_182, n_2129, n_727);
  nand g1987 (n_2130, n_725, n_726);
  nand g1988 (n_2131, n_727, n_726);
  nand g1989 (n_2132, n_725, n_727);
  nand g1990 (n_100, n_2130, n_2131, n_2132);
  xor g1991 (n_2133, A[43], A[41]);
  xor g1992 (n_732, n_2133, A[37]);
  nand g1993 (n_2134, A[43], A[41]);
  nand g1994 (n_2135, A[37], A[41]);
  nand g1995 (n_2136, A[43], A[37]);
  nand g1996 (n_742, n_2134, n_2135, n_2136);
  xor g1998 (n_733, n_1685, A[35]);
  nand g2000 (n_2139, A[35], A[27]);
  nand g2002 (n_743, n_1686, n_2139, n_1880);
  xor g2003 (n_2141, A[25], A[39]);
  xor g2004 (n_731, n_2141, A[33]);
  nand g2005 (n_2142, A[25], A[39]);
  nand g2008 (n_744, n_2142, n_2008, n_2075);
  xor g2009 (n_2145, A[31], n_728);
  xor g2010 (n_735, n_2145, n_729);
  nand g2011 (n_2146, A[31], n_728);
  nand g2012 (n_2147, n_729, n_728);
  nand g2013 (n_2148, A[31], n_729);
  nand g2014 (n_748, n_2146, n_2147, n_2148);
  xor g2015 (n_2149, n_730, n_731);
  xor g2016 (n_737, n_2149, n_732);
  nand g2017 (n_2150, n_730, n_731);
  nand g2018 (n_2151, n_732, n_731);
  nand g2019 (n_2152, n_730, n_732);
  nand g2020 (n_750, n_2150, n_2151, n_2152);
  xor g2021 (n_2153, n_733, n_734);
  xor g2022 (n_739, n_2153, n_735);
  nand g2023 (n_2154, n_733, n_734);
  nand g2024 (n_2155, n_735, n_734);
  nand g2025 (n_2156, n_733, n_735);
  nand g2026 (n_752, n_2154, n_2155, n_2156);
  xor g2027 (n_2157, n_736, n_737);
  xor g2028 (n_740, n_2157, n_738);
  nand g2029 (n_2158, n_736, n_737);
  nand g2030 (n_2159, n_738, n_737);
  nand g2031 (n_2160, n_736, n_738);
  nand g2032 (n_755, n_2158, n_2159, n_2160);
  xor g2033 (n_2161, n_739, n_740);
  xor g2034 (n_181, n_2161, n_741);
  nand g2035 (n_2162, n_739, n_740);
  nand g2036 (n_2163, n_741, n_740);
  nand g2037 (n_2164, n_739, n_741);
  nand g2038 (n_99, n_2162, n_2163, n_2164);
  xor g2039 (n_2165, A[44], A[42]);
  xor g2040 (n_746, n_2165, A[38]);
  nand g2041 (n_2166, A[44], A[42]);
  nand g2042 (n_2167, A[38], A[42]);
  nand g2043 (n_2168, A[44], A[38]);
  nand g2044 (n_756, n_2166, n_2167, n_2168);
  xor g2046 (n_747, n_1717, A[36]);
  nand g2048 (n_2171, A[36], A[28]);
  nand g2050 (n_757, n_1718, n_2171, n_1912);
  xor g2051 (n_2173, A[26], A[40]);
  xor g2052 (n_745, n_2173, A[34]);
  nand g2053 (n_2174, A[26], A[40]);
  nand g2056 (n_758, n_2174, n_2040, n_2107);
  xor g2057 (n_2177, A[32], n_742);
  xor g2058 (n_749, n_2177, n_743);
  nand g2059 (n_2178, A[32], n_742);
  nand g2060 (n_2179, n_743, n_742);
  nand g2061 (n_2180, A[32], n_743);
  nand g2062 (n_762, n_2178, n_2179, n_2180);
  xor g2063 (n_2181, n_744, n_745);
  xor g2064 (n_751, n_2181, n_746);
  nand g2065 (n_2182, n_744, n_745);
  nand g2066 (n_2183, n_746, n_745);
  nand g2067 (n_2184, n_744, n_746);
  nand g2068 (n_764, n_2182, n_2183, n_2184);
  xor g2069 (n_2185, n_747, n_748);
  xor g2070 (n_753, n_2185, n_749);
  nand g2071 (n_2186, n_747, n_748);
  nand g2072 (n_2187, n_749, n_748);
  nand g2073 (n_2188, n_747, n_749);
  nand g2074 (n_766, n_2186, n_2187, n_2188);
  xor g2075 (n_2189, n_750, n_751);
  xor g2076 (n_754, n_2189, n_752);
  nand g2077 (n_2190, n_750, n_751);
  nand g2078 (n_2191, n_752, n_751);
  nand g2079 (n_2192, n_750, n_752);
  nand g2080 (n_769, n_2190, n_2191, n_2192);
  xor g2081 (n_2193, n_753, n_754);
  xor g2082 (n_180, n_2193, n_755);
  nand g2083 (n_2194, n_753, n_754);
  nand g2084 (n_2195, n_755, n_754);
  nand g2085 (n_2196, n_753, n_755);
  nand g2086 (n_98, n_2194, n_2195, n_2196);
  xor g2087 (n_2197, A[45], A[43]);
  xor g2088 (n_760, n_2197, A[39]);
  nand g2089 (n_2198, A[45], A[43]);
  nand g2090 (n_2199, A[39], A[43]);
  nand g2091 (n_2200, A[45], A[39]);
  nand g2092 (n_770, n_2198, n_2199, n_2200);
  xor g2094 (n_761, n_1749, A[37]);
  nand g2096 (n_2203, A[37], A[29]);
  nand g2098 (n_771, n_1750, n_2203, n_1944);
  xor g2099 (n_2205, A[27], A[41]);
  xor g2100 (n_759, n_2205, A[35]);
  nand g2101 (n_2206, A[27], A[41]);
  nand g2104 (n_772, n_2206, n_2072, n_2139);
  xor g2105 (n_2209, A[33], n_756);
  xor g2106 (n_763, n_2209, n_757);
  nand g2107 (n_2210, A[33], n_756);
  nand g2108 (n_2211, n_757, n_756);
  nand g2109 (n_2212, A[33], n_757);
  nand g2110 (n_776, n_2210, n_2211, n_2212);
  xor g2111 (n_2213, n_758, n_759);
  xor g2112 (n_765, n_2213, n_760);
  nand g2113 (n_2214, n_758, n_759);
  nand g2114 (n_2215, n_760, n_759);
  nand g2115 (n_2216, n_758, n_760);
  nand g2116 (n_778, n_2214, n_2215, n_2216);
  xor g2117 (n_2217, n_761, n_762);
  xor g2118 (n_767, n_2217, n_763);
  nand g2119 (n_2218, n_761, n_762);
  nand g2120 (n_2219, n_763, n_762);
  nand g2121 (n_2220, n_761, n_763);
  nand g2122 (n_780, n_2218, n_2219, n_2220);
  xor g2123 (n_2221, n_764, n_765);
  xor g2124 (n_768, n_2221, n_766);
  nand g2125 (n_2222, n_764, n_765);
  nand g2126 (n_2223, n_766, n_765);
  nand g2127 (n_2224, n_764, n_766);
  nand g2128 (n_783, n_2222, n_2223, n_2224);
  xor g2129 (n_2225, n_767, n_768);
  xor g2130 (n_179, n_2225, n_769);
  nand g2131 (n_2226, n_767, n_768);
  nand g2132 (n_2227, n_769, n_768);
  nand g2133 (n_2228, n_767, n_769);
  nand g2134 (n_97, n_2226, n_2227, n_2228);
  xor g2135 (n_2229, A[46], A[44]);
  xor g2136 (n_774, n_2229, A[40]);
  nand g2137 (n_2230, A[46], A[44]);
  nand g2138 (n_2231, A[40], A[44]);
  nand g2139 (n_2232, A[46], A[40]);
  nand g2140 (n_784, n_2230, n_2231, n_2232);
  xor g2142 (n_775, n_1781, A[38]);
  nand g2144 (n_2235, A[38], A[30]);
  nand g2146 (n_785, n_1782, n_2235, n_1976);
  xor g2147 (n_2237, A[28], A[42]);
  xor g2148 (n_773, n_2237, A[36]);
  nand g2149 (n_2238, A[28], A[42]);
  nand g2152 (n_786, n_2238, n_2104, n_2171);
  xor g2153 (n_2241, A[34], n_770);
  xor g2154 (n_777, n_2241, n_771);
  nand g2155 (n_2242, A[34], n_770);
  nand g2156 (n_2243, n_771, n_770);
  nand g2157 (n_2244, A[34], n_771);
  nand g2158 (n_790, n_2242, n_2243, n_2244);
  xor g2159 (n_2245, n_772, n_773);
  xor g2160 (n_779, n_2245, n_774);
  nand g2161 (n_2246, n_772, n_773);
  nand g2162 (n_2247, n_774, n_773);
  nand g2163 (n_2248, n_772, n_774);
  nand g2164 (n_792, n_2246, n_2247, n_2248);
  xor g2165 (n_2249, n_775, n_776);
  xor g2166 (n_781, n_2249, n_777);
  nand g2167 (n_2250, n_775, n_776);
  nand g2168 (n_2251, n_777, n_776);
  nand g2169 (n_2252, n_775, n_777);
  nand g2170 (n_794, n_2250, n_2251, n_2252);
  xor g2171 (n_2253, n_778, n_779);
  xor g2172 (n_782, n_2253, n_780);
  nand g2173 (n_2254, n_778, n_779);
  nand g2174 (n_2255, n_780, n_779);
  nand g2175 (n_2256, n_778, n_780);
  nand g2176 (n_797, n_2254, n_2255, n_2256);
  xor g2177 (n_2257, n_781, n_782);
  xor g2178 (n_178, n_2257, n_783);
  nand g2179 (n_2258, n_781, n_782);
  nand g2180 (n_2259, n_783, n_782);
  nand g2181 (n_2260, n_781, n_783);
  nand g2182 (n_96, n_2258, n_2259, n_2260);
  xor g2183 (n_2261, A[47], A[45]);
  xor g2184 (n_788, n_2261, A[41]);
  nand g2185 (n_2262, A[47], A[45]);
  nand g2186 (n_2263, A[41], A[45]);
  nand g2187 (n_2264, A[47], A[41]);
  nand g2188 (n_798, n_2262, n_2263, n_2264);
  xor g2190 (n_789, n_1813, A[39]);
  nand g2192 (n_2267, A[39], A[31]);
  nand g2194 (n_799, n_1814, n_2267, n_2008);
  xor g2195 (n_2269, A[29], A[43]);
  xor g2196 (n_787, n_2269, A[37]);
  nand g2197 (n_2270, A[29], A[43]);
  nand g2200 (n_800, n_2270, n_2136, n_2203);
  xor g2201 (n_2273, A[35], n_784);
  xor g2202 (n_791, n_2273, n_785);
  nand g2203 (n_2274, A[35], n_784);
  nand g2204 (n_2275, n_785, n_784);
  nand g2205 (n_2276, A[35], n_785);
  nand g2206 (n_804, n_2274, n_2275, n_2276);
  xor g2207 (n_2277, n_786, n_787);
  xor g2208 (n_793, n_2277, n_788);
  nand g2209 (n_2278, n_786, n_787);
  nand g2210 (n_2279, n_788, n_787);
  nand g2211 (n_2280, n_786, n_788);
  nand g2212 (n_806, n_2278, n_2279, n_2280);
  xor g2213 (n_2281, n_789, n_790);
  xor g2214 (n_795, n_2281, n_791);
  nand g2215 (n_2282, n_789, n_790);
  nand g2216 (n_2283, n_791, n_790);
  nand g2217 (n_2284, n_789, n_791);
  nand g2218 (n_808, n_2282, n_2283, n_2284);
  xor g2219 (n_2285, n_792, n_793);
  xor g2220 (n_796, n_2285, n_794);
  nand g2221 (n_2286, n_792, n_793);
  nand g2222 (n_2287, n_794, n_793);
  nand g2223 (n_2288, n_792, n_794);
  nand g2224 (n_811, n_2286, n_2287, n_2288);
  xor g2225 (n_2289, n_795, n_796);
  xor g2226 (n_177, n_2289, n_797);
  nand g2227 (n_2290, n_795, n_796);
  nand g2228 (n_2291, n_797, n_796);
  nand g2229 (n_2292, n_795, n_797);
  nand g2230 (n_95, n_2290, n_2291, n_2292);
  xor g2231 (n_2293, A[48], A[46]);
  xor g2232 (n_802, n_2293, A[42]);
  nand g2233 (n_2294, A[48], A[46]);
  nand g2234 (n_2295, A[42], A[46]);
  nand g2235 (n_2296, A[48], A[42]);
  nand g2236 (n_812, n_2294, n_2295, n_2296);
  xor g2238 (n_803, n_1845, A[40]);
  nand g2240 (n_2299, A[40], A[32]);
  nand g2242 (n_813, n_1846, n_2299, n_2040);
  xor g2243 (n_2301, A[30], A[44]);
  xor g2244 (n_801, n_2301, A[38]);
  nand g2245 (n_2302, A[30], A[44]);
  nand g2248 (n_814, n_2302, n_2168, n_2235);
  xor g2249 (n_2305, A[36], n_798);
  xor g2250 (n_805, n_2305, n_799);
  nand g2251 (n_2306, A[36], n_798);
  nand g2252 (n_2307, n_799, n_798);
  nand g2253 (n_2308, A[36], n_799);
  nand g2254 (n_818, n_2306, n_2307, n_2308);
  xor g2255 (n_2309, n_800, n_801);
  xor g2256 (n_807, n_2309, n_802);
  nand g2257 (n_2310, n_800, n_801);
  nand g2258 (n_2311, n_802, n_801);
  nand g2259 (n_2312, n_800, n_802);
  nand g2260 (n_820, n_2310, n_2311, n_2312);
  xor g2261 (n_2313, n_803, n_804);
  xor g2262 (n_809, n_2313, n_805);
  nand g2263 (n_2314, n_803, n_804);
  nand g2264 (n_2315, n_805, n_804);
  nand g2265 (n_2316, n_803, n_805);
  nand g2266 (n_822, n_2314, n_2315, n_2316);
  xor g2267 (n_2317, n_806, n_807);
  xor g2268 (n_810, n_2317, n_808);
  nand g2269 (n_2318, n_806, n_807);
  nand g2270 (n_2319, n_808, n_807);
  nand g2271 (n_2320, n_806, n_808);
  nand g2272 (n_825, n_2318, n_2319, n_2320);
  xor g2273 (n_2321, n_809, n_810);
  xor g2274 (n_176, n_2321, n_811);
  nand g2275 (n_2322, n_809, n_810);
  nand g2276 (n_2323, n_811, n_810);
  nand g2277 (n_2324, n_809, n_811);
  nand g2278 (n_94, n_2322, n_2323, n_2324);
  xor g2279 (n_2325, A[49], A[47]);
  xor g2280 (n_816, n_2325, A[43]);
  nand g2281 (n_2326, A[49], A[47]);
  nand g2282 (n_2327, A[43], A[47]);
  nand g2283 (n_2328, A[49], A[43]);
  nand g2284 (n_826, n_2326, n_2327, n_2328);
  xor g2286 (n_817, n_1877, A[41]);
  nand g2288 (n_2331, A[41], A[33]);
  nand g2290 (n_827, n_1878, n_2331, n_2072);
  xor g2291 (n_2333, A[31], A[45]);
  xor g2292 (n_815, n_2333, A[39]);
  nand g2293 (n_2334, A[31], A[45]);
  nand g2296 (n_828, n_2334, n_2200, n_2267);
  xor g2297 (n_2337, A[37], n_812);
  xor g2298 (n_819, n_2337, n_813);
  nand g2299 (n_2338, A[37], n_812);
  nand g2300 (n_2339, n_813, n_812);
  nand g2301 (n_2340, A[37], n_813);
  nand g2302 (n_832, n_2338, n_2339, n_2340);
  xor g2303 (n_2341, n_814, n_815);
  xor g2304 (n_821, n_2341, n_816);
  nand g2305 (n_2342, n_814, n_815);
  nand g2306 (n_2343, n_816, n_815);
  nand g2307 (n_2344, n_814, n_816);
  nand g2308 (n_834, n_2342, n_2343, n_2344);
  xor g2309 (n_2345, n_817, n_818);
  xor g2310 (n_823, n_2345, n_819);
  nand g2311 (n_2346, n_817, n_818);
  nand g2312 (n_2347, n_819, n_818);
  nand g2313 (n_2348, n_817, n_819);
  nand g2314 (n_836, n_2346, n_2347, n_2348);
  xor g2315 (n_2349, n_820, n_821);
  xor g2316 (n_824, n_2349, n_822);
  nand g2317 (n_2350, n_820, n_821);
  nand g2318 (n_2351, n_822, n_821);
  nand g2319 (n_2352, n_820, n_822);
  nand g2320 (n_839, n_2350, n_2351, n_2352);
  xor g2321 (n_2353, n_823, n_824);
  xor g2322 (n_175, n_2353, n_825);
  nand g2323 (n_2354, n_823, n_824);
  nand g2324 (n_2355, n_825, n_824);
  nand g2325 (n_2356, n_823, n_825);
  nand g2326 (n_93, n_2354, n_2355, n_2356);
  xor g2327 (n_2357, A[50], A[48]);
  xor g2328 (n_830, n_2357, A[44]);
  nand g2329 (n_2358, A[50], A[48]);
  nand g2330 (n_2359, A[44], A[48]);
  nand g2331 (n_2360, A[50], A[44]);
  nand g2332 (n_840, n_2358, n_2359, n_2360);
  xor g2334 (n_831, n_1909, A[42]);
  nand g2336 (n_2363, A[42], A[34]);
  nand g2338 (n_841, n_1910, n_2363, n_2104);
  xor g2339 (n_2365, A[32], A[46]);
  xor g2340 (n_829, n_2365, A[40]);
  nand g2341 (n_2366, A[32], A[46]);
  nand g2344 (n_842, n_2366, n_2232, n_2299);
  xor g2345 (n_2369, A[38], n_826);
  xor g2346 (n_833, n_2369, n_827);
  nand g2347 (n_2370, A[38], n_826);
  nand g2348 (n_2371, n_827, n_826);
  nand g2349 (n_2372, A[38], n_827);
  nand g2350 (n_846, n_2370, n_2371, n_2372);
  xor g2351 (n_2373, n_828, n_829);
  xor g2352 (n_835, n_2373, n_830);
  nand g2353 (n_2374, n_828, n_829);
  nand g2354 (n_2375, n_830, n_829);
  nand g2355 (n_2376, n_828, n_830);
  nand g2356 (n_848, n_2374, n_2375, n_2376);
  xor g2357 (n_2377, n_831, n_832);
  xor g2358 (n_837, n_2377, n_833);
  nand g2359 (n_2378, n_831, n_832);
  nand g2360 (n_2379, n_833, n_832);
  nand g2361 (n_2380, n_831, n_833);
  nand g2362 (n_850, n_2378, n_2379, n_2380);
  xor g2363 (n_2381, n_834, n_835);
  xor g2364 (n_838, n_2381, n_836);
  nand g2365 (n_2382, n_834, n_835);
  nand g2366 (n_2383, n_836, n_835);
  nand g2367 (n_2384, n_834, n_836);
  nand g2368 (n_853, n_2382, n_2383, n_2384);
  xor g2369 (n_2385, n_837, n_838);
  xor g2370 (n_174, n_2385, n_839);
  nand g2371 (n_2386, n_837, n_838);
  nand g2372 (n_2387, n_839, n_838);
  nand g2373 (n_2388, n_837, n_839);
  nand g2374 (n_92, n_2386, n_2387, n_2388);
  xor g2375 (n_2389, A[51], A[49]);
  xor g2376 (n_844, n_2389, A[45]);
  nand g2377 (n_2390, A[51], A[49]);
  nand g2378 (n_2391, A[45], A[49]);
  nand g2379 (n_2392, A[51], A[45]);
  nand g2380 (n_854, n_2390, n_2391, n_2392);
  xor g2382 (n_845, n_1941, A[43]);
  nand g2384 (n_2395, A[43], A[35]);
  nand g2386 (n_855, n_1942, n_2395, n_2136);
  xor g2387 (n_2397, A[33], A[47]);
  xor g2388 (n_843, n_2397, A[41]);
  nand g2389 (n_2398, A[33], A[47]);
  nand g2392 (n_856, n_2398, n_2264, n_2331);
  xor g2393 (n_2401, A[39], n_840);
  xor g2394 (n_847, n_2401, n_841);
  nand g2395 (n_2402, A[39], n_840);
  nand g2396 (n_2403, n_841, n_840);
  nand g2397 (n_2404, A[39], n_841);
  nand g2398 (n_860, n_2402, n_2403, n_2404);
  xor g2399 (n_2405, n_842, n_843);
  xor g2400 (n_849, n_2405, n_844);
  nand g2401 (n_2406, n_842, n_843);
  nand g2402 (n_2407, n_844, n_843);
  nand g2403 (n_2408, n_842, n_844);
  nand g2404 (n_862, n_2406, n_2407, n_2408);
  xor g2405 (n_2409, n_845, n_846);
  xor g2406 (n_851, n_2409, n_847);
  nand g2407 (n_2410, n_845, n_846);
  nand g2408 (n_2411, n_847, n_846);
  nand g2409 (n_2412, n_845, n_847);
  nand g2410 (n_864, n_2410, n_2411, n_2412);
  xor g2411 (n_2413, n_848, n_849);
  xor g2412 (n_852, n_2413, n_850);
  nand g2413 (n_2414, n_848, n_849);
  nand g2414 (n_2415, n_850, n_849);
  nand g2415 (n_2416, n_848, n_850);
  nand g2416 (n_867, n_2414, n_2415, n_2416);
  xor g2417 (n_2417, n_851, n_852);
  xor g2418 (n_173, n_2417, n_853);
  nand g2419 (n_2418, n_851, n_852);
  nand g2420 (n_2419, n_853, n_852);
  nand g2421 (n_2420, n_851, n_853);
  nand g2422 (n_91, n_2418, n_2419, n_2420);
  xor g2423 (n_2421, A[52], A[50]);
  xor g2424 (n_858, n_2421, A[46]);
  nand g2425 (n_2422, A[52], A[50]);
  nand g2426 (n_2423, A[46], A[50]);
  nand g2427 (n_2424, A[52], A[46]);
  nand g2428 (n_868, n_2422, n_2423, n_2424);
  xor g2430 (n_859, n_1973, A[44]);
  nand g2432 (n_2427, A[44], A[36]);
  nand g2434 (n_869, n_1974, n_2427, n_2168);
  xor g2435 (n_2429, A[34], A[48]);
  xor g2436 (n_857, n_2429, A[42]);
  nand g2437 (n_2430, A[34], A[48]);
  nand g2440 (n_870, n_2430, n_2296, n_2363);
  xor g2441 (n_2433, A[40], n_854);
  xor g2442 (n_861, n_2433, n_855);
  nand g2443 (n_2434, A[40], n_854);
  nand g2444 (n_2435, n_855, n_854);
  nand g2445 (n_2436, A[40], n_855);
  nand g2446 (n_874, n_2434, n_2435, n_2436);
  xor g2447 (n_2437, n_856, n_857);
  xor g2448 (n_863, n_2437, n_858);
  nand g2449 (n_2438, n_856, n_857);
  nand g2450 (n_2439, n_858, n_857);
  nand g2451 (n_2440, n_856, n_858);
  nand g2452 (n_876, n_2438, n_2439, n_2440);
  xor g2453 (n_2441, n_859, n_860);
  xor g2454 (n_865, n_2441, n_861);
  nand g2455 (n_2442, n_859, n_860);
  nand g2456 (n_2443, n_861, n_860);
  nand g2457 (n_2444, n_859, n_861);
  nand g2458 (n_878, n_2442, n_2443, n_2444);
  xor g2459 (n_2445, n_862, n_863);
  xor g2460 (n_866, n_2445, n_864);
  nand g2461 (n_2446, n_862, n_863);
  nand g2462 (n_2447, n_864, n_863);
  nand g2463 (n_2448, n_862, n_864);
  nand g2464 (n_881, n_2446, n_2447, n_2448);
  xor g2465 (n_2449, n_865, n_866);
  xor g2466 (n_172, n_2449, n_867);
  nand g2467 (n_2450, n_865, n_866);
  nand g2468 (n_2451, n_867, n_866);
  nand g2469 (n_2452, n_865, n_867);
  nand g2470 (n_90, n_2450, n_2451, n_2452);
  xor g2471 (n_2453, A[53], A[51]);
  xor g2472 (n_872, n_2453, A[47]);
  nand g2473 (n_2454, A[53], A[51]);
  nand g2474 (n_2455, A[47], A[51]);
  nand g2475 (n_2456, A[53], A[47]);
  nand g2476 (n_882, n_2454, n_2455, n_2456);
  xor g2478 (n_873, n_2005, A[45]);
  nand g2480 (n_2459, A[45], A[37]);
  nand g2482 (n_883, n_2006, n_2459, n_2200);
  xor g2483 (n_2461, A[35], A[49]);
  xor g2484 (n_871, n_2461, A[43]);
  nand g2485 (n_2462, A[35], A[49]);
  nand g2488 (n_884, n_2462, n_2328, n_2395);
  xor g2489 (n_2465, A[41], n_868);
  xor g2490 (n_875, n_2465, n_869);
  nand g2491 (n_2466, A[41], n_868);
  nand g2492 (n_2467, n_869, n_868);
  nand g2493 (n_2468, A[41], n_869);
  nand g2494 (n_888, n_2466, n_2467, n_2468);
  xor g2495 (n_2469, n_870, n_871);
  xor g2496 (n_877, n_2469, n_872);
  nand g2497 (n_2470, n_870, n_871);
  nand g2498 (n_2471, n_872, n_871);
  nand g2499 (n_2472, n_870, n_872);
  nand g2500 (n_890, n_2470, n_2471, n_2472);
  xor g2501 (n_2473, n_873, n_874);
  xor g2502 (n_879, n_2473, n_875);
  nand g2503 (n_2474, n_873, n_874);
  nand g2504 (n_2475, n_875, n_874);
  nand g2505 (n_2476, n_873, n_875);
  nand g2506 (n_892, n_2474, n_2475, n_2476);
  xor g2507 (n_2477, n_876, n_877);
  xor g2508 (n_880, n_2477, n_878);
  nand g2509 (n_2478, n_876, n_877);
  nand g2510 (n_2479, n_878, n_877);
  nand g2511 (n_2480, n_876, n_878);
  nand g2512 (n_895, n_2478, n_2479, n_2480);
  xor g2513 (n_2481, n_879, n_880);
  xor g2514 (n_171, n_2481, n_881);
  nand g2515 (n_2482, n_879, n_880);
  nand g2516 (n_2483, n_881, n_880);
  nand g2517 (n_2484, n_879, n_881);
  nand g2518 (n_89, n_2482, n_2483, n_2484);
  xor g2519 (n_2485, A[54], A[52]);
  xor g2520 (n_886, n_2485, A[48]);
  nand g2521 (n_2486, A[54], A[52]);
  nand g2522 (n_2487, A[48], A[52]);
  nand g2523 (n_2488, A[54], A[48]);
  nand g2524 (n_896, n_2486, n_2487, n_2488);
  xor g2526 (n_887, n_2037, A[46]);
  nand g2528 (n_2491, A[46], A[38]);
  nand g2530 (n_897, n_2038, n_2491, n_2232);
  xor g2531 (n_2493, A[36], A[50]);
  xor g2532 (n_885, n_2493, A[44]);
  nand g2533 (n_2494, A[36], A[50]);
  nand g2536 (n_898, n_2494, n_2360, n_2427);
  xor g2537 (n_2497, A[42], n_882);
  xor g2538 (n_889, n_2497, n_883);
  nand g2539 (n_2498, A[42], n_882);
  nand g2540 (n_2499, n_883, n_882);
  nand g2541 (n_2500, A[42], n_883);
  nand g2542 (n_902, n_2498, n_2499, n_2500);
  xor g2543 (n_2501, n_884, n_885);
  xor g2544 (n_891, n_2501, n_886);
  nand g2545 (n_2502, n_884, n_885);
  nand g2546 (n_2503, n_886, n_885);
  nand g2547 (n_2504, n_884, n_886);
  nand g2548 (n_904, n_2502, n_2503, n_2504);
  xor g2549 (n_2505, n_887, n_888);
  xor g2550 (n_893, n_2505, n_889);
  nand g2551 (n_2506, n_887, n_888);
  nand g2552 (n_2507, n_889, n_888);
  nand g2553 (n_2508, n_887, n_889);
  nand g2554 (n_906, n_2506, n_2507, n_2508);
  xor g2555 (n_2509, n_890, n_891);
  xor g2556 (n_894, n_2509, n_892);
  nand g2557 (n_2510, n_890, n_891);
  nand g2558 (n_2511, n_892, n_891);
  nand g2559 (n_2512, n_890, n_892);
  nand g2560 (n_909, n_2510, n_2511, n_2512);
  xor g2561 (n_2513, n_893, n_894);
  xor g2562 (n_170, n_2513, n_895);
  nand g2563 (n_2514, n_893, n_894);
  nand g2564 (n_2515, n_895, n_894);
  nand g2565 (n_2516, n_893, n_895);
  nand g2566 (n_88, n_2514, n_2515, n_2516);
  xor g2567 (n_2517, A[55], A[53]);
  xor g2568 (n_900, n_2517, A[49]);
  nand g2569 (n_2518, A[55], A[53]);
  nand g2570 (n_2519, A[49], A[53]);
  nand g2571 (n_2520, A[55], A[49]);
  nand g2572 (n_910, n_2518, n_2519, n_2520);
  xor g2574 (n_901, n_2069, A[47]);
  nand g2576 (n_2523, A[47], A[39]);
  nand g2578 (n_911, n_2070, n_2523, n_2264);
  xor g2579 (n_2525, A[37], A[51]);
  xor g2580 (n_899, n_2525, A[45]);
  nand g2581 (n_2526, A[37], A[51]);
  nand g2584 (n_912, n_2526, n_2392, n_2459);
  xor g2585 (n_2529, A[43], n_896);
  xor g2586 (n_903, n_2529, n_897);
  nand g2587 (n_2530, A[43], n_896);
  nand g2588 (n_2531, n_897, n_896);
  nand g2589 (n_2532, A[43], n_897);
  nand g2590 (n_916, n_2530, n_2531, n_2532);
  xor g2591 (n_2533, n_898, n_899);
  xor g2592 (n_905, n_2533, n_900);
  nand g2593 (n_2534, n_898, n_899);
  nand g2594 (n_2535, n_900, n_899);
  nand g2595 (n_2536, n_898, n_900);
  nand g2596 (n_918, n_2534, n_2535, n_2536);
  xor g2597 (n_2537, n_901, n_902);
  xor g2598 (n_907, n_2537, n_903);
  nand g2599 (n_2538, n_901, n_902);
  nand g2600 (n_2539, n_903, n_902);
  nand g2601 (n_2540, n_901, n_903);
  nand g2602 (n_920, n_2538, n_2539, n_2540);
  xor g2603 (n_2541, n_904, n_905);
  xor g2604 (n_908, n_2541, n_906);
  nand g2605 (n_2542, n_904, n_905);
  nand g2606 (n_2543, n_906, n_905);
  nand g2607 (n_2544, n_904, n_906);
  nand g2608 (n_923, n_2542, n_2543, n_2544);
  xor g2609 (n_2545, n_907, n_908);
  xor g2610 (n_169, n_2545, n_909);
  nand g2611 (n_2546, n_907, n_908);
  nand g2612 (n_2547, n_909, n_908);
  nand g2613 (n_2548, n_907, n_909);
  nand g2614 (n_87, n_2546, n_2547, n_2548);
  xor g2615 (n_2549, A[56], A[54]);
  xor g2616 (n_914, n_2549, A[50]);
  nand g2617 (n_2550, A[56], A[54]);
  nand g2618 (n_2551, A[50], A[54]);
  nand g2619 (n_2552, A[56], A[50]);
  nand g2620 (n_924, n_2550, n_2551, n_2552);
  xor g2622 (n_915, n_2101, A[48]);
  nand g2624 (n_2555, A[48], A[40]);
  nand g2626 (n_925, n_2102, n_2555, n_2296);
  xor g2627 (n_2557, A[38], A[52]);
  xor g2628 (n_913, n_2557, A[46]);
  nand g2629 (n_2558, A[38], A[52]);
  nand g2632 (n_926, n_2558, n_2424, n_2491);
  xor g2633 (n_2561, A[44], n_910);
  xor g2634 (n_917, n_2561, n_911);
  nand g2635 (n_2562, A[44], n_910);
  nand g2636 (n_2563, n_911, n_910);
  nand g2637 (n_2564, A[44], n_911);
  nand g2638 (n_930, n_2562, n_2563, n_2564);
  xor g2639 (n_2565, n_912, n_913);
  xor g2640 (n_919, n_2565, n_914);
  nand g2641 (n_2566, n_912, n_913);
  nand g2642 (n_2567, n_914, n_913);
  nand g2643 (n_2568, n_912, n_914);
  nand g2644 (n_932, n_2566, n_2567, n_2568);
  xor g2645 (n_2569, n_915, n_916);
  xor g2646 (n_921, n_2569, n_917);
  nand g2647 (n_2570, n_915, n_916);
  nand g2648 (n_2571, n_917, n_916);
  nand g2649 (n_2572, n_915, n_917);
  nand g2650 (n_934, n_2570, n_2571, n_2572);
  xor g2651 (n_2573, n_918, n_919);
  xor g2652 (n_922, n_2573, n_920);
  nand g2653 (n_2574, n_918, n_919);
  nand g2654 (n_2575, n_920, n_919);
  nand g2655 (n_2576, n_918, n_920);
  nand g2656 (n_937, n_2574, n_2575, n_2576);
  xor g2657 (n_2577, n_921, n_922);
  xor g2658 (n_168, n_2577, n_923);
  nand g2659 (n_2578, n_921, n_922);
  nand g2660 (n_2579, n_923, n_922);
  nand g2661 (n_2580, n_921, n_923);
  nand g2662 (n_86, n_2578, n_2579, n_2580);
  xor g2663 (n_2581, A[57], A[55]);
  xor g2664 (n_928, n_2581, A[51]);
  nand g2665 (n_2582, A[57], A[55]);
  nand g2666 (n_2583, A[51], A[55]);
  nand g2667 (n_2584, A[57], A[51]);
  nand g2668 (n_938, n_2582, n_2583, n_2584);
  xor g2670 (n_929, n_2133, A[49]);
  nand g2672 (n_2587, A[49], A[41]);
  nand g2674 (n_939, n_2134, n_2587, n_2328);
  xor g2675 (n_2589, A[39], A[53]);
  xor g2676 (n_927, n_2589, A[47]);
  nand g2677 (n_2590, A[39], A[53]);
  nand g2680 (n_940, n_2590, n_2456, n_2523);
  xor g2681 (n_2593, A[45], n_924);
  xor g2682 (n_931, n_2593, n_925);
  nand g2683 (n_2594, A[45], n_924);
  nand g2684 (n_2595, n_925, n_924);
  nand g2685 (n_2596, A[45], n_925);
  nand g2686 (n_944, n_2594, n_2595, n_2596);
  xor g2687 (n_2597, n_926, n_927);
  xor g2688 (n_933, n_2597, n_928);
  nand g2689 (n_2598, n_926, n_927);
  nand g2690 (n_2599, n_928, n_927);
  nand g2691 (n_2600, n_926, n_928);
  nand g2692 (n_946, n_2598, n_2599, n_2600);
  xor g2693 (n_2601, n_929, n_930);
  xor g2694 (n_935, n_2601, n_931);
  nand g2695 (n_2602, n_929, n_930);
  nand g2696 (n_2603, n_931, n_930);
  nand g2697 (n_2604, n_929, n_931);
  nand g2698 (n_948, n_2602, n_2603, n_2604);
  xor g2699 (n_2605, n_932, n_933);
  xor g2700 (n_936, n_2605, n_934);
  nand g2701 (n_2606, n_932, n_933);
  nand g2702 (n_2607, n_934, n_933);
  nand g2703 (n_2608, n_932, n_934);
  nand g2704 (n_951, n_2606, n_2607, n_2608);
  xor g2705 (n_2609, n_935, n_936);
  xor g2706 (n_167, n_2609, n_937);
  nand g2707 (n_2610, n_935, n_936);
  nand g2708 (n_2611, n_937, n_936);
  nand g2709 (n_2612, n_935, n_937);
  nand g2710 (n_85, n_2610, n_2611, n_2612);
  xor g2711 (n_2613, A[58], A[56]);
  xor g2712 (n_942, n_2613, A[52]);
  nand g2713 (n_2614, A[58], A[56]);
  nand g2714 (n_2615, A[52], A[56]);
  nand g2715 (n_2616, A[58], A[52]);
  nand g2716 (n_952, n_2614, n_2615, n_2616);
  xor g2718 (n_943, n_2165, A[50]);
  nand g2720 (n_2619, A[50], A[42]);
  nand g2722 (n_953, n_2166, n_2619, n_2360);
  xor g2723 (n_2621, A[40], A[54]);
  xor g2724 (n_941, n_2621, A[48]);
  nand g2725 (n_2622, A[40], A[54]);
  nand g2728 (n_954, n_2622, n_2488, n_2555);
  xor g2729 (n_2625, A[46], n_938);
  xor g2730 (n_945, n_2625, n_939);
  nand g2731 (n_2626, A[46], n_938);
  nand g2732 (n_2627, n_939, n_938);
  nand g2733 (n_2628, A[46], n_939);
  nand g2734 (n_958, n_2626, n_2627, n_2628);
  xor g2735 (n_2629, n_940, n_941);
  xor g2736 (n_947, n_2629, n_942);
  nand g2737 (n_2630, n_940, n_941);
  nand g2738 (n_2631, n_942, n_941);
  nand g2739 (n_2632, n_940, n_942);
  nand g2740 (n_960, n_2630, n_2631, n_2632);
  xor g2741 (n_2633, n_943, n_944);
  xor g2742 (n_949, n_2633, n_945);
  nand g2743 (n_2634, n_943, n_944);
  nand g2744 (n_2635, n_945, n_944);
  nand g2745 (n_2636, n_943, n_945);
  nand g2746 (n_962, n_2634, n_2635, n_2636);
  xor g2747 (n_2637, n_946, n_947);
  xor g2748 (n_950, n_2637, n_948);
  nand g2749 (n_2638, n_946, n_947);
  nand g2750 (n_2639, n_948, n_947);
  nand g2751 (n_2640, n_946, n_948);
  nand g2752 (n_965, n_2638, n_2639, n_2640);
  xor g2753 (n_2641, n_949, n_950);
  xor g2754 (n_166, n_2641, n_951);
  nand g2755 (n_2642, n_949, n_950);
  nand g2756 (n_2643, n_951, n_950);
  nand g2757 (n_2644, n_949, n_951);
  nand g2758 (n_84, n_2642, n_2643, n_2644);
  xor g2759 (n_2645, A[59], A[57]);
  xor g2760 (n_956, n_2645, A[53]);
  nand g2761 (n_2646, A[59], A[57]);
  nand g2762 (n_2647, A[53], A[57]);
  nand g2763 (n_2648, A[59], A[53]);
  nand g2764 (n_966, n_2646, n_2647, n_2648);
  xor g2766 (n_957, n_2197, A[51]);
  nand g2768 (n_2651, A[51], A[43]);
  nand g2770 (n_967, n_2198, n_2651, n_2392);
  xor g2771 (n_2653, A[41], A[55]);
  xor g2772 (n_955, n_2653, A[49]);
  nand g2773 (n_2654, A[41], A[55]);
  nand g2776 (n_968, n_2654, n_2520, n_2587);
  xor g2777 (n_2657, A[47], n_952);
  xor g2778 (n_959, n_2657, n_953);
  nand g2779 (n_2658, A[47], n_952);
  nand g2780 (n_2659, n_953, n_952);
  nand g2781 (n_2660, A[47], n_953);
  nand g2782 (n_972, n_2658, n_2659, n_2660);
  xor g2783 (n_2661, n_954, n_955);
  xor g2784 (n_961, n_2661, n_956);
  nand g2785 (n_2662, n_954, n_955);
  nand g2786 (n_2663, n_956, n_955);
  nand g2787 (n_2664, n_954, n_956);
  nand g2788 (n_974, n_2662, n_2663, n_2664);
  xor g2789 (n_2665, n_957, n_958);
  xor g2790 (n_963, n_2665, n_959);
  nand g2791 (n_2666, n_957, n_958);
  nand g2792 (n_2667, n_959, n_958);
  nand g2793 (n_2668, n_957, n_959);
  nand g2794 (n_976, n_2666, n_2667, n_2668);
  xor g2795 (n_2669, n_960, n_961);
  xor g2796 (n_964, n_2669, n_962);
  nand g2797 (n_2670, n_960, n_961);
  nand g2798 (n_2671, n_962, n_961);
  nand g2799 (n_2672, n_960, n_962);
  nand g2800 (n_979, n_2670, n_2671, n_2672);
  xor g2801 (n_2673, n_963, n_964);
  xor g2802 (n_165, n_2673, n_965);
  nand g2803 (n_2674, n_963, n_964);
  nand g2804 (n_2675, n_965, n_964);
  nand g2805 (n_2676, n_963, n_965);
  nand g2806 (n_83, n_2674, n_2675, n_2676);
  xor g2807 (n_2677, A[60], A[58]);
  xor g2808 (n_970, n_2677, A[54]);
  nand g2809 (n_2678, A[60], A[58]);
  nand g2810 (n_2679, A[54], A[58]);
  nand g2811 (n_2680, A[60], A[54]);
  nand g2812 (n_983, n_2678, n_2679, n_2680);
  xor g2814 (n_971, n_2229, A[52]);
  nand g2816 (n_2683, A[52], A[44]);
  nand g2818 (n_984, n_2230, n_2683, n_2424);
  xor g2819 (n_2685, A[42], A[56]);
  xor g2820 (n_969, n_2685, A[50]);
  nand g2821 (n_2686, A[42], A[56]);
  nand g2824 (n_982, n_2686, n_2552, n_2619);
  xor g2825 (n_2689, A[48], n_966);
  xor g2826 (n_973, n_2689, n_967);
  nand g2827 (n_2690, A[48], n_966);
  nand g2828 (n_2691, n_967, n_966);
  nand g2829 (n_2692, A[48], n_967);
  nand g2830 (n_988, n_2690, n_2691, n_2692);
  xor g2831 (n_2693, n_968, n_969);
  xor g2832 (n_975, n_2693, n_970);
  nand g2833 (n_2694, n_968, n_969);
  nand g2834 (n_2695, n_970, n_969);
  nand g2835 (n_2696, n_968, n_970);
  nand g2836 (n_990, n_2694, n_2695, n_2696);
  xor g2837 (n_2697, n_971, n_972);
  xor g2838 (n_977, n_2697, n_973);
  nand g2839 (n_2698, n_971, n_972);
  nand g2840 (n_2699, n_973, n_972);
  nand g2841 (n_2700, n_971, n_973);
  nand g2842 (n_992, n_2698, n_2699, n_2700);
  xor g2843 (n_2701, n_974, n_975);
  xor g2844 (n_978, n_2701, n_976);
  nand g2845 (n_2702, n_974, n_975);
  nand g2846 (n_2703, n_976, n_975);
  nand g2847 (n_2704, n_974, n_976);
  nand g2848 (n_995, n_2702, n_2703, n_2704);
  xor g2849 (n_2705, n_977, n_978);
  xor g2850 (n_164, n_2705, n_979);
  nand g2851 (n_2706, n_977, n_978);
  nand g2852 (n_2707, n_979, n_978);
  nand g2853 (n_2708, n_977, n_979);
  nand g2854 (n_82, n_2706, n_2707, n_2708);
  xor g2857 (n_2709, A[61], A[55]);
  xor g2858 (n_986, n_2709, A[47]);
  nand g2859 (n_2710, A[61], A[55]);
  nand g2860 (n_2711, A[47], A[55]);
  nand g2861 (n_2712, A[61], A[47]);
  nand g2862 (n_1000, n_2710, n_2711, n_2712);
  xor g2863 (n_2713, A[45], A[59]);
  xor g2864 (n_987, n_2713, A[43]);
  nand g2865 (n_2714, A[45], A[59]);
  nand g2866 (n_2715, A[43], A[59]);
  nand g2868 (n_1001, n_2714, n_2715, n_2198);
  xor g2869 (n_2717, A[53], A[57]);
  xor g2870 (n_985, n_2717, A[51]);
  nand g2874 (n_999, n_2647, n_2584, n_2454);
  xor g2875 (n_2721, A[49], n_982);
  xor g2876 (n_989, n_2721, n_983);
  nand g2877 (n_2722, A[49], n_982);
  nand g2878 (n_2723, n_983, n_982);
  nand g2879 (n_2724, A[49], n_983);
  nand g2880 (n_1005, n_2722, n_2723, n_2724);
  xor g2881 (n_2725, n_984, n_985);
  xor g2882 (n_991, n_2725, n_986);
  nand g2883 (n_2726, n_984, n_985);
  nand g2884 (n_2727, n_986, n_985);
  nand g2885 (n_2728, n_984, n_986);
  nand g2886 (n_1007, n_2726, n_2727, n_2728);
  xor g2887 (n_2729, n_987, n_988);
  xor g2888 (n_993, n_2729, n_989);
  nand g2889 (n_2730, n_987, n_988);
  nand g2890 (n_2731, n_989, n_988);
  nand g2891 (n_2732, n_987, n_989);
  nand g2892 (n_1009, n_2730, n_2731, n_2732);
  xor g2893 (n_2733, n_990, n_991);
  xor g2894 (n_994, n_2733, n_992);
  nand g2895 (n_2734, n_990, n_991);
  nand g2896 (n_2735, n_992, n_991);
  nand g2897 (n_2736, n_990, n_992);
  nand g2898 (n_1012, n_2734, n_2735, n_2736);
  xor g2899 (n_2737, n_993, n_994);
  xor g2900 (n_163, n_2737, n_995);
  nand g2901 (n_2738, n_993, n_994);
  nand g2902 (n_2739, n_995, n_994);
  nand g2903 (n_2740, n_993, n_995);
  nand g2904 (n_81, n_2738, n_2739, n_2740);
  xor g2907 (n_2741, A[54], A[46]);
  xor g2908 (n_1003, n_2741, A[44]);
  nand g2909 (n_2742, A[54], A[46]);
  nand g2911 (n_2744, A[54], A[44]);
  nand g2912 (n_1014, n_2742, n_2230, n_2744);
  xor g2913 (n_2745, A[61], A[60]);
  xor g2914 (n_1004, n_2745, A[52]);
  nand g2915 (n_2746, A[61], A[60]);
  nand g2916 (n_2747, A[52], A[60]);
  nand g2917 (n_2748, A[61], A[52]);
  nand g2918 (n_1015, n_2746, n_2747, n_2748);
  xor g2920 (n_1002, n_2613, A[50]);
  nand g2923 (n_2752, A[58], A[50]);
  nand g2924 (n_1016, n_2614, n_2552, n_2752);
  xor g2925 (n_2753, A[48], n_999);
  xor g2926 (n_1006, n_2753, n_1000);
  nand g2927 (n_2754, A[48], n_999);
  nand g2928 (n_2755, n_1000, n_999);
  nand g2929 (n_2756, A[48], n_1000);
  nand g2930 (n_1020, n_2754, n_2755, n_2756);
  xor g2931 (n_2757, n_1001, n_1002);
  xor g2932 (n_1008, n_2757, n_1003);
  nand g2933 (n_2758, n_1001, n_1002);
  nand g2934 (n_2759, n_1003, n_1002);
  nand g2935 (n_2760, n_1001, n_1003);
  nand g2936 (n_1022, n_2758, n_2759, n_2760);
  xor g2937 (n_2761, n_1004, n_1005);
  xor g2938 (n_1010, n_2761, n_1006);
  nand g2939 (n_2762, n_1004, n_1005);
  nand g2940 (n_2763, n_1006, n_1005);
  nand g2941 (n_2764, n_1004, n_1006);
  nand g2942 (n_1024, n_2762, n_2763, n_2764);
  xor g2943 (n_2765, n_1007, n_1008);
  xor g2944 (n_1011, n_2765, n_1009);
  nand g2945 (n_2766, n_1007, n_1008);
  nand g2946 (n_2767, n_1009, n_1008);
  nand g2947 (n_2768, n_1007, n_1009);
  nand g2948 (n_1027, n_2766, n_2767, n_2768);
  xor g2949 (n_2769, n_1010, n_1011);
  xor g2950 (n_162, n_2769, n_1012);
  nand g2951 (n_2770, n_1010, n_1011);
  nand g2952 (n_2771, n_1012, n_1011);
  nand g2953 (n_2772, n_1010, n_1012);
  nand g2954 (n_80, n_2770, n_2771, n_2772);
  xor g2956 (n_1018, n_2773, A[55]);
  nand g2958 (n_2775, A[55], A[59]);
  nand g2960 (n_1030, n_2774, n_2775, n_2776);
  xor g2962 (n_1019, n_2261, A[53]);
  nand g2964 (n_2779, A[53], A[45]);
  nand g2966 (n_1031, n_2262, n_2779, n_2456);
  xor g2968 (n_1017, n_2781, A[51]);
  nand g2972 (n_1032, n_2782, n_2584, n_2784);
  xor g2973 (n_2785, A[49], n_1014);
  xor g2974 (n_1021, n_2785, n_1015);
  nand g2975 (n_2786, A[49], n_1014);
  nand g2976 (n_2787, n_1015, n_1014);
  nand g2977 (n_2788, A[49], n_1015);
  nand g2978 (n_1036, n_2786, n_2787, n_2788);
  xor g2979 (n_2789, n_1016, n_1017);
  xor g2980 (n_1023, n_2789, n_1018);
  nand g2981 (n_2790, n_1016, n_1017);
  nand g2982 (n_2791, n_1018, n_1017);
  nand g2983 (n_2792, n_1016, n_1018);
  nand g2984 (n_1038, n_2790, n_2791, n_2792);
  xor g2985 (n_2793, n_1019, n_1020);
  xor g2986 (n_1025, n_2793, n_1021);
  nand g2987 (n_2794, n_1019, n_1020);
  nand g2988 (n_2795, n_1021, n_1020);
  nand g2989 (n_2796, n_1019, n_1021);
  nand g2990 (n_1040, n_2794, n_2795, n_2796);
  xor g2991 (n_2797, n_1022, n_1023);
  xor g2992 (n_1026, n_2797, n_1024);
  nand g2993 (n_2798, n_1022, n_1023);
  nand g2994 (n_2799, n_1024, n_1023);
  nand g2995 (n_2800, n_1022, n_1024);
  nand g2996 (n_1042, n_2798, n_2799, n_2800);
  xor g2997 (n_2801, n_1025, n_1026);
  xor g2998 (n_161, n_2801, n_1027);
  nand g2999 (n_2802, n_1025, n_1026);
  nand g3000 (n_2803, n_1027, n_1026);
  nand g3001 (n_2804, n_1025, n_1027);
  nand g3002 (n_79, n_2802, n_2803, n_2804);
  xor g3005 (n_2805, A[58], A[46]);
  xor g3006 (n_1034, n_2805, A[54]);
  nand g3007 (n_2806, A[58], A[46]);
  nand g3010 (n_1045, n_2806, n_2742, n_2679);
  xor g3011 (n_2809, A[52], A[56]);
  xor g3012 (n_1033, n_2809, A[50]);
  nand g3016 (n_1044, n_2615, n_2552, n_2422);
  xor g3018 (n_1035, n_2813, n_1030);
  nand g3021 (n_2816, A[48], n_1030);
  nand g3022 (n_1049, n_2814, n_2815, n_2816);
  xor g3023 (n_2817, n_1031, n_1032);
  xor g3024 (n_1037, n_2817, n_1033);
  nand g3025 (n_2818, n_1031, n_1032);
  nand g3026 (n_2819, n_1033, n_1032);
  nand g3027 (n_2820, n_1031, n_1033);
  nand g3028 (n_1051, n_2818, n_2819, n_2820);
  xor g3029 (n_2821, n_1034, n_1035);
  xor g3030 (n_1039, n_2821, n_1036);
  nand g3031 (n_2822, n_1034, n_1035);
  nand g3032 (n_2823, n_1036, n_1035);
  nand g3033 (n_2824, n_1034, n_1036);
  nand g3034 (n_1052, n_2822, n_2823, n_2824);
  xor g3035 (n_2825, n_1037, n_1038);
  xor g3036 (n_1041, n_2825, n_1039);
  nand g3037 (n_2826, n_1037, n_1038);
  nand g3038 (n_2827, n_1039, n_1038);
  nand g3039 (n_2828, n_1037, n_1039);
  nand g3040 (n_1055, n_2826, n_2827, n_2828);
  xor g3041 (n_2829, n_1040, n_1041);
  xor g3042 (n_160, n_2829, n_1042);
  nand g3043 (n_2830, n_1040, n_1041);
  nand g3044 (n_2831, n_1042, n_1041);
  nand g3045 (n_2832, n_1040, n_1042);
  nand g3046 (n_78, n_2830, n_2831, n_2832);
  xor g3053 (n_2837, A[47], A[53]);
  xor g3054 (n_1047, n_2837, A[57]);
  nand g3057 (n_2840, A[47], A[57]);
  nand g3058 (n_1059, n_2456, n_2647, n_2840);
  xor g3060 (n_1048, n_2389, A[60]);
  nand g3062 (n_2843, A[60], A[49]);
  nand g3063 (n_2844, A[51], A[60]);
  nand g3064 (n_1062, n_2390, n_2843, n_2844);
  xor g3065 (n_2845, n_1044, n_1045);
  xor g3066 (n_1050, n_2845, n_1018);
  nand g3067 (n_2846, n_1044, n_1045);
  nand g3068 (n_2847, n_1018, n_1045);
  nand g3069 (n_2848, n_1044, n_1018);
  nand g3070 (n_1064, n_2846, n_2847, n_2848);
  xor g3071 (n_2849, n_1047, n_1048);
  xor g3072 (n_1053, n_2849, n_1049);
  nand g3073 (n_2850, n_1047, n_1048);
  nand g3074 (n_2851, n_1049, n_1048);
  nand g3075 (n_2852, n_1047, n_1049);
  nand g3076 (n_1066, n_2850, n_2851, n_2852);
  xor g3077 (n_2853, n_1050, n_1051);
  xor g3078 (n_1054, n_2853, n_1052);
  nand g3079 (n_2854, n_1050, n_1051);
  nand g3080 (n_2855, n_1052, n_1051);
  nand g3081 (n_2856, n_1050, n_1052);
  nand g3082 (n_1068, n_2854, n_2855, n_2856);
  xor g3083 (n_2857, n_1053, n_1054);
  xor g3084 (n_159, n_2857, n_1055);
  nand g3085 (n_2858, n_1053, n_1054);
  nand g3086 (n_2859, n_1055, n_1054);
  nand g3087 (n_2860, n_1053, n_1055);
  nand g3088 (n_158, n_2858, n_2859, n_2860);
  xor g3091 (n_2861, A[58], A[54]);
  xor g3092 (n_1061, n_2861, A[52]);
  nand g3096 (n_1070, n_2679, n_2486, n_2616);
  xor g3097 (n_2865, A[56], A[50]);
  xor g3098 (n_1060, n_2865, A[48]);
  nand g3101 (n_2868, A[56], A[48]);
  nand g3102 (n_1071, n_2552, n_2358, n_2868);
  xor g3104 (n_1063, n_2869, n_1059);
  nand g3106 (n_2871, n_1059, n_1030);
  nand g3108 (n_1075, n_2815, n_2871, n_2872);
  xor g3109 (n_2873, n_1060, n_1061);
  xor g3110 (n_1065, n_2873, n_1062);
  nand g3111 (n_2874, n_1060, n_1061);
  nand g3112 (n_2875, n_1062, n_1061);
  nand g3113 (n_2876, n_1060, n_1062);
  nand g3114 (n_1076, n_2874, n_2875, n_2876);
  xor g3115 (n_2877, n_1063, n_1064);
  xor g3116 (n_1067, n_2877, n_1065);
  nand g3117 (n_2878, n_1063, n_1064);
  nand g3118 (n_2879, n_1065, n_1064);
  nand g3119 (n_2880, n_1063, n_1065);
  nand g3120 (n_1079, n_2878, n_2879, n_2880);
  xor g3121 (n_2881, n_1066, n_1067);
  xor g3122 (n_77, n_2881, n_1068);
  nand g3123 (n_2882, n_1066, n_1067);
  nand g3124 (n_2883, n_1068, n_1067);
  nand g3125 (n_2884, n_1066, n_1068);
  nand g3126 (n_76, n_2882, n_2883, n_2884);
  xor g3139 (n_2893, A[49], A[60]);
  xor g3140 (n_1074, n_2893, n_1070);
  nand g3142 (n_2895, n_1070, A[60]);
  nand g3143 (n_2896, A[49], n_1070);
  nand g3144 (n_1086, n_2843, n_2895, n_2896);
  xor g3145 (n_2897, n_1071, n_985);
  xor g3146 (n_1077, n_2897, n_1018);
  nand g3147 (n_2898, n_1071, n_985);
  nand g3148 (n_2899, n_1018, n_985);
  nand g3149 (n_2900, n_1071, n_1018);
  nand g3150 (n_1087, n_2898, n_2899, n_2900);
  xor g3151 (n_2901, n_1074, n_1075);
  xor g3152 (n_1078, n_2901, n_1076);
  nand g3153 (n_2902, n_1074, n_1075);
  nand g3154 (n_2903, n_1076, n_1075);
  nand g3155 (n_2904, n_1074, n_1076);
  nand g3156 (n_1090, n_2902, n_2903, n_2904);
  xor g3157 (n_2905, n_1077, n_1078);
  xor g3158 (n_157, n_2905, n_1079);
  nand g3159 (n_2906, n_1077, n_1078);
  nand g3160 (n_2907, n_1079, n_1078);
  nand g3161 (n_2908, n_1077, n_1079);
  nand g3162 (n_75, n_2906, n_2907, n_2908);
  xor g3166 (n_1084, n_2485, A[60]);
  nand g3170 (n_1092, n_2486, n_2747, n_2680);
  nand g3176 (n_1095, n_2552, n_2915, n_2916);
  xor g3177 (n_2917, n_999, n_1030);
  xor g3178 (n_1088, n_2917, n_1084);
  nand g3179 (n_2918, n_999, n_1030);
  nand g3180 (n_2919, n_1084, n_1030);
  nand g3181 (n_2920, n_999, n_1084);
  nand g3182 (n_1097, n_2918, n_2919, n_2920);
  xor g3183 (n_2921, n_1085, n_1086);
  xor g3184 (n_1089, n_2921, n_1087);
  nand g3185 (n_2922, n_1085, n_1086);
  nand g3186 (n_2923, n_1087, n_1086);
  nand g3187 (n_2924, n_1085, n_1087);
  nand g3188 (n_1099, n_2922, n_2923, n_2924);
  xor g3189 (n_2925, n_1088, n_1089);
  xor g3190 (n_156, n_2925, n_1090);
  nand g3191 (n_2926, n_1088, n_1089);
  nand g3192 (n_2927, n_1090, n_1089);
  nand g3193 (n_2928, n_1088, n_1090);
  nand g3194 (n_74, n_2926, n_2927, n_2928);
  xor g3207 (n_2937, A[58], n_1092);
  xor g3208 (n_1096, n_2937, n_985);
  nand g3209 (n_2938, A[58], n_1092);
  nand g3210 (n_2939, n_985, n_1092);
  nand g3211 (n_2940, A[58], n_985);
  nand g3212 (n_1106, n_2938, n_2939, n_2940);
  xor g3213 (n_2941, n_1018, n_1095);
  xor g3214 (n_1098, n_2941, n_1096);
  nand g3215 (n_2942, n_1018, n_1095);
  nand g3216 (n_2943, n_1096, n_1095);
  nand g3217 (n_2944, n_1018, n_1096);
  nand g3218 (n_1108, n_2942, n_2943, n_2944);
  xor g3219 (n_2945, n_1097, n_1098);
  xor g3220 (n_155, n_2945, n_1099);
  nand g3221 (n_2946, n_1097, n_1098);
  nand g3222 (n_2947, n_1099, n_1098);
  nand g3223 (n_2948, n_1097, n_1099);
  nand g3224 (n_73, n_2946, n_2947, n_2948);
  nand g3237 (n_2956, A[56], n_999);
  nand g3238 (n_1113, n_2915, n_2955, n_2956);
  xor g3239 (n_2957, n_1030, n_1084);
  xor g3240 (n_1107, n_2957, n_1105);
  nand g3242 (n_2959, n_1105, n_1084);
  nand g3243 (n_2960, n_1030, n_1105);
  nand g3244 (n_1115, n_2919, n_2959, n_2960);
  xor g3245 (n_2961, n_1106, n_1107);
  xor g3246 (n_154, n_2961, n_1108);
  nand g3247 (n_2962, n_1106, n_1107);
  nand g3248 (n_2963, n_1108, n_1107);
  nand g3249 (n_2964, n_1106, n_1108);
  nand g3250 (n_153, n_2962, n_2963, n_2964);
  xor g3258 (n_1112, n_2717, A[58]);
  nand g3260 (n_2971, A[58], A[57]);
  nand g3261 (n_2972, A[53], A[58]);
  nand g3262 (n_1120, n_2647, n_2971, n_2972);
  xor g3263 (n_2973, n_1092, n_1018);
  xor g3264 (n_1114, n_2973, n_1112);
  nand g3265 (n_2974, n_1092, n_1018);
  nand g3266 (n_2975, n_1112, n_1018);
  nand g3267 (n_2976, n_1092, n_1112);
  nand g3268 (n_1122, n_2974, n_2975, n_2976);
  xor g3269 (n_2977, n_1113, n_1114);
  xor g3270 (n_72, n_2977, n_1115);
  nand g3271 (n_2978, n_1113, n_1114);
  nand g3272 (n_2979, n_1115, n_1114);
  nand g3273 (n_2980, n_1113, n_1115);
  nand g3274 (n_152, n_2978, n_2979, n_2980);
  xor g3278 (n_1119, n_2861, A[56]);
  nand g3282 (n_1124, n_2679, n_2614, n_2550);
  xor g3284 (n_1121, n_2869, n_1119);
  nand g3286 (n_2987, n_1119, n_1030);
  nand g3288 (n_1127, n_2815, n_2987, n_2988);
  xor g3289 (n_2989, n_1120, n_1121);
  xor g3290 (n_71, n_2989, n_1122);
  nand g3291 (n_2990, n_1120, n_1121);
  nand g3292 (n_2991, n_1122, n_1121);
  nand g3293 (n_2992, n_1120, n_1122);
  nand g3294 (n_151, n_2990, n_2991, n_2992);
  xor g3301 (n_2997, A[57], A[60]);
  xor g3302 (n_1126, n_2997, n_1124);
  nand g3303 (n_2998, A[57], A[60]);
  nand g3304 (n_2999, n_1124, A[60]);
  nand g3305 (n_3000, A[57], n_1124);
  nand g3306 (n_1132, n_2998, n_2999, n_3000);
  xor g3307 (n_3001, n_1018, n_1126);
  xor g3308 (n_70, n_3001, n_1127);
  nand g3309 (n_3002, n_1018, n_1126);
  nand g3310 (n_3003, n_1127, n_1126);
  nand g3311 (n_3004, n_1018, n_1127);
  nand g3312 (n_150, n_3002, n_3003, n_3004);
  nand g3320 (n_1135, n_2614, n_3007, n_3008);
  xor g3321 (n_3009, n_1030, n_1131);
  xor g3322 (n_69, n_3009, n_1132);
  nand g3323 (n_3010, n_1030, n_1131);
  nand g3324 (n_3011, n_1132, n_1131);
  nand g3325 (n_3012, n_1030, n_1132);
  nand g3326 (n_149, n_3010, n_3011, n_3012);
  xor g3328 (n_1134, n_2773, A[57]);
  nand g3332 (n_1138, n_2774, n_2646, n_2782);
  xor g3333 (n_3017, A[60], n_1134);
  xor g3334 (n_68, n_3017, n_1135);
  nand g3335 (n_3018, A[60], n_1134);
  nand g3336 (n_3019, n_1135, n_1134);
  nand g3337 (n_3020, A[60], n_1135);
  nand g3338 (n_148, n_3018, n_3019, n_3020);
  nand g3345 (n_3024, A[60], n_1138);
  nand g3346 (n_147, n_3022, n_3023, n_3024);
  xor g3348 (n_66, n_2773, A[58]);
  nand g3350 (n_3027, A[58], A[59]);
  nand g3352 (n_146, n_2774, n_3027, n_3028);
  nor g11 (n_3044, A[2], A[0]);
  nor g13 (n_3040, A[3], A[1]);
  nor g15 (n_3050, A[2], n_220);
  nand g16 (n_3045, A[2], n_220);
  nor g17 (n_3046, n_138, n_219);
  nand g18 (n_3047, n_138, n_219);
  nor g19 (n_3056, n_137, n_218);
  nand g20 (n_3051, n_137, n_218);
  nor g21 (n_3052, n_136, n_217);
  nand g22 (n_3053, n_136, n_217);
  nor g23 (n_3062, n_135, n_216);
  nand g24 (n_3057, n_135, n_216);
  nor g25 (n_3058, n_134, n_215);
  nand g26 (n_3059, n_134, n_215);
  nor g27 (n_3068, n_133, n_214);
  nand g28 (n_3063, n_133, n_214);
  nor g29 (n_3064, n_132, n_213);
  nand g30 (n_3065, n_132, n_213);
  nor g31 (n_3074, n_131, n_212);
  nand g32 (n_3069, n_131, n_212);
  nor g33 (n_3070, n_130, n_211);
  nand g34 (n_3071, n_130, n_211);
  nor g35 (n_3080, n_129, n_210);
  nand g36 (n_3075, n_129, n_210);
  nor g37 (n_3076, n_128, n_209);
  nand g38 (n_3077, n_128, n_209);
  nor g39 (n_3086, n_127, n_208);
  nand g40 (n_3081, n_127, n_208);
  nor g41 (n_3082, n_126, n_207);
  nand g42 (n_3083, n_126, n_207);
  nor g43 (n_3092, n_125, n_206);
  nand g44 (n_3087, n_125, n_206);
  nor g45 (n_3088, n_124, n_205);
  nand g46 (n_3089, n_124, n_205);
  nor g47 (n_3098, n_123, n_204);
  nand g48 (n_3093, n_123, n_204);
  nor g49 (n_3094, n_122, n_203);
  nand g50 (n_3095, n_122, n_203);
  nor g51 (n_3104, n_121, n_202);
  nand g52 (n_3099, n_121, n_202);
  nor g53 (n_3100, n_120, n_201);
  nand g54 (n_3101, n_120, n_201);
  nor g55 (n_3110, n_119, n_200);
  nand g56 (n_3105, n_119, n_200);
  nor g57 (n_3106, n_118, n_199);
  nand g58 (n_3107, n_118, n_199);
  nor g59 (n_3116, n_117, n_198);
  nand g60 (n_3111, n_117, n_198);
  nor g61 (n_3112, n_116, n_197);
  nand g62 (n_3113, n_116, n_197);
  nor g63 (n_3122, n_115, n_196);
  nand g64 (n_3117, n_115, n_196);
  nor g65 (n_3118, n_114, n_195);
  nand g66 (n_3119, n_114, n_195);
  nor g67 (n_3128, n_113, n_194);
  nand g68 (n_3123, n_113, n_194);
  nor g69 (n_3124, n_112, n_193);
  nand g70 (n_3125, n_112, n_193);
  nor g71 (n_3134, n_111, n_192);
  nand g72 (n_3129, n_111, n_192);
  nor g73 (n_3130, n_110, n_191);
  nand g74 (n_3131, n_110, n_191);
  nor g75 (n_3140, n_109, n_190);
  nand g76 (n_3135, n_109, n_190);
  nor g77 (n_3136, n_108, n_189);
  nand g78 (n_3137, n_108, n_189);
  nor g79 (n_3146, n_107, n_188);
  nand g80 (n_3141, n_107, n_188);
  nor g81 (n_3142, n_106, n_187);
  nand g82 (n_3143, n_106, n_187);
  nor g83 (n_3152, n_105, n_186);
  nand g84 (n_3147, n_105, n_186);
  nor g85 (n_3148, n_104, n_185);
  nand g86 (n_3149, n_104, n_185);
  nor g87 (n_3158, n_103, n_184);
  nand g88 (n_3153, n_103, n_184);
  nor g89 (n_3154, n_102, n_183);
  nand g90 (n_3155, n_102, n_183);
  nor g91 (n_3164, n_101, n_182);
  nand g92 (n_3159, n_101, n_182);
  nor g93 (n_3160, n_100, n_181);
  nand g94 (n_3161, n_100, n_181);
  nor g95 (n_3170, n_99, n_180);
  nand g96 (n_3165, n_99, n_180);
  nor g97 (n_3166, n_98, n_179);
  nand g98 (n_3167, n_98, n_179);
  nor g99 (n_3176, n_97, n_178);
  nand g100 (n_3171, n_97, n_178);
  nor g101 (n_3172, n_96, n_177);
  nand g102 (n_3173, n_96, n_177);
  nor g103 (n_3182, n_95, n_176);
  nand g104 (n_3177, n_95, n_176);
  nor g105 (n_3178, n_94, n_175);
  nand g106 (n_3179, n_94, n_175);
  nor g107 (n_3188, n_93, n_174);
  nand g108 (n_3183, n_93, n_174);
  nor g109 (n_3184, n_92, n_173);
  nand g110 (n_3185, n_92, n_173);
  nor g111 (n_3194, n_91, n_172);
  nand g112 (n_3189, n_91, n_172);
  nor g113 (n_3190, n_90, n_171);
  nand g114 (n_3191, n_90, n_171);
  nor g115 (n_3200, n_89, n_170);
  nand g116 (n_3195, n_89, n_170);
  nor g117 (n_3196, n_88, n_169);
  nand g118 (n_3197, n_88, n_169);
  nor g119 (n_3206, n_87, n_168);
  nand g120 (n_3201, n_87, n_168);
  nor g121 (n_3202, n_86, n_167);
  nand g122 (n_3203, n_86, n_167);
  nor g123 (n_3212, n_85, n_166);
  nand g124 (n_3207, n_85, n_166);
  nor g125 (n_3208, n_84, n_165);
  nand g126 (n_3209, n_84, n_165);
  nor g127 (n_3218, n_83, n_164);
  nand g128 (n_3213, n_83, n_164);
  nor g129 (n_3214, n_82, n_163);
  nand g130 (n_3215, n_82, n_163);
  nor g131 (n_3224, n_81, n_162);
  nand g132 (n_3219, n_81, n_162);
  nor g133 (n_3220, n_80, n_161);
  nand g134 (n_3221, n_80, n_161);
  nor g135 (n_3230, n_79, n_160);
  nand g136 (n_3225, n_79, n_160);
  nor g137 (n_3226, n_78, n_159);
  nand g138 (n_3227, n_78, n_159);
  nor g139 (n_3236, n_77, n_158);
  nand g140 (n_3231, n_77, n_158);
  nor g141 (n_3232, n_76, n_157);
  nand g142 (n_3233, n_76, n_157);
  nor g143 (n_3242, n_75, n_156);
  nand g144 (n_3237, n_75, n_156);
  nor g145 (n_3238, n_74, n_155);
  nand g146 (n_3239, n_74, n_155);
  nor g147 (n_3248, n_73, n_154);
  nand g148 (n_3243, n_73, n_154);
  nor g149 (n_3244, n_72, n_153);
  nand g150 (n_3245, n_72, n_153);
  nor g151 (n_3254, n_71, n_152);
  nand g152 (n_3249, n_71, n_152);
  nor g153 (n_3250, n_70, n_151);
  nand g154 (n_3251, n_70, n_151);
  nor g155 (n_3260, n_69, n_150);
  nand g156 (n_3255, n_69, n_150);
  nor g157 (n_3256, n_68, n_149);
  nand g158 (n_3257, n_68, n_149);
  nor g159 (n_3266, n_67, n_148);
  nand g160 (n_3261, n_67, n_148);
  nor g161 (n_3262, n_66, n_147);
  nand g162 (n_3263, n_66, n_147);
  nor g172 (n_3042, n_1146, n_3040);
  nor g176 (n_3048, n_3045, n_3046);
  nor g179 (n_3283, n_3050, n_3046);
  nor g180 (n_3054, n_3051, n_3052);
  nor g183 (n_3277, n_3056, n_3052);
  nor g184 (n_3060, n_3057, n_3058);
  nor g187 (n_3290, n_3062, n_3058);
  nor g188 (n_3066, n_3063, n_3064);
  nor g191 (n_3284, n_3068, n_3064);
  nor g192 (n_3072, n_3069, n_3070);
  nor g195 (n_3297, n_3074, n_3070);
  nor g196 (n_3078, n_3075, n_3076);
  nor g199 (n_3291, n_3080, n_3076);
  nor g200 (n_3084, n_3081, n_3082);
  nor g203 (n_3304, n_3086, n_3082);
  nor g204 (n_3090, n_3087, n_3088);
  nor g207 (n_3298, n_3092, n_3088);
  nor g208 (n_3096, n_3093, n_3094);
  nor g211 (n_3311, n_3098, n_3094);
  nor g212 (n_3102, n_3099, n_3100);
  nor g215 (n_3305, n_3104, n_3100);
  nor g216 (n_3108, n_3105, n_3106);
  nor g219 (n_3318, n_3110, n_3106);
  nor g220 (n_3114, n_3111, n_3112);
  nor g223 (n_3312, n_3116, n_3112);
  nor g224 (n_3120, n_3117, n_3118);
  nor g227 (n_3325, n_3122, n_3118);
  nor g228 (n_3126, n_3123, n_3124);
  nor g231 (n_3319, n_3128, n_3124);
  nor g232 (n_3132, n_3129, n_3130);
  nor g235 (n_3332, n_3134, n_3130);
  nor g236 (n_3138, n_3135, n_3136);
  nor g239 (n_3326, n_3140, n_3136);
  nor g240 (n_3144, n_3141, n_3142);
  nor g243 (n_3339, n_3146, n_3142);
  nor g244 (n_3150, n_3147, n_3148);
  nor g247 (n_3333, n_3152, n_3148);
  nor g248 (n_3156, n_3153, n_3154);
  nor g251 (n_3346, n_3158, n_3154);
  nor g252 (n_3162, n_3159, n_3160);
  nor g255 (n_3340, n_3164, n_3160);
  nor g256 (n_3168, n_3165, n_3166);
  nor g259 (n_3353, n_3170, n_3166);
  nor g260 (n_3174, n_3171, n_3172);
  nor g263 (n_3347, n_3176, n_3172);
  nor g264 (n_3180, n_3177, n_3178);
  nor g267 (n_3360, n_3182, n_3178);
  nor g268 (n_3186, n_3183, n_3184);
  nor g271 (n_3354, n_3188, n_3184);
  nor g272 (n_3192, n_3189, n_3190);
  nor g275 (n_3367, n_3194, n_3190);
  nor g276 (n_3198, n_3195, n_3196);
  nor g279 (n_3361, n_3200, n_3196);
  nor g280 (n_3204, n_3201, n_3202);
  nor g283 (n_3374, n_3206, n_3202);
  nor g284 (n_3210, n_3207, n_3208);
  nor g287 (n_3368, n_3212, n_3208);
  nor g288 (n_3216, n_3213, n_3214);
  nor g291 (n_3381, n_3218, n_3214);
  nor g292 (n_3222, n_3219, n_3220);
  nor g295 (n_3375, n_3224, n_3220);
  nor g296 (n_3228, n_3225, n_3226);
  nor g299 (n_3388, n_3230, n_3226);
  nor g300 (n_3234, n_3231, n_3232);
  nor g303 (n_3382, n_3236, n_3232);
  nor g304 (n_3240, n_3237, n_3238);
  nor g307 (n_3395, n_3242, n_3238);
  nor g308 (n_3246, n_3243, n_3244);
  nor g311 (n_3389, n_3248, n_3244);
  nor g312 (n_3252, n_3249, n_3250);
  nor g315 (n_3402, n_3254, n_3250);
  nor g316 (n_3258, n_3255, n_3256);
  nor g319 (n_3396, n_3260, n_3256);
  nor g320 (n_3264, n_3261, n_3262);
  nor g323 (n_3409, n_3266, n_3262);
  nor g324 (n_3270, n_3267, n_3268);
  nor g327 (n_3403, n_3272, n_3268);
  nand g334 (n_3410, n_3283, n_3277);
  nand g339 (n_3420, n_3290, n_3284);
  nand g344 (n_3415, n_3297, n_3291);
  nand g349 (n_3426, n_3304, n_3298);
  nand g354 (n_3421, n_3311, n_3305);
  nand g359 (n_3432, n_3318, n_3312);
  nand g364 (n_3427, n_3325, n_3319);
  nand g369 (n_3438, n_3332, n_3326);
  nand g374 (n_3433, n_3339, n_3333);
  nand g379 (n_3444, n_3346, n_3340);
  nand g384 (n_3439, n_3353, n_3347);
  nand g389 (n_3450, n_3360, n_3354);
  nand g394 (n_3445, n_3367, n_3361);
  nand g399 (n_3456, n_3374, n_3368);
  nand g404 (n_3451, n_3381, n_3375);
  nand g409 (n_3462, n_3388, n_3382);
  nand g414 (n_3457, n_3395, n_3389);
  nand g419 (n_3468, n_3402, n_3396);
  nand g424 (n_3463, n_3409, n_3403);
  nand g427 (n_3470, n_3413, n_3414);
  nor g428 (n_3418, n_3415, n_3416);
  nor g431 (n_3469, n_3420, n_3415);
  nor g432 (n_3424, n_3421, n_3422);
  nor g435 (n_3479, n_3426, n_3421);
  nor g436 (n_3430, n_3427, n_3428);
  nor g439 (n_3473, n_3432, n_3427);
  nor g440 (n_3436, n_3433, n_3434);
  nor g443 (n_3486, n_3438, n_3433);
  nor g444 (n_3442, n_3439, n_3440);
  nor g447 (n_3480, n_3444, n_3439);
  nor g448 (n_3448, n_3445, n_3446);
  nor g451 (n_3493, n_3450, n_3445);
  nor g452 (n_3454, n_3451, n_3452);
  nor g455 (n_3487, n_3456, n_3451);
  nor g456 (n_3460, n_3457, n_3458);
  nor g459 (n_3500, n_3462, n_3457);
  nor g460 (n_3466, n_3463, n_3464);
  nor g463 (n_3494, n_3468, n_3463);
  nand g464 (n_3472, n_3469, n_3470);
  nand g465 (n_3502, n_3471, n_3472);
  nand g470 (n_3501, n_3479, n_3473);
  nand g475 (n_3511, n_3486, n_3480);
  nand g480 (n_3506, n_3493, n_3487);
  nand g485 (n_3518, n_3500, n_3494);
  nand g488 (n_3513, n_3504, n_3505);
  nor g489 (n_3509, n_3506, n_3507);
  nor g3360 (n_3512, n_3511, n_3506);
  nand g3361 (n_3515, n_3512, n_3513);
  nand g3362 (n_3519, n_3514, n_3515);
  nand g3365 (n_3525, n_3507, n_3517);
  nand g3368 (n_3676, n_3521, n_3522);
  nand g3369 (n_3523, n_3479, n_3502);
  nand g3370 (n_3532, n_3474, n_3523);
  nand g3371 (n_3524, n_3486, n_3513);
  nand g3372 (n_3537, n_3481, n_3524);
  nand g3373 (n_3526, n_3493, n_3525);
  nand g3374 (n_3542, n_3488, n_3526);
  nand g3375 (n_3527, n_3500, n_3519);
  nand g3376 (n_3547, n_3495, n_3527);
  nand g3379 (n_3552, n_3416, n_3529);
  nand g3382 (n_3555, n_3422, n_3531);
  nand g3385 (n_3558, n_3428, n_3534);
  nand g3388 (n_3561, n_3434, n_3536);
  nand g3391 (n_3564, n_3440, n_3539);
  nand g3394 (n_3567, n_3446, n_3541);
  nand g3397 (n_3570, n_3452, n_3544);
  nand g3400 (n_3573, n_3458, n_3546);
  nand g3403 (n_3576, n_3464, n_3549);
  nand g3405 (n_3582, n_3278, n_3550);
  nand g3406 (n_3551, n_3290, n_3470);
  nand g3407 (n_3587, n_3285, n_3551);
  nand g3408 (n_3553, n_3297, n_3552);
  nand g3409 (n_3592, n_3292, n_3553);
  nand g3410 (n_3554, n_3304, n_3502);
  nand g3411 (n_3597, n_3299, n_3554);
  nand g3412 (n_3556, n_3311, n_3555);
  nand g3413 (n_3602, n_3306, n_3556);
  nand g3414 (n_3557, n_3318, n_3532);
  nand g3415 (n_3607, n_3313, n_3557);
  nand g3416 (n_3559, n_3325, n_3558);
  nand g3417 (n_3612, n_3320, n_3559);
  nand g3418 (n_3560, n_3332, n_3513);
  nand g3419 (n_3617, n_3327, n_3560);
  nand g3420 (n_3562, n_3339, n_3561);
  nand g3421 (n_3622, n_3334, n_3562);
  nand g3422 (n_3563, n_3346, n_3537);
  nand g3423 (n_3627, n_3341, n_3563);
  nand g3424 (n_3565, n_3353, n_3564);
  nand g3425 (n_3632, n_3348, n_3565);
  nand g3426 (n_3566, n_3360, n_3525);
  nand g3427 (n_3637, n_3355, n_3566);
  nand g3428 (n_3568, n_3367, n_3567);
  nand g3429 (n_3642, n_3362, n_3568);
  nand g3430 (n_3569, n_3374, n_3542);
  nand g3431 (n_3647, n_3369, n_3569);
  nand g3432 (n_3571, n_3381, n_3570);
  nand g3433 (n_3652, n_3376, n_3571);
  nand g3434 (n_3572, n_3388, n_3519);
  nand g3435 (n_3657, n_3383, n_3572);
  nand g3436 (n_3574, n_3395, n_3573);
  nand g3437 (n_3662, n_3390, n_3574);
  nand g3438 (n_3575, n_3402, n_3547);
  nand g3439 (n_3667, n_3397, n_3575);
  nand g3440 (n_3577, n_3409, n_3576);
  nand g3441 (n_3672, n_3404, n_3577);
  nand g3447 (n_3686, n_3045, n_3581);
  nand g3450 (n_3690, n_3051, n_3584);
  nand g3453 (n_3694, n_3057, n_3586);
  nand g3456 (n_3698, n_3063, n_3589);
  nand g3459 (n_3702, n_3069, n_3591);
  nand g3462 (n_3706, n_3075, n_3594);
  nand g3465 (n_3710, n_3081, n_3596);
  nand g3468 (n_3714, n_3087, n_3599);
  nand g3471 (n_3718, n_3093, n_3601);
  nand g3474 (n_3722, n_3099, n_3604);
  nand g3477 (n_3726, n_3105, n_3606);
  nand g3480 (n_3730, n_3111, n_3609);
  nand g3483 (n_3734, n_3117, n_3611);
  nand g3486 (n_3738, n_3123, n_3614);
  nand g3489 (n_3742, n_3129, n_3616);
  nand g3492 (n_3746, n_3135, n_3619);
  nand g3495 (n_3750, n_3141, n_3621);
  nand g3498 (n_3754, n_3147, n_3624);
  nand g3501 (n_3758, n_3153, n_3626);
  nand g3504 (n_3762, n_3159, n_3629);
  nand g3507 (n_3766, n_3165, n_3631);
  nand g3510 (n_3770, n_3171, n_3634);
  nand g3513 (n_3774, n_3177, n_3636);
  nand g3516 (n_3778, n_3183, n_3639);
  nand g3519 (n_3782, n_3189, n_3641);
  nand g3522 (n_3786, n_3195, n_3644);
  nand g3525 (n_3790, n_3201, n_3646);
  nand g3528 (n_3794, n_3207, n_3649);
  nand g3531 (n_3798, n_3213, n_3651);
  nand g3534 (n_3802, n_3219, n_3654);
  nand g3537 (n_3806, n_3225, n_3656);
  nand g3540 (n_3810, n_3231, n_3659);
  nand g3543 (n_3814, n_3237, n_3661);
  nand g3546 (n_3818, n_3243, n_3664);
  nand g3549 (n_3822, n_3249, n_3666);
  nand g3552 (n_3826, n_3255, n_3669);
  nand g3555 (n_3830, n_3261, n_3671);
  nand g3558 (n_3834, n_3267, n_3674);
  xnor g3571 (Z[5], n_3686, n_3687);
  xnor g3573 (Z[6], n_3582, n_3688);
  xnor g3576 (Z[7], n_3690, n_3691);
  xnor g3578 (Z[8], n_3470, n_3692);
  xnor g3581 (Z[9], n_3694, n_3695);
  xnor g3583 (Z[10], n_3587, n_3696);
  xnor g3586 (Z[11], n_3698, n_3699);
  xnor g3588 (Z[12], n_3552, n_3700);
  xnor g3591 (Z[13], n_3702, n_3703);
  xnor g3593 (Z[14], n_3592, n_3704);
  xnor g3596 (Z[15], n_3706, n_3707);
  xnor g3598 (Z[16], n_3502, n_3708);
  xnor g3601 (Z[17], n_3710, n_3711);
  xnor g3603 (Z[18], n_3597, n_3712);
  xnor g3606 (Z[19], n_3714, n_3715);
  xnor g3608 (Z[20], n_3555, n_3716);
  xnor g3611 (Z[21], n_3718, n_3719);
  xnor g3613 (Z[22], n_3602, n_3720);
  xnor g3616 (Z[23], n_3722, n_3723);
  xnor g3618 (Z[24], n_3532, n_3724);
  xnor g3621 (Z[25], n_3726, n_3727);
  xnor g3623 (Z[26], n_3607, n_3728);
  xnor g3626 (Z[27], n_3730, n_3731);
  xnor g3628 (Z[28], n_3558, n_3732);
  xnor g3631 (Z[29], n_3734, n_3735);
  xnor g3633 (Z[30], n_3612, n_3736);
  xnor g3636 (Z[31], n_3738, n_3739);
  xnor g3638 (Z[32], n_3513, n_3740);
  xnor g3641 (Z[33], n_3742, n_3743);
  xnor g3643 (Z[34], n_3617, n_3744);
  xnor g3646 (Z[35], n_3746, n_3747);
  xnor g3648 (Z[36], n_3561, n_3748);
  xnor g3651 (Z[37], n_3750, n_3751);
  xnor g3653 (Z[38], n_3622, n_3752);
  xnor g3656 (Z[39], n_3754, n_3755);
  xnor g3658 (Z[40], n_3537, n_3756);
  xnor g3661 (Z[41], n_3758, n_3759);
  xnor g3663 (Z[42], n_3627, n_3760);
  xnor g3666 (Z[43], n_3762, n_3763);
  xnor g3668 (Z[44], n_3564, n_3764);
  xnor g3671 (Z[45], n_3766, n_3767);
  xnor g3673 (Z[46], n_3632, n_3768);
  xnor g3676 (Z[47], n_3770, n_3771);
  xnor g3678 (Z[48], n_3525, n_3772);
  xnor g3681 (Z[49], n_3774, n_3775);
  xnor g3683 (Z[50], n_3637, n_3776);
  xnor g3686 (Z[51], n_3778, n_3779);
  xnor g3688 (Z[52], n_3567, n_3780);
  xnor g3691 (Z[53], n_3782, n_3783);
  xnor g3693 (Z[54], n_3642, n_3784);
  xnor g3696 (Z[55], n_3786, n_3787);
  xnor g3698 (Z[56], n_3542, n_3788);
  xnor g3701 (Z[57], n_3790, n_3791);
  xnor g3703 (Z[58], n_3647, n_3792);
  xnor g3706 (Z[59], n_3794, n_3795);
  xnor g3708 (Z[60], n_3570, n_3796);
  xnor g3711 (Z[61], n_3798, n_3799);
  xnor g3713 (Z[62], n_3652, n_3800);
  xnor g3716 (Z[63], n_3802, n_3803);
  xnor g3718 (Z[64], n_3519, n_3804);
  xnor g3721 (Z[65], n_3806, n_3807);
  xnor g3723 (Z[66], n_3657, n_3808);
  xnor g3726 (Z[67], n_3810, n_3811);
  xnor g3728 (Z[68], n_3573, n_3812);
  xnor g3731 (Z[69], n_3814, n_3815);
  xnor g3733 (Z[70], n_3662, n_3816);
  xnor g3736 (Z[71], n_3818, n_3819);
  xnor g3738 (Z[72], n_3547, n_3820);
  xnor g3741 (Z[73], n_3822, n_3823);
  xnor g3743 (Z[74], n_3667, n_3824);
  xnor g3746 (Z[75], n_3826, n_3827);
  xnor g3748 (Z[76], n_3576, n_3828);
  xnor g3751 (Z[77], n_3830, n_3831);
  xnor g3753 (Z[78], n_3672, n_3832);
  xnor g3756 (Z[79], n_3834, n_3835);
  or g3771 (n_314, wc, wc0, n_138);
  not gc0 (wc0, n_1146);
  not gc (wc, n_1160);
  or g3772 (n_323, wc1, wc2, n_308);
  not gc2 (wc2, n_1160);
  not gc1 (wc1, n_1179);
  or g3773 (n_336, wc3, n_313, n_308);
  not gc3 (wc3, n_1207);
  or g3774 (n_353, wc4, wc5, n_313);
  not gc5 (wc5, n_1242);
  not gc4 (wc4, n_1243);
  or g3775 (n_375, wc6, wc7, n_313);
  not gc7 (wc7, n_1290);
  not gc6 (wc6, n_1291);
  or g3776 (n_423, wc8, wc9, n_308);
  not gc9 (wc9, n_1291);
  not gc8 (wc8, n_1338);
  or g3777 (n_451, wc10, wc11, n_313);
  not gc11 (wc11, n_1467);
  not gc10 (wc10, n_1468);
  or g3778 (n_479, wc12, wc13, n_322);
  not gc13 (wc13, n_1407);
  not gc12 (wc12, n_1531);
  or g3779 (n_505, wc14, wc15, n_335);
  not gc15 (wc15, n_1471);
  not gc14 (wc14, n_1595);
  or g3780 (n_533, wc16, wc17, n_352);
  not gc17 (wc17, n_1400);
  not gc16 (wc16, n_1659);
  or g3781 (n_561, wc18, wc19, n_373);
  not gc19 (wc19, n_1464);
  not gc18 (wc18, n_1723);
  or g3782 (n_589, wc20, wc21, n_398);
  not gc21 (wc21, n_1528);
  not gc20 (wc20, n_1787);
  xnor g3783 (n_2773, A[61], A[59]);
  or g3784 (n_2774, wc22, A[61]);
  not gc22 (wc22, A[59]);
  or g3785 (n_2776, wc23, A[61]);
  not gc23 (wc23, A[55]);
  xnor g3786 (n_2813, A[60], A[48]);
  or g3787 (n_2814, wc24, A[60]);
  not gc24 (wc24, A[48]);
  xnor g3788 (n_1085, n_2865, A[58]);
  or g3789 (n_2915, wc25, A[58]);
  not gc25 (wc25, A[56]);
  or g3790 (n_2916, wc26, A[58]);
  not gc26 (wc26, A[50]);
  xnor g3792 (n_1131, n_2613, A[60]);
  or g3793 (n_3007, wc27, A[60]);
  not gc27 (wc27, A[56]);
  or g3794 (n_3008, wc28, A[60]);
  not gc28 (wc28, A[58]);
  or g3795 (n_2782, wc29, A[61]);
  not gc29 (wc29, A[57]);
  or g3797 (n_3022, A[58], wc30);
  not gc30 (wc30, A[60]);
  or g3798 (n_3028, wc31, A[61]);
  not gc31 (wc31, A[58]);
  and g3799 (n_3268, wc32, A[61]);
  not gc32 (wc32, A[60]);
  or g3800 (n_3269, wc33, A[61]);
  not gc33 (wc33, A[60]);
  or g3801 (n_404, wc34, wc35, n_313);
  not gc35 (wc35, n_1347);
  not gc34 (wc34, n_1348);
  or g3802 (n_2872, A[60], wc36);
  not gc36 (wc36, n_1059);
  xnor g3803 (n_1105, n_2613, n_999);
  or g3804 (n_2955, A[58], wc37);
  not gc37 (wc37, n_999);
  or g3805 (n_2988, A[60], wc38);
  not gc38 (wc38, n_1119);
  and g3806 (n_3275, wc39, n_1143);
  not gc39 (wc39, n_3042);
  or g3808 (n_3680, n_3044, wc40);
  not gc40 (wc40, n_1146);
  or g3809 (n_3683, n_3040, wc41);
  not gc41 (wc41, n_1143);
  xnor g3810 (n_2781, A[61], A[57]);
  or g3811 (n_2784, wc42, A[61]);
  not gc42 (wc42, A[51]);
  or g3812 (n_2815, A[60], wc43);
  not gc43 (wc43, n_1030);
  xnor g3813 (n_2869, n_1030, A[60]);
  xnor g3814 (n_67, n_2677, n_1138);
  or g3815 (n_3023, A[58], wc44);
  not gc44 (wc44, n_1138);
  and g3816 (n_3272, A[60], wc45);
  not gc45 (wc45, n_146);
  or g3817 (n_3267, A[60], wc46);
  not gc46 (wc46, n_146);
  or g3818 (n_3684, wc47, n_3050);
  not gc47 (wc47, n_3045);
  or g3819 (n_3835, wc48, n_3268);
  not gc48 (wc48, n_3269);
  and g3820 (n_3278, wc49, n_3047);
  not gc49 (wc49, n_3048);
  not g3821 (Z[2], n_3680);
  or g3822 (n_3687, wc50, n_3046);
  not gc50 (wc50, n_3047);
  or g3823 (n_3688, wc51, n_3056);
  not gc51 (wc51, n_3051);
  and g3824 (n_3280, wc52, n_3053);
  not gc52 (wc52, n_3054);
  and g3825 (n_3406, n_3269, wc53);
  not gc53 (wc53, n_3270);
  or g3828 (n_3691, wc54, n_3052);
  not gc54 (wc54, n_3053);
  or g3829 (n_3832, wc55, n_3272);
  not gc55 (wc55, n_3267);
  and g3830 (n_3285, wc56, n_3059);
  not gc56 (wc56, n_3060);
  and g3831 (n_3281, wc57, n_3277);
  not gc57 (wc57, n_3278);
  or g3832 (n_3550, n_3275, wc58);
  not gc58 (wc58, n_3283);
  or g3833 (n_3581, n_3050, n_3275);
  xor g3834 (Z[3], n_1146, n_3683);
  xor g3835 (Z[4], n_3275, n_3684);
  or g3836 (n_3692, wc59, n_3062);
  not gc59 (wc59, n_3057);
  or g3837 (n_3695, wc60, n_3058);
  not gc60 (wc60, n_3059);
  and g3838 (n_3404, wc61, n_3263);
  not gc61 (wc61, n_3264);
  and g3839 (n_3413, wc62, n_3280);
  not gc62 (wc62, n_3281);
  or g3840 (n_3414, n_3410, n_3275);
  or g3841 (n_3696, wc63, n_3068);
  not gc63 (wc63, n_3063);
  or g3842 (n_3828, wc64, n_3266);
  not gc64 (wc64, n_3261);
  or g3843 (n_3831, wc65, n_3262);
  not gc65 (wc65, n_3263);
  and g3844 (n_3287, wc66, n_3065);
  not gc66 (wc66, n_3066);
  and g3845 (n_3292, wc67, n_3071);
  not gc67 (wc67, n_3072);
  and g3846 (n_3407, wc68, n_3403);
  not gc68 (wc68, n_3404);
  or g3847 (n_3584, wc69, n_3056);
  not gc69 (wc69, n_3582);
  or g3848 (n_3699, wc70, n_3064);
  not gc70 (wc70, n_3065);
  or g3849 (n_3700, wc71, n_3074);
  not gc71 (wc71, n_3069);
  or g3850 (n_3703, wc72, n_3070);
  not gc72 (wc72, n_3071);
  or g3851 (n_3827, wc73, n_3256);
  not gc73 (wc73, n_3257);
  and g3852 (n_3294, wc74, n_3077);
  not gc74 (wc74, n_3078);
  and g3853 (n_3397, wc75, n_3251);
  not gc75 (wc75, n_3252);
  and g3854 (n_3399, wc76, n_3257);
  not gc76 (wc76, n_3258);
  and g3855 (n_3288, wc77, n_3284);
  not gc77 (wc77, n_3285);
  and g3856 (n_3465, wc78, n_3406);
  not gc78 (wc78, n_3407);
  or g3857 (n_3586, wc79, n_3062);
  not gc79 (wc79, n_3470);
  or g3858 (n_3704, wc80, n_3080);
  not gc80 (wc80, n_3075);
  or g3859 (n_3707, wc81, n_3076);
  not gc81 (wc81, n_3077);
  or g3860 (n_3820, wc82, n_3254);
  not gc82 (wc82, n_3249);
  or g3861 (n_3823, wc83, n_3250);
  not gc83 (wc83, n_3251);
  or g3862 (n_3824, wc84, n_3260);
  not gc84 (wc84, n_3255);
  and g3863 (n_3299, wc85, n_3083);
  not gc85 (wc85, n_3084);
  and g3864 (n_3301, wc86, n_3089);
  not gc86 (wc86, n_3090);
  and g3865 (n_3416, wc87, n_3287);
  not gc87 (wc87, n_3288);
  and g3866 (n_3295, wc88, n_3291);
  not gc88 (wc88, n_3292);
  and g3867 (n_3400, wc89, n_3396);
  not gc89 (wc89, n_3397);
  or g3868 (n_3529, wc90, n_3420);
  not gc90 (wc90, n_3470);
  or g3869 (n_3708, wc91, n_3086);
  not gc91 (wc91, n_3081);
  or g3870 (n_3711, wc92, n_3082);
  not gc92 (wc92, n_3083);
  or g3871 (n_3712, wc93, n_3092);
  not gc93 (wc93, n_3087);
  or g3872 (n_3715, wc94, n_3088);
  not gc94 (wc94, n_3089);
  or g3873 (n_3716, wc95, n_3098);
  not gc95 (wc95, n_3093);
  or g3874 (n_3819, wc96, n_3244);
  not gc96 (wc96, n_3245);
  and g3875 (n_3306, wc97, n_3095);
  not gc97 (wc97, n_3096);
  and g3876 (n_3390, wc98, n_3239);
  not gc98 (wc98, n_3240);
  and g3877 (n_3392, wc99, n_3245);
  not gc99 (wc99, n_3246);
  and g3878 (n_3417, wc100, n_3294);
  not gc100 (wc100, n_3295);
  and g3879 (n_3302, wc101, n_3298);
  not gc101 (wc101, n_3299);
  and g3880 (n_3464, wc102, n_3399);
  not gc102 (wc102, n_3400);
  or g3881 (n_3589, wc103, n_3068);
  not gc103 (wc103, n_3587);
  or g3882 (n_3719, wc104, n_3094);
  not gc104 (wc104, n_3095);
  or g3883 (n_3720, wc105, n_3104);
  not gc105 (wc105, n_3099);
  or g3884 (n_3812, wc106, n_3242);
  not gc106 (wc106, n_3237);
  or g3885 (n_3815, wc107, n_3238);
  not gc107 (wc107, n_3239);
  or g3886 (n_3816, wc108, n_3248);
  not gc108 (wc108, n_3243);
  and g3887 (n_3308, wc109, n_3101);
  not gc109 (wc109, n_3102);
  and g3888 (n_3313, wc110, n_3107);
  not gc110 (wc110, n_3108);
  and g3889 (n_3315, wc111, n_3113);
  not gc111 (wc111, n_3114);
  and g3890 (n_3320, wc112, n_3119);
  not gc112 (wc112, n_3120);
  and g3891 (n_3322, wc113, n_3125);
  not gc113 (wc113, n_3126);
  and g3892 (n_3327, wc114, n_3131);
  not gc114 (wc114, n_3132);
  and g3893 (n_3329, wc115, n_3137);
  not gc115 (wc115, n_3138);
  and g3894 (n_3334, wc116, n_3143);
  not gc116 (wc116, n_3144);
  and g3895 (n_3336, wc117, n_3149);
  not gc117 (wc117, n_3150);
  and g3896 (n_3341, wc118, n_3155);
  not gc118 (wc118, n_3156);
  and g3897 (n_3343, wc119, n_3161);
  not gc119 (wc119, n_3162);
  and g3898 (n_3348, wc120, n_3167);
  not gc120 (wc120, n_3168);
  and g3899 (n_3350, wc121, n_3173);
  not gc121 (wc121, n_3174);
  and g3900 (n_3355, wc122, n_3179);
  not gc122 (wc122, n_3180);
  and g3901 (n_3357, wc123, n_3185);
  not gc123 (wc123, n_3186);
  and g3902 (n_3362, wc124, n_3191);
  not gc124 (wc124, n_3192);
  and g3903 (n_3364, wc125, n_3197);
  not gc125 (wc125, n_3198);
  and g3904 (n_3369, wc126, n_3203);
  not gc126 (wc126, n_3204);
  and g3905 (n_3371, wc127, n_3209);
  not gc127 (wc127, n_3210);
  and g3906 (n_3376, wc128, n_3215);
  not gc128 (wc128, n_3216);
  and g3907 (n_3422, wc129, n_3301);
  not gc129 (wc129, n_3302);
  and g3908 (n_3393, wc130, n_3389);
  not gc130 (wc130, n_3390);
  or g3909 (n_3591, wc131, n_3074);
  not gc131 (wc131, n_3552);
  or g3910 (n_3723, wc132, n_3100);
  not gc132 (wc132, n_3101);
  or g3911 (n_3724, wc133, n_3110);
  not gc133 (wc133, n_3105);
  or g3912 (n_3727, wc134, n_3106);
  not gc134 (wc134, n_3107);
  or g3913 (n_3728, wc135, n_3116);
  not gc135 (wc135, n_3111);
  or g3914 (n_3731, wc136, n_3112);
  not gc136 (wc136, n_3113);
  or g3915 (n_3732, wc137, n_3122);
  not gc137 (wc137, n_3117);
  or g3916 (n_3735, wc138, n_3118);
  not gc138 (wc138, n_3119);
  or g3917 (n_3736, wc139, n_3128);
  not gc139 (wc139, n_3123);
  or g3918 (n_3739, wc140, n_3124);
  not gc140 (wc140, n_3125);
  or g3919 (n_3740, wc141, n_3134);
  not gc141 (wc141, n_3129);
  or g3920 (n_3743, wc142, n_3130);
  not gc142 (wc142, n_3131);
  or g3921 (n_3744, wc143, n_3140);
  not gc143 (wc143, n_3135);
  or g3922 (n_3747, wc144, n_3136);
  not gc144 (wc144, n_3137);
  or g3923 (n_3748, wc145, n_3146);
  not gc145 (wc145, n_3141);
  or g3924 (n_3751, wc146, n_3142);
  not gc146 (wc146, n_3143);
  or g3925 (n_3752, wc147, n_3152);
  not gc147 (wc147, n_3147);
  or g3926 (n_3755, wc148, n_3148);
  not gc148 (wc148, n_3149);
  or g3927 (n_3756, wc149, n_3158);
  not gc149 (wc149, n_3153);
  or g3928 (n_3759, wc150, n_3154);
  not gc150 (wc150, n_3155);
  or g3929 (n_3760, wc151, n_3164);
  not gc151 (wc151, n_3159);
  or g3930 (n_3763, wc152, n_3160);
  not gc152 (wc152, n_3161);
  or g3931 (n_3764, wc153, n_3170);
  not gc153 (wc153, n_3165);
  or g3932 (n_3767, wc154, n_3166);
  not gc154 (wc154, n_3167);
  or g3933 (n_3768, wc155, n_3176);
  not gc155 (wc155, n_3171);
  or g3934 (n_3771, wc156, n_3172);
  not gc156 (wc156, n_3173);
  or g3935 (n_3772, wc157, n_3182);
  not gc157 (wc157, n_3177);
  or g3936 (n_3775, wc158, n_3178);
  not gc158 (wc158, n_3179);
  or g3937 (n_3776, wc159, n_3188);
  not gc159 (wc159, n_3183);
  or g3938 (n_3779, wc160, n_3184);
  not gc160 (wc160, n_3185);
  or g3939 (n_3780, wc161, n_3194);
  not gc161 (wc161, n_3189);
  or g3940 (n_3783, wc162, n_3190);
  not gc162 (wc162, n_3191);
  or g3941 (n_3784, wc163, n_3200);
  not gc163 (wc163, n_3195);
  or g3942 (n_3787, wc164, n_3196);
  not gc164 (wc164, n_3197);
  or g3943 (n_3788, wc165, n_3206);
  not gc165 (wc165, n_3201);
  or g3944 (n_3791, wc166, n_3202);
  not gc166 (wc166, n_3203);
  or g3945 (n_3792, wc167, n_3212);
  not gc167 (wc167, n_3207);
  or g3946 (n_3795, wc168, n_3208);
  not gc168 (wc168, n_3209);
  or g3947 (n_3796, wc169, n_3218);
  not gc169 (wc169, n_3213);
  or g3948 (n_3799, wc170, n_3214);
  not gc170 (wc170, n_3215);
  or g3949 (n_3800, wc171, n_3224);
  not gc171 (wc171, n_3219);
  and g3950 (n_3378, wc172, n_3221);
  not gc172 (wc172, n_3222);
  and g3951 (n_3309, wc173, n_3305);
  not gc173 (wc173, n_3306);
  and g3952 (n_3316, wc174, n_3312);
  not gc174 (wc174, n_3313);
  and g3953 (n_3323, wc175, n_3319);
  not gc175 (wc175, n_3320);
  and g3954 (n_3330, wc176, n_3326);
  not gc176 (wc176, n_3327);
  and g3955 (n_3337, wc177, n_3333);
  not gc177 (wc177, n_3334);
  and g3956 (n_3344, wc178, n_3340);
  not gc178 (wc178, n_3341);
  and g3957 (n_3351, wc179, n_3347);
  not gc179 (wc179, n_3348);
  and g3958 (n_3358, wc180, n_3354);
  not gc180 (wc180, n_3355);
  and g3959 (n_3365, wc181, n_3361);
  not gc181 (wc181, n_3362);
  and g3960 (n_3372, wc182, n_3368);
  not gc182 (wc182, n_3369);
  and g3961 (n_3459, wc183, n_3392);
  not gc183 (wc183, n_3393);
  and g3962 (n_3471, n_3417, wc184);
  not gc184 (wc184, n_3418);
  and g3963 (n_3497, n_3465, wc185);
  not gc185 (wc185, n_3466);
  or g3964 (n_3803, wc186, n_3220);
  not gc186 (wc186, n_3221);
  or g3965 (n_3804, wc187, n_3230);
  not gc187 (wc187, n_3225);
  and g3966 (n_3383, wc188, n_3227);
  not gc188 (wc188, n_3228);
  and g3967 (n_3423, wc189, n_3308);
  not gc189 (wc189, n_3309);
  and g3968 (n_3428, wc190, n_3315);
  not gc190 (wc190, n_3316);
  and g3969 (n_3429, wc191, n_3322);
  not gc191 (wc191, n_3323);
  and g3970 (n_3434, wc192, n_3329);
  not gc192 (wc192, n_3330);
  and g3971 (n_3435, wc193, n_3336);
  not gc193 (wc193, n_3337);
  and g3972 (n_3440, wc194, n_3343);
  not gc194 (wc194, n_3344);
  and g3973 (n_3441, wc195, n_3350);
  not gc195 (wc195, n_3351);
  and g3974 (n_3446, wc196, n_3357);
  not gc196 (wc196, n_3358);
  and g3975 (n_3447, wc197, n_3364);
  not gc197 (wc197, n_3365);
  and g3976 (n_3452, wc198, n_3371);
  not gc198 (wc198, n_3372);
  and g3977 (n_3379, wc199, n_3375);
  not gc199 (wc199, n_3376);
  or g3978 (n_3594, wc200, n_3080);
  not gc200 (wc200, n_3592);
  or g3979 (n_3807, wc201, n_3226);
  not gc201 (wc201, n_3227);
  or g3980 (n_3808, wc202, n_3236);
  not gc202 (wc202, n_3231);
  and g3981 (n_3385, wc203, n_3233);
  not gc203 (wc203, n_3234);
  and g3982 (n_3453, wc204, n_3378);
  not gc204 (wc204, n_3379);
  or g3983 (n_3531, wc205, n_3426);
  not gc205 (wc205, n_3502);
  or g3984 (n_3596, wc206, n_3086);
  not gc206 (wc206, n_3502);
  or g3985 (n_3811, wc207, n_3232);
  not gc207 (wc207, n_3233);
  and g3986 (n_3386, wc208, n_3382);
  not gc208 (wc208, n_3383);
  and g3987 (n_3474, n_3423, wc209);
  not gc209 (wc209, n_3424);
  and g3988 (n_3476, n_3429, wc210);
  not gc210 (wc210, n_3430);
  and g3989 (n_3481, n_3435, wc211);
  not gc211 (wc211, n_3436);
  and g3990 (n_3483, n_3441, wc212);
  not gc212 (wc212, n_3442);
  and g3991 (n_3488, n_3447, wc213);
  not gc213 (wc213, n_3448);
  or g3992 (n_3505, n_3501, wc214);
  not gc214 (wc214, n_3502);
  and g3993 (n_3458, wc215, n_3385);
  not gc215 (wc215, n_3386);
  and g3994 (n_3490, n_3453, wc216);
  not gc216 (wc216, n_3454);
  and g3995 (n_3477, wc217, n_3473);
  not gc217 (wc217, n_3474);
  and g3996 (n_3484, wc218, n_3480);
  not gc218 (wc218, n_3481);
  and g3997 (n_3491, wc219, n_3487);
  not gc219 (wc219, n_3488);
  or g3998 (n_3599, wc220, n_3092);
  not gc220 (wc220, n_3597);
  or g3999 (n_3601, wc221, n_3098);
  not gc221 (wc221, n_3555);
  and g4000 (n_3504, wc222, n_3476);
  not gc222 (wc222, n_3477);
  and g4001 (n_3507, wc223, n_3483);
  not gc223 (wc223, n_3484);
  or g4002 (n_3534, wc224, n_3432);
  not gc224 (wc224, n_3532);
  or g4003 (n_3606, wc225, n_3110);
  not gc225 (wc225, n_3532);
  and g4004 (n_3495, n_3459, wc226);
  not gc226 (wc226, n_3460);
  and g4005 (n_3508, wc227, n_3490);
  not gc227 (wc227, n_3491);
  or g4006 (n_3604, wc228, n_3104);
  not gc228 (wc228, n_3602);
  and g4007 (n_3498, wc229, n_3494);
  not gc229 (wc229, n_3495);
  or g4008 (n_3517, wc230, n_3511);
  not gc230 (wc230, n_3513);
  or g4009 (n_3536, wc231, n_3438);
  not gc231 (wc231, n_3513);
  or g4010 (n_3609, wc232, n_3116);
  not gc232 (wc232, n_3607);
  or g4011 (n_3611, wc233, n_3122);
  not gc233 (wc233, n_3558);
  or g4012 (n_3616, wc234, n_3134);
  not gc234 (wc234, n_3513);
  and g4013 (n_3521, wc235, n_3497);
  not gc235 (wc235, n_3498);
  and g4014 (n_3514, n_3508, wc236);
  not gc236 (wc236, n_3509);
  or g4015 (n_3539, wc237, n_3444);
  not gc237 (wc237, n_3537);
  or g4016 (n_3541, wc238, n_3450);
  not gc238 (wc238, n_3525);
  or g4017 (n_3614, wc239, n_3128);
  not gc239 (wc239, n_3612);
  or g4018 (n_3619, wc240, n_3140);
  not gc240 (wc240, n_3617);
  or g4019 (n_3621, wc241, n_3146);
  not gc241 (wc241, n_3561);
  or g4020 (n_3626, wc242, n_3158);
  not gc242 (wc242, n_3537);
  or g4021 (n_3636, wc243, n_3182);
  not gc243 (wc243, n_3525);
  or g4022 (n_3522, wc244, n_3518);
  not gc244 (wc244, n_3519);
  or g4023 (n_3546, wc245, n_3462);
  not gc245 (wc245, n_3519);
  or g4024 (n_3656, wc246, n_3230);
  not gc246 (wc246, n_3519);
  or g4025 (n_3544, wc247, n_3456);
  not gc247 (wc247, n_3542);
  or g4026 (n_3624, wc248, n_3152);
  not gc248 (wc248, n_3622);
  or g4027 (n_3629, wc249, n_3164);
  not gc249 (wc249, n_3627);
  or g4028 (n_3631, wc250, n_3170);
  not gc250 (wc250, n_3564);
  or g4029 (n_3639, wc251, n_3188);
  not gc251 (wc251, n_3637);
  or g4030 (n_3641, wc252, n_3194);
  not gc252 (wc252, n_3567);
  or g4031 (n_3646, wc253, n_3206);
  not gc253 (wc253, n_3542);
  or g4032 (n_3549, wc254, n_3468);
  not gc254 (wc254, n_3547);
  or g4033 (n_3659, wc255, n_3236);
  not gc255 (wc255, n_3657);
  or g4034 (n_3661, wc256, n_3242);
  not gc256 (wc256, n_3573);
  or g4035 (n_3666, wc257, n_3254);
  not gc257 (wc257, n_3547);
  not g4036 (Z[80], n_3676);
  or g4037 (n_3634, wc258, n_3176);
  not gc258 (wc258, n_3632);
  or g4038 (n_3644, wc259, n_3200);
  not gc259 (wc259, n_3642);
  or g4039 (n_3649, wc260, n_3212);
  not gc260 (wc260, n_3647);
  or g4040 (n_3651, wc261, n_3218);
  not gc261 (wc261, n_3570);
  or g4041 (n_3664, wc262, n_3248);
  not gc262 (wc262, n_3662);
  or g4042 (n_3669, wc263, n_3260);
  not gc263 (wc263, n_3667);
  or g4043 (n_3671, wc264, n_3266);
  not gc264 (wc264, n_3576);
  or g4044 (n_3654, wc265, n_3224);
  not gc265 (wc265, n_3652);
  or g4045 (n_3674, n_3272, wc266);
  not gc266 (wc266, n_3672);
endmodule

module mult_signed_const_14732_GENERIC(A, Z);
  input [61:0] A;
  output [80:0] Z;
  wire [61:0] A;
  wire [80:0] Z;
  mult_signed_const_14732_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_15239_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [63:0] A;
  output [82:0] Z;
  wire [63:0] A;
  wire [82:0] Z;
  wire n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213;
  wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_315;
  wire n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323;
  wire n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331;
  wire n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339;
  wire n_340, n_341, n_342, n_343, n_344, n_345, n_346, n_347;
  wire n_348, n_349, n_350, n_351, n_352, n_353, n_354, n_355;
  wire n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371;
  wire n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395;
  wire n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403;
  wire n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411;
  wire n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419;
  wire n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476;
  wire n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484;
  wire n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492;
  wire n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500;
  wire n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508;
  wire n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516;
  wire n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524;
  wire n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_532;
  wire n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540;
  wire n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548;
  wire n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_556;
  wire n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564;
  wire n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572;
  wire n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580;
  wire n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588;
  wire n_589, n_590, n_591, n_592, n_593, n_594, n_595, n_596;
  wire n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604;
  wire n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612;
  wire n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620;
  wire n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628;
  wire n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636;
  wire n_637, n_638, n_639, n_640, n_641, n_642, n_643, n_644;
  wire n_645, n_646, n_647, n_648, n_649, n_650, n_651, n_652;
  wire n_653, n_654, n_655, n_656, n_657, n_658, n_659, n_660;
  wire n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668;
  wire n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676;
  wire n_677, n_678, n_679, n_680, n_681, n_682, n_683, n_684;
  wire n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692;
  wire n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700;
  wire n_701, n_702, n_703, n_704, n_705, n_706, n_707, n_708;
  wire n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716;
  wire n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724;
  wire n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732;
  wire n_733, n_734, n_735, n_736, n_737, n_738, n_739, n_740;
  wire n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748;
  wire n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756;
  wire n_757, n_758, n_759, n_760, n_761, n_762, n_763, n_764;
  wire n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772;
  wire n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780;
  wire n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788;
  wire n_789, n_790, n_791, n_792, n_793, n_794, n_795, n_796;
  wire n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804;
  wire n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812;
  wire n_813, n_814, n_815, n_816, n_817, n_818, n_819, n_820;
  wire n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828;
  wire n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836;
  wire n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844;
  wire n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860;
  wire n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868;
  wire n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876;
  wire n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884;
  wire n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892;
  wire n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900;
  wire n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908;
  wire n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932;
  wire n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940;
  wire n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948;
  wire n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956;
  wire n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964;
  wire n_965, n_966, n_967, n_968, n_969, n_970, n_971, n_972;
  wire n_973, n_974, n_975, n_976, n_977, n_978, n_979, n_980;
  wire n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988;
  wire n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996;
  wire n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004;
  wire n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012;
  wire n_1013, n_1014, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022;
  wire n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030;
  wire n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041;
  wire n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1049, n_1050;
  wire n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058;
  wire n_1059, n_1060, n_1061, n_1062, n_1065, n_1066, n_1067, n_1068;
  wire n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
  wire n_1077, n_1079, n_1080, n_1082, n_1083, n_1084, n_1085, n_1086;
  wire n_1087, n_1088, n_1089, n_1090, n_1094, n_1096, n_1097, n_1098;
  wire n_1099, n_1100, n_1101, n_1102, n_1103, n_1105, n_1109, n_1110;
  wire n_1111, n_1112, n_1113, n_1114, n_1119, n_1120, n_1121, n_1122;
  wire n_1123, n_1124, n_1125, n_1127, n_1130, n_1131, n_1132, n_1133;
  wire n_1134, n_1140, n_1141, n_1142, n_1143, n_1147, n_1148, n_1149;
  wire n_1150, n_1154, n_1155, n_1156, n_1157, n_1159, n_1161, n_1162;
  wire n_1166, n_1167, n_1169, n_1170, n_1173, n_1176, n_1177, n_1178;
  wire n_1179, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1188;
  wire n_1189, n_1190, n_1191, n_1195, n_1196, n_1197, n_1198, n_1199;
  wire n_1200, n_1201, n_1202, n_1204, n_1206, n_1207, n_1208, n_1209;
  wire n_1210, n_1211, n_1212, n_1214, n_1216, n_1217, n_1218, n_1219;
  wire n_1220, n_1221, n_1222, n_1223, n_1226, n_1228, n_1229, n_1230;
  wire n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238;
  wire n_1239, n_1242, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251;
  wire n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1260, n_1261;
  wire n_1262, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270;
  wire n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278;
  wire n_1280, n_1281, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288;
  wire n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1298, n_1299, n_1300, n_1301, n_1303, n_1304, n_1306;
  wire n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314;
  wire n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1323, n_1324;
  wire n_1325, n_1326, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333;
  wire n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341;
  wire n_1342, n_1343, n_1344, n_1345, n_1346, n_1352, n_1353, n_1356;
  wire n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364;
  wire n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372;
  wire n_1373, n_1375, n_1376, n_1378, n_1379, n_1382, n_1383, n_1384;
  wire n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392;
  wire n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400;
  wire n_1401, n_1402, n_1406, n_1407, n_1408, n_1409, n_1410, n_1412;
  wire n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420;
  wire n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428;
  wire n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1440;
  wire n_1441, n_1442, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449;
  wire n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457;
  wire n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465;
  wire n_1466, n_1467, n_1472, n_1474, n_1476, n_1477, n_1478, n_1479;
  wire n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487;
  wire n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495;
  wire n_1496, n_1497, n_1498, n_1499, n_1502, n_1503, n_1504, n_1505;
  wire n_1506, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514;
  wire n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522;
  wire n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530;
  wire n_1531, n_1534, n_1536, n_1537, n_1540, n_1541, n_1542, n_1543;
  wire n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551;
  wire n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559;
  wire n_1560, n_1561, n_1562, n_1563, n_1566, n_1568, n_1569, n_1572;
  wire n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580;
  wire n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588;
  wire n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596;
  wire n_1598, n_1600, n_1601, n_1604, n_1605, n_1606, n_1607, n_1608;
  wire n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616;
  wire n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624;
  wire n_1625, n_1626, n_1627, n_1630, n_1632, n_1633, n_1636, n_1637;
  wire n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645;
  wire n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653;
  wire n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661;
  wire n_1662, n_1664, n_1665, n_1668, n_1669, n_1670, n_1671, n_1672;
  wire n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680;
  wire n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688;
  wire n_1689, n_1690, n_1691, n_1694, n_1696, n_1697, n_1700, n_1701;
  wire n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709;
  wire n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717;
  wire n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1726;
  wire n_1728, n_1729, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737;
  wire n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745;
  wire n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753;
  wire n_1754, n_1755, n_1758, n_1760, n_1761, n_1764, n_1765, n_1766;
  wire n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774;
  wire n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782;
  wire n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1790, n_1792;
  wire n_1793, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802;
  wire n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810;
  wire n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818;
  wire n_1819, n_1822, n_1824, n_1825, n_1828, n_1829, n_1830, n_1831;
  wire n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839;
  wire n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847;
  wire n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1856;
  wire n_1857, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866;
  wire n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874;
  wire n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882;
  wire n_1883, n_1886, n_1888, n_1889, n_1892, n_1893, n_1894, n_1895;
  wire n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903;
  wire n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911;
  wire n_1912, n_1913, n_1914, n_1915, n_1918, n_1920, n_1921, n_1924;
  wire n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932;
  wire n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940;
  wire n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1950;
  wire n_1952, n_1953, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961;
  wire n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969;
  wire n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977;
  wire n_1978, n_1979, n_1982, n_1984, n_1985, n_1988, n_1989, n_1990;
  wire n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998;
  wire n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006;
  wire n_2007, n_2008, n_2009, n_2010, n_2011, n_2014, n_2016, n_2017;
  wire n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027;
  wire n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035;
  wire n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043;
  wire n_2046, n_2048, n_2049, n_2052, n_2053, n_2054, n_2055, n_2056;
  wire n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064;
  wire n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072;
  wire n_2073, n_2074, n_2075, n_2078, n_2080, n_2081, n_2084, n_2085;
  wire n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093;
  wire n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101;
  wire n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2110, n_2112;
  wire n_2113, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122;
  wire n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130;
  wire n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138;
  wire n_2139, n_2142, n_2144, n_2145, n_2148, n_2149, n_2150, n_2151;
  wire n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159;
  wire n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167;
  wire n_2168, n_2169, n_2170, n_2171, n_2174, n_2176, n_2177, n_2180;
  wire n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188;
  wire n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196;
  wire n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2206;
  wire n_2208, n_2209, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217;
  wire n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225;
  wire n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233;
  wire n_2234, n_2235, n_2238, n_2240, n_2241, n_2244, n_2245, n_2246;
  wire n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254;
  wire n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262;
  wire n_2263, n_2264, n_2265, n_2266, n_2267, n_2270, n_2272, n_2273;
  wire n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283;
  wire n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291;
  wire n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299;
  wire n_2302, n_2304, n_2305, n_2308, n_2309, n_2310, n_2311, n_2312;
  wire n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320;
  wire n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328;
  wire n_2329, n_2330, n_2331, n_2334, n_2336, n_2337, n_2340, n_2341;
  wire n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349;
  wire n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357;
  wire n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2366, n_2368;
  wire n_2369, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378;
  wire n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386;
  wire n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394;
  wire n_2395, n_2398, n_2400, n_2401, n_2404, n_2405, n_2406, n_2407;
  wire n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415;
  wire n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423;
  wire n_2424, n_2425, n_2426, n_2427, n_2430, n_2432, n_2433, n_2436;
  wire n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444;
  wire n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452;
  wire n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2462;
  wire n_2464, n_2465, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473;
  wire n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481;
  wire n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489;
  wire n_2490, n_2491, n_2494, n_2496, n_2497, n_2500, n_2501, n_2502;
  wire n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510;
  wire n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518;
  wire n_2519, n_2520, n_2521, n_2522, n_2523, n_2526, n_2528, n_2529;
  wire n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539;
  wire n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547;
  wire n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555;
  wire n_2558, n_2560, n_2561, n_2564, n_2565, n_2566, n_2567, n_2568;
  wire n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576;
  wire n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584;
  wire n_2585, n_2586, n_2587, n_2590, n_2592, n_2593, n_2596, n_2597;
  wire n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605;
  wire n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613;
  wire n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2622, n_2624;
  wire n_2625, n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634;
  wire n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642;
  wire n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650;
  wire n_2651, n_2654, n_2656, n_2657, n_2660, n_2661, n_2662, n_2663;
  wire n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671;
  wire n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679;
  wire n_2680, n_2681, n_2682, n_2683, n_2686, n_2688, n_2689, n_2692;
  wire n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700;
  wire n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708;
  wire n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2718;
  wire n_2720, n_2721, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729;
  wire n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737;
  wire n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745;
  wire n_2746, n_2747, n_2750, n_2752, n_2753, n_2756, n_2757, n_2758;
  wire n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766;
  wire n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774;
  wire n_2775, n_2776, n_2777, n_2778, n_2779, n_2782, n_2784, n_2785;
  wire n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, n_2795;
  wire n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803;
  wire n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811;
  wire n_2812, n_2813, n_2814, n_2816, n_2820, n_2821, n_2822, n_2823;
  wire n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831;
  wire n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839;
  wire n_2840, n_2841, n_2843, n_2844, n_2845, n_2848, n_2851, n_2852;
  wire n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860;
  wire n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868;
  wire n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, n_2878;
  wire n_2880, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889;
  wire n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897;
  wire n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905;
  wire n_2908, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918;
  wire n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926;
  wire n_2927, n_2928, n_2929, n_2930, n_2931, n_2936, n_2939, n_2942;
  wire n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950;
  wire n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958;
  wire n_2959, n_2960, n_2968, n_2970, n_2971, n_2972, n_2973, n_2974;
  wire n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982;
  wire n_2983, n_2992, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999;
  wire n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007;
  wire n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021;
  wire n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3036, n_3037;
  wire n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045;
  wire n_3046, n_3047, n_3054, n_3055, n_3056, n_3058, n_3059, n_3060;
  wire n_3061, n_3062, n_3063, n_3070, n_3071, n_3072, n_3073, n_3074;
  wire n_3075, n_3076, n_3077, n_3078, n_3079, n_3086, n_3087, n_3088;
  wire n_3089, n_3090, n_3091, n_3096, n_3097, n_3098, n_3099, n_3100;
  wire n_3101, n_3102, n_3103, n_3106, n_3107, n_3108, n_3109, n_3110;
  wire n_3111, n_3115, n_3116, n_3117, n_3118, n_3119, n_3121, n_3122;
  wire n_3123, n_3126, n_3127, n_3146, n_3147, n_3149, n_3150, n_3151;
  wire n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159;
  wire n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167;
  wire n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175;
  wire n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183;
  wire n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191;
  wire n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199;
  wire n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207;
  wire n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215;
  wire n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, n_3222, n_3223;
  wire n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, n_3231;
  wire n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239;
  wire n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247;
  wire n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255;
  wire n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3263;
  wire n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271;
  wire n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279;
  wire n_3280, n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287;
  wire n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, n_3294, n_3295;
  wire n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, n_3303;
  wire n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311;
  wire n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319;
  wire n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327;
  wire n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335;
  wire n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343;
  wire n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351;
  wire n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359;
  wire n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, n_3366, n_3367;
  wire n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, n_3375;
  wire n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383;
  wire n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391;
  wire n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399;
  wire n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, n_3407;
  wire n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415;
  wire n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423;
  wire n_3424, n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431;
  wire n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, n_3438, n_3439;
  wire n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, n_3447;
  wire n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455;
  wire n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463;
  wire n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471;
  wire n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, n_3479;
  wire n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487;
  wire n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495;
  wire n_3496, n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503;
  wire n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, n_3510, n_3511;
  wire n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3519;
  wire n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527;
  wire n_3528, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535;
  wire n_3536, n_3537, n_3538, n_3539;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g508 (n_226, A[4], A[0]);
  and g2 (n_142, A[4], A[0]);
  xor g509 (n_1176, A[1], A[3]);
  xor g510 (n_225, n_1176, A[5]);
  nand g3 (n_1177, A[1], A[3]);
  nand g511 (n_1178, A[5], A[3]);
  nand g512 (n_1179, A[1], A[5]);
  nand g513 (n_141, n_1177, n_1178, n_1179);
  xor g514 (n_315, A[6], A[4]);
  and g515 (n_316, A[6], A[4]);
  xor g516 (Z[2], A[0], A[2]);
  xor g517 (n_224, Z[2], n_315);
  nand g518 (n_1181, A[0], A[2]);
  nand g4 (n_1182, n_315, A[2]);
  nand g5 (n_1183, A[0], n_315);
  nand g519 (n_140, n_1181, n_1182, n_1183);
  xor g520 (n_1184, A[1], A[7]);
  xor g521 (n_317, n_1184, A[5]);
  nand g522 (n_1185, A[1], A[7]);
  nand g523 (n_1186, A[5], A[7]);
  nand g6 (n_319, n_1185, n_1186, n_1179);
  xor g525 (n_1188, A[3], n_316);
  xor g526 (n_223, n_1188, n_317);
  nand g527 (n_1189, A[3], n_316);
  nand g528 (n_1190, n_317, n_316);
  nand g529 (n_1191, A[3], n_317);
  nand g530 (n_139, n_1189, n_1190, n_1191);
  xor g531 (n_318, A[8], A[6]);
  and g532 (n_321, A[8], A[6]);
  xor g534 (n_320, Z[2], A[4]);
  nand g537 (n_1195, A[2], A[4]);
  xor g539 (n_1196, n_318, n_319);
  xor g540 (n_222, n_1196, n_320);
  nand g541 (n_1197, n_318, n_319);
  nand g542 (n_1198, n_320, n_319);
  nand g543 (n_1199, n_318, n_320);
  nand g544 (n_138, n_1197, n_1198, n_1199);
  xor g545 (n_1200, A[1], A[9]);
  xor g546 (n_323, n_1200, A[3]);
  nand g547 (n_1201, A[1], A[9]);
  nand g548 (n_1202, A[3], A[9]);
  nand g550 (n_326, n_1201, n_1202, n_1177);
  xor g551 (n_1204, A[7], A[5]);
  xor g552 (n_324, n_1204, n_321);
  nand g554 (n_1206, n_321, A[5]);
  nand g555 (n_1207, A[7], n_321);
  nand g556 (n_328, n_1186, n_1206, n_1207);
  xor g557 (n_1208, n_322, n_323);
  xor g558 (n_221, n_1208, n_324);
  nand g559 (n_1209, n_322, n_323);
  nand g560 (n_1210, n_324, n_323);
  nand g561 (n_1211, n_322, n_324);
  nand g562 (n_137, n_1209, n_1210, n_1211);
  xor g563 (n_325, A[10], A[8]);
  and g564 (n_330, A[10], A[8]);
  xor g565 (n_1212, A[4], A[2]);
  xor g566 (n_327, n_1212, A[6]);
  nand g568 (n_1214, A[6], A[2]);
  xor g571 (n_1216, A[0], n_325);
  xor g572 (n_329, n_1216, n_326);
  nand g573 (n_1217, A[0], n_325);
  nand g574 (n_1218, n_326, n_325);
  nand g575 (n_1219, A[0], n_326);
  nand g576 (n_334, n_1217, n_1218, n_1219);
  xor g577 (n_1220, n_327, n_328);
  xor g578 (n_220, n_1220, n_329);
  nand g579 (n_1221, n_327, n_328);
  nand g580 (n_1222, n_329, n_328);
  nand g581 (n_1223, n_327, n_329);
  nand g582 (n_136, n_1221, n_1222, n_1223);
  xor g584 (n_332, n_1200, A[5]);
  nand g586 (n_1226, A[5], A[9]);
  nand g588 (n_337, n_1201, n_1226, n_1179);
  xor g589 (n_1228, A[3], A[11]);
  xor g590 (n_333, n_1228, A[7]);
  nand g591 (n_1229, A[3], A[11]);
  nand g592 (n_1230, A[7], A[11]);
  nand g593 (n_1231, A[3], A[7]);
  nand g594 (n_338, n_1229, n_1230, n_1231);
  xor g595 (n_1232, n_330, n_331);
  xor g596 (n_335, n_1232, n_332);
  nand g597 (n_1233, n_330, n_331);
  nand g598 (n_1234, n_332, n_331);
  nand g599 (n_1235, n_330, n_332);
  nand g600 (n_342, n_1233, n_1234, n_1235);
  xor g601 (n_1236, n_333, n_334);
  xor g602 (n_219, n_1236, n_335);
  nand g603 (n_1237, n_333, n_334);
  nand g604 (n_1238, n_335, n_334);
  nand g605 (n_1239, n_333, n_335);
  nand g606 (n_135, n_1237, n_1238, n_1239);
  xor g607 (n_336, A[12], A[10]);
  and g608 (n_343, A[12], A[10]);
  xor g610 (n_339, n_315, A[8]);
  nand g612 (n_1242, A[8], A[4]);
  xor g616 (n_340, Z[2], n_336);
  nand g618 (n_1246, n_336, A[0]);
  nand g619 (n_1247, A[2], n_336);
  nand g620 (n_347, n_1181, n_1246, n_1247);
  xor g621 (n_1248, n_337, n_338);
  xor g622 (n_341, n_1248, n_339);
  nand g623 (n_1249, n_337, n_338);
  nand g624 (n_1250, n_339, n_338);
  nand g625 (n_1251, n_337, n_339);
  nand g626 (n_349, n_1249, n_1250, n_1251);
  xor g627 (n_1252, n_340, n_341);
  xor g628 (n_218, n_1252, n_342);
  nand g629 (n_1253, n_340, n_341);
  nand g630 (n_1254, n_342, n_341);
  nand g631 (n_1255, n_340, n_342);
  nand g632 (n_134, n_1253, n_1254, n_1255);
  xor g633 (n_1256, A[1], A[11]);
  xor g634 (n_346, n_1256, A[7]);
  nand g635 (n_1257, A[1], A[11]);
  nand g638 (n_352, n_1257, n_1230, n_1185);
  xor g639 (n_1260, A[5], A[13]);
  xor g640 (n_345, n_1260, A[3]);
  nand g641 (n_1261, A[5], A[13]);
  nand g642 (n_1262, A[3], A[13]);
  nand g644 (n_353, n_1261, n_1262, n_1178);
  xor g645 (n_1264, A[9], n_343);
  xor g646 (n_348, n_1264, n_344);
  nand g647 (n_1265, A[9], n_343);
  nand g648 (n_1266, n_344, n_343);
  nand g649 (n_1267, A[9], n_344);
  nand g650 (n_356, n_1265, n_1266, n_1267);
  xor g651 (n_1268, n_345, n_346);
  xor g652 (n_350, n_1268, n_347);
  nand g653 (n_1269, n_345, n_346);
  nand g654 (n_1270, n_347, n_346);
  nand g655 (n_1271, n_345, n_347);
  nand g656 (n_358, n_1269, n_1270, n_1271);
  xor g657 (n_1272, n_348, n_349);
  xor g658 (n_217, n_1272, n_350);
  nand g659 (n_1273, n_348, n_349);
  nand g660 (n_1274, n_350, n_349);
  nand g661 (n_1275, n_348, n_350);
  nand g662 (n_133, n_1273, n_1274, n_1275);
  xor g663 (n_351, A[14], A[12]);
  and g664 (n_360, A[14], A[12]);
  xor g665 (n_1276, A[8], A[0]);
  xor g666 (n_355, n_1276, A[6]);
  nand g667 (n_1277, A[8], A[0]);
  nand g668 (n_1278, A[6], A[0]);
  xor g671 (n_1280, A[10], A[4]);
  xor g672 (n_354, n_1280, A[2]);
  nand g673 (n_1281, A[10], A[4]);
  nand g675 (n_1283, A[10], A[2]);
  nand g676 (n_362, n_1281, n_1195, n_1283);
  xor g677 (n_1284, n_351, n_352);
  xor g678 (n_357, n_1284, n_353);
  nand g679 (n_1285, n_351, n_352);
  nand g680 (n_1286, n_353, n_352);
  nand g681 (n_1287, n_351, n_353);
  nand g682 (n_366, n_1285, n_1286, n_1287);
  xor g683 (n_1288, n_354, n_355);
  xor g684 (n_359, n_1288, n_356);
  nand g685 (n_1289, n_354, n_355);
  nand g686 (n_1290, n_356, n_355);
  nand g687 (n_1291, n_354, n_356);
  nand g688 (n_369, n_1289, n_1290, n_1291);
  xor g689 (n_1292, n_357, n_358);
  xor g690 (n_216, n_1292, n_359);
  nand g691 (n_1293, n_357, n_358);
  nand g692 (n_1294, n_359, n_358);
  nand g693 (n_1295, n_357, n_359);
  nand g694 (n_132, n_1293, n_1294, n_1295);
  xor g695 (n_1296, A[1], A[15]);
  xor g696 (n_363, n_1296, A[13]);
  nand g697 (n_1297, A[1], A[15]);
  nand g698 (n_1298, A[13], A[15]);
  nand g699 (n_1299, A[1], A[13]);
  nand g700 (n_371, n_1297, n_1298, n_1299);
  xor g701 (n_1300, A[9], A[7]);
  xor g702 (n_364, n_1300, A[11]);
  nand g703 (n_1301, A[9], A[7]);
  nand g705 (n_1303, A[9], A[11]);
  nand g706 (n_372, n_1301, n_1230, n_1303);
  xor g707 (n_1304, A[5], A[3]);
  xor g708 (n_365, n_1304, n_360);
  nand g710 (n_1306, n_360, A[3]);
  nand g711 (n_1307, A[5], n_360);
  nand g712 (n_375, n_1178, n_1306, n_1307);
  xor g713 (n_1308, n_361, n_362);
  xor g714 (n_367, n_1308, n_363);
  nand g715 (n_1309, n_361, n_362);
  nand g716 (n_1310, n_363, n_362);
  nand g717 (n_1311, n_361, n_363);
  nand g718 (n_377, n_1309, n_1310, n_1311);
  xor g719 (n_1312, n_364, n_365);
  xor g720 (n_368, n_1312, n_366);
  nand g721 (n_1313, n_364, n_365);
  nand g722 (n_1314, n_366, n_365);
  nand g723 (n_1315, n_364, n_366);
  nand g724 (n_379, n_1313, n_1314, n_1315);
  xor g725 (n_1316, n_367, n_368);
  xor g726 (n_215, n_1316, n_369);
  nand g727 (n_1317, n_367, n_368);
  nand g728 (n_1318, n_369, n_368);
  nand g729 (n_1319, n_367, n_369);
  nand g730 (n_131, n_1317, n_1318, n_1319);
  xor g731 (n_370, A[16], A[14]);
  and g732 (n_381, A[16], A[14]);
  xor g733 (n_1320, A[10], A[2]);
  xor g734 (n_374, n_1320, A[0]);
  nand g737 (n_1323, A[10], A[0]);
  nand g738 (n_382, n_1283, n_1181, n_1323);
  xor g739 (n_1324, A[8], A[12]);
  xor g740 (n_373, n_1324, A[6]);
  nand g741 (n_1325, A[8], A[12]);
  nand g742 (n_1326, A[6], A[12]);
  xor g745 (n_1328, A[4], n_370);
  xor g746 (n_376, n_1328, n_371);
  nand g747 (n_1329, A[4], n_370);
  nand g748 (n_1330, n_371, n_370);
  nand g749 (n_1331, A[4], n_371);
  nand g750 (n_387, n_1329, n_1330, n_1331);
  xor g751 (n_1332, n_372, n_373);
  xor g752 (n_378, n_1332, n_374);
  nand g753 (n_1333, n_372, n_373);
  nand g754 (n_1334, n_374, n_373);
  nand g755 (n_1335, n_372, n_374);
  nand g756 (n_389, n_1333, n_1334, n_1335);
  xor g757 (n_1336, n_375, n_376);
  xor g758 (n_380, n_1336, n_377);
  nand g759 (n_1337, n_375, n_376);
  nand g760 (n_1338, n_377, n_376);
  nand g761 (n_1339, n_375, n_377);
  nand g762 (n_391, n_1337, n_1338, n_1339);
  xor g763 (n_1340, n_378, n_379);
  xor g764 (n_214, n_1340, n_380);
  nand g765 (n_1341, n_378, n_379);
  nand g766 (n_1342, n_380, n_379);
  nand g767 (n_1343, n_378, n_380);
  nand g768 (n_130, n_1341, n_1342, n_1343);
  xor g769 (n_1344, A[1], A[17]);
  xor g770 (n_385, n_1344, A[15]);
  nand g771 (n_1345, A[1], A[17]);
  nand g772 (n_1346, A[15], A[17]);
  nand g774 (n_394, n_1345, n_1346, n_1297);
  xor g776 (n_386, n_1228, A[9]);
  nand g780 (n_396, n_1229, n_1303, n_1202);
  xor g781 (n_1352, A[13], A[7]);
  xor g782 (n_384, n_1352, A[5]);
  nand g783 (n_1353, A[13], A[7]);
  nand g786 (n_395, n_1353, n_1186, n_1261);
  xor g787 (n_1356, n_381, n_382);
  xor g788 (n_388, n_1356, n_383);
  nand g789 (n_1357, n_381, n_382);
  nand g790 (n_1358, n_383, n_382);
  nand g791 (n_1359, n_381, n_383);
  nand g792 (n_400, n_1357, n_1358, n_1359);
  xor g793 (n_1360, n_384, n_385);
  xor g794 (n_390, n_1360, n_386);
  nand g795 (n_1361, n_384, n_385);
  nand g796 (n_1362, n_386, n_385);
  nand g797 (n_1363, n_384, n_386);
  nand g798 (n_402, n_1361, n_1362, n_1363);
  xor g799 (n_1364, n_387, n_388);
  xor g800 (n_392, n_1364, n_389);
  nand g801 (n_1365, n_387, n_388);
  nand g802 (n_1366, n_389, n_388);
  nand g803 (n_1367, n_387, n_389);
  nand g804 (n_404, n_1365, n_1366, n_1367);
  xor g805 (n_1368, n_390, n_391);
  xor g806 (n_213, n_1368, n_392);
  nand g807 (n_1369, n_390, n_391);
  nand g808 (n_1370, n_392, n_391);
  nand g809 (n_1371, n_390, n_392);
  nand g810 (n_129, n_1369, n_1370, n_1371);
  xor g811 (n_393, A[18], A[16]);
  and g812 (n_406, A[18], A[16]);
  xor g813 (n_1372, A[12], A[4]);
  xor g814 (n_397, n_1372, A[2]);
  nand g815 (n_1373, A[12], A[4]);
  nand g817 (n_1375, A[12], A[2]);
  nand g818 (n_407, n_1373, n_1195, n_1375);
  xor g819 (n_1376, A[10], A[0]);
  xor g820 (n_398, n_1376, A[14]);
  nand g822 (n_1378, A[14], A[0]);
  nand g823 (n_1379, A[10], A[14]);
  nand g824 (n_408, n_1323, n_1378, n_1379);
  xor g826 (n_399, n_318, n_393);
  nand g828 (n_1382, n_393, A[6]);
  nand g829 (n_1383, A[8], n_393);
  xor g831 (n_1384, n_394, n_395);
  xor g832 (n_401, n_1384, n_396);
  nand g833 (n_1385, n_394, n_395);
  nand g834 (n_1386, n_396, n_395);
  nand g835 (n_1387, n_394, n_396);
  nand g836 (n_414, n_1385, n_1386, n_1387);
  xor g837 (n_1388, n_397, n_398);
  xor g838 (n_403, n_1388, n_399);
  nand g839 (n_1389, n_397, n_398);
  nand g840 (n_1390, n_399, n_398);
  nand g841 (n_1391, n_397, n_399);
  nand g842 (n_415, n_1389, n_1390, n_1391);
  xor g843 (n_1392, n_400, n_401);
  xor g844 (n_405, n_1392, n_402);
  nand g845 (n_1393, n_400, n_401);
  nand g846 (n_1394, n_402, n_401);
  nand g847 (n_1395, n_400, n_402);
  nand g848 (n_418, n_1393, n_1394, n_1395);
  xor g849 (n_1396, n_403, n_404);
  xor g850 (n_212, n_1396, n_405);
  nand g851 (n_1397, n_403, n_404);
  nand g852 (n_1398, n_405, n_404);
  nand g853 (n_1399, n_403, n_405);
  nand g854 (n_128, n_1397, n_1398, n_1399);
  xor g855 (n_1400, A[1], A[19]);
  xor g856 (n_410, n_1400, A[13]);
  nand g857 (n_1401, A[1], A[19]);
  nand g858 (n_1402, A[13], A[19]);
  nand g860 (n_420, n_1401, n_1402, n_1299);
  xor g862 (n_411, n_1304, A[17]);
  nand g864 (n_1406, A[17], A[3]);
  nand g865 (n_1407, A[5], A[17]);
  nand g866 (n_421, n_1178, n_1406, n_1407);
  xor g867 (n_1408, A[11], A[15]);
  xor g868 (n_409, n_1408, A[9]);
  nand g869 (n_1409, A[11], A[15]);
  nand g870 (n_1410, A[9], A[15]);
  nand g872 (n_422, n_1409, n_1410, n_1303);
  xor g873 (n_1412, A[7], n_406);
  xor g874 (n_413, n_1412, n_407);
  nand g875 (n_1413, A[7], n_406);
  nand g876 (n_1414, n_407, n_406);
  nand g877 (n_1415, A[7], n_407);
  nand g878 (n_426, n_1413, n_1414, n_1415);
  xor g879 (n_1416, n_408, n_409);
  xor g880 (n_416, n_1416, n_410);
  nand g881 (n_1417, n_408, n_409);
  nand g882 (n_1418, n_410, n_409);
  nand g883 (n_1419, n_408, n_410);
  nand g884 (n_428, n_1417, n_1418, n_1419);
  xor g885 (n_1420, n_411, n_412);
  xor g886 (n_417, n_1420, n_413);
  nand g887 (n_1421, n_411, n_412);
  nand g888 (n_1422, n_413, n_412);
  nand g889 (n_1423, n_411, n_413);
  nand g890 (n_430, n_1421, n_1422, n_1423);
  xor g891 (n_1424, n_414, n_415);
  xor g892 (n_419, n_1424, n_416);
  nand g893 (n_1425, n_414, n_415);
  nand g894 (n_1426, n_416, n_415);
  nand g895 (n_1427, n_414, n_416);
  nand g896 (n_432, n_1425, n_1426, n_1427);
  xor g897 (n_1428, n_417, n_418);
  xor g898 (n_211, n_1428, n_419);
  nand g899 (n_1429, n_417, n_418);
  nand g900 (n_1430, n_419, n_418);
  nand g901 (n_1431, n_417, n_419);
  nand g902 (n_127, n_1429, n_1430, n_1431);
  xor g903 (n_1432, A[20], A[18]);
  xor g904 (n_424, n_1432, A[14]);
  nand g905 (n_1433, A[20], A[18]);
  nand g906 (n_1434, A[14], A[18]);
  nand g907 (n_1435, A[20], A[14]);
  nand g908 (n_143, n_1433, n_1434, n_1435);
  xor g910 (n_425, n_315, A[12]);
  xor g915 (n_1440, A[2], A[16]);
  xor g916 (n_423, n_1440, A[10]);
  nand g917 (n_1441, A[2], A[16]);
  nand g918 (n_1442, A[10], A[16]);
  nand g920 (n_145, n_1441, n_1442, n_1283);
  xor g921 (n_1444, A[8], n_420);
  xor g922 (n_427, n_1444, n_421);
  nand g923 (n_1445, A[8], n_420);
  nand g924 (n_1446, n_421, n_420);
  nand g925 (n_1447, A[8], n_421);
  nand g926 (n_435, n_1445, n_1446, n_1447);
  xor g927 (n_1448, n_422, n_423);
  xor g928 (n_429, n_1448, n_424);
  nand g929 (n_1449, n_422, n_423);
  nand g930 (n_1450, n_424, n_423);
  nand g931 (n_1451, n_422, n_424);
  nand g932 (n_437, n_1449, n_1450, n_1451);
  xor g933 (n_1452, n_425, n_426);
  xor g934 (n_431, n_1452, n_427);
  nand g935 (n_1453, n_425, n_426);
  nand g936 (n_1454, n_427, n_426);
  nand g937 (n_1455, n_425, n_427);
  nand g938 (n_439, n_1453, n_1454, n_1455);
  xor g939 (n_1456, n_428, n_429);
  xor g940 (n_433, n_1456, n_430);
  nand g941 (n_1457, n_428, n_429);
  nand g942 (n_1458, n_430, n_429);
  nand g943 (n_1459, n_428, n_430);
  nand g944 (n_441, n_1457, n_1458, n_1459);
  xor g945 (n_1460, n_431, n_432);
  xor g946 (n_210, n_1460, n_433);
  nand g947 (n_1461, n_431, n_432);
  nand g948 (n_1462, n_433, n_432);
  nand g949 (n_1463, n_431, n_433);
  nand g950 (n_126, n_1461, n_1462, n_1463);
  xor g951 (n_1464, A[21], A[19]);
  xor g952 (n_147, n_1464, A[15]);
  nand g953 (n_1465, A[21], A[19]);
  nand g954 (n_1466, A[15], A[19]);
  nand g955 (n_1467, A[21], A[15]);
  nand g956 (n_443, n_1465, n_1466, n_1467);
  xor g958 (n_434, n_1204, A[13]);
  xor g963 (n_1472, A[3], A[17]);
  xor g964 (n_146, n_1472, A[11]);
  nand g966 (n_1474, A[11], A[17]);
  nand g968 (n_445, n_1406, n_1474, n_1229);
  xor g969 (n_1476, A[9], n_143);
  xor g970 (n_436, n_1476, n_144);
  nand g971 (n_1477, A[9], n_143);
  nand g972 (n_1478, n_144, n_143);
  nand g973 (n_1479, A[9], n_144);
  nand g974 (n_449, n_1477, n_1478, n_1479);
  xor g975 (n_1480, n_145, n_146);
  xor g976 (n_438, n_1480, n_147);
  nand g977 (n_1481, n_145, n_146);
  nand g978 (n_1482, n_147, n_146);
  nand g979 (n_1483, n_145, n_147);
  nand g980 (n_451, n_1481, n_1482, n_1483);
  xor g981 (n_1484, n_434, n_435);
  xor g982 (n_440, n_1484, n_436);
  nand g983 (n_1485, n_434, n_435);
  nand g984 (n_1486, n_436, n_435);
  nand g985 (n_1487, n_434, n_436);
  nand g986 (n_453, n_1485, n_1486, n_1487);
  xor g987 (n_1488, n_437, n_438);
  xor g988 (n_442, n_1488, n_439);
  nand g989 (n_1489, n_437, n_438);
  nand g990 (n_1490, n_439, n_438);
  nand g991 (n_1491, n_437, n_439);
  nand g992 (n_456, n_1489, n_1490, n_1491);
  xor g993 (n_1492, n_440, n_441);
  xor g994 (n_209, n_1492, n_442);
  nand g995 (n_1493, n_440, n_441);
  nand g996 (n_1494, n_442, n_441);
  nand g997 (n_1495, n_440, n_442);
  nand g998 (n_125, n_1493, n_1494, n_1495);
  xor g999 (n_1496, A[22], A[20]);
  xor g1000 (n_447, n_1496, A[16]);
  nand g1001 (n_1497, A[22], A[20]);
  nand g1002 (n_1498, A[16], A[20]);
  nand g1003 (n_1499, A[22], A[16]);
  nand g1004 (n_457, n_1497, n_1498, n_1499);
  xor g1006 (n_448, n_318, A[14]);
  nand g1008 (n_1502, A[14], A[6]);
  nand g1009 (n_1503, A[8], A[14]);
  xor g1011 (n_1504, A[4], A[18]);
  xor g1012 (n_446, n_1504, A[12]);
  nand g1013 (n_1505, A[4], A[18]);
  nand g1014 (n_1506, A[12], A[18]);
  nand g1016 (n_459, n_1505, n_1506, n_1373);
  xor g1017 (n_1508, A[10], n_443);
  xor g1018 (n_450, n_1508, n_395);
  nand g1019 (n_1509, A[10], n_443);
  nand g1020 (n_1510, n_395, n_443);
  nand g1021 (n_1511, A[10], n_395);
  nand g1022 (n_463, n_1509, n_1510, n_1511);
  xor g1023 (n_1512, n_445, n_446);
  xor g1024 (n_452, n_1512, n_447);
  nand g1025 (n_1513, n_445, n_446);
  nand g1026 (n_1514, n_447, n_446);
  nand g1027 (n_1515, n_445, n_447);
  nand g1028 (n_465, n_1513, n_1514, n_1515);
  xor g1029 (n_1516, n_448, n_449);
  xor g1030 (n_454, n_1516, n_450);
  nand g1031 (n_1517, n_448, n_449);
  nand g1032 (n_1518, n_450, n_449);
  nand g1033 (n_1519, n_448, n_450);
  nand g1034 (n_467, n_1517, n_1518, n_1519);
  xor g1035 (n_1520, n_451, n_452);
  xor g1036 (n_455, n_1520, n_453);
  nand g1037 (n_1521, n_451, n_452);
  nand g1038 (n_1522, n_453, n_452);
  nand g1039 (n_1523, n_451, n_453);
  nand g1040 (n_470, n_1521, n_1522, n_1523);
  xor g1041 (n_1524, n_454, n_455);
  xor g1042 (n_208, n_1524, n_456);
  nand g1043 (n_1525, n_454, n_455);
  nand g1044 (n_1526, n_456, n_455);
  nand g1045 (n_1527, n_454, n_456);
  nand g1046 (n_124, n_1525, n_1526, n_1527);
  xor g1047 (n_1528, A[23], A[21]);
  xor g1048 (n_461, n_1528, A[17]);
  nand g1049 (n_1529, A[23], A[21]);
  nand g1050 (n_1530, A[17], A[21]);
  nand g1051 (n_1531, A[23], A[17]);
  nand g1052 (n_471, n_1529, n_1530, n_1531);
  xor g1054 (n_462, n_1300, A[15]);
  nand g1056 (n_1534, A[15], A[7]);
  nand g1058 (n_472, n_1301, n_1534, n_1410);
  xor g1059 (n_1536, A[5], A[19]);
  xor g1060 (n_460, n_1536, A[13]);
  nand g1061 (n_1537, A[5], A[19]);
  nand g1064 (n_473, n_1537, n_1402, n_1261);
  xor g1065 (n_1540, A[11], n_457);
  xor g1066 (n_464, n_1540, n_458);
  nand g1067 (n_1541, A[11], n_457);
  nand g1068 (n_1542, n_458, n_457);
  nand g1069 (n_1543, A[11], n_458);
  nand g1070 (n_477, n_1541, n_1542, n_1543);
  xor g1071 (n_1544, n_459, n_460);
  xor g1072 (n_466, n_1544, n_461);
  nand g1073 (n_1545, n_459, n_460);
  nand g1074 (n_1546, n_461, n_460);
  nand g1075 (n_1547, n_459, n_461);
  nand g1076 (n_479, n_1545, n_1546, n_1547);
  xor g1077 (n_1548, n_462, n_463);
  xor g1078 (n_468, n_1548, n_464);
  nand g1079 (n_1549, n_462, n_463);
  nand g1080 (n_1550, n_464, n_463);
  nand g1081 (n_1551, n_462, n_464);
  nand g1082 (n_481, n_1549, n_1550, n_1551);
  xor g1083 (n_1552, n_465, n_466);
  xor g1084 (n_469, n_1552, n_467);
  nand g1085 (n_1553, n_465, n_466);
  nand g1086 (n_1554, n_467, n_466);
  nand g1087 (n_1555, n_465, n_467);
  nand g1088 (n_484, n_1553, n_1554, n_1555);
  xor g1089 (n_1556, n_468, n_469);
  xor g1090 (n_207, n_1556, n_470);
  nand g1091 (n_1557, n_468, n_469);
  nand g1092 (n_1558, n_470, n_469);
  nand g1093 (n_1559, n_468, n_470);
  nand g1094 (n_123, n_1557, n_1558, n_1559);
  xor g1095 (n_1560, A[24], A[22]);
  xor g1096 (n_475, n_1560, A[18]);
  nand g1097 (n_1561, A[24], A[22]);
  nand g1098 (n_1562, A[18], A[22]);
  nand g1099 (n_1563, A[24], A[18]);
  nand g1100 (n_485, n_1561, n_1562, n_1563);
  xor g1102 (n_476, n_325, A[16]);
  nand g1104 (n_1566, A[16], A[8]);
  xor g1107 (n_1568, A[6], A[20]);
  xor g1108 (n_474, n_1568, A[14]);
  nand g1109 (n_1569, A[6], A[20]);
  nand g1112 (n_487, n_1569, n_1435, n_1502);
  xor g1113 (n_1572, A[12], n_471);
  xor g1114 (n_478, n_1572, n_472);
  nand g1115 (n_1573, A[12], n_471);
  nand g1116 (n_1574, n_472, n_471);
  nand g1117 (n_1575, A[12], n_472);
  nand g1118 (n_491, n_1573, n_1574, n_1575);
  xor g1119 (n_1576, n_473, n_474);
  xor g1120 (n_480, n_1576, n_475);
  nand g1121 (n_1577, n_473, n_474);
  nand g1122 (n_1578, n_475, n_474);
  nand g1123 (n_1579, n_473, n_475);
  nand g1124 (n_493, n_1577, n_1578, n_1579);
  xor g1125 (n_1580, n_476, n_477);
  xor g1126 (n_482, n_1580, n_478);
  nand g1127 (n_1581, n_476, n_477);
  nand g1128 (n_1582, n_478, n_477);
  nand g1129 (n_1583, n_476, n_478);
  nand g1130 (n_495, n_1581, n_1582, n_1583);
  xor g1131 (n_1584, n_479, n_480);
  xor g1132 (n_483, n_1584, n_481);
  nand g1133 (n_1585, n_479, n_480);
  nand g1134 (n_1586, n_481, n_480);
  nand g1135 (n_1587, n_479, n_481);
  nand g1136 (n_498, n_1585, n_1586, n_1587);
  xor g1137 (n_1588, n_482, n_483);
  xor g1138 (n_206, n_1588, n_484);
  nand g1139 (n_1589, n_482, n_483);
  nand g1140 (n_1590, n_484, n_483);
  nand g1141 (n_1591, n_482, n_484);
  nand g1142 (n_122, n_1589, n_1590, n_1591);
  xor g1143 (n_1592, A[25], A[23]);
  xor g1144 (n_489, n_1592, A[19]);
  nand g1145 (n_1593, A[25], A[23]);
  nand g1146 (n_1594, A[19], A[23]);
  nand g1147 (n_1595, A[25], A[19]);
  nand g1148 (n_499, n_1593, n_1594, n_1595);
  xor g1149 (n_1596, A[11], A[9]);
  xor g1150 (n_490, n_1596, A[17]);
  nand g1152 (n_1598, A[17], A[9]);
  nand g1154 (n_500, n_1303, n_1598, n_1474);
  xor g1155 (n_1600, A[7], A[21]);
  xor g1156 (n_488, n_1600, A[15]);
  nand g1157 (n_1601, A[7], A[21]);
  nand g1160 (n_501, n_1601, n_1467, n_1534);
  xor g1161 (n_1604, A[13], n_485);
  xor g1162 (n_492, n_1604, n_486);
  nand g1163 (n_1605, A[13], n_485);
  nand g1164 (n_1606, n_486, n_485);
  nand g1165 (n_1607, A[13], n_486);
  nand g1166 (n_505, n_1605, n_1606, n_1607);
  xor g1167 (n_1608, n_487, n_488);
  xor g1168 (n_494, n_1608, n_489);
  nand g1169 (n_1609, n_487, n_488);
  nand g1170 (n_1610, n_489, n_488);
  nand g1171 (n_1611, n_487, n_489);
  nand g1172 (n_507, n_1609, n_1610, n_1611);
  xor g1173 (n_1612, n_490, n_491);
  xor g1174 (n_496, n_1612, n_492);
  nand g1175 (n_1613, n_490, n_491);
  nand g1176 (n_1614, n_492, n_491);
  nand g1177 (n_1615, n_490, n_492);
  nand g1178 (n_228, n_1613, n_1614, n_1615);
  xor g1179 (n_1616, n_493, n_494);
  xor g1180 (n_497, n_1616, n_495);
  nand g1181 (n_1617, n_493, n_494);
  nand g1182 (n_1618, n_495, n_494);
  nand g1183 (n_1619, n_493, n_495);
  nand g1184 (n_510, n_1617, n_1618, n_1619);
  xor g1185 (n_1620, n_496, n_497);
  xor g1186 (n_205, n_1620, n_498);
  nand g1187 (n_1621, n_496, n_497);
  nand g1188 (n_1622, n_498, n_497);
  nand g1189 (n_1623, n_496, n_498);
  nand g1190 (n_121, n_1621, n_1622, n_1623);
  xor g1191 (n_1624, A[26], A[24]);
  xor g1192 (n_503, n_1624, A[20]);
  nand g1193 (n_1625, A[26], A[24]);
  nand g1194 (n_1626, A[20], A[24]);
  nand g1195 (n_1627, A[26], A[20]);
  nand g1196 (n_511, n_1625, n_1626, n_1627);
  xor g1198 (n_504, n_336, A[18]);
  nand g1200 (n_1630, A[18], A[10]);
  xor g1203 (n_1632, A[8], A[22]);
  xor g1204 (n_502, n_1632, A[16]);
  nand g1205 (n_1633, A[8], A[22]);
  nand g1208 (n_513, n_1633, n_1499, n_1566);
  xor g1209 (n_1636, A[14], n_499);
  xor g1210 (n_506, n_1636, n_500);
  nand g1211 (n_1637, A[14], n_499);
  nand g1212 (n_1638, n_500, n_499);
  nand g1213 (n_1639, A[14], n_500);
  nand g1214 (n_517, n_1637, n_1638, n_1639);
  xor g1215 (n_1640, n_501, n_502);
  xor g1216 (n_227, n_1640, n_503);
  nand g1217 (n_1641, n_501, n_502);
  nand g1218 (n_1642, n_503, n_502);
  nand g1219 (n_1643, n_501, n_503);
  nand g1220 (n_519, n_1641, n_1642, n_1643);
  xor g1221 (n_1644, n_504, n_505);
  xor g1222 (n_508, n_1644, n_506);
  nand g1223 (n_1645, n_504, n_505);
  nand g1224 (n_1646, n_506, n_505);
  nand g1225 (n_1647, n_504, n_506);
  nand g1226 (n_521, n_1645, n_1646, n_1647);
  xor g1227 (n_1648, n_507, n_227);
  xor g1228 (n_509, n_1648, n_228);
  nand g1229 (n_1649, n_507, n_227);
  nand g1230 (n_1650, n_228, n_227);
  nand g1231 (n_1651, n_507, n_228);
  nand g1232 (n_524, n_1649, n_1650, n_1651);
  xor g1233 (n_1652, n_508, n_509);
  xor g1234 (n_204, n_1652, n_510);
  nand g1235 (n_1653, n_508, n_509);
  nand g1236 (n_1654, n_510, n_509);
  nand g1237 (n_1655, n_508, n_510);
  nand g1238 (n_120, n_1653, n_1654, n_1655);
  xor g1239 (n_1656, A[27], A[25]);
  xor g1240 (n_515, n_1656, A[21]);
  nand g1241 (n_1657, A[27], A[25]);
  nand g1242 (n_1658, A[21], A[25]);
  nand g1243 (n_1659, A[27], A[21]);
  nand g1244 (n_525, n_1657, n_1658, n_1659);
  xor g1245 (n_1660, A[13], A[11]);
  xor g1246 (n_516, n_1660, A[19]);
  nand g1247 (n_1661, A[13], A[11]);
  nand g1248 (n_1662, A[19], A[11]);
  nand g1250 (n_526, n_1661, n_1662, n_1402);
  xor g1251 (n_1664, A[9], A[23]);
  xor g1252 (n_514, n_1664, A[17]);
  nand g1253 (n_1665, A[9], A[23]);
  nand g1256 (n_527, n_1665, n_1531, n_1598);
  xor g1257 (n_1668, A[15], n_511);
  xor g1258 (n_518, n_1668, n_512);
  nand g1259 (n_1669, A[15], n_511);
  nand g1260 (n_1670, n_512, n_511);
  nand g1261 (n_1671, A[15], n_512);
  nand g1262 (n_531, n_1669, n_1670, n_1671);
  xor g1263 (n_1672, n_513, n_514);
  xor g1264 (n_520, n_1672, n_515);
  nand g1265 (n_1673, n_513, n_514);
  nand g1266 (n_1674, n_515, n_514);
  nand g1267 (n_1675, n_513, n_515);
  nand g1268 (n_533, n_1673, n_1674, n_1675);
  xor g1269 (n_1676, n_516, n_517);
  xor g1270 (n_522, n_1676, n_518);
  nand g1271 (n_1677, n_516, n_517);
  nand g1272 (n_1678, n_518, n_517);
  nand g1273 (n_1679, n_516, n_518);
  nand g1274 (n_535, n_1677, n_1678, n_1679);
  xor g1275 (n_1680, n_519, n_520);
  xor g1276 (n_523, n_1680, n_521);
  nand g1277 (n_1681, n_519, n_520);
  nand g1278 (n_1682, n_521, n_520);
  nand g1279 (n_1683, n_519, n_521);
  nand g1280 (n_538, n_1681, n_1682, n_1683);
  xor g1281 (n_1684, n_522, n_523);
  xor g1282 (n_203, n_1684, n_524);
  nand g1283 (n_1685, n_522, n_523);
  nand g1284 (n_1686, n_524, n_523);
  nand g1285 (n_1687, n_522, n_524);
  nand g1286 (n_119, n_1685, n_1686, n_1687);
  xor g1287 (n_1688, A[28], A[26]);
  xor g1288 (n_529, n_1688, A[22]);
  nand g1289 (n_1689, A[28], A[26]);
  nand g1290 (n_1690, A[22], A[26]);
  nand g1291 (n_1691, A[28], A[22]);
  nand g1292 (n_539, n_1689, n_1690, n_1691);
  xor g1294 (n_530, n_351, A[20]);
  nand g1296 (n_1694, A[20], A[12]);
  xor g1299 (n_1696, A[10], A[24]);
  xor g1300 (n_528, n_1696, A[18]);
  nand g1301 (n_1697, A[10], A[24]);
  nand g1304 (n_541, n_1697, n_1563, n_1630);
  xor g1305 (n_1700, A[16], n_525);
  xor g1306 (n_532, n_1700, n_526);
  nand g1307 (n_1701, A[16], n_525);
  nand g1308 (n_1702, n_526, n_525);
  nand g1309 (n_1703, A[16], n_526);
  nand g1310 (n_545, n_1701, n_1702, n_1703);
  xor g1311 (n_1704, n_527, n_528);
  xor g1312 (n_534, n_1704, n_529);
  nand g1313 (n_1705, n_527, n_528);
  nand g1314 (n_1706, n_529, n_528);
  nand g1315 (n_1707, n_527, n_529);
  nand g1316 (n_547, n_1705, n_1706, n_1707);
  xor g1317 (n_1708, n_530, n_531);
  xor g1318 (n_536, n_1708, n_532);
  nand g1319 (n_1709, n_530, n_531);
  nand g1320 (n_1710, n_532, n_531);
  nand g1321 (n_1711, n_530, n_532);
  nand g1322 (n_549, n_1709, n_1710, n_1711);
  xor g1323 (n_1712, n_533, n_534);
  xor g1324 (n_537, n_1712, n_535);
  nand g1325 (n_1713, n_533, n_534);
  nand g1326 (n_1714, n_535, n_534);
  nand g1327 (n_1715, n_533, n_535);
  nand g1328 (n_552, n_1713, n_1714, n_1715);
  xor g1329 (n_1716, n_536, n_537);
  xor g1330 (n_202, n_1716, n_538);
  nand g1331 (n_1717, n_536, n_537);
  nand g1332 (n_1718, n_538, n_537);
  nand g1333 (n_1719, n_536, n_538);
  nand g1334 (n_118, n_1717, n_1718, n_1719);
  xor g1335 (n_1720, A[29], A[27]);
  xor g1336 (n_543, n_1720, A[23]);
  nand g1337 (n_1721, A[29], A[27]);
  nand g1338 (n_1722, A[23], A[27]);
  nand g1339 (n_1723, A[29], A[23]);
  nand g1340 (n_553, n_1721, n_1722, n_1723);
  xor g1341 (n_1724, A[15], A[13]);
  xor g1342 (n_544, n_1724, A[21]);
  nand g1344 (n_1726, A[21], A[13]);
  nand g1346 (n_554, n_1298, n_1726, n_1467);
  xor g1347 (n_1728, A[11], A[25]);
  xor g1348 (n_542, n_1728, A[19]);
  nand g1349 (n_1729, A[11], A[25]);
  nand g1352 (n_555, n_1729, n_1595, n_1662);
  xor g1353 (n_1732, A[17], n_539);
  xor g1354 (n_546, n_1732, n_540);
  nand g1355 (n_1733, A[17], n_539);
  nand g1356 (n_1734, n_540, n_539);
  nand g1357 (n_1735, A[17], n_540);
  nand g1358 (n_559, n_1733, n_1734, n_1735);
  xor g1359 (n_1736, n_541, n_542);
  xor g1360 (n_548, n_1736, n_543);
  nand g1361 (n_1737, n_541, n_542);
  nand g1362 (n_1738, n_543, n_542);
  nand g1363 (n_1739, n_541, n_543);
  nand g1364 (n_561, n_1737, n_1738, n_1739);
  xor g1365 (n_1740, n_544, n_545);
  xor g1366 (n_550, n_1740, n_546);
  nand g1367 (n_1741, n_544, n_545);
  nand g1368 (n_1742, n_546, n_545);
  nand g1369 (n_1743, n_544, n_546);
  nand g1370 (n_563, n_1741, n_1742, n_1743);
  xor g1371 (n_1744, n_547, n_548);
  xor g1372 (n_551, n_1744, n_549);
  nand g1373 (n_1745, n_547, n_548);
  nand g1374 (n_1746, n_549, n_548);
  nand g1375 (n_1747, n_547, n_549);
  nand g1376 (n_566, n_1745, n_1746, n_1747);
  xor g1377 (n_1748, n_550, n_551);
  xor g1378 (n_201, n_1748, n_552);
  nand g1379 (n_1749, n_550, n_551);
  nand g1380 (n_1750, n_552, n_551);
  nand g1381 (n_1751, n_550, n_552);
  nand g1382 (n_117, n_1749, n_1750, n_1751);
  xor g1383 (n_1752, A[30], A[28]);
  xor g1384 (n_557, n_1752, A[24]);
  nand g1385 (n_1753, A[30], A[28]);
  nand g1386 (n_1754, A[24], A[28]);
  nand g1387 (n_1755, A[30], A[24]);
  nand g1388 (n_567, n_1753, n_1754, n_1755);
  xor g1390 (n_558, n_370, A[22]);
  nand g1392 (n_1758, A[22], A[14]);
  xor g1395 (n_1760, A[12], A[26]);
  xor g1396 (n_556, n_1760, A[20]);
  nand g1397 (n_1761, A[12], A[26]);
  nand g1400 (n_569, n_1761, n_1627, n_1694);
  xor g1401 (n_1764, A[18], n_553);
  xor g1402 (n_560, n_1764, n_554);
  nand g1403 (n_1765, A[18], n_553);
  nand g1404 (n_1766, n_554, n_553);
  nand g1405 (n_1767, A[18], n_554);
  nand g1406 (n_573, n_1765, n_1766, n_1767);
  xor g1407 (n_1768, n_555, n_556);
  xor g1408 (n_562, n_1768, n_557);
  nand g1409 (n_1769, n_555, n_556);
  nand g1410 (n_1770, n_557, n_556);
  nand g1411 (n_1771, n_555, n_557);
  nand g1412 (n_575, n_1769, n_1770, n_1771);
  xor g1413 (n_1772, n_558, n_559);
  xor g1414 (n_564, n_1772, n_560);
  nand g1415 (n_1773, n_558, n_559);
  nand g1416 (n_1774, n_560, n_559);
  nand g1417 (n_1775, n_558, n_560);
  nand g1418 (n_577, n_1773, n_1774, n_1775);
  xor g1419 (n_1776, n_561, n_562);
  xor g1420 (n_565, n_1776, n_563);
  nand g1421 (n_1777, n_561, n_562);
  nand g1422 (n_1778, n_563, n_562);
  nand g1423 (n_1779, n_561, n_563);
  nand g1424 (n_580, n_1777, n_1778, n_1779);
  xor g1425 (n_1780, n_564, n_565);
  xor g1426 (n_200, n_1780, n_566);
  nand g1427 (n_1781, n_564, n_565);
  nand g1428 (n_1782, n_566, n_565);
  nand g1429 (n_1783, n_564, n_566);
  nand g1430 (n_116, n_1781, n_1782, n_1783);
  xor g1431 (n_1784, A[31], A[29]);
  xor g1432 (n_571, n_1784, A[25]);
  nand g1433 (n_1785, A[31], A[29]);
  nand g1434 (n_1786, A[25], A[29]);
  nand g1435 (n_1787, A[31], A[25]);
  nand g1436 (n_581, n_1785, n_1786, n_1787);
  xor g1437 (n_1788, A[17], A[15]);
  xor g1438 (n_572, n_1788, A[23]);
  nand g1440 (n_1790, A[23], A[15]);
  nand g1442 (n_582, n_1346, n_1790, n_1531);
  xor g1443 (n_1792, A[13], A[27]);
  xor g1444 (n_570, n_1792, A[21]);
  nand g1445 (n_1793, A[13], A[27]);
  nand g1448 (n_583, n_1793, n_1659, n_1726);
  xor g1449 (n_1796, A[19], n_567);
  xor g1450 (n_574, n_1796, n_568);
  nand g1451 (n_1797, A[19], n_567);
  nand g1452 (n_1798, n_568, n_567);
  nand g1453 (n_1799, A[19], n_568);
  nand g1454 (n_587, n_1797, n_1798, n_1799);
  xor g1455 (n_1800, n_569, n_570);
  xor g1456 (n_576, n_1800, n_571);
  nand g1457 (n_1801, n_569, n_570);
  nand g1458 (n_1802, n_571, n_570);
  nand g1459 (n_1803, n_569, n_571);
  nand g1460 (n_589, n_1801, n_1802, n_1803);
  xor g1461 (n_1804, n_572, n_573);
  xor g1462 (n_578, n_1804, n_574);
  nand g1463 (n_1805, n_572, n_573);
  nand g1464 (n_1806, n_574, n_573);
  nand g1465 (n_1807, n_572, n_574);
  nand g1466 (n_591, n_1805, n_1806, n_1807);
  xor g1467 (n_1808, n_575, n_576);
  xor g1468 (n_579, n_1808, n_577);
  nand g1469 (n_1809, n_575, n_576);
  nand g1470 (n_1810, n_577, n_576);
  nand g1471 (n_1811, n_575, n_577);
  nand g1472 (n_594, n_1809, n_1810, n_1811);
  xor g1473 (n_1812, n_578, n_579);
  xor g1474 (n_199, n_1812, n_580);
  nand g1475 (n_1813, n_578, n_579);
  nand g1476 (n_1814, n_580, n_579);
  nand g1477 (n_1815, n_578, n_580);
  nand g1478 (n_115, n_1813, n_1814, n_1815);
  xor g1479 (n_1816, A[32], A[30]);
  xor g1480 (n_585, n_1816, A[26]);
  nand g1481 (n_1817, A[32], A[30]);
  nand g1482 (n_1818, A[26], A[30]);
  nand g1483 (n_1819, A[32], A[26]);
  nand g1484 (n_595, n_1817, n_1818, n_1819);
  xor g1486 (n_586, n_393, A[24]);
  nand g1488 (n_1822, A[24], A[16]);
  xor g1491 (n_1824, A[14], A[28]);
  xor g1492 (n_584, n_1824, A[22]);
  nand g1493 (n_1825, A[14], A[28]);
  nand g1496 (n_597, n_1825, n_1691, n_1758);
  xor g1497 (n_1828, A[20], n_581);
  xor g1498 (n_588, n_1828, n_582);
  nand g1499 (n_1829, A[20], n_581);
  nand g1500 (n_1830, n_582, n_581);
  nand g1501 (n_1831, A[20], n_582);
  nand g1502 (n_601, n_1829, n_1830, n_1831);
  xor g1503 (n_1832, n_583, n_584);
  xor g1504 (n_590, n_1832, n_585);
  nand g1505 (n_1833, n_583, n_584);
  nand g1506 (n_1834, n_585, n_584);
  nand g1507 (n_1835, n_583, n_585);
  nand g1508 (n_603, n_1833, n_1834, n_1835);
  xor g1509 (n_1836, n_586, n_587);
  xor g1510 (n_592, n_1836, n_588);
  nand g1511 (n_1837, n_586, n_587);
  nand g1512 (n_1838, n_588, n_587);
  nand g1513 (n_1839, n_586, n_588);
  nand g1514 (n_605, n_1837, n_1838, n_1839);
  xor g1515 (n_1840, n_589, n_590);
  xor g1516 (n_593, n_1840, n_591);
  nand g1517 (n_1841, n_589, n_590);
  nand g1518 (n_1842, n_591, n_590);
  nand g1519 (n_1843, n_589, n_591);
  nand g1520 (n_608, n_1841, n_1842, n_1843);
  xor g1521 (n_1844, n_592, n_593);
  xor g1522 (n_198, n_1844, n_594);
  nand g1523 (n_1845, n_592, n_593);
  nand g1524 (n_1846, n_594, n_593);
  nand g1525 (n_1847, n_592, n_594);
  nand g1526 (n_114, n_1845, n_1846, n_1847);
  xor g1527 (n_1848, A[33], A[31]);
  xor g1528 (n_599, n_1848, A[27]);
  nand g1529 (n_1849, A[33], A[31]);
  nand g1530 (n_1850, A[27], A[31]);
  nand g1531 (n_1851, A[33], A[27]);
  nand g1532 (n_609, n_1849, n_1850, n_1851);
  xor g1533 (n_1852, A[19], A[17]);
  xor g1534 (n_600, n_1852, A[25]);
  nand g1535 (n_1853, A[19], A[17]);
  nand g1536 (n_1854, A[25], A[17]);
  nand g1538 (n_610, n_1853, n_1854, n_1595);
  xor g1539 (n_1856, A[15], A[29]);
  xor g1540 (n_598, n_1856, A[23]);
  nand g1541 (n_1857, A[15], A[29]);
  nand g1544 (n_611, n_1857, n_1723, n_1790);
  xor g1545 (n_1860, A[21], n_595);
  xor g1546 (n_602, n_1860, n_596);
  nand g1547 (n_1861, A[21], n_595);
  nand g1548 (n_1862, n_596, n_595);
  nand g1549 (n_1863, A[21], n_596);
  nand g1550 (n_615, n_1861, n_1862, n_1863);
  xor g1551 (n_1864, n_597, n_598);
  xor g1552 (n_604, n_1864, n_599);
  nand g1553 (n_1865, n_597, n_598);
  nand g1554 (n_1866, n_599, n_598);
  nand g1555 (n_1867, n_597, n_599);
  nand g1556 (n_617, n_1865, n_1866, n_1867);
  xor g1557 (n_1868, n_600, n_601);
  xor g1558 (n_606, n_1868, n_602);
  nand g1559 (n_1869, n_600, n_601);
  nand g1560 (n_1870, n_602, n_601);
  nand g1561 (n_1871, n_600, n_602);
  nand g1562 (n_619, n_1869, n_1870, n_1871);
  xor g1563 (n_1872, n_603, n_604);
  xor g1564 (n_607, n_1872, n_605);
  nand g1565 (n_1873, n_603, n_604);
  nand g1566 (n_1874, n_605, n_604);
  nand g1567 (n_1875, n_603, n_605);
  nand g1568 (n_622, n_1873, n_1874, n_1875);
  xor g1569 (n_1876, n_606, n_607);
  xor g1570 (n_197, n_1876, n_608);
  nand g1571 (n_1877, n_606, n_607);
  nand g1572 (n_1878, n_608, n_607);
  nand g1573 (n_1879, n_606, n_608);
  nand g1574 (n_113, n_1877, n_1878, n_1879);
  xor g1575 (n_1880, A[34], A[32]);
  xor g1576 (n_613, n_1880, A[28]);
  nand g1577 (n_1881, A[34], A[32]);
  nand g1578 (n_1882, A[28], A[32]);
  nand g1579 (n_1883, A[34], A[28]);
  nand g1580 (n_623, n_1881, n_1882, n_1883);
  xor g1582 (n_614, n_1432, A[26]);
  nand g1584 (n_1886, A[26], A[18]);
  nand g1586 (n_624, n_1433, n_1886, n_1627);
  xor g1587 (n_1888, A[16], A[30]);
  xor g1588 (n_612, n_1888, A[24]);
  nand g1589 (n_1889, A[16], A[30]);
  nand g1592 (n_625, n_1889, n_1755, n_1822);
  xor g1593 (n_1892, A[22], n_609);
  xor g1594 (n_616, n_1892, n_610);
  nand g1595 (n_1893, A[22], n_609);
  nand g1596 (n_1894, n_610, n_609);
  nand g1597 (n_1895, A[22], n_610);
  nand g1598 (n_629, n_1893, n_1894, n_1895);
  xor g1599 (n_1896, n_611, n_612);
  xor g1600 (n_618, n_1896, n_613);
  nand g1601 (n_1897, n_611, n_612);
  nand g1602 (n_1898, n_613, n_612);
  nand g1603 (n_1899, n_611, n_613);
  nand g1604 (n_631, n_1897, n_1898, n_1899);
  xor g1605 (n_1900, n_614, n_615);
  xor g1606 (n_620, n_1900, n_616);
  nand g1607 (n_1901, n_614, n_615);
  nand g1608 (n_1902, n_616, n_615);
  nand g1609 (n_1903, n_614, n_616);
  nand g1610 (n_633, n_1901, n_1902, n_1903);
  xor g1611 (n_1904, n_617, n_618);
  xor g1612 (n_621, n_1904, n_619);
  nand g1613 (n_1905, n_617, n_618);
  nand g1614 (n_1906, n_619, n_618);
  nand g1615 (n_1907, n_617, n_619);
  nand g1616 (n_636, n_1905, n_1906, n_1907);
  xor g1617 (n_1908, n_620, n_621);
  xor g1618 (n_196, n_1908, n_622);
  nand g1619 (n_1909, n_620, n_621);
  nand g1620 (n_1910, n_622, n_621);
  nand g1621 (n_1911, n_620, n_622);
  nand g1622 (n_112, n_1909, n_1910, n_1911);
  xor g1623 (n_1912, A[35], A[33]);
  xor g1624 (n_627, n_1912, A[29]);
  nand g1625 (n_1913, A[35], A[33]);
  nand g1626 (n_1914, A[29], A[33]);
  nand g1627 (n_1915, A[35], A[29]);
  nand g1628 (n_637, n_1913, n_1914, n_1915);
  xor g1630 (n_628, n_1464, A[27]);
  nand g1632 (n_1918, A[27], A[19]);
  nand g1634 (n_638, n_1465, n_1918, n_1659);
  xor g1635 (n_1920, A[17], A[31]);
  xor g1636 (n_626, n_1920, A[25]);
  nand g1637 (n_1921, A[17], A[31]);
  nand g1640 (n_639, n_1921, n_1787, n_1854);
  xor g1641 (n_1924, A[23], n_623);
  xor g1642 (n_630, n_1924, n_624);
  nand g1643 (n_1925, A[23], n_623);
  nand g1644 (n_1926, n_624, n_623);
  nand g1645 (n_1927, A[23], n_624);
  nand g1646 (n_643, n_1925, n_1926, n_1927);
  xor g1647 (n_1928, n_625, n_626);
  xor g1648 (n_632, n_1928, n_627);
  nand g1649 (n_1929, n_625, n_626);
  nand g1650 (n_1930, n_627, n_626);
  nand g1651 (n_1931, n_625, n_627);
  nand g1652 (n_645, n_1929, n_1930, n_1931);
  xor g1653 (n_1932, n_628, n_629);
  xor g1654 (n_634, n_1932, n_630);
  nand g1655 (n_1933, n_628, n_629);
  nand g1656 (n_1934, n_630, n_629);
  nand g1657 (n_1935, n_628, n_630);
  nand g1658 (n_647, n_1933, n_1934, n_1935);
  xor g1659 (n_1936, n_631, n_632);
  xor g1660 (n_635, n_1936, n_633);
  nand g1661 (n_1937, n_631, n_632);
  nand g1662 (n_1938, n_633, n_632);
  nand g1663 (n_1939, n_631, n_633);
  nand g1664 (n_650, n_1937, n_1938, n_1939);
  xor g1665 (n_1940, n_634, n_635);
  xor g1666 (n_195, n_1940, n_636);
  nand g1667 (n_1941, n_634, n_635);
  nand g1668 (n_1942, n_636, n_635);
  nand g1669 (n_1943, n_634, n_636);
  nand g1670 (n_111, n_1941, n_1942, n_1943);
  xor g1671 (n_1944, A[36], A[34]);
  xor g1672 (n_641, n_1944, A[30]);
  nand g1673 (n_1945, A[36], A[34]);
  nand g1674 (n_1946, A[30], A[34]);
  nand g1675 (n_1947, A[36], A[30]);
  nand g1676 (n_651, n_1945, n_1946, n_1947);
  xor g1678 (n_642, n_1496, A[28]);
  nand g1680 (n_1950, A[28], A[20]);
  nand g1682 (n_652, n_1497, n_1950, n_1691);
  xor g1683 (n_1952, A[18], A[32]);
  xor g1684 (n_640, n_1952, A[26]);
  nand g1685 (n_1953, A[18], A[32]);
  nand g1688 (n_653, n_1953, n_1819, n_1886);
  xor g1689 (n_1956, A[24], n_637);
  xor g1690 (n_644, n_1956, n_638);
  nand g1691 (n_1957, A[24], n_637);
  nand g1692 (n_1958, n_638, n_637);
  nand g1693 (n_1959, A[24], n_638);
  nand g1694 (n_657, n_1957, n_1958, n_1959);
  xor g1695 (n_1960, n_639, n_640);
  xor g1696 (n_646, n_1960, n_641);
  nand g1697 (n_1961, n_639, n_640);
  nand g1698 (n_1962, n_641, n_640);
  nand g1699 (n_1963, n_639, n_641);
  nand g1700 (n_659, n_1961, n_1962, n_1963);
  xor g1701 (n_1964, n_642, n_643);
  xor g1702 (n_648, n_1964, n_644);
  nand g1703 (n_1965, n_642, n_643);
  nand g1704 (n_1966, n_644, n_643);
  nand g1705 (n_1967, n_642, n_644);
  nand g1706 (n_661, n_1965, n_1966, n_1967);
  xor g1707 (n_1968, n_645, n_646);
  xor g1708 (n_649, n_1968, n_647);
  nand g1709 (n_1969, n_645, n_646);
  nand g1710 (n_1970, n_647, n_646);
  nand g1711 (n_1971, n_645, n_647);
  nand g1712 (n_664, n_1969, n_1970, n_1971);
  xor g1713 (n_1972, n_648, n_649);
  xor g1714 (n_194, n_1972, n_650);
  nand g1715 (n_1973, n_648, n_649);
  nand g1716 (n_1974, n_650, n_649);
  nand g1717 (n_1975, n_648, n_650);
  nand g1718 (n_110, n_1973, n_1974, n_1975);
  xor g1719 (n_1976, A[37], A[35]);
  xor g1720 (n_655, n_1976, A[31]);
  nand g1721 (n_1977, A[37], A[35]);
  nand g1722 (n_1978, A[31], A[35]);
  nand g1723 (n_1979, A[37], A[31]);
  nand g1724 (n_665, n_1977, n_1978, n_1979);
  xor g1726 (n_656, n_1528, A[29]);
  nand g1728 (n_1982, A[29], A[21]);
  nand g1730 (n_666, n_1529, n_1982, n_1723);
  xor g1731 (n_1984, A[19], A[33]);
  xor g1732 (n_654, n_1984, A[27]);
  nand g1733 (n_1985, A[19], A[33]);
  nand g1736 (n_667, n_1985, n_1851, n_1918);
  xor g1737 (n_1988, A[25], n_651);
  xor g1738 (n_658, n_1988, n_652);
  nand g1739 (n_1989, A[25], n_651);
  nand g1740 (n_1990, n_652, n_651);
  nand g1741 (n_1991, A[25], n_652);
  nand g1742 (n_671, n_1989, n_1990, n_1991);
  xor g1743 (n_1992, n_653, n_654);
  xor g1744 (n_660, n_1992, n_655);
  nand g1745 (n_1993, n_653, n_654);
  nand g1746 (n_1994, n_655, n_654);
  nand g1747 (n_1995, n_653, n_655);
  nand g1748 (n_673, n_1993, n_1994, n_1995);
  xor g1749 (n_1996, n_656, n_657);
  xor g1750 (n_662, n_1996, n_658);
  nand g1751 (n_1997, n_656, n_657);
  nand g1752 (n_1998, n_658, n_657);
  nand g1753 (n_1999, n_656, n_658);
  nand g1754 (n_675, n_1997, n_1998, n_1999);
  xor g1755 (n_2000, n_659, n_660);
  xor g1756 (n_663, n_2000, n_661);
  nand g1757 (n_2001, n_659, n_660);
  nand g1758 (n_2002, n_661, n_660);
  nand g1759 (n_2003, n_659, n_661);
  nand g1760 (n_678, n_2001, n_2002, n_2003);
  xor g1761 (n_2004, n_662, n_663);
  xor g1762 (n_193, n_2004, n_664);
  nand g1763 (n_2005, n_662, n_663);
  nand g1764 (n_2006, n_664, n_663);
  nand g1765 (n_2007, n_662, n_664);
  nand g1766 (n_109, n_2005, n_2006, n_2007);
  xor g1767 (n_2008, A[38], A[36]);
  xor g1768 (n_669, n_2008, A[32]);
  nand g1769 (n_2009, A[38], A[36]);
  nand g1770 (n_2010, A[32], A[36]);
  nand g1771 (n_2011, A[38], A[32]);
  nand g1772 (n_679, n_2009, n_2010, n_2011);
  xor g1774 (n_670, n_1560, A[30]);
  nand g1776 (n_2014, A[30], A[22]);
  nand g1778 (n_680, n_1561, n_2014, n_1755);
  xor g1779 (n_2016, A[20], A[34]);
  xor g1780 (n_668, n_2016, A[28]);
  nand g1781 (n_2017, A[20], A[34]);
  nand g1784 (n_681, n_2017, n_1883, n_1950);
  xor g1785 (n_2020, A[26], n_665);
  xor g1786 (n_672, n_2020, n_666);
  nand g1787 (n_2021, A[26], n_665);
  nand g1788 (n_2022, n_666, n_665);
  nand g1789 (n_2023, A[26], n_666);
  nand g1790 (n_685, n_2021, n_2022, n_2023);
  xor g1791 (n_2024, n_667, n_668);
  xor g1792 (n_674, n_2024, n_669);
  nand g1793 (n_2025, n_667, n_668);
  nand g1794 (n_2026, n_669, n_668);
  nand g1795 (n_2027, n_667, n_669);
  nand g1796 (n_687, n_2025, n_2026, n_2027);
  xor g1797 (n_2028, n_670, n_671);
  xor g1798 (n_676, n_2028, n_672);
  nand g1799 (n_2029, n_670, n_671);
  nand g1800 (n_2030, n_672, n_671);
  nand g1801 (n_2031, n_670, n_672);
  nand g1802 (n_689, n_2029, n_2030, n_2031);
  xor g1803 (n_2032, n_673, n_674);
  xor g1804 (n_677, n_2032, n_675);
  nand g1805 (n_2033, n_673, n_674);
  nand g1806 (n_2034, n_675, n_674);
  nand g1807 (n_2035, n_673, n_675);
  nand g1808 (n_692, n_2033, n_2034, n_2035);
  xor g1809 (n_2036, n_676, n_677);
  xor g1810 (n_192, n_2036, n_678);
  nand g1811 (n_2037, n_676, n_677);
  nand g1812 (n_2038, n_678, n_677);
  nand g1813 (n_2039, n_676, n_678);
  nand g1814 (n_108, n_2037, n_2038, n_2039);
  xor g1815 (n_2040, A[39], A[37]);
  xor g1816 (n_683, n_2040, A[33]);
  nand g1817 (n_2041, A[39], A[37]);
  nand g1818 (n_2042, A[33], A[37]);
  nand g1819 (n_2043, A[39], A[33]);
  nand g1820 (n_693, n_2041, n_2042, n_2043);
  xor g1822 (n_684, n_1592, A[31]);
  nand g1824 (n_2046, A[31], A[23]);
  nand g1826 (n_694, n_1593, n_2046, n_1787);
  xor g1827 (n_2048, A[21], A[35]);
  xor g1828 (n_682, n_2048, A[29]);
  nand g1829 (n_2049, A[21], A[35]);
  nand g1832 (n_695, n_2049, n_1915, n_1982);
  xor g1833 (n_2052, A[27], n_679);
  xor g1834 (n_686, n_2052, n_680);
  nand g1835 (n_2053, A[27], n_679);
  nand g1836 (n_2054, n_680, n_679);
  nand g1837 (n_2055, A[27], n_680);
  nand g1838 (n_699, n_2053, n_2054, n_2055);
  xor g1839 (n_2056, n_681, n_682);
  xor g1840 (n_688, n_2056, n_683);
  nand g1841 (n_2057, n_681, n_682);
  nand g1842 (n_2058, n_683, n_682);
  nand g1843 (n_2059, n_681, n_683);
  nand g1844 (n_701, n_2057, n_2058, n_2059);
  xor g1845 (n_2060, n_684, n_685);
  xor g1846 (n_690, n_2060, n_686);
  nand g1847 (n_2061, n_684, n_685);
  nand g1848 (n_2062, n_686, n_685);
  nand g1849 (n_2063, n_684, n_686);
  nand g1850 (n_703, n_2061, n_2062, n_2063);
  xor g1851 (n_2064, n_687, n_688);
  xor g1852 (n_691, n_2064, n_689);
  nand g1853 (n_2065, n_687, n_688);
  nand g1854 (n_2066, n_689, n_688);
  nand g1855 (n_2067, n_687, n_689);
  nand g1856 (n_706, n_2065, n_2066, n_2067);
  xor g1857 (n_2068, n_690, n_691);
  xor g1858 (n_191, n_2068, n_692);
  nand g1859 (n_2069, n_690, n_691);
  nand g1860 (n_2070, n_692, n_691);
  nand g1861 (n_2071, n_690, n_692);
  nand g1862 (n_107, n_2069, n_2070, n_2071);
  xor g1863 (n_2072, A[40], A[38]);
  xor g1864 (n_697, n_2072, A[34]);
  nand g1865 (n_2073, A[40], A[38]);
  nand g1866 (n_2074, A[34], A[38]);
  nand g1867 (n_2075, A[40], A[34]);
  nand g1868 (n_707, n_2073, n_2074, n_2075);
  xor g1870 (n_698, n_1624, A[32]);
  nand g1872 (n_2078, A[32], A[24]);
  nand g1874 (n_708, n_1625, n_2078, n_1819);
  xor g1875 (n_2080, A[22], A[36]);
  xor g1876 (n_696, n_2080, A[30]);
  nand g1877 (n_2081, A[22], A[36]);
  nand g1880 (n_709, n_2081, n_1947, n_2014);
  xor g1881 (n_2084, A[28], n_693);
  xor g1882 (n_700, n_2084, n_694);
  nand g1883 (n_2085, A[28], n_693);
  nand g1884 (n_2086, n_694, n_693);
  nand g1885 (n_2087, A[28], n_694);
  nand g1886 (n_713, n_2085, n_2086, n_2087);
  xor g1887 (n_2088, n_695, n_696);
  xor g1888 (n_702, n_2088, n_697);
  nand g1889 (n_2089, n_695, n_696);
  nand g1890 (n_2090, n_697, n_696);
  nand g1891 (n_2091, n_695, n_697);
  nand g1892 (n_715, n_2089, n_2090, n_2091);
  xor g1893 (n_2092, n_698, n_699);
  xor g1894 (n_704, n_2092, n_700);
  nand g1895 (n_2093, n_698, n_699);
  nand g1896 (n_2094, n_700, n_699);
  nand g1897 (n_2095, n_698, n_700);
  nand g1898 (n_717, n_2093, n_2094, n_2095);
  xor g1899 (n_2096, n_701, n_702);
  xor g1900 (n_705, n_2096, n_703);
  nand g1901 (n_2097, n_701, n_702);
  nand g1902 (n_2098, n_703, n_702);
  nand g1903 (n_2099, n_701, n_703);
  nand g1904 (n_720, n_2097, n_2098, n_2099);
  xor g1905 (n_2100, n_704, n_705);
  xor g1906 (n_190, n_2100, n_706);
  nand g1907 (n_2101, n_704, n_705);
  nand g1908 (n_2102, n_706, n_705);
  nand g1909 (n_2103, n_704, n_706);
  nand g1910 (n_106, n_2101, n_2102, n_2103);
  xor g1911 (n_2104, A[41], A[39]);
  xor g1912 (n_711, n_2104, A[35]);
  nand g1913 (n_2105, A[41], A[39]);
  nand g1914 (n_2106, A[35], A[39]);
  nand g1915 (n_2107, A[41], A[35]);
  nand g1916 (n_721, n_2105, n_2106, n_2107);
  xor g1918 (n_712, n_1656, A[33]);
  nand g1920 (n_2110, A[33], A[25]);
  nand g1922 (n_722, n_1657, n_2110, n_1851);
  xor g1923 (n_2112, A[23], A[37]);
  xor g1924 (n_710, n_2112, A[31]);
  nand g1925 (n_2113, A[23], A[37]);
  nand g1928 (n_723, n_2113, n_1979, n_2046);
  xor g1929 (n_2116, A[29], n_707);
  xor g1930 (n_714, n_2116, n_708);
  nand g1931 (n_2117, A[29], n_707);
  nand g1932 (n_2118, n_708, n_707);
  nand g1933 (n_2119, A[29], n_708);
  nand g1934 (n_727, n_2117, n_2118, n_2119);
  xor g1935 (n_2120, n_709, n_710);
  xor g1936 (n_716, n_2120, n_711);
  nand g1937 (n_2121, n_709, n_710);
  nand g1938 (n_2122, n_711, n_710);
  nand g1939 (n_2123, n_709, n_711);
  nand g1940 (n_729, n_2121, n_2122, n_2123);
  xor g1941 (n_2124, n_712, n_713);
  xor g1942 (n_718, n_2124, n_714);
  nand g1943 (n_2125, n_712, n_713);
  nand g1944 (n_2126, n_714, n_713);
  nand g1945 (n_2127, n_712, n_714);
  nand g1946 (n_731, n_2125, n_2126, n_2127);
  xor g1947 (n_2128, n_715, n_716);
  xor g1948 (n_719, n_2128, n_717);
  nand g1949 (n_2129, n_715, n_716);
  nand g1950 (n_2130, n_717, n_716);
  nand g1951 (n_2131, n_715, n_717);
  nand g1952 (n_734, n_2129, n_2130, n_2131);
  xor g1953 (n_2132, n_718, n_719);
  xor g1954 (n_189, n_2132, n_720);
  nand g1955 (n_2133, n_718, n_719);
  nand g1956 (n_2134, n_720, n_719);
  nand g1957 (n_2135, n_718, n_720);
  nand g1958 (n_105, n_2133, n_2134, n_2135);
  xor g1959 (n_2136, A[42], A[40]);
  xor g1960 (n_725, n_2136, A[36]);
  nand g1961 (n_2137, A[42], A[40]);
  nand g1962 (n_2138, A[36], A[40]);
  nand g1963 (n_2139, A[42], A[36]);
  nand g1964 (n_735, n_2137, n_2138, n_2139);
  xor g1966 (n_726, n_1688, A[34]);
  nand g1968 (n_2142, A[34], A[26]);
  nand g1970 (n_736, n_1689, n_2142, n_1883);
  xor g1971 (n_2144, A[24], A[38]);
  xor g1972 (n_724, n_2144, A[32]);
  nand g1973 (n_2145, A[24], A[38]);
  nand g1976 (n_737, n_2145, n_2011, n_2078);
  xor g1977 (n_2148, A[30], n_721);
  xor g1978 (n_728, n_2148, n_722);
  nand g1979 (n_2149, A[30], n_721);
  nand g1980 (n_2150, n_722, n_721);
  nand g1981 (n_2151, A[30], n_722);
  nand g1982 (n_741, n_2149, n_2150, n_2151);
  xor g1983 (n_2152, n_723, n_724);
  xor g1984 (n_730, n_2152, n_725);
  nand g1985 (n_2153, n_723, n_724);
  nand g1986 (n_2154, n_725, n_724);
  nand g1987 (n_2155, n_723, n_725);
  nand g1988 (n_743, n_2153, n_2154, n_2155);
  xor g1989 (n_2156, n_726, n_727);
  xor g1990 (n_732, n_2156, n_728);
  nand g1991 (n_2157, n_726, n_727);
  nand g1992 (n_2158, n_728, n_727);
  nand g1993 (n_2159, n_726, n_728);
  nand g1994 (n_745, n_2157, n_2158, n_2159);
  xor g1995 (n_2160, n_729, n_730);
  xor g1996 (n_733, n_2160, n_731);
  nand g1997 (n_2161, n_729, n_730);
  nand g1998 (n_2162, n_731, n_730);
  nand g1999 (n_2163, n_729, n_731);
  nand g2000 (n_748, n_2161, n_2162, n_2163);
  xor g2001 (n_2164, n_732, n_733);
  xor g2002 (n_188, n_2164, n_734);
  nand g2003 (n_2165, n_732, n_733);
  nand g2004 (n_2166, n_734, n_733);
  nand g2005 (n_2167, n_732, n_734);
  nand g2006 (n_104, n_2165, n_2166, n_2167);
  xor g2007 (n_2168, A[43], A[41]);
  xor g2008 (n_739, n_2168, A[37]);
  nand g2009 (n_2169, A[43], A[41]);
  nand g2010 (n_2170, A[37], A[41]);
  nand g2011 (n_2171, A[43], A[37]);
  nand g2012 (n_749, n_2169, n_2170, n_2171);
  xor g2014 (n_740, n_1720, A[35]);
  nand g2016 (n_2174, A[35], A[27]);
  nand g2018 (n_750, n_1721, n_2174, n_1915);
  xor g2019 (n_2176, A[25], A[39]);
  xor g2020 (n_738, n_2176, A[33]);
  nand g2021 (n_2177, A[25], A[39]);
  nand g2024 (n_751, n_2177, n_2043, n_2110);
  xor g2025 (n_2180, A[31], n_735);
  xor g2026 (n_742, n_2180, n_736);
  nand g2027 (n_2181, A[31], n_735);
  nand g2028 (n_2182, n_736, n_735);
  nand g2029 (n_2183, A[31], n_736);
  nand g2030 (n_755, n_2181, n_2182, n_2183);
  xor g2031 (n_2184, n_737, n_738);
  xor g2032 (n_744, n_2184, n_739);
  nand g2033 (n_2185, n_737, n_738);
  nand g2034 (n_2186, n_739, n_738);
  nand g2035 (n_2187, n_737, n_739);
  nand g2036 (n_757, n_2185, n_2186, n_2187);
  xor g2037 (n_2188, n_740, n_741);
  xor g2038 (n_746, n_2188, n_742);
  nand g2039 (n_2189, n_740, n_741);
  nand g2040 (n_2190, n_742, n_741);
  nand g2041 (n_2191, n_740, n_742);
  nand g2042 (n_759, n_2189, n_2190, n_2191);
  xor g2043 (n_2192, n_743, n_744);
  xor g2044 (n_747, n_2192, n_745);
  nand g2045 (n_2193, n_743, n_744);
  nand g2046 (n_2194, n_745, n_744);
  nand g2047 (n_2195, n_743, n_745);
  nand g2048 (n_762, n_2193, n_2194, n_2195);
  xor g2049 (n_2196, n_746, n_747);
  xor g2050 (n_187, n_2196, n_748);
  nand g2051 (n_2197, n_746, n_747);
  nand g2052 (n_2198, n_748, n_747);
  nand g2053 (n_2199, n_746, n_748);
  nand g2054 (n_103, n_2197, n_2198, n_2199);
  xor g2055 (n_2200, A[44], A[42]);
  xor g2056 (n_753, n_2200, A[38]);
  nand g2057 (n_2201, A[44], A[42]);
  nand g2058 (n_2202, A[38], A[42]);
  nand g2059 (n_2203, A[44], A[38]);
  nand g2060 (n_763, n_2201, n_2202, n_2203);
  xor g2062 (n_754, n_1752, A[36]);
  nand g2064 (n_2206, A[36], A[28]);
  nand g2066 (n_764, n_1753, n_2206, n_1947);
  xor g2067 (n_2208, A[26], A[40]);
  xor g2068 (n_752, n_2208, A[34]);
  nand g2069 (n_2209, A[26], A[40]);
  nand g2072 (n_765, n_2209, n_2075, n_2142);
  xor g2073 (n_2212, A[32], n_749);
  xor g2074 (n_756, n_2212, n_750);
  nand g2075 (n_2213, A[32], n_749);
  nand g2076 (n_2214, n_750, n_749);
  nand g2077 (n_2215, A[32], n_750);
  nand g2078 (n_769, n_2213, n_2214, n_2215);
  xor g2079 (n_2216, n_751, n_752);
  xor g2080 (n_758, n_2216, n_753);
  nand g2081 (n_2217, n_751, n_752);
  nand g2082 (n_2218, n_753, n_752);
  nand g2083 (n_2219, n_751, n_753);
  nand g2084 (n_771, n_2217, n_2218, n_2219);
  xor g2085 (n_2220, n_754, n_755);
  xor g2086 (n_760, n_2220, n_756);
  nand g2087 (n_2221, n_754, n_755);
  nand g2088 (n_2222, n_756, n_755);
  nand g2089 (n_2223, n_754, n_756);
  nand g2090 (n_773, n_2221, n_2222, n_2223);
  xor g2091 (n_2224, n_757, n_758);
  xor g2092 (n_761, n_2224, n_759);
  nand g2093 (n_2225, n_757, n_758);
  nand g2094 (n_2226, n_759, n_758);
  nand g2095 (n_2227, n_757, n_759);
  nand g2096 (n_776, n_2225, n_2226, n_2227);
  xor g2097 (n_2228, n_760, n_761);
  xor g2098 (n_186, n_2228, n_762);
  nand g2099 (n_2229, n_760, n_761);
  nand g2100 (n_2230, n_762, n_761);
  nand g2101 (n_2231, n_760, n_762);
  nand g2102 (n_102, n_2229, n_2230, n_2231);
  xor g2103 (n_2232, A[45], A[43]);
  xor g2104 (n_767, n_2232, A[39]);
  nand g2105 (n_2233, A[45], A[43]);
  nand g2106 (n_2234, A[39], A[43]);
  nand g2107 (n_2235, A[45], A[39]);
  nand g2108 (n_777, n_2233, n_2234, n_2235);
  xor g2110 (n_768, n_1784, A[37]);
  nand g2112 (n_2238, A[37], A[29]);
  nand g2114 (n_778, n_1785, n_2238, n_1979);
  xor g2115 (n_2240, A[27], A[41]);
  xor g2116 (n_766, n_2240, A[35]);
  nand g2117 (n_2241, A[27], A[41]);
  nand g2120 (n_779, n_2241, n_2107, n_2174);
  xor g2121 (n_2244, A[33], n_763);
  xor g2122 (n_770, n_2244, n_764);
  nand g2123 (n_2245, A[33], n_763);
  nand g2124 (n_2246, n_764, n_763);
  nand g2125 (n_2247, A[33], n_764);
  nand g2126 (n_783, n_2245, n_2246, n_2247);
  xor g2127 (n_2248, n_765, n_766);
  xor g2128 (n_772, n_2248, n_767);
  nand g2129 (n_2249, n_765, n_766);
  nand g2130 (n_2250, n_767, n_766);
  nand g2131 (n_2251, n_765, n_767);
  nand g2132 (n_785, n_2249, n_2250, n_2251);
  xor g2133 (n_2252, n_768, n_769);
  xor g2134 (n_774, n_2252, n_770);
  nand g2135 (n_2253, n_768, n_769);
  nand g2136 (n_2254, n_770, n_769);
  nand g2137 (n_2255, n_768, n_770);
  nand g2138 (n_787, n_2253, n_2254, n_2255);
  xor g2139 (n_2256, n_771, n_772);
  xor g2140 (n_775, n_2256, n_773);
  nand g2141 (n_2257, n_771, n_772);
  nand g2142 (n_2258, n_773, n_772);
  nand g2143 (n_2259, n_771, n_773);
  nand g2144 (n_790, n_2257, n_2258, n_2259);
  xor g2145 (n_2260, n_774, n_775);
  xor g2146 (n_185, n_2260, n_776);
  nand g2147 (n_2261, n_774, n_775);
  nand g2148 (n_2262, n_776, n_775);
  nand g2149 (n_2263, n_774, n_776);
  nand g2150 (n_101, n_2261, n_2262, n_2263);
  xor g2151 (n_2264, A[46], A[44]);
  xor g2152 (n_781, n_2264, A[40]);
  nand g2153 (n_2265, A[46], A[44]);
  nand g2154 (n_2266, A[40], A[44]);
  nand g2155 (n_2267, A[46], A[40]);
  nand g2156 (n_791, n_2265, n_2266, n_2267);
  xor g2158 (n_782, n_1816, A[38]);
  nand g2160 (n_2270, A[38], A[30]);
  nand g2162 (n_792, n_1817, n_2270, n_2011);
  xor g2163 (n_2272, A[28], A[42]);
  xor g2164 (n_780, n_2272, A[36]);
  nand g2165 (n_2273, A[28], A[42]);
  nand g2168 (n_793, n_2273, n_2139, n_2206);
  xor g2169 (n_2276, A[34], n_777);
  xor g2170 (n_784, n_2276, n_778);
  nand g2171 (n_2277, A[34], n_777);
  nand g2172 (n_2278, n_778, n_777);
  nand g2173 (n_2279, A[34], n_778);
  nand g2174 (n_797, n_2277, n_2278, n_2279);
  xor g2175 (n_2280, n_779, n_780);
  xor g2176 (n_786, n_2280, n_781);
  nand g2177 (n_2281, n_779, n_780);
  nand g2178 (n_2282, n_781, n_780);
  nand g2179 (n_2283, n_779, n_781);
  nand g2180 (n_799, n_2281, n_2282, n_2283);
  xor g2181 (n_2284, n_782, n_783);
  xor g2182 (n_788, n_2284, n_784);
  nand g2183 (n_2285, n_782, n_783);
  nand g2184 (n_2286, n_784, n_783);
  nand g2185 (n_2287, n_782, n_784);
  nand g2186 (n_801, n_2285, n_2286, n_2287);
  xor g2187 (n_2288, n_785, n_786);
  xor g2188 (n_789, n_2288, n_787);
  nand g2189 (n_2289, n_785, n_786);
  nand g2190 (n_2290, n_787, n_786);
  nand g2191 (n_2291, n_785, n_787);
  nand g2192 (n_804, n_2289, n_2290, n_2291);
  xor g2193 (n_2292, n_788, n_789);
  xor g2194 (n_184, n_2292, n_790);
  nand g2195 (n_2293, n_788, n_789);
  nand g2196 (n_2294, n_790, n_789);
  nand g2197 (n_2295, n_788, n_790);
  nand g2198 (n_100, n_2293, n_2294, n_2295);
  xor g2199 (n_2296, A[47], A[45]);
  xor g2200 (n_795, n_2296, A[41]);
  nand g2201 (n_2297, A[47], A[45]);
  nand g2202 (n_2298, A[41], A[45]);
  nand g2203 (n_2299, A[47], A[41]);
  nand g2204 (n_805, n_2297, n_2298, n_2299);
  xor g2206 (n_796, n_1848, A[39]);
  nand g2208 (n_2302, A[39], A[31]);
  nand g2210 (n_806, n_1849, n_2302, n_2043);
  xor g2211 (n_2304, A[29], A[43]);
  xor g2212 (n_794, n_2304, A[37]);
  nand g2213 (n_2305, A[29], A[43]);
  nand g2216 (n_807, n_2305, n_2171, n_2238);
  xor g2217 (n_2308, A[35], n_791);
  xor g2218 (n_798, n_2308, n_792);
  nand g2219 (n_2309, A[35], n_791);
  nand g2220 (n_2310, n_792, n_791);
  nand g2221 (n_2311, A[35], n_792);
  nand g2222 (n_811, n_2309, n_2310, n_2311);
  xor g2223 (n_2312, n_793, n_794);
  xor g2224 (n_800, n_2312, n_795);
  nand g2225 (n_2313, n_793, n_794);
  nand g2226 (n_2314, n_795, n_794);
  nand g2227 (n_2315, n_793, n_795);
  nand g2228 (n_813, n_2313, n_2314, n_2315);
  xor g2229 (n_2316, n_796, n_797);
  xor g2230 (n_802, n_2316, n_798);
  nand g2231 (n_2317, n_796, n_797);
  nand g2232 (n_2318, n_798, n_797);
  nand g2233 (n_2319, n_796, n_798);
  nand g2234 (n_815, n_2317, n_2318, n_2319);
  xor g2235 (n_2320, n_799, n_800);
  xor g2236 (n_803, n_2320, n_801);
  nand g2237 (n_2321, n_799, n_800);
  nand g2238 (n_2322, n_801, n_800);
  nand g2239 (n_2323, n_799, n_801);
  nand g2240 (n_818, n_2321, n_2322, n_2323);
  xor g2241 (n_2324, n_802, n_803);
  xor g2242 (n_183, n_2324, n_804);
  nand g2243 (n_2325, n_802, n_803);
  nand g2244 (n_2326, n_804, n_803);
  nand g2245 (n_2327, n_802, n_804);
  nand g2246 (n_99, n_2325, n_2326, n_2327);
  xor g2247 (n_2328, A[48], A[46]);
  xor g2248 (n_809, n_2328, A[42]);
  nand g2249 (n_2329, A[48], A[46]);
  nand g2250 (n_2330, A[42], A[46]);
  nand g2251 (n_2331, A[48], A[42]);
  nand g2252 (n_819, n_2329, n_2330, n_2331);
  xor g2254 (n_810, n_1880, A[40]);
  nand g2256 (n_2334, A[40], A[32]);
  nand g2258 (n_820, n_1881, n_2334, n_2075);
  xor g2259 (n_2336, A[30], A[44]);
  xor g2260 (n_808, n_2336, A[38]);
  nand g2261 (n_2337, A[30], A[44]);
  nand g2264 (n_821, n_2337, n_2203, n_2270);
  xor g2265 (n_2340, A[36], n_805);
  xor g2266 (n_812, n_2340, n_806);
  nand g2267 (n_2341, A[36], n_805);
  nand g2268 (n_2342, n_806, n_805);
  nand g2269 (n_2343, A[36], n_806);
  nand g2270 (n_825, n_2341, n_2342, n_2343);
  xor g2271 (n_2344, n_807, n_808);
  xor g2272 (n_814, n_2344, n_809);
  nand g2273 (n_2345, n_807, n_808);
  nand g2274 (n_2346, n_809, n_808);
  nand g2275 (n_2347, n_807, n_809);
  nand g2276 (n_827, n_2345, n_2346, n_2347);
  xor g2277 (n_2348, n_810, n_811);
  xor g2278 (n_816, n_2348, n_812);
  nand g2279 (n_2349, n_810, n_811);
  nand g2280 (n_2350, n_812, n_811);
  nand g2281 (n_2351, n_810, n_812);
  nand g2282 (n_829, n_2349, n_2350, n_2351);
  xor g2283 (n_2352, n_813, n_814);
  xor g2284 (n_817, n_2352, n_815);
  nand g2285 (n_2353, n_813, n_814);
  nand g2286 (n_2354, n_815, n_814);
  nand g2287 (n_2355, n_813, n_815);
  nand g2288 (n_832, n_2353, n_2354, n_2355);
  xor g2289 (n_2356, n_816, n_817);
  xor g2290 (n_182, n_2356, n_818);
  nand g2291 (n_2357, n_816, n_817);
  nand g2292 (n_2358, n_818, n_817);
  nand g2293 (n_2359, n_816, n_818);
  nand g2294 (n_98, n_2357, n_2358, n_2359);
  xor g2295 (n_2360, A[49], A[47]);
  xor g2296 (n_823, n_2360, A[43]);
  nand g2297 (n_2361, A[49], A[47]);
  nand g2298 (n_2362, A[43], A[47]);
  nand g2299 (n_2363, A[49], A[43]);
  nand g2300 (n_833, n_2361, n_2362, n_2363);
  xor g2302 (n_824, n_1912, A[41]);
  nand g2304 (n_2366, A[41], A[33]);
  nand g2306 (n_834, n_1913, n_2366, n_2107);
  xor g2307 (n_2368, A[31], A[45]);
  xor g2308 (n_822, n_2368, A[39]);
  nand g2309 (n_2369, A[31], A[45]);
  nand g2312 (n_835, n_2369, n_2235, n_2302);
  xor g2313 (n_2372, A[37], n_819);
  xor g2314 (n_826, n_2372, n_820);
  nand g2315 (n_2373, A[37], n_819);
  nand g2316 (n_2374, n_820, n_819);
  nand g2317 (n_2375, A[37], n_820);
  nand g2318 (n_839, n_2373, n_2374, n_2375);
  xor g2319 (n_2376, n_821, n_822);
  xor g2320 (n_828, n_2376, n_823);
  nand g2321 (n_2377, n_821, n_822);
  nand g2322 (n_2378, n_823, n_822);
  nand g2323 (n_2379, n_821, n_823);
  nand g2324 (n_841, n_2377, n_2378, n_2379);
  xor g2325 (n_2380, n_824, n_825);
  xor g2326 (n_830, n_2380, n_826);
  nand g2327 (n_2381, n_824, n_825);
  nand g2328 (n_2382, n_826, n_825);
  nand g2329 (n_2383, n_824, n_826);
  nand g2330 (n_843, n_2381, n_2382, n_2383);
  xor g2331 (n_2384, n_827, n_828);
  xor g2332 (n_831, n_2384, n_829);
  nand g2333 (n_2385, n_827, n_828);
  nand g2334 (n_2386, n_829, n_828);
  nand g2335 (n_2387, n_827, n_829);
  nand g2336 (n_846, n_2385, n_2386, n_2387);
  xor g2337 (n_2388, n_830, n_831);
  xor g2338 (n_181, n_2388, n_832);
  nand g2339 (n_2389, n_830, n_831);
  nand g2340 (n_2390, n_832, n_831);
  nand g2341 (n_2391, n_830, n_832);
  nand g2342 (n_97, n_2389, n_2390, n_2391);
  xor g2343 (n_2392, A[50], A[48]);
  xor g2344 (n_837, n_2392, A[44]);
  nand g2345 (n_2393, A[50], A[48]);
  nand g2346 (n_2394, A[44], A[48]);
  nand g2347 (n_2395, A[50], A[44]);
  nand g2348 (n_847, n_2393, n_2394, n_2395);
  xor g2350 (n_838, n_1944, A[42]);
  nand g2352 (n_2398, A[42], A[34]);
  nand g2354 (n_848, n_1945, n_2398, n_2139);
  xor g2355 (n_2400, A[32], A[46]);
  xor g2356 (n_836, n_2400, A[40]);
  nand g2357 (n_2401, A[32], A[46]);
  nand g2360 (n_849, n_2401, n_2267, n_2334);
  xor g2361 (n_2404, A[38], n_833);
  xor g2362 (n_840, n_2404, n_834);
  nand g2363 (n_2405, A[38], n_833);
  nand g2364 (n_2406, n_834, n_833);
  nand g2365 (n_2407, A[38], n_834);
  nand g2366 (n_853, n_2405, n_2406, n_2407);
  xor g2367 (n_2408, n_835, n_836);
  xor g2368 (n_842, n_2408, n_837);
  nand g2369 (n_2409, n_835, n_836);
  nand g2370 (n_2410, n_837, n_836);
  nand g2371 (n_2411, n_835, n_837);
  nand g2372 (n_855, n_2409, n_2410, n_2411);
  xor g2373 (n_2412, n_838, n_839);
  xor g2374 (n_844, n_2412, n_840);
  nand g2375 (n_2413, n_838, n_839);
  nand g2376 (n_2414, n_840, n_839);
  nand g2377 (n_2415, n_838, n_840);
  nand g2378 (n_857, n_2413, n_2414, n_2415);
  xor g2379 (n_2416, n_841, n_842);
  xor g2380 (n_845, n_2416, n_843);
  nand g2381 (n_2417, n_841, n_842);
  nand g2382 (n_2418, n_843, n_842);
  nand g2383 (n_2419, n_841, n_843);
  nand g2384 (n_860, n_2417, n_2418, n_2419);
  xor g2385 (n_2420, n_844, n_845);
  xor g2386 (n_180, n_2420, n_846);
  nand g2387 (n_2421, n_844, n_845);
  nand g2388 (n_2422, n_846, n_845);
  nand g2389 (n_2423, n_844, n_846);
  nand g2390 (n_96, n_2421, n_2422, n_2423);
  xor g2391 (n_2424, A[51], A[49]);
  xor g2392 (n_851, n_2424, A[45]);
  nand g2393 (n_2425, A[51], A[49]);
  nand g2394 (n_2426, A[45], A[49]);
  nand g2395 (n_2427, A[51], A[45]);
  nand g2396 (n_861, n_2425, n_2426, n_2427);
  xor g2398 (n_852, n_1976, A[43]);
  nand g2400 (n_2430, A[43], A[35]);
  nand g2402 (n_862, n_1977, n_2430, n_2171);
  xor g2403 (n_2432, A[33], A[47]);
  xor g2404 (n_850, n_2432, A[41]);
  nand g2405 (n_2433, A[33], A[47]);
  nand g2408 (n_863, n_2433, n_2299, n_2366);
  xor g2409 (n_2436, A[39], n_847);
  xor g2410 (n_854, n_2436, n_848);
  nand g2411 (n_2437, A[39], n_847);
  nand g2412 (n_2438, n_848, n_847);
  nand g2413 (n_2439, A[39], n_848);
  nand g2414 (n_867, n_2437, n_2438, n_2439);
  xor g2415 (n_2440, n_849, n_850);
  xor g2416 (n_856, n_2440, n_851);
  nand g2417 (n_2441, n_849, n_850);
  nand g2418 (n_2442, n_851, n_850);
  nand g2419 (n_2443, n_849, n_851);
  nand g2420 (n_869, n_2441, n_2442, n_2443);
  xor g2421 (n_2444, n_852, n_853);
  xor g2422 (n_858, n_2444, n_854);
  nand g2423 (n_2445, n_852, n_853);
  nand g2424 (n_2446, n_854, n_853);
  nand g2425 (n_2447, n_852, n_854);
  nand g2426 (n_871, n_2445, n_2446, n_2447);
  xor g2427 (n_2448, n_855, n_856);
  xor g2428 (n_859, n_2448, n_857);
  nand g2429 (n_2449, n_855, n_856);
  nand g2430 (n_2450, n_857, n_856);
  nand g2431 (n_2451, n_855, n_857);
  nand g2432 (n_874, n_2449, n_2450, n_2451);
  xor g2433 (n_2452, n_858, n_859);
  xor g2434 (n_179, n_2452, n_860);
  nand g2435 (n_2453, n_858, n_859);
  nand g2436 (n_2454, n_860, n_859);
  nand g2437 (n_2455, n_858, n_860);
  nand g2438 (n_95, n_2453, n_2454, n_2455);
  xor g2439 (n_2456, A[52], A[50]);
  xor g2440 (n_865, n_2456, A[46]);
  nand g2441 (n_2457, A[52], A[50]);
  nand g2442 (n_2458, A[46], A[50]);
  nand g2443 (n_2459, A[52], A[46]);
  nand g2444 (n_875, n_2457, n_2458, n_2459);
  xor g2446 (n_866, n_2008, A[44]);
  nand g2448 (n_2462, A[44], A[36]);
  nand g2450 (n_876, n_2009, n_2462, n_2203);
  xor g2451 (n_2464, A[34], A[48]);
  xor g2452 (n_864, n_2464, A[42]);
  nand g2453 (n_2465, A[34], A[48]);
  nand g2456 (n_877, n_2465, n_2331, n_2398);
  xor g2457 (n_2468, A[40], n_861);
  xor g2458 (n_868, n_2468, n_862);
  nand g2459 (n_2469, A[40], n_861);
  nand g2460 (n_2470, n_862, n_861);
  nand g2461 (n_2471, A[40], n_862);
  nand g2462 (n_881, n_2469, n_2470, n_2471);
  xor g2463 (n_2472, n_863, n_864);
  xor g2464 (n_870, n_2472, n_865);
  nand g2465 (n_2473, n_863, n_864);
  nand g2466 (n_2474, n_865, n_864);
  nand g2467 (n_2475, n_863, n_865);
  nand g2468 (n_883, n_2473, n_2474, n_2475);
  xor g2469 (n_2476, n_866, n_867);
  xor g2470 (n_872, n_2476, n_868);
  nand g2471 (n_2477, n_866, n_867);
  nand g2472 (n_2478, n_868, n_867);
  nand g2473 (n_2479, n_866, n_868);
  nand g2474 (n_885, n_2477, n_2478, n_2479);
  xor g2475 (n_2480, n_869, n_870);
  xor g2476 (n_873, n_2480, n_871);
  nand g2477 (n_2481, n_869, n_870);
  nand g2478 (n_2482, n_871, n_870);
  nand g2479 (n_2483, n_869, n_871);
  nand g2480 (n_888, n_2481, n_2482, n_2483);
  xor g2481 (n_2484, n_872, n_873);
  xor g2482 (n_178, n_2484, n_874);
  nand g2483 (n_2485, n_872, n_873);
  nand g2484 (n_2486, n_874, n_873);
  nand g2485 (n_2487, n_872, n_874);
  nand g2486 (n_94, n_2485, n_2486, n_2487);
  xor g2487 (n_2488, A[53], A[51]);
  xor g2488 (n_879, n_2488, A[47]);
  nand g2489 (n_2489, A[53], A[51]);
  nand g2490 (n_2490, A[47], A[51]);
  nand g2491 (n_2491, A[53], A[47]);
  nand g2492 (n_889, n_2489, n_2490, n_2491);
  xor g2494 (n_880, n_2040, A[45]);
  nand g2496 (n_2494, A[45], A[37]);
  nand g2498 (n_890, n_2041, n_2494, n_2235);
  xor g2499 (n_2496, A[35], A[49]);
  xor g2500 (n_878, n_2496, A[43]);
  nand g2501 (n_2497, A[35], A[49]);
  nand g2504 (n_891, n_2497, n_2363, n_2430);
  xor g2505 (n_2500, A[41], n_875);
  xor g2506 (n_882, n_2500, n_876);
  nand g2507 (n_2501, A[41], n_875);
  nand g2508 (n_2502, n_876, n_875);
  nand g2509 (n_2503, A[41], n_876);
  nand g2510 (n_895, n_2501, n_2502, n_2503);
  xor g2511 (n_2504, n_877, n_878);
  xor g2512 (n_884, n_2504, n_879);
  nand g2513 (n_2505, n_877, n_878);
  nand g2514 (n_2506, n_879, n_878);
  nand g2515 (n_2507, n_877, n_879);
  nand g2516 (n_897, n_2505, n_2506, n_2507);
  xor g2517 (n_2508, n_880, n_881);
  xor g2518 (n_886, n_2508, n_882);
  nand g2519 (n_2509, n_880, n_881);
  nand g2520 (n_2510, n_882, n_881);
  nand g2521 (n_2511, n_880, n_882);
  nand g2522 (n_899, n_2509, n_2510, n_2511);
  xor g2523 (n_2512, n_883, n_884);
  xor g2524 (n_887, n_2512, n_885);
  nand g2525 (n_2513, n_883, n_884);
  nand g2526 (n_2514, n_885, n_884);
  nand g2527 (n_2515, n_883, n_885);
  nand g2528 (n_902, n_2513, n_2514, n_2515);
  xor g2529 (n_2516, n_886, n_887);
  xor g2530 (n_177, n_2516, n_888);
  nand g2531 (n_2517, n_886, n_887);
  nand g2532 (n_2518, n_888, n_887);
  nand g2533 (n_2519, n_886, n_888);
  nand g2534 (n_93, n_2517, n_2518, n_2519);
  xor g2535 (n_2520, A[54], A[52]);
  xor g2536 (n_893, n_2520, A[48]);
  nand g2537 (n_2521, A[54], A[52]);
  nand g2538 (n_2522, A[48], A[52]);
  nand g2539 (n_2523, A[54], A[48]);
  nand g2540 (n_903, n_2521, n_2522, n_2523);
  xor g2542 (n_894, n_2072, A[46]);
  nand g2544 (n_2526, A[46], A[38]);
  nand g2546 (n_904, n_2073, n_2526, n_2267);
  xor g2547 (n_2528, A[36], A[50]);
  xor g2548 (n_892, n_2528, A[44]);
  nand g2549 (n_2529, A[36], A[50]);
  nand g2552 (n_905, n_2529, n_2395, n_2462);
  xor g2553 (n_2532, A[42], n_889);
  xor g2554 (n_896, n_2532, n_890);
  nand g2555 (n_2533, A[42], n_889);
  nand g2556 (n_2534, n_890, n_889);
  nand g2557 (n_2535, A[42], n_890);
  nand g2558 (n_909, n_2533, n_2534, n_2535);
  xor g2559 (n_2536, n_891, n_892);
  xor g2560 (n_898, n_2536, n_893);
  nand g2561 (n_2537, n_891, n_892);
  nand g2562 (n_2538, n_893, n_892);
  nand g2563 (n_2539, n_891, n_893);
  nand g2564 (n_911, n_2537, n_2538, n_2539);
  xor g2565 (n_2540, n_894, n_895);
  xor g2566 (n_900, n_2540, n_896);
  nand g2567 (n_2541, n_894, n_895);
  nand g2568 (n_2542, n_896, n_895);
  nand g2569 (n_2543, n_894, n_896);
  nand g2570 (n_913, n_2541, n_2542, n_2543);
  xor g2571 (n_2544, n_897, n_898);
  xor g2572 (n_901, n_2544, n_899);
  nand g2573 (n_2545, n_897, n_898);
  nand g2574 (n_2546, n_899, n_898);
  nand g2575 (n_2547, n_897, n_899);
  nand g2576 (n_916, n_2545, n_2546, n_2547);
  xor g2577 (n_2548, n_900, n_901);
  xor g2578 (n_176, n_2548, n_902);
  nand g2579 (n_2549, n_900, n_901);
  nand g2580 (n_2550, n_902, n_901);
  nand g2581 (n_2551, n_900, n_902);
  nand g2582 (n_92, n_2549, n_2550, n_2551);
  xor g2583 (n_2552, A[55], A[53]);
  xor g2584 (n_907, n_2552, A[49]);
  nand g2585 (n_2553, A[55], A[53]);
  nand g2586 (n_2554, A[49], A[53]);
  nand g2587 (n_2555, A[55], A[49]);
  nand g2588 (n_917, n_2553, n_2554, n_2555);
  xor g2590 (n_908, n_2104, A[47]);
  nand g2592 (n_2558, A[47], A[39]);
  nand g2594 (n_918, n_2105, n_2558, n_2299);
  xor g2595 (n_2560, A[37], A[51]);
  xor g2596 (n_906, n_2560, A[45]);
  nand g2597 (n_2561, A[37], A[51]);
  nand g2600 (n_919, n_2561, n_2427, n_2494);
  xor g2601 (n_2564, A[43], n_903);
  xor g2602 (n_910, n_2564, n_904);
  nand g2603 (n_2565, A[43], n_903);
  nand g2604 (n_2566, n_904, n_903);
  nand g2605 (n_2567, A[43], n_904);
  nand g2606 (n_923, n_2565, n_2566, n_2567);
  xor g2607 (n_2568, n_905, n_906);
  xor g2608 (n_912, n_2568, n_907);
  nand g2609 (n_2569, n_905, n_906);
  nand g2610 (n_2570, n_907, n_906);
  nand g2611 (n_2571, n_905, n_907);
  nand g2612 (n_925, n_2569, n_2570, n_2571);
  xor g2613 (n_2572, n_908, n_909);
  xor g2614 (n_914, n_2572, n_910);
  nand g2615 (n_2573, n_908, n_909);
  nand g2616 (n_2574, n_910, n_909);
  nand g2617 (n_2575, n_908, n_910);
  nand g2618 (n_927, n_2573, n_2574, n_2575);
  xor g2619 (n_2576, n_911, n_912);
  xor g2620 (n_915, n_2576, n_913);
  nand g2621 (n_2577, n_911, n_912);
  nand g2622 (n_2578, n_913, n_912);
  nand g2623 (n_2579, n_911, n_913);
  nand g2624 (n_930, n_2577, n_2578, n_2579);
  xor g2625 (n_2580, n_914, n_915);
  xor g2626 (n_175, n_2580, n_916);
  nand g2627 (n_2581, n_914, n_915);
  nand g2628 (n_2582, n_916, n_915);
  nand g2629 (n_2583, n_914, n_916);
  nand g2630 (n_91, n_2581, n_2582, n_2583);
  xor g2631 (n_2584, A[56], A[54]);
  xor g2632 (n_921, n_2584, A[50]);
  nand g2633 (n_2585, A[56], A[54]);
  nand g2634 (n_2586, A[50], A[54]);
  nand g2635 (n_2587, A[56], A[50]);
  nand g2636 (n_931, n_2585, n_2586, n_2587);
  xor g2638 (n_922, n_2136, A[48]);
  nand g2640 (n_2590, A[48], A[40]);
  nand g2642 (n_932, n_2137, n_2590, n_2331);
  xor g2643 (n_2592, A[38], A[52]);
  xor g2644 (n_920, n_2592, A[46]);
  nand g2645 (n_2593, A[38], A[52]);
  nand g2648 (n_933, n_2593, n_2459, n_2526);
  xor g2649 (n_2596, A[44], n_917);
  xor g2650 (n_924, n_2596, n_918);
  nand g2651 (n_2597, A[44], n_917);
  nand g2652 (n_2598, n_918, n_917);
  nand g2653 (n_2599, A[44], n_918);
  nand g2654 (n_937, n_2597, n_2598, n_2599);
  xor g2655 (n_2600, n_919, n_920);
  xor g2656 (n_926, n_2600, n_921);
  nand g2657 (n_2601, n_919, n_920);
  nand g2658 (n_2602, n_921, n_920);
  nand g2659 (n_2603, n_919, n_921);
  nand g2660 (n_939, n_2601, n_2602, n_2603);
  xor g2661 (n_2604, n_922, n_923);
  xor g2662 (n_928, n_2604, n_924);
  nand g2663 (n_2605, n_922, n_923);
  nand g2664 (n_2606, n_924, n_923);
  nand g2665 (n_2607, n_922, n_924);
  nand g2666 (n_941, n_2605, n_2606, n_2607);
  xor g2667 (n_2608, n_925, n_926);
  xor g2668 (n_929, n_2608, n_927);
  nand g2669 (n_2609, n_925, n_926);
  nand g2670 (n_2610, n_927, n_926);
  nand g2671 (n_2611, n_925, n_927);
  nand g2672 (n_944, n_2609, n_2610, n_2611);
  xor g2673 (n_2612, n_928, n_929);
  xor g2674 (n_174, n_2612, n_930);
  nand g2675 (n_2613, n_928, n_929);
  nand g2676 (n_2614, n_930, n_929);
  nand g2677 (n_2615, n_928, n_930);
  nand g2678 (n_90, n_2613, n_2614, n_2615);
  xor g2679 (n_2616, A[57], A[55]);
  xor g2680 (n_935, n_2616, A[51]);
  nand g2681 (n_2617, A[57], A[55]);
  nand g2682 (n_2618, A[51], A[55]);
  nand g2683 (n_2619, A[57], A[51]);
  nand g2684 (n_945, n_2617, n_2618, n_2619);
  xor g2686 (n_936, n_2168, A[49]);
  nand g2688 (n_2622, A[49], A[41]);
  nand g2690 (n_946, n_2169, n_2622, n_2363);
  xor g2691 (n_2624, A[39], A[53]);
  xor g2692 (n_934, n_2624, A[47]);
  nand g2693 (n_2625, A[39], A[53]);
  nand g2696 (n_947, n_2625, n_2491, n_2558);
  xor g2697 (n_2628, A[45], n_931);
  xor g2698 (n_938, n_2628, n_932);
  nand g2699 (n_2629, A[45], n_931);
  nand g2700 (n_2630, n_932, n_931);
  nand g2701 (n_2631, A[45], n_932);
  nand g2702 (n_951, n_2629, n_2630, n_2631);
  xor g2703 (n_2632, n_933, n_934);
  xor g2704 (n_940, n_2632, n_935);
  nand g2705 (n_2633, n_933, n_934);
  nand g2706 (n_2634, n_935, n_934);
  nand g2707 (n_2635, n_933, n_935);
  nand g2708 (n_953, n_2633, n_2634, n_2635);
  xor g2709 (n_2636, n_936, n_937);
  xor g2710 (n_942, n_2636, n_938);
  nand g2711 (n_2637, n_936, n_937);
  nand g2712 (n_2638, n_938, n_937);
  nand g2713 (n_2639, n_936, n_938);
  nand g2714 (n_955, n_2637, n_2638, n_2639);
  xor g2715 (n_2640, n_939, n_940);
  xor g2716 (n_943, n_2640, n_941);
  nand g2717 (n_2641, n_939, n_940);
  nand g2718 (n_2642, n_941, n_940);
  nand g2719 (n_2643, n_939, n_941);
  nand g2720 (n_958, n_2641, n_2642, n_2643);
  xor g2721 (n_2644, n_942, n_943);
  xor g2722 (n_173, n_2644, n_944);
  nand g2723 (n_2645, n_942, n_943);
  nand g2724 (n_2646, n_944, n_943);
  nand g2725 (n_2647, n_942, n_944);
  nand g2726 (n_89, n_2645, n_2646, n_2647);
  xor g2727 (n_2648, A[58], A[56]);
  xor g2728 (n_949, n_2648, A[52]);
  nand g2729 (n_2649, A[58], A[56]);
  nand g2730 (n_2650, A[52], A[56]);
  nand g2731 (n_2651, A[58], A[52]);
  nand g2732 (n_959, n_2649, n_2650, n_2651);
  xor g2734 (n_950, n_2200, A[50]);
  nand g2736 (n_2654, A[50], A[42]);
  nand g2738 (n_960, n_2201, n_2654, n_2395);
  xor g2739 (n_2656, A[40], A[54]);
  xor g2740 (n_948, n_2656, A[48]);
  nand g2741 (n_2657, A[40], A[54]);
  nand g2744 (n_961, n_2657, n_2523, n_2590);
  xor g2745 (n_2660, A[46], n_945);
  xor g2746 (n_952, n_2660, n_946);
  nand g2747 (n_2661, A[46], n_945);
  nand g2748 (n_2662, n_946, n_945);
  nand g2749 (n_2663, A[46], n_946);
  nand g2750 (n_965, n_2661, n_2662, n_2663);
  xor g2751 (n_2664, n_947, n_948);
  xor g2752 (n_954, n_2664, n_949);
  nand g2753 (n_2665, n_947, n_948);
  nand g2754 (n_2666, n_949, n_948);
  nand g2755 (n_2667, n_947, n_949);
  nand g2756 (n_967, n_2665, n_2666, n_2667);
  xor g2757 (n_2668, n_950, n_951);
  xor g2758 (n_956, n_2668, n_952);
  nand g2759 (n_2669, n_950, n_951);
  nand g2760 (n_2670, n_952, n_951);
  nand g2761 (n_2671, n_950, n_952);
  nand g2762 (n_969, n_2669, n_2670, n_2671);
  xor g2763 (n_2672, n_953, n_954);
  xor g2764 (n_957, n_2672, n_955);
  nand g2765 (n_2673, n_953, n_954);
  nand g2766 (n_2674, n_955, n_954);
  nand g2767 (n_2675, n_953, n_955);
  nand g2768 (n_972, n_2673, n_2674, n_2675);
  xor g2769 (n_2676, n_956, n_957);
  xor g2770 (n_172, n_2676, n_958);
  nand g2771 (n_2677, n_956, n_957);
  nand g2772 (n_2678, n_958, n_957);
  nand g2773 (n_2679, n_956, n_958);
  nand g2774 (n_88, n_2677, n_2678, n_2679);
  xor g2775 (n_2680, A[59], A[57]);
  xor g2776 (n_963, n_2680, A[53]);
  nand g2777 (n_2681, A[59], A[57]);
  nand g2778 (n_2682, A[53], A[57]);
  nand g2779 (n_2683, A[59], A[53]);
  nand g2780 (n_973, n_2681, n_2682, n_2683);
  xor g2782 (n_964, n_2232, A[51]);
  nand g2784 (n_2686, A[51], A[43]);
  nand g2786 (n_974, n_2233, n_2686, n_2427);
  xor g2787 (n_2688, A[41], A[55]);
  xor g2788 (n_962, n_2688, A[49]);
  nand g2789 (n_2689, A[41], A[55]);
  nand g2792 (n_975, n_2689, n_2555, n_2622);
  xor g2793 (n_2692, A[47], n_959);
  xor g2794 (n_966, n_2692, n_960);
  nand g2795 (n_2693, A[47], n_959);
  nand g2796 (n_2694, n_960, n_959);
  nand g2797 (n_2695, A[47], n_960);
  nand g2798 (n_979, n_2693, n_2694, n_2695);
  xor g2799 (n_2696, n_961, n_962);
  xor g2800 (n_968, n_2696, n_963);
  nand g2801 (n_2697, n_961, n_962);
  nand g2802 (n_2698, n_963, n_962);
  nand g2803 (n_2699, n_961, n_963);
  nand g2804 (n_981, n_2697, n_2698, n_2699);
  xor g2805 (n_2700, n_964, n_965);
  xor g2806 (n_970, n_2700, n_966);
  nand g2807 (n_2701, n_964, n_965);
  nand g2808 (n_2702, n_966, n_965);
  nand g2809 (n_2703, n_964, n_966);
  nand g2810 (n_983, n_2701, n_2702, n_2703);
  xor g2811 (n_2704, n_967, n_968);
  xor g2812 (n_971, n_2704, n_969);
  nand g2813 (n_2705, n_967, n_968);
  nand g2814 (n_2706, n_969, n_968);
  nand g2815 (n_2707, n_967, n_969);
  nand g2816 (n_986, n_2705, n_2706, n_2707);
  xor g2817 (n_2708, n_970, n_971);
  xor g2818 (n_171, n_2708, n_972);
  nand g2819 (n_2709, n_970, n_971);
  nand g2820 (n_2710, n_972, n_971);
  nand g2821 (n_2711, n_970, n_972);
  nand g2822 (n_87, n_2709, n_2710, n_2711);
  xor g2823 (n_2712, A[60], A[58]);
  xor g2824 (n_977, n_2712, A[54]);
  nand g2825 (n_2713, A[60], A[58]);
  nand g2826 (n_2714, A[54], A[58]);
  nand g2827 (n_2715, A[60], A[54]);
  nand g2828 (n_987, n_2713, n_2714, n_2715);
  xor g2830 (n_978, n_2264, A[52]);
  nand g2832 (n_2718, A[52], A[44]);
  nand g2834 (n_988, n_2265, n_2718, n_2459);
  xor g2835 (n_2720, A[42], A[56]);
  xor g2836 (n_976, n_2720, A[50]);
  nand g2837 (n_2721, A[42], A[56]);
  nand g2840 (n_989, n_2721, n_2587, n_2654);
  xor g2841 (n_2724, A[48], n_973);
  xor g2842 (n_980, n_2724, n_974);
  nand g2843 (n_2725, A[48], n_973);
  nand g2844 (n_2726, n_974, n_973);
  nand g2845 (n_2727, A[48], n_974);
  nand g2846 (n_993, n_2725, n_2726, n_2727);
  xor g2847 (n_2728, n_975, n_976);
  xor g2848 (n_982, n_2728, n_977);
  nand g2849 (n_2729, n_975, n_976);
  nand g2850 (n_2730, n_977, n_976);
  nand g2851 (n_2731, n_975, n_977);
  nand g2852 (n_995, n_2729, n_2730, n_2731);
  xor g2853 (n_2732, n_978, n_979);
  xor g2854 (n_984, n_2732, n_980);
  nand g2855 (n_2733, n_978, n_979);
  nand g2856 (n_2734, n_980, n_979);
  nand g2857 (n_2735, n_978, n_980);
  nand g2858 (n_997, n_2733, n_2734, n_2735);
  xor g2859 (n_2736, n_981, n_982);
  xor g2860 (n_985, n_2736, n_983);
  nand g2861 (n_2737, n_981, n_982);
  nand g2862 (n_2738, n_983, n_982);
  nand g2863 (n_2739, n_981, n_983);
  nand g2864 (n_1000, n_2737, n_2738, n_2739);
  xor g2865 (n_2740, n_984, n_985);
  xor g2866 (n_170, n_2740, n_986);
  nand g2867 (n_2741, n_984, n_985);
  nand g2868 (n_2742, n_986, n_985);
  nand g2869 (n_2743, n_984, n_986);
  nand g2870 (n_86, n_2741, n_2742, n_2743);
  xor g2871 (n_2744, A[61], A[59]);
  xor g2872 (n_991, n_2744, A[55]);
  nand g2873 (n_2745, A[61], A[59]);
  nand g2874 (n_2746, A[55], A[59]);
  nand g2875 (n_2747, A[61], A[55]);
  nand g2876 (n_1001, n_2745, n_2746, n_2747);
  xor g2878 (n_992, n_2296, A[53]);
  nand g2880 (n_2750, A[53], A[45]);
  nand g2882 (n_1002, n_2297, n_2750, n_2491);
  xor g2883 (n_2752, A[43], A[57]);
  xor g2884 (n_990, n_2752, A[51]);
  nand g2885 (n_2753, A[43], A[57]);
  nand g2888 (n_1003, n_2753, n_2619, n_2686);
  xor g2889 (n_2756, A[49], n_987);
  xor g2890 (n_994, n_2756, n_988);
  nand g2891 (n_2757, A[49], n_987);
  nand g2892 (n_2758, n_988, n_987);
  nand g2893 (n_2759, A[49], n_988);
  nand g2894 (n_1007, n_2757, n_2758, n_2759);
  xor g2895 (n_2760, n_989, n_990);
  xor g2896 (n_996, n_2760, n_991);
  nand g2897 (n_2761, n_989, n_990);
  nand g2898 (n_2762, n_991, n_990);
  nand g2899 (n_2763, n_989, n_991);
  nand g2900 (n_1009, n_2761, n_2762, n_2763);
  xor g2901 (n_2764, n_992, n_993);
  xor g2902 (n_998, n_2764, n_994);
  nand g2903 (n_2765, n_992, n_993);
  nand g2904 (n_2766, n_994, n_993);
  nand g2905 (n_2767, n_992, n_994);
  nand g2906 (n_1011, n_2765, n_2766, n_2767);
  xor g2907 (n_2768, n_995, n_996);
  xor g2908 (n_999, n_2768, n_997);
  nand g2909 (n_2769, n_995, n_996);
  nand g2910 (n_2770, n_997, n_996);
  nand g2911 (n_2771, n_995, n_997);
  nand g2912 (n_1014, n_2769, n_2770, n_2771);
  xor g2913 (n_2772, n_998, n_999);
  xor g2914 (n_169, n_2772, n_1000);
  nand g2915 (n_2773, n_998, n_999);
  nand g2916 (n_2774, n_1000, n_999);
  nand g2917 (n_2775, n_998, n_1000);
  nand g2918 (n_85, n_2773, n_2774, n_2775);
  xor g2919 (n_2776, A[62], A[60]);
  xor g2920 (n_1005, n_2776, A[56]);
  nand g2921 (n_2777, A[62], A[60]);
  nand g2922 (n_2778, A[56], A[60]);
  nand g2923 (n_2779, A[62], A[56]);
  nand g2924 (n_1018, n_2777, n_2778, n_2779);
  xor g2926 (n_1006, n_2328, A[54]);
  nand g2928 (n_2782, A[54], A[46]);
  nand g2930 (n_1019, n_2329, n_2782, n_2523);
  xor g2931 (n_2784, A[44], A[58]);
  xor g2932 (n_1004, n_2784, A[52]);
  nand g2933 (n_2785, A[44], A[58]);
  nand g2936 (n_1017, n_2785, n_2651, n_2718);
  xor g2937 (n_2788, A[50], n_1001);
  xor g2938 (n_1008, n_2788, n_1002);
  nand g2939 (n_2789, A[50], n_1001);
  nand g2940 (n_2790, n_1002, n_1001);
  nand g2941 (n_2791, A[50], n_1002);
  nand g2942 (n_1023, n_2789, n_2790, n_2791);
  xor g2943 (n_2792, n_1003, n_1004);
  xor g2944 (n_1010, n_2792, n_1005);
  nand g2945 (n_2793, n_1003, n_1004);
  nand g2946 (n_2794, n_1005, n_1004);
  nand g2947 (n_2795, n_1003, n_1005);
  nand g2948 (n_1025, n_2793, n_2794, n_2795);
  xor g2949 (n_2796, n_1006, n_1007);
  xor g2950 (n_1012, n_2796, n_1008);
  nand g2951 (n_2797, n_1006, n_1007);
  nand g2952 (n_2798, n_1008, n_1007);
  nand g2953 (n_2799, n_1006, n_1008);
  nand g2954 (n_1027, n_2797, n_2798, n_2799);
  xor g2955 (n_2800, n_1009, n_1010);
  xor g2956 (n_1013, n_2800, n_1011);
  nand g2957 (n_2801, n_1009, n_1010);
  nand g2958 (n_2802, n_1011, n_1010);
  nand g2959 (n_2803, n_1009, n_1011);
  nand g2960 (n_1030, n_2801, n_2802, n_2803);
  xor g2961 (n_2804, n_1012, n_1013);
  xor g2962 (n_168, n_2804, n_1014);
  nand g2963 (n_2805, n_1012, n_1013);
  nand g2964 (n_2806, n_1014, n_1013);
  nand g2965 (n_2807, n_1012, n_1014);
  nand g2966 (n_84, n_2805, n_2806, n_2807);
  xor g2969 (n_2808, A[63], A[57]);
  xor g2970 (n_1021, n_2808, A[49]);
  nand g2971 (n_2809, A[63], A[57]);
  nand g2972 (n_2810, A[49], A[57]);
  nand g2973 (n_2811, A[63], A[49]);
  nand g2974 (n_1034, n_2809, n_2810, n_2811);
  xor g2975 (n_2812, A[47], A[61]);
  xor g2976 (n_1022, n_2812, A[45]);
  nand g2977 (n_2813, A[47], A[61]);
  nand g2978 (n_2814, A[45], A[61]);
  nand g2980 (n_1035, n_2813, n_2814, n_2297);
  xor g2981 (n_2816, A[55], A[59]);
  xor g2982 (n_1020, n_2816, A[53]);
  nand g2986 (n_1036, n_2746, n_2683, n_2553);
  xor g2987 (n_2820, A[51], n_1017);
  xor g2988 (n_1024, n_2820, n_1018);
  nand g2989 (n_2821, A[51], n_1017);
  nand g2990 (n_2822, n_1018, n_1017);
  nand g2991 (n_2823, A[51], n_1018);
  nand g2992 (n_1040, n_2821, n_2822, n_2823);
  xor g2993 (n_2824, n_1019, n_1020);
  xor g2994 (n_1026, n_2824, n_1021);
  nand g2995 (n_2825, n_1019, n_1020);
  nand g2996 (n_2826, n_1021, n_1020);
  nand g2997 (n_2827, n_1019, n_1021);
  nand g2998 (n_1042, n_2825, n_2826, n_2827);
  xor g2999 (n_2828, n_1022, n_1023);
  xor g3000 (n_1028, n_2828, n_1024);
  nand g3001 (n_2829, n_1022, n_1023);
  nand g3002 (n_2830, n_1024, n_1023);
  nand g3003 (n_2831, n_1022, n_1024);
  nand g3004 (n_1045, n_2829, n_2830, n_2831);
  xor g3005 (n_2832, n_1025, n_1026);
  xor g3006 (n_1029, n_2832, n_1027);
  nand g3007 (n_2833, n_1025, n_1026);
  nand g3008 (n_2834, n_1027, n_1026);
  nand g3009 (n_2835, n_1025, n_1027);
  nand g3010 (n_1047, n_2833, n_2834, n_2835);
  xor g3011 (n_2836, n_1028, n_1029);
  xor g3012 (n_167, n_2836, n_1030);
  nand g3013 (n_2837, n_1028, n_1029);
  nand g3014 (n_2838, n_1030, n_1029);
  nand g3015 (n_2839, n_1028, n_1030);
  nand g3016 (n_83, n_2837, n_2838, n_2839);
  xor g3019 (n_2840, A[56], A[48]);
  xor g3020 (n_1038, n_2840, A[46]);
  nand g3021 (n_2841, A[56], A[48]);
  nand g3023 (n_2843, A[56], A[46]);
  nand g3024 (n_1049, n_2841, n_2329, n_2843);
  xor g3025 (n_2844, A[62], A[54]);
  xor g3026 (n_1039, n_2844, A[60]);
  nand g3027 (n_2845, A[62], A[54]);
  nand g3030 (n_1051, n_2845, n_2715, n_2777);
  xor g3031 (n_2848, A[58], A[52]);
  xor g3032 (n_1037, n_2848, A[50]);
  nand g3035 (n_2851, A[58], A[50]);
  nand g3036 (n_1050, n_2651, n_2457, n_2851);
  xor g3037 (n_2852, A[63], n_1034);
  xor g3038 (n_1041, n_2852, n_1035);
  nand g3039 (n_2853, A[63], n_1034);
  nand g3040 (n_2854, n_1035, n_1034);
  nand g3041 (n_2855, A[63], n_1035);
  nand g3042 (n_1055, n_2853, n_2854, n_2855);
  xor g3043 (n_2856, n_1036, n_1037);
  xor g3044 (n_1043, n_2856, n_1038);
  nand g3045 (n_2857, n_1036, n_1037);
  nand g3046 (n_2858, n_1038, n_1037);
  nand g3047 (n_2859, n_1036, n_1038);
  nand g3048 (n_1057, n_2857, n_2858, n_2859);
  xor g3049 (n_2860, n_1039, n_1040);
  xor g3050 (n_1044, n_2860, n_1041);
  nand g3051 (n_2861, n_1039, n_1040);
  nand g3052 (n_2862, n_1041, n_1040);
  nand g3053 (n_2863, n_1039, n_1041);
  nand g3054 (n_1060, n_2861, n_2862, n_2863);
  xor g3055 (n_2864, n_1042, n_1043);
  xor g3056 (n_1046, n_2864, n_1044);
  nand g3057 (n_2865, n_1042, n_1043);
  nand g3058 (n_2866, n_1044, n_1043);
  nand g3059 (n_2867, n_1042, n_1044);
  nand g3060 (n_1062, n_2865, n_2866, n_2867);
  xor g3061 (n_2868, n_1045, n_1046);
  xor g3062 (n_166, n_2868, n_1047);
  nand g3063 (n_2869, n_1045, n_1046);
  nand g3064 (n_2870, n_1047, n_1046);
  nand g3065 (n_2871, n_1045, n_1047);
  nand g3066 (n_82, n_2869, n_2870, n_2871);
  xor g3068 (n_1053, n_2872, A[57]);
  nand g3070 (n_2874, A[57], A[61]);
  nand g3072 (n_1065, n_2873, n_2874, n_2875);
  xor g3074 (n_1054, n_2360, A[55]);
  nand g3076 (n_2878, A[55], A[47]);
  nand g3078 (n_1066, n_2361, n_2878, n_2555);
  xor g3079 (n_2880, A[59], A[53]);
  xor g3080 (n_1052, n_2880, A[51]);
  nand g3083 (n_2883, A[59], A[51]);
  nand g3084 (n_1067, n_2683, n_2489, n_2883);
  xor g3086 (n_1056, n_2884, n_1050);
  nand g3088 (n_2886, n_1050, n_1049);
  nand g3090 (n_1071, n_2885, n_2886, n_2887);
  xor g3091 (n_2888, n_1051, n_1052);
  xor g3092 (n_1058, n_2888, n_1053);
  nand g3093 (n_2889, n_1051, n_1052);
  nand g3094 (n_2890, n_1053, n_1052);
  nand g3095 (n_2891, n_1051, n_1053);
  nand g3096 (n_1073, n_2889, n_2890, n_2891);
  xor g3097 (n_2892, n_1054, n_1055);
  xor g3098 (n_1059, n_2892, n_1056);
  nand g3099 (n_2893, n_1054, n_1055);
  nand g3100 (n_2894, n_1056, n_1055);
  nand g3101 (n_2895, n_1054, n_1056);
  nand g3102 (n_1075, n_2893, n_2894, n_2895);
  xor g3103 (n_2896, n_1057, n_1058);
  xor g3104 (n_1061, n_2896, n_1059);
  nand g3105 (n_2897, n_1057, n_1058);
  nand g3106 (n_2898, n_1059, n_1058);
  nand g3107 (n_2899, n_1057, n_1059);
  nand g3108 (n_1077, n_2897, n_2898, n_2899);
  xor g3109 (n_2900, n_1060, n_1061);
  xor g3110 (n_165, n_2900, n_1062);
  nand g3111 (n_2901, n_1060, n_1061);
  nand g3112 (n_2902, n_1062, n_1061);
  nand g3113 (n_2903, n_1060, n_1062);
  nand g3114 (n_81, n_2901, n_2902, n_2903);
  xor g3117 (n_2904, A[60], A[48]);
  xor g3118 (n_1069, n_2904, A[56]);
  nand g3119 (n_2905, A[60], A[48]);
  nand g3122 (n_1080, n_2905, n_2841, n_2778);
  xor g3123 (n_2908, A[54], A[58]);
  xor g3124 (n_1068, n_2908, A[52]);
  nand g3128 (n_1079, n_2714, n_2651, n_2521);
  xor g3130 (n_1070, n_2912, n_1065);
  nand g3133 (n_2915, A[50], n_1065);
  nand g3134 (n_1084, n_2913, n_2914, n_2915);
  xor g3135 (n_2916, n_1066, n_1067);
  xor g3136 (n_1072, n_2916, n_1068);
  nand g3137 (n_2917, n_1066, n_1067);
  nand g3138 (n_2918, n_1068, n_1067);
  nand g3139 (n_2919, n_1066, n_1068);
  nand g3140 (n_1086, n_2917, n_2918, n_2919);
  xor g3141 (n_2920, n_1069, n_1070);
  xor g3142 (n_1074, n_2920, n_1071);
  nand g3143 (n_2921, n_1069, n_1070);
  nand g3144 (n_2922, n_1071, n_1070);
  nand g3145 (n_2923, n_1069, n_1071);
  nand g3146 (n_1087, n_2921, n_2922, n_2923);
  xor g3147 (n_2924, n_1072, n_1073);
  xor g3148 (n_1076, n_2924, n_1074);
  nand g3149 (n_2925, n_1072, n_1073);
  nand g3150 (n_2926, n_1074, n_1073);
  nand g3151 (n_2927, n_1072, n_1074);
  nand g3152 (n_1090, n_2925, n_2926, n_2927);
  xor g3153 (n_2928, n_1075, n_1076);
  xor g3154 (n_164, n_2928, n_1077);
  nand g3155 (n_2929, n_1075, n_1076);
  nand g3156 (n_2930, n_1077, n_1076);
  nand g3157 (n_2931, n_1075, n_1077);
  nand g3158 (n_80, n_2929, n_2930, n_2931);
  xor g3165 (n_2936, A[49], A[55]);
  xor g3166 (n_1082, n_2936, A[59]);
  nand g3169 (n_2939, A[49], A[59]);
  nand g3170 (n_1094, n_2555, n_2746, n_2939);
  xor g3172 (n_1083, n_2488, A[62]);
  nand g3174 (n_2942, A[62], A[51]);
  nand g3175 (n_2943, A[53], A[62]);
  nand g3176 (n_1097, n_2489, n_2942, n_2943);
  xor g3177 (n_2944, n_1079, n_1080);
  xor g3178 (n_1085, n_2944, n_1053);
  nand g3179 (n_2945, n_1079, n_1080);
  nand g3180 (n_2946, n_1053, n_1080);
  nand g3181 (n_2947, n_1079, n_1053);
  nand g3182 (n_1099, n_2945, n_2946, n_2947);
  xor g3183 (n_2948, n_1082, n_1083);
  xor g3184 (n_1088, n_2948, n_1084);
  nand g3185 (n_2949, n_1082, n_1083);
  nand g3186 (n_2950, n_1084, n_1083);
  nand g3187 (n_2951, n_1082, n_1084);
  nand g3188 (n_1101, n_2949, n_2950, n_2951);
  xor g3189 (n_2952, n_1085, n_1086);
  xor g3190 (n_1089, n_2952, n_1087);
  nand g3191 (n_2953, n_1085, n_1086);
  nand g3192 (n_2954, n_1087, n_1086);
  nand g3193 (n_2955, n_1085, n_1087);
  nand g3194 (n_1103, n_2953, n_2954, n_2955);
  xor g3195 (n_2956, n_1088, n_1089);
  xor g3196 (n_163, n_2956, n_1090);
  nand g3197 (n_2957, n_1088, n_1089);
  nand g3198 (n_2958, n_1090, n_1089);
  nand g3199 (n_2959, n_1088, n_1090);
  nand g3200 (n_162, n_2957, n_2958, n_2959);
  xor g3203 (n_2960, A[60], A[56]);
  xor g3204 (n_1096, n_2960, A[54]);
  nand g3208 (n_1105, n_2778, n_2585, n_2715);
  xor g3216 (n_1098, n_2968, n_1094);
  nand g3218 (n_2970, n_1094, n_1065);
  nand g3220 (n_1110, n_2914, n_2970, n_2971);
  xor g3221 (n_2972, n_1037, n_1096);
  xor g3222 (n_1100, n_2972, n_1097);
  nand g3223 (n_2973, n_1037, n_1096);
  nand g3224 (n_2974, n_1097, n_1096);
  nand g3225 (n_2975, n_1037, n_1097);
  nand g3226 (n_1111, n_2973, n_2974, n_2975);
  xor g3227 (n_2976, n_1098, n_1099);
  xor g3228 (n_1102, n_2976, n_1100);
  nand g3229 (n_2977, n_1098, n_1099);
  nand g3230 (n_2978, n_1100, n_1099);
  nand g3231 (n_2979, n_1098, n_1100);
  nand g3232 (n_1114, n_2977, n_2978, n_2979);
  xor g3233 (n_2980, n_1101, n_1102);
  xor g3234 (n_79, n_2980, n_1103);
  nand g3235 (n_2981, n_1101, n_1102);
  nand g3236 (n_2982, n_1103, n_1102);
  nand g3237 (n_2983, n_1101, n_1103);
  nand g3238 (n_78, n_2981, n_2982, n_2983);
  xor g3251 (n_2992, A[51], A[62]);
  xor g3252 (n_1109, n_2992, n_1105);
  nand g3254 (n_2994, n_1105, A[62]);
  nand g3255 (n_2995, A[51], n_1105);
  nand g3256 (n_1121, n_2942, n_2994, n_2995);
  xor g3257 (n_2996, n_1050, n_1020);
  xor g3258 (n_1112, n_2996, n_1053);
  nand g3259 (n_2997, n_1050, n_1020);
  nand g3260 (n_2998, n_1053, n_1020);
  nand g3261 (n_2999, n_1050, n_1053);
  nand g3262 (n_1122, n_2997, n_2998, n_2999);
  xor g3263 (n_3000, n_1109, n_1110);
  xor g3264 (n_1113, n_3000, n_1111);
  nand g3265 (n_3001, n_1109, n_1110);
  nand g3266 (n_3002, n_1111, n_1110);
  nand g3267 (n_3003, n_1109, n_1111);
  nand g3268 (n_1125, n_3001, n_3002, n_3003);
  xor g3269 (n_3004, n_1112, n_1113);
  xor g3270 (n_161, n_3004, n_1114);
  nand g3271 (n_3005, n_1112, n_1113);
  nand g3272 (n_3006, n_1114, n_1113);
  nand g3273 (n_3007, n_1112, n_1114);
  nand g3274 (n_77, n_3005, n_3006, n_3007);
  xor g3278 (n_1119, n_2584, A[62]);
  nand g3282 (n_1127, n_2585, n_2845, n_2779);
  nand g3288 (n_1130, n_2651, n_3014, n_3015);
  xor g3289 (n_3016, n_1036, n_1065);
  xor g3290 (n_1123, n_3016, n_1119);
  nand g3291 (n_3017, n_1036, n_1065);
  nand g3292 (n_3018, n_1119, n_1065);
  nand g3293 (n_3019, n_1036, n_1119);
  nand g3294 (n_1132, n_3017, n_3018, n_3019);
  xor g3295 (n_3020, n_1120, n_1121);
  xor g3296 (n_1124, n_3020, n_1122);
  nand g3297 (n_3021, n_1120, n_1121);
  nand g3298 (n_3022, n_1122, n_1121);
  nand g3299 (n_3023, n_1120, n_1122);
  nand g3300 (n_1134, n_3021, n_3022, n_3023);
  xor g3301 (n_3024, n_1123, n_1124);
  xor g3302 (n_160, n_3024, n_1125);
  nand g3303 (n_3025, n_1123, n_1124);
  nand g3304 (n_3026, n_1125, n_1124);
  nand g3305 (n_3027, n_1123, n_1125);
  nand g3306 (n_76, n_3025, n_3026, n_3027);
  xor g3319 (n_3036, A[60], n_1127);
  xor g3320 (n_1131, n_3036, n_1020);
  nand g3321 (n_3037, A[60], n_1127);
  nand g3322 (n_3038, n_1020, n_1127);
  nand g3323 (n_3039, A[60], n_1020);
  nand g3324 (n_1141, n_3037, n_3038, n_3039);
  xor g3325 (n_3040, n_1053, n_1130);
  xor g3326 (n_1133, n_3040, n_1131);
  nand g3327 (n_3041, n_1053, n_1130);
  nand g3328 (n_3042, n_1131, n_1130);
  nand g3329 (n_3043, n_1053, n_1131);
  nand g3330 (n_1143, n_3041, n_3042, n_3043);
  xor g3331 (n_3044, n_1132, n_1133);
  xor g3332 (n_159, n_3044, n_1134);
  nand g3333 (n_3045, n_1132, n_1133);
  nand g3334 (n_3046, n_1134, n_1133);
  nand g3335 (n_3047, n_1132, n_1134);
  nand g3336 (n_75, n_3045, n_3046, n_3047);
  nand g3349 (n_3055, A[58], n_1036);
  nand g3350 (n_1148, n_3014, n_3054, n_3055);
  xor g3351 (n_3056, n_1065, n_1119);
  xor g3352 (n_1142, n_3056, n_1140);
  nand g3354 (n_3058, n_1140, n_1119);
  nand g3355 (n_3059, n_1065, n_1140);
  nand g3356 (n_1150, n_3018, n_3058, n_3059);
  xor g3357 (n_3060, n_1141, n_1142);
  xor g3358 (n_158, n_3060, n_1143);
  nand g3359 (n_3061, n_1141, n_1142);
  nand g3360 (n_3062, n_1143, n_1142);
  nand g3361 (n_3063, n_1141, n_1143);
  nand g3362 (n_157, n_3061, n_3062, n_3063);
  xor g3370 (n_1147, n_2816, A[60]);
  nand g3372 (n_3070, A[60], A[59]);
  nand g3373 (n_3071, A[55], A[60]);
  nand g3374 (n_1155, n_2746, n_3070, n_3071);
  xor g3375 (n_3072, n_1127, n_1053);
  xor g3376 (n_1149, n_3072, n_1147);
  nand g3377 (n_3073, n_1127, n_1053);
  nand g3378 (n_3074, n_1147, n_1053);
  nand g3379 (n_3075, n_1127, n_1147);
  nand g3380 (n_1157, n_3073, n_3074, n_3075);
  xor g3381 (n_3076, n_1148, n_1149);
  xor g3382 (n_74, n_3076, n_1150);
  nand g3383 (n_3077, n_1148, n_1149);
  nand g3384 (n_3078, n_1150, n_1149);
  nand g3385 (n_3079, n_1148, n_1150);
  nand g3386 (n_156, n_3077, n_3078, n_3079);
  xor g3390 (n_1154, n_2960, A[58]);
  nand g3394 (n_1159, n_2778, n_2713, n_2649);
  xor g3396 (n_1156, n_2968, n_1154);
  nand g3398 (n_3086, n_1154, n_1065);
  nand g3400 (n_1162, n_2914, n_3086, n_3087);
  xor g3401 (n_3088, n_1155, n_1156);
  xor g3402 (n_73, n_3088, n_1157);
  nand g3403 (n_3089, n_1155, n_1156);
  nand g3404 (n_3090, n_1157, n_1156);
  nand g3405 (n_3091, n_1155, n_1157);
  nand g3406 (n_155, n_3089, n_3090, n_3091);
  xor g3413 (n_3096, A[59], A[62]);
  xor g3414 (n_1161, n_3096, n_1159);
  nand g3415 (n_3097, A[59], A[62]);
  nand g3416 (n_3098, n_1159, A[62]);
  nand g3417 (n_3099, A[59], n_1159);
  nand g3418 (n_1167, n_3097, n_3098, n_3099);
  xor g3419 (n_3100, n_1053, n_1161);
  xor g3420 (n_72, n_3100, n_1162);
  nand g3421 (n_3101, n_1053, n_1161);
  nand g3422 (n_3102, n_1162, n_1161);
  nand g3423 (n_3103, n_1053, n_1162);
  nand g3424 (n_154, n_3101, n_3102, n_3103);
  nand g3432 (n_1170, n_2713, n_3106, n_3107);
  xor g3433 (n_3108, n_1065, n_1166);
  xor g3434 (n_71, n_3108, n_1167);
  nand g3435 (n_3109, n_1065, n_1166);
  nand g3436 (n_3110, n_1167, n_1166);
  nand g3437 (n_3111, n_1065, n_1167);
  nand g3438 (n_153, n_3109, n_3110, n_3111);
  xor g3440 (n_1169, n_2872, A[59]);
  nand g3444 (n_1173, n_2873, n_2745, n_3115);
  xor g3445 (n_3116, A[62], n_1169);
  xor g3446 (n_70, n_3116, n_1170);
  nand g3447 (n_3117, A[62], n_1169);
  nand g3448 (n_3118, n_1170, n_1169);
  nand g3449 (n_3119, A[62], n_1170);
  nand g3450 (n_152, n_3117, n_3118, n_3119);
  nand g3457 (n_3123, A[62], n_1173);
  nand g3458 (n_151, n_3121, n_3122, n_3123);
  xor g3460 (n_68, n_2872, A[60]);
  nand g3462 (n_3126, A[60], A[61]);
  nand g3464 (n_150, n_2873, n_3126, n_3127);
  nand g25 (n_3149, n_1177, n_3146, n_3147);
  nand g28 (n_3150, A[2], n_226);
  nand g29 (n_3151, A[2], n_3149);
  nand g30 (n_3152, n_226, n_3149);
  nand g31 (n_3154, n_3150, n_3151, n_3152);
  xor g32 (n_3153, A[2], n_226);
  xor g33 (Z[4], n_3149, n_3153);
  nand g34 (n_3155, n_142, n_225);
  nand g35 (n_3156, n_142, n_3154);
  nand g36 (n_3157, n_225, n_3154);
  nand g37 (n_3159, n_3155, n_3156, n_3157);
  xor g38 (n_3158, n_142, n_225);
  xor g39 (Z[5], n_3154, n_3158);
  nand g40 (n_3160, n_141, n_224);
  nand g41 (n_3161, n_141, n_3159);
  nand g42 (n_3162, n_224, n_3159);
  nand g43 (n_3164, n_3160, n_3161, n_3162);
  xor g44 (n_3163, n_141, n_224);
  xor g45 (Z[6], n_3159, n_3163);
  nand g46 (n_3165, n_140, n_223);
  nand g47 (n_3166, n_140, n_3164);
  nand g48 (n_3167, n_223, n_3164);
  nand g49 (n_3169, n_3165, n_3166, n_3167);
  xor g50 (n_3168, n_140, n_223);
  xor g51 (Z[7], n_3164, n_3168);
  nand g52 (n_3170, n_139, n_222);
  nand g53 (n_3171, n_139, n_3169);
  nand g54 (n_3172, n_222, n_3169);
  nand g55 (n_3174, n_3170, n_3171, n_3172);
  xor g56 (n_3173, n_139, n_222);
  xor g57 (Z[8], n_3169, n_3173);
  nand g58 (n_3175, n_138, n_221);
  nand g59 (n_3176, n_138, n_3174);
  nand g60 (n_3177, n_221, n_3174);
  nand g61 (n_3179, n_3175, n_3176, n_3177);
  xor g62 (n_3178, n_138, n_221);
  xor g63 (Z[9], n_3174, n_3178);
  nand g64 (n_3180, n_137, n_220);
  nand g65 (n_3181, n_137, n_3179);
  nand g66 (n_3182, n_220, n_3179);
  nand g67 (n_3184, n_3180, n_3181, n_3182);
  xor g68 (n_3183, n_137, n_220);
  xor g69 (Z[10], n_3179, n_3183);
  nand g70 (n_3185, n_136, n_219);
  nand g71 (n_3186, n_136, n_3184);
  nand g72 (n_3187, n_219, n_3184);
  nand g73 (n_3189, n_3185, n_3186, n_3187);
  xor g74 (n_3188, n_136, n_219);
  xor g75 (Z[11], n_3184, n_3188);
  nand g76 (n_3190, n_135, n_218);
  nand g77 (n_3191, n_135, n_3189);
  nand g78 (n_3192, n_218, n_3189);
  nand g79 (n_3194, n_3190, n_3191, n_3192);
  xor g80 (n_3193, n_135, n_218);
  xor g81 (Z[12], n_3189, n_3193);
  nand g82 (n_3195, n_134, n_217);
  nand g83 (n_3196, n_134, n_3194);
  nand g84 (n_3197, n_217, n_3194);
  nand g85 (n_3199, n_3195, n_3196, n_3197);
  xor g86 (n_3198, n_134, n_217);
  xor g87 (Z[13], n_3194, n_3198);
  nand g88 (n_3200, n_133, n_216);
  nand g89 (n_3201, n_133, n_3199);
  nand g90 (n_3202, n_216, n_3199);
  nand g91 (n_3204, n_3200, n_3201, n_3202);
  xor g92 (n_3203, n_133, n_216);
  xor g93 (Z[14], n_3199, n_3203);
  nand g94 (n_3205, n_132, n_215);
  nand g95 (n_3206, n_132, n_3204);
  nand g96 (n_3207, n_215, n_3204);
  nand g97 (n_3209, n_3205, n_3206, n_3207);
  xor g98 (n_3208, n_132, n_215);
  xor g99 (Z[15], n_3204, n_3208);
  nand g100 (n_3210, n_131, n_214);
  nand g101 (n_3211, n_131, n_3209);
  nand g102 (n_3212, n_214, n_3209);
  nand g103 (n_3214, n_3210, n_3211, n_3212);
  xor g104 (n_3213, n_131, n_214);
  xor g105 (Z[16], n_3209, n_3213);
  nand g106 (n_3215, n_130, n_213);
  nand g107 (n_3216, n_130, n_3214);
  nand g108 (n_3217, n_213, n_3214);
  nand g109 (n_3219, n_3215, n_3216, n_3217);
  xor g110 (n_3218, n_130, n_213);
  xor g111 (Z[17], n_3214, n_3218);
  nand g112 (n_3220, n_129, n_212);
  nand g113 (n_3221, n_129, n_3219);
  nand g114 (n_3222, n_212, n_3219);
  nand g115 (n_3224, n_3220, n_3221, n_3222);
  xor g116 (n_3223, n_129, n_212);
  xor g117 (Z[18], n_3219, n_3223);
  nand g118 (n_3225, n_128, n_211);
  nand g119 (n_3226, n_128, n_3224);
  nand g120 (n_3227, n_211, n_3224);
  nand g121 (n_3229, n_3225, n_3226, n_3227);
  xor g122 (n_3228, n_128, n_211);
  xor g123 (Z[19], n_3224, n_3228);
  nand g124 (n_3230, n_127, n_210);
  nand g125 (n_3231, n_127, n_3229);
  nand g126 (n_3232, n_210, n_3229);
  nand g127 (n_3234, n_3230, n_3231, n_3232);
  xor g128 (n_3233, n_127, n_210);
  xor g129 (Z[20], n_3229, n_3233);
  nand g130 (n_3235, n_126, n_209);
  nand g131 (n_3236, n_126, n_3234);
  nand g132 (n_3237, n_209, n_3234);
  nand g133 (n_3239, n_3235, n_3236, n_3237);
  xor g134 (n_3238, n_126, n_209);
  xor g135 (Z[21], n_3234, n_3238);
  nand g136 (n_3240, n_125, n_208);
  nand g137 (n_3241, n_125, n_3239);
  nand g138 (n_3242, n_208, n_3239);
  nand g139 (n_3244, n_3240, n_3241, n_3242);
  xor g140 (n_3243, n_125, n_208);
  xor g141 (Z[22], n_3239, n_3243);
  nand g142 (n_3245, n_124, n_207);
  nand g143 (n_3246, n_124, n_3244);
  nand g144 (n_3247, n_207, n_3244);
  nand g145 (n_3249, n_3245, n_3246, n_3247);
  xor g146 (n_3248, n_124, n_207);
  xor g147 (Z[23], n_3244, n_3248);
  nand g148 (n_3250, n_123, n_206);
  nand g149 (n_3251, n_123, n_3249);
  nand g150 (n_3252, n_206, n_3249);
  nand g151 (n_3254, n_3250, n_3251, n_3252);
  xor g152 (n_3253, n_123, n_206);
  xor g153 (Z[24], n_3249, n_3253);
  nand g154 (n_3255, n_122, n_205);
  nand g155 (n_3256, n_122, n_3254);
  nand g156 (n_3257, n_205, n_3254);
  nand g157 (n_3259, n_3255, n_3256, n_3257);
  xor g158 (n_3258, n_122, n_205);
  xor g159 (Z[25], n_3254, n_3258);
  nand g160 (n_3260, n_121, n_204);
  nand g161 (n_3261, n_121, n_3259);
  nand g162 (n_3262, n_204, n_3259);
  nand g163 (n_3264, n_3260, n_3261, n_3262);
  xor g164 (n_3263, n_121, n_204);
  xor g165 (Z[26], n_3259, n_3263);
  nand g166 (n_3265, n_120, n_203);
  nand g167 (n_3266, n_120, n_3264);
  nand g168 (n_3267, n_203, n_3264);
  nand g169 (n_3269, n_3265, n_3266, n_3267);
  xor g170 (n_3268, n_120, n_203);
  xor g171 (Z[27], n_3264, n_3268);
  nand g172 (n_3270, n_119, n_202);
  nand g173 (n_3271, n_119, n_3269);
  nand g174 (n_3272, n_202, n_3269);
  nand g175 (n_3274, n_3270, n_3271, n_3272);
  xor g176 (n_3273, n_119, n_202);
  xor g177 (Z[28], n_3269, n_3273);
  nand g178 (n_3275, n_118, n_201);
  nand g179 (n_3276, n_118, n_3274);
  nand g180 (n_3277, n_201, n_3274);
  nand g181 (n_3279, n_3275, n_3276, n_3277);
  xor g182 (n_3278, n_118, n_201);
  xor g183 (Z[29], n_3274, n_3278);
  nand g184 (n_3280, n_117, n_200);
  nand g185 (n_3281, n_117, n_3279);
  nand g186 (n_3282, n_200, n_3279);
  nand g187 (n_3284, n_3280, n_3281, n_3282);
  xor g188 (n_3283, n_117, n_200);
  xor g189 (Z[30], n_3279, n_3283);
  nand g190 (n_3285, n_116, n_199);
  nand g191 (n_3286, n_116, n_3284);
  nand g192 (n_3287, n_199, n_3284);
  nand g193 (n_3289, n_3285, n_3286, n_3287);
  xor g194 (n_3288, n_116, n_199);
  xor g195 (Z[31], n_3284, n_3288);
  nand g196 (n_3290, n_115, n_198);
  nand g197 (n_3291, n_115, n_3289);
  nand g198 (n_3292, n_198, n_3289);
  nand g199 (n_3294, n_3290, n_3291, n_3292);
  xor g200 (n_3293, n_115, n_198);
  xor g201 (Z[32], n_3289, n_3293);
  nand g202 (n_3295, n_114, n_197);
  nand g203 (n_3296, n_114, n_3294);
  nand g204 (n_3297, n_197, n_3294);
  nand g205 (n_3299, n_3295, n_3296, n_3297);
  xor g206 (n_3298, n_114, n_197);
  xor g207 (Z[33], n_3294, n_3298);
  nand g208 (n_3300, n_113, n_196);
  nand g209 (n_3301, n_113, n_3299);
  nand g210 (n_3302, n_196, n_3299);
  nand g211 (n_3304, n_3300, n_3301, n_3302);
  xor g212 (n_3303, n_113, n_196);
  xor g213 (Z[34], n_3299, n_3303);
  nand g214 (n_3305, n_112, n_195);
  nand g215 (n_3306, n_112, n_3304);
  nand g216 (n_3307, n_195, n_3304);
  nand g217 (n_3309, n_3305, n_3306, n_3307);
  xor g218 (n_3308, n_112, n_195);
  xor g219 (Z[35], n_3304, n_3308);
  nand g220 (n_3310, n_111, n_194);
  nand g221 (n_3311, n_111, n_3309);
  nand g222 (n_3312, n_194, n_3309);
  nand g223 (n_3314, n_3310, n_3311, n_3312);
  xor g224 (n_3313, n_111, n_194);
  xor g225 (Z[36], n_3309, n_3313);
  nand g226 (n_3315, n_110, n_193);
  nand g227 (n_3316, n_110, n_3314);
  nand g228 (n_3317, n_193, n_3314);
  nand g229 (n_3319, n_3315, n_3316, n_3317);
  xor g230 (n_3318, n_110, n_193);
  xor g231 (Z[37], n_3314, n_3318);
  nand g232 (n_3320, n_109, n_192);
  nand g233 (n_3321, n_109, n_3319);
  nand g234 (n_3322, n_192, n_3319);
  nand g235 (n_3324, n_3320, n_3321, n_3322);
  xor g236 (n_3323, n_109, n_192);
  xor g237 (Z[38], n_3319, n_3323);
  nand g238 (n_3325, n_108, n_191);
  nand g239 (n_3326, n_108, n_3324);
  nand g240 (n_3327, n_191, n_3324);
  nand g241 (n_3329, n_3325, n_3326, n_3327);
  xor g242 (n_3328, n_108, n_191);
  xor g243 (Z[39], n_3324, n_3328);
  nand g244 (n_3330, n_107, n_190);
  nand g245 (n_3331, n_107, n_3329);
  nand g246 (n_3332, n_190, n_3329);
  nand g247 (n_3334, n_3330, n_3331, n_3332);
  xor g248 (n_3333, n_107, n_190);
  xor g249 (Z[40], n_3329, n_3333);
  nand g250 (n_3335, n_106, n_189);
  nand g251 (n_3336, n_106, n_3334);
  nand g252 (n_3337, n_189, n_3334);
  nand g253 (n_3339, n_3335, n_3336, n_3337);
  xor g254 (n_3338, n_106, n_189);
  xor g255 (Z[41], n_3334, n_3338);
  nand g256 (n_3340, n_105, n_188);
  nand g257 (n_3341, n_105, n_3339);
  nand g258 (n_3342, n_188, n_3339);
  nand g259 (n_3344, n_3340, n_3341, n_3342);
  xor g260 (n_3343, n_105, n_188);
  xor g261 (Z[42], n_3339, n_3343);
  nand g262 (n_3345, n_104, n_187);
  nand g263 (n_3346, n_104, n_3344);
  nand g264 (n_3347, n_187, n_3344);
  nand g265 (n_3349, n_3345, n_3346, n_3347);
  xor g266 (n_3348, n_104, n_187);
  xor g267 (Z[43], n_3344, n_3348);
  nand g268 (n_3350, n_103, n_186);
  nand g269 (n_3351, n_103, n_3349);
  nand g270 (n_3352, n_186, n_3349);
  nand g271 (n_3354, n_3350, n_3351, n_3352);
  xor g272 (n_3353, n_103, n_186);
  xor g273 (Z[44], n_3349, n_3353);
  nand g274 (n_3355, n_102, n_185);
  nand g275 (n_3356, n_102, n_3354);
  nand g276 (n_3357, n_185, n_3354);
  nand g277 (n_3359, n_3355, n_3356, n_3357);
  xor g278 (n_3358, n_102, n_185);
  xor g279 (Z[45], n_3354, n_3358);
  nand g280 (n_3360, n_101, n_184);
  nand g281 (n_3361, n_101, n_3359);
  nand g282 (n_3362, n_184, n_3359);
  nand g283 (n_3364, n_3360, n_3361, n_3362);
  xor g284 (n_3363, n_101, n_184);
  xor g285 (Z[46], n_3359, n_3363);
  nand g286 (n_3365, n_100, n_183);
  nand g287 (n_3366, n_100, n_3364);
  nand g288 (n_3367, n_183, n_3364);
  nand g289 (n_3369, n_3365, n_3366, n_3367);
  xor g290 (n_3368, n_100, n_183);
  xor g291 (Z[47], n_3364, n_3368);
  nand g292 (n_3370, n_99, n_182);
  nand g293 (n_3371, n_99, n_3369);
  nand g294 (n_3372, n_182, n_3369);
  nand g295 (n_3374, n_3370, n_3371, n_3372);
  xor g296 (n_3373, n_99, n_182);
  xor g297 (Z[48], n_3369, n_3373);
  nand g298 (n_3375, n_98, n_181);
  nand g299 (n_3376, n_98, n_3374);
  nand g300 (n_3377, n_181, n_3374);
  nand g301 (n_3379, n_3375, n_3376, n_3377);
  xor g302 (n_3378, n_98, n_181);
  xor g303 (Z[49], n_3374, n_3378);
  nand g304 (n_3380, n_97, n_180);
  nand g305 (n_3381, n_97, n_3379);
  nand g306 (n_3382, n_180, n_3379);
  nand g307 (n_3384, n_3380, n_3381, n_3382);
  xor g308 (n_3383, n_97, n_180);
  xor g309 (Z[50], n_3379, n_3383);
  nand g310 (n_3385, n_96, n_179);
  nand g311 (n_3386, n_96, n_3384);
  nand g312 (n_3387, n_179, n_3384);
  nand g313 (n_3389, n_3385, n_3386, n_3387);
  xor g314 (n_3388, n_96, n_179);
  xor g315 (Z[51], n_3384, n_3388);
  nand g316 (n_3390, n_95, n_178);
  nand g317 (n_3391, n_95, n_3389);
  nand g318 (n_3392, n_178, n_3389);
  nand g319 (n_3394, n_3390, n_3391, n_3392);
  xor g320 (n_3393, n_95, n_178);
  xor g321 (Z[52], n_3389, n_3393);
  nand g322 (n_3395, n_94, n_177);
  nand g323 (n_3396, n_94, n_3394);
  nand g324 (n_3397, n_177, n_3394);
  nand g325 (n_3399, n_3395, n_3396, n_3397);
  xor g326 (n_3398, n_94, n_177);
  xor g327 (Z[53], n_3394, n_3398);
  nand g328 (n_3400, n_93, n_176);
  nand g329 (n_3401, n_93, n_3399);
  nand g330 (n_3402, n_176, n_3399);
  nand g331 (n_3404, n_3400, n_3401, n_3402);
  xor g332 (n_3403, n_93, n_176);
  xor g333 (Z[54], n_3399, n_3403);
  nand g334 (n_3405, n_92, n_175);
  nand g335 (n_3406, n_92, n_3404);
  nand g336 (n_3407, n_175, n_3404);
  nand g337 (n_3409, n_3405, n_3406, n_3407);
  xor g338 (n_3408, n_92, n_175);
  xor g339 (Z[55], n_3404, n_3408);
  nand g340 (n_3410, n_91, n_174);
  nand g341 (n_3411, n_91, n_3409);
  nand g342 (n_3412, n_174, n_3409);
  nand g343 (n_3414, n_3410, n_3411, n_3412);
  xor g344 (n_3413, n_91, n_174);
  xor g345 (Z[56], n_3409, n_3413);
  nand g346 (n_3415, n_90, n_173);
  nand g347 (n_3416, n_90, n_3414);
  nand g348 (n_3417, n_173, n_3414);
  nand g349 (n_3419, n_3415, n_3416, n_3417);
  xor g350 (n_3418, n_90, n_173);
  xor g351 (Z[57], n_3414, n_3418);
  nand g352 (n_3420, n_89, n_172);
  nand g353 (n_3421, n_89, n_3419);
  nand g354 (n_3422, n_172, n_3419);
  nand g355 (n_3424, n_3420, n_3421, n_3422);
  xor g356 (n_3423, n_89, n_172);
  xor g357 (Z[58], n_3419, n_3423);
  nand g358 (n_3425, n_88, n_171);
  nand g359 (n_3426, n_88, n_3424);
  nand g360 (n_3427, n_171, n_3424);
  nand g361 (n_3429, n_3425, n_3426, n_3427);
  xor g362 (n_3428, n_88, n_171);
  xor g363 (Z[59], n_3424, n_3428);
  nand g364 (n_3430, n_87, n_170);
  nand g365 (n_3431, n_87, n_3429);
  nand g366 (n_3432, n_170, n_3429);
  nand g367 (n_3434, n_3430, n_3431, n_3432);
  xor g368 (n_3433, n_87, n_170);
  xor g369 (Z[60], n_3429, n_3433);
  nand g370 (n_3435, n_86, n_169);
  nand g371 (n_3436, n_86, n_3434);
  nand g372 (n_3437, n_169, n_3434);
  nand g373 (n_3439, n_3435, n_3436, n_3437);
  xor g374 (n_3438, n_86, n_169);
  xor g375 (Z[61], n_3434, n_3438);
  nand g376 (n_3440, n_85, n_168);
  nand g377 (n_3441, n_85, n_3439);
  nand g378 (n_3442, n_168, n_3439);
  nand g379 (n_3444, n_3440, n_3441, n_3442);
  xor g380 (n_3443, n_85, n_168);
  xor g381 (Z[62], n_3439, n_3443);
  nand g382 (n_3445, n_84, n_167);
  nand g383 (n_3446, n_84, n_3444);
  nand g384 (n_3447, n_167, n_3444);
  nand g385 (n_3449, n_3445, n_3446, n_3447);
  xor g386 (n_3448, n_84, n_167);
  xor g387 (Z[63], n_3444, n_3448);
  nand g388 (n_3450, n_83, n_166);
  nand g389 (n_3451, n_83, n_3449);
  nand g390 (n_3452, n_166, n_3449);
  nand g391 (n_3454, n_3450, n_3451, n_3452);
  xor g392 (n_3453, n_83, n_166);
  xor g393 (Z[64], n_3449, n_3453);
  nand g394 (n_3455, n_82, n_165);
  nand g395 (n_3456, n_82, n_3454);
  nand g396 (n_3457, n_165, n_3454);
  nand g397 (n_3459, n_3455, n_3456, n_3457);
  xor g398 (n_3458, n_82, n_165);
  xor g399 (Z[65], n_3454, n_3458);
  nand g400 (n_3460, n_81, n_164);
  nand g401 (n_3461, n_81, n_3459);
  nand g402 (n_3462, n_164, n_3459);
  nand g403 (n_3464, n_3460, n_3461, n_3462);
  xor g404 (n_3463, n_81, n_164);
  xor g405 (Z[66], n_3459, n_3463);
  nand g406 (n_3465, n_80, n_163);
  nand g407 (n_3466, n_80, n_3464);
  nand g408 (n_3467, n_163, n_3464);
  nand g409 (n_3469, n_3465, n_3466, n_3467);
  xor g410 (n_3468, n_80, n_163);
  xor g411 (Z[67], n_3464, n_3468);
  nand g412 (n_3470, n_79, n_162);
  nand g413 (n_3471, n_79, n_3469);
  nand g414 (n_3472, n_162, n_3469);
  nand g415 (n_3474, n_3470, n_3471, n_3472);
  xor g416 (n_3473, n_79, n_162);
  xor g417 (Z[68], n_3469, n_3473);
  nand g418 (n_3475, n_78, n_161);
  nand g419 (n_3476, n_78, n_3474);
  nand g420 (n_3477, n_161, n_3474);
  nand g421 (n_3479, n_3475, n_3476, n_3477);
  xor g422 (n_3478, n_78, n_161);
  xor g423 (Z[69], n_3474, n_3478);
  nand g424 (n_3480, n_77, n_160);
  nand g425 (n_3481, n_77, n_3479);
  nand g426 (n_3482, n_160, n_3479);
  nand g427 (n_3484, n_3480, n_3481, n_3482);
  xor g428 (n_3483, n_77, n_160);
  xor g429 (Z[70], n_3479, n_3483);
  nand g430 (n_3485, n_76, n_159);
  nand g431 (n_3486, n_76, n_3484);
  nand g432 (n_3487, n_159, n_3484);
  nand g433 (n_3489, n_3485, n_3486, n_3487);
  xor g434 (n_3488, n_76, n_159);
  xor g435 (Z[71], n_3484, n_3488);
  nand g436 (n_3490, n_75, n_158);
  nand g437 (n_3491, n_75, n_3489);
  nand g438 (n_3492, n_158, n_3489);
  nand g439 (n_3494, n_3490, n_3491, n_3492);
  xor g440 (n_3493, n_75, n_158);
  xor g441 (Z[72], n_3489, n_3493);
  nand g442 (n_3495, n_74, n_157);
  nand g443 (n_3496, n_74, n_3494);
  nand g444 (n_3497, n_157, n_3494);
  nand g445 (n_3499, n_3495, n_3496, n_3497);
  xor g446 (n_3498, n_74, n_157);
  xor g447 (Z[73], n_3494, n_3498);
  nand g448 (n_3500, n_73, n_156);
  nand g449 (n_3501, n_73, n_3499);
  nand g450 (n_3502, n_156, n_3499);
  nand g451 (n_3504, n_3500, n_3501, n_3502);
  xor g452 (n_3503, n_73, n_156);
  xor g453 (Z[74], n_3499, n_3503);
  nand g454 (n_3505, n_72, n_155);
  nand g455 (n_3506, n_72, n_3504);
  nand g456 (n_3507, n_155, n_3504);
  nand g457 (n_3509, n_3505, n_3506, n_3507);
  xor g458 (n_3508, n_72, n_155);
  xor g459 (Z[75], n_3504, n_3508);
  nand g460 (n_3510, n_71, n_154);
  nand g461 (n_3511, n_71, n_3509);
  nand g462 (n_3512, n_154, n_3509);
  nand g463 (n_3514, n_3510, n_3511, n_3512);
  xor g464 (n_3513, n_71, n_154);
  xor g465 (Z[76], n_3509, n_3513);
  nand g466 (n_3515, n_70, n_153);
  nand g467 (n_3516, n_70, n_3514);
  nand g468 (n_3517, n_153, n_3514);
  nand g469 (n_3519, n_3515, n_3516, n_3517);
  xor g470 (n_3518, n_70, n_153);
  xor g471 (Z[77], n_3514, n_3518);
  nand g472 (n_3520, n_69, n_152);
  nand g473 (n_3521, n_69, n_3519);
  nand g474 (n_3522, n_152, n_3519);
  nand g475 (n_3524, n_3520, n_3521, n_3522);
  xor g476 (n_3523, n_69, n_152);
  xor g477 (Z[78], n_3519, n_3523);
  nand g478 (n_3525, n_68, n_151);
  nand g479 (n_3526, n_68, n_3524);
  nand g480 (n_3527, n_151, n_3524);
  nand g481 (n_3529, n_3525, n_3526, n_3527);
  xor g482 (n_3528, n_68, n_151);
  xor g483 (Z[79], n_3524, n_3528);
  nand g486 (n_3532, n_150, n_3529);
  nand g487 (n_3534, n_3530, n_3531, n_3532);
  xor g489 (Z[80], n_3529, n_3533);
  nand g492 (n_3537, A[62], n_3534);
  nand g493 (n_3539, n_3535, n_3536, n_3537);
  xor g495 (Z[81], n_3534, n_3538);
  or g3482 (n_322, wc, wc0, n_142);
  not gc0 (wc0, n_1181);
  not gc (wc, n_1195);
  or g3483 (n_331, wc1, wc2, n_316);
  not gc2 (wc2, n_1195);
  not gc1 (wc1, n_1214);
  or g3484 (n_344, wc3, n_321, n_316);
  not gc3 (wc3, n_1242);
  or g3485 (n_361, wc4, wc5, n_321);
  not gc5 (wc5, n_1277);
  not gc4 (wc4, n_1278);
  or g3486 (n_383, wc6, wc7, n_321);
  not gc7 (wc7, n_1325);
  not gc6 (wc6, n_1326);
  or g3487 (n_144, wc8, wc9, n_316);
  not gc9 (wc9, n_1326);
  not gc8 (wc8, n_1373);
  or g3488 (n_458, wc10, wc11, n_321);
  not gc11 (wc11, n_1502);
  not gc10 (wc10, n_1503);
  or g3489 (n_486, wc12, wc13, n_330);
  not gc13 (wc13, n_1442);
  not gc12 (wc12, n_1566);
  or g3490 (n_512, wc14, wc15, n_343);
  not gc15 (wc15, n_1506);
  not gc14 (wc14, n_1630);
  or g3491 (n_540, wc16, wc17, n_360);
  not gc17 (wc17, n_1435);
  not gc16 (wc16, n_1694);
  or g3492 (n_568, wc18, wc19, n_381);
  not gc19 (wc19, n_1499);
  not gc18 (wc18, n_1758);
  or g3493 (n_596, wc20, wc21, n_406);
  not gc21 (wc21, n_1563);
  not gc20 (wc20, n_1822);
  xnor g3494 (n_2872, A[63], A[61]);
  or g3495 (n_2873, wc22, A[63]);
  not gc22 (wc22, A[61]);
  or g3496 (n_2875, wc23, A[63]);
  not gc23 (wc23, A[57]);
  xnor g3497 (n_2912, A[62], A[50]);
  or g3498 (n_2913, wc24, A[62]);
  not gc24 (wc24, A[50]);
  xnor g3499 (n_1120, n_2848, A[60]);
  or g3500 (n_3014, wc25, A[60]);
  not gc25 (wc25, A[58]);
  or g3501 (n_3015, wc26, A[60]);
  not gc26 (wc26, A[52]);
  xnor g3503 (n_1166, n_2712, A[62]);
  or g3504 (n_3106, wc27, A[62]);
  not gc27 (wc27, A[58]);
  or g3505 (n_3107, wc28, A[62]);
  not gc28 (wc28, A[60]);
  or g3506 (n_3115, wc29, A[63]);
  not gc29 (wc29, A[59]);
  or g3508 (n_3121, A[60], wc30);
  not gc30 (wc30, A[62]);
  or g3509 (n_3127, wc31, A[63]);
  not gc31 (wc31, A[60]);
  or g3510 (n_3535, wc32, A[63]);
  not gc32 (wc32, A[62]);
  xnor g3511 (n_3538, A[63], A[62]);
  or g3512 (n_412, wc33, wc34, n_321);
  not gc34 (wc34, n_1382);
  not gc33 (wc33, n_1383);
  or g3513 (n_2971, A[62], wc35);
  not gc35 (wc35, n_1094);
  xnor g3514 (n_1140, n_2712, n_1036);
  or g3515 (n_3054, A[60], wc36);
  not gc36 (wc36, n_1036);
  or g3516 (n_3087, A[62], wc37);
  not gc37 (wc37, n_1154);
  xnor g3517 (n_2884, n_1049, A[63]);
  or g3518 (n_2885, A[63], wc38);
  not gc38 (wc38, n_1049);
  or g3519 (n_2887, A[63], wc39);
  not gc39 (wc39, n_1050);
  or g3520 (n_2914, A[62], wc40);
  not gc40 (wc40, n_1065);
  xnor g3521 (n_2968, n_1065, A[62]);
  xnor g3522 (n_69, n_2776, n_1173);
  or g3523 (n_3122, A[60], wc41);
  not gc41 (wc41, n_1173);
  or g3524 (n_3530, A[62], wc42);
  not gc42 (wc42, n_150);
  xnor g3525 (n_3533, n_150, A[62]);
  or g3527 (n_3146, wc43, n_1181);
  not gc43 (wc43, A[1]);
  or g3528 (n_3147, wc44, n_1181);
  not gc44 (wc44, A[3]);
  xnor g3529 (Z[3], n_1176, n_1181);
  or g3530 (n_3531, A[62], wc45);
  not gc45 (wc45, n_3529);
  or g3531 (n_3536, A[63], wc46);
  not gc46 (wc46, n_3534);
  not g3532 (Z[82], n_3539);
endmodule

module mult_signed_const_15239_GENERIC(A, Z);
  input [63:0] A;
  output [82:0] Z;
  wire [63:0] A;
  wire [82:0] Z;
  mult_signed_const_15239_GENERIC_REAL g1(.A ({A[63:2], A[0], A[0]}),
       .Z (Z));
endmodule

module mult_signed_const_15762_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [65:0] A;
  output [84:0] Z;
  wire [65:0] A;
  wire [84:0] Z;
  wire n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77;
  wire n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85;
  wire n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93;
  wire n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101;
  wire n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109;
  wire n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117;
  wire n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125;
  wire n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133;
  wire n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150, n_151, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231;
  wire n_232, n_233, n_234, n_323, n_324, n_325, n_326, n_327;
  wire n_328, n_329, n_330, n_331, n_332, n_333, n_334, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351;
  wire n_352, n_353, n_354, n_355, n_356, n_357, n_358, n_359;
  wire n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367;
  wire n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431;
  wire n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439;
  wire n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447;
  wire n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455;
  wire n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463;
  wire n_464, n_465, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538;
  wire n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562;
  wire n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_577, n_578, n_579;
  wire n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587;
  wire n_588, n_589, n_590, n_591, n_592, n_593, n_594, n_595;
  wire n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603;
  wire n_605, n_606, n_607, n_608, n_609, n_610, n_611, n_612;
  wire n_613, n_614, n_615, n_616, n_617, n_618, n_619, n_620;
  wire n_621, n_622, n_623, n_624, n_625, n_626, n_627, n_628;
  wire n_629, n_630, n_631, n_633, n_634, n_635, n_636, n_637;
  wire n_638, n_639, n_640, n_641, n_642, n_643, n_644, n_645;
  wire n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
  wire n_654, n_655, n_656, n_657, n_658, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669;
  wire n_670, n_671, n_672, n_673, n_674, n_675, n_676, n_677;
  wire n_678, n_679, n_680, n_681, n_682, n_683, n_684, n_685;
  wire n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693;
  wire n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701;
  wire n_702, n_703, n_704, n_705, n_706, n_707, n_708, n_709;
  wire n_710, n_711, n_712, n_713, n_714, n_715, n_716, n_717;
  wire n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725;
  wire n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733;
  wire n_734, n_735, n_736, n_737, n_738, n_739, n_740, n_741;
  wire n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749;
  wire n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757;
  wire n_758, n_759, n_760, n_761, n_762, n_763, n_764, n_765;
  wire n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_779, n_780, n_781;
  wire n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789;
  wire n_790, n_791, n_792, n_793, n_794, n_795, n_796, n_797;
  wire n_798, n_799, n_801, n_802, n_803, n_804, n_805, n_806;
  wire n_807, n_808, n_809, n_810, n_811, n_812, n_813, n_815;
  wire n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823;
  wire n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831;
  wire n_832, n_833, n_834, n_835, n_836, n_837, n_838, n_839;
  wire n_840, n_841, n_842, n_843, n_844, n_845, n_846, n_847;
  wire n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855;
  wire n_857, n_858, n_859, n_860, n_861, n_862, n_863, n_864;
  wire n_865, n_866, n_867, n_868, n_869, n_871, n_872, n_873;
  wire n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897;
  wire n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905;
  wire n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913;
  wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
  wire n_922, n_923, n_924, n_925, n_927, n_928, n_929, n_930;
  wire n_931, n_932, n_933, n_934, n_935, n_936, n_937, n_938;
  wire n_941, n_942, n_943, n_944, n_945, n_946, n_947, n_948;
  wire n_949, n_950, n_951, n_952, n_955, n_956, n_957, n_958;
  wire n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966;
  wire n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976;
  wire n_977, n_978, n_979, n_980, n_982, n_983, n_984, n_985;
  wire n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993;
  wire n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001;
  wire n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1010;
  wire n_1011, n_1012, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019;
  wire n_1020, n_1021, n_1022, n_1025, n_1028, n_1029, n_1030, n_1031;
  wire n_1032, n_1033, n_1034, n_1035, n_1036, n_1038, n_1040, n_1041;
  wire n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049;
  wire n_1050, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059;
  wire n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1070;
  wire n_1071, n_1072, n_1073, n_1075, n_1076, n_1077, n_1078, n_1079;
  wire n_1080, n_1081, n_1082, n_1083, n_1086, n_1087, n_1088, n_1089;
  wire n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097;
  wire n_1098, n_1101, n_1102, n_1103, n_1105, n_1106, n_1107, n_1108;
  wire n_1109, n_1110, n_1111, n_1112, n_1113, n_1116, n_1118, n_1119;
  wire n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1130;
  wire n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138;
  wire n_1139, n_1141, n_1142, n_1143, n_1145, n_1146, n_1147, n_1148;
  wire n_1149, n_1150, n_1153, n_1155, n_1156, n_1157, n_1158, n_1159;
  wire n_1160, n_1161, n_1163, n_1166, n_1167, n_1168, n_1169, n_1170;
  wire n_1176, n_1177, n_1178, n_1179, n_1183, n_1184, n_1185, n_1186;
  wire n_1190, n_1191, n_1192, n_1193, n_1195, n_1197, n_1198, n_1202;
  wire n_1203, n_1205, n_1206, n_1209, n_1212, n_1213, n_1214, n_1215;
  wire n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1224, n_1225;
  wire n_1226, n_1227, n_1230, n_1232, n_1233, n_1234, n_1235, n_1236;
  wire n_1237, n_1238, n_1240, n_1242, n_1243, n_1244, n_1245, n_1246;
  wire n_1247, n_1250, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257;
  wire n_1258, n_1259, n_1262, n_1264, n_1265, n_1266, n_1267, n_1268;
  wire n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276;
  wire n_1277, n_1278, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285;
  wire n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293;
  wire n_1296, n_1297, n_1298, n_1300, n_1301, n_1302, n_1303, n_1304;
  wire n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312;
  wire n_1315, n_1316, n_1317, n_1320, n_1321, n_1322, n_1323, n_1324;
  wire n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332;
  wire n_1333, n_1334, n_1335, n_1336, n_1339, n_1342, n_1343, n_1344;
  wire n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352;
  wire n_1353, n_1354, n_1355, n_1356, n_1363, n_1364, n_1365, n_1366;
  wire n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374;
  wire n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382;
  wire n_1384, n_1387, n_1388, n_1392, n_1393, n_1394, n_1395, n_1396;
  wire n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404;
  wire n_1405, n_1406, n_1407, n_1408, n_1409, n_1415, n_1418, n_1419;
  wire n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427;
  wire n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435;
  wire n_1436, n_1437, n_1438, n_1440, n_1441, n_1442, n_1443, n_1444;
  wire n_1445, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453;
  wire n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461;
  wire n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469;
  wire n_1470, n_1471, n_1474, n_1475, n_1478, n_1479, n_1480, n_1481;
  wire n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489;
  wire n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
  wire n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1507, n_1508;
  wire n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518;
  wire n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526;
  wire n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534;
  wire n_1535, n_1540, n_1541, n_1542, n_1544, n_1545, n_1546, n_1547;
  wire n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555;
  wire n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563;
  wire n_1564, n_1565, n_1566, n_1567, n_1572, n_1573, n_1576, n_1577;
  wire n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585;
  wire n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593;
  wire n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1602, n_1603;
  wire n_1604, n_1605, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613;
  wire n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621;
  wire n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629;
  wire n_1630, n_1631, n_1636, n_1637, n_1640, n_1641, n_1642, n_1643;
  wire n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651;
  wire n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659;
  wire n_1660, n_1661, n_1662, n_1663, n_1664, n_1666, n_1668, n_1671;
  wire n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679;
  wire n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687;
  wire n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695;
  wire n_1696, n_1698, n_1700, n_1701, n_1704, n_1705, n_1706, n_1707;
  wire n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715;
  wire n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723;
  wire n_1724, n_1725, n_1726, n_1727, n_1728, n_1730, n_1731, n_1732;
  wire n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742;
  wire n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750;
  wire n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758;
  wire n_1759, n_1760, n_1762, n_1764, n_1765, n_1768, n_1769, n_1770;
  wire n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778;
  wire n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786;
  wire n_1787, n_1788, n_1789, n_1790, n_1791, n_1796, n_1799, n_1800;
  wire n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1826, n_1828, n_1829, n_1832, n_1833, n_1834, n_1835, n_1836;
  wire n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844;
  wire n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852;
  wire n_1853, n_1854, n_1855, n_1860, n_1861, n_1864, n_1865, n_1866;
  wire n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874;
  wire n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882;
  wire n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890;
  wire n_1892, n_1893, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901;
  wire n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909;
  wire n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917;
  wire n_1918, n_1919, n_1924, n_1925, n_1928, n_1929, n_1930, n_1931;
  wire n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939;
  wire n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947;
  wire n_1948, n_1949, n_1950, n_1951, n_1954, n_1956, n_1957, n_1960;
  wire n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968;
  wire n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976;
  wire n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1986;
  wire n_1988, n_1989, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997;
  wire n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005;
  wire n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013;
  wire n_2014, n_2015, n_2018, n_2020, n_2021, n_2024, n_2025, n_2026;
  wire n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034;
  wire n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042;
  wire n_2043, n_2044, n_2045, n_2046, n_2047, n_2050, n_2052, n_2053;
  wire n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063;
  wire n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071;
  wire n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079;
  wire n_2082, n_2084, n_2085, n_2088, n_2089, n_2090, n_2091, n_2092;
  wire n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100;
  wire n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108;
  wire n_2109, n_2110, n_2111, n_2114, n_2116, n_2117, n_2120, n_2121;
  wire n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129;
  wire n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137;
  wire n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2146, n_2148;
  wire n_2149, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158;
  wire n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166;
  wire n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174;
  wire n_2175, n_2176, n_2177, n_2178, n_2180, n_2183, n_2184, n_2185;
  wire n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193;
  wire n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201;
  wire n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209;
  wire n_2210, n_2212, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220;
  wire n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228;
  wire n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236;
  wire n_2237, n_2239, n_2240, n_2242, n_2244, n_2247, n_2248, n_2249;
  wire n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257;
  wire n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265;
  wire n_2266, n_2267, n_2268, n_2269, n_2271, n_2272, n_2274, n_2276;
  wire n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286;
  wire n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294;
  wire n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302;
  wire n_2303, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318;
  wire n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326;
  wire n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334;
  wire n_2335, n_2344, n_2345, n_2346, n_2348, n_2349, n_2350, n_2351;
  wire n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359;
  wire n_2360, n_2361, n_2362, n_2363, n_2364, n_2367, n_2371, n_2374;
  wire n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382;
  wire n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390;
  wire n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2399, n_2403;
  wire n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413;
  wire n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421;
  wire n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2430, n_2431;
  wire n_2436, n_2437, n_2438, n_2440, n_2441, n_2442, n_2443, n_2444;
  wire n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452;
  wire n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2462;
  wire n_2463, n_2468, n_2469, n_2470, n_2472, n_2473, n_2474, n_2475;
  wire n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483;
  wire n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491;
  wire n_2495, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506;
  wire n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514;
  wire n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522;
  wire n_2523, n_2527, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537;
  wire n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545;
  wire n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553;
  wire n_2554, n_2555, n_2560, n_2562, n_2563, n_2564, n_2565, n_2567;
  wire n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575;
  wire n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583;
  wire n_2584, n_2585, n_2586, n_2587, n_2592, n_2594, n_2595, n_2596;
  wire n_2597, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605;
  wire n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613;
  wire n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2624, n_2625;
  wire n_2626, n_2627, n_2628, n_2629, n_2630, n_2632, n_2633, n_2634;
  wire n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642;
  wire n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650;
  wire n_2651, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662;
  wire n_2664, n_2665, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672;
  wire n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680;
  wire n_2681, n_2682, n_2683, n_2688, n_2689, n_2691, n_2692, n_2693;
  wire n_2694, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702;
  wire n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710;
  wire n_2711, n_2712, n_2713, n_2714, n_2715, n_2720, n_2721, n_2723;
  wire n_2724, n_2725, n_2726, n_2728, n_2729, n_2730, n_2731, n_2732;
  wire n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740;
  wire n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2750;
  wire n_2751, n_2752, n_2753, n_2754, n_2756, n_2758, n_2762, n_2763;
  wire n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771;
  wire n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779;
  wire n_2782, n_2783, n_2784, n_2785, n_2786, n_2788, n_2790, n_2792;
  wire n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800;
  wire n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808;
  wire n_2809, n_2810, n_2811, n_2816, n_2817, n_2818, n_2819, n_2824;
  wire n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832;
  wire n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, n_2840;
  wire n_2841, n_2842, n_2843, n_2848, n_2849, n_2850, n_2851, n_2856;
  wire n_2857, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865;
  wire n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873;
  wire n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2883, n_2884;
  wire n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892;
  wire n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900;
  wire n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908;
  wire n_2909, n_2910, n_2911, n_2915, n_2916, n_2917, n_2918, n_2919;
  wire n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927;
  wire n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935;
  wire n_2936, n_2937, n_2938, n_2939, n_2945, n_2946, n_2947, n_2948;
  wire n_2949, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, n_2957;
  wire n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965;
  wire n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973;
  wire n_2974, n_2975, n_2980, n_2981, n_2983, n_2984, n_2985, n_2986;
  wire n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994;
  wire n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, n_3002;
  wire n_3003, n_3004, n_3007, n_3012, n_3013, n_3014, n_3015, n_3016;
  wire n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024;
  wire n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3036;
  wire n_3038, n_3039, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047;
  wire n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055;
  wire n_3056, n_3057, n_3058, n_3059, n_3060, n_3062, n_3064, n_3067;
  wire n_3068, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076;
  wire n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3088;
  wire n_3091, n_3092, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099;
  wire n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107;
  wire n_3108, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120;
  wire n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3136;
  wire n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144;
  wire n_3145, n_3146, n_3147, n_3154, n_3155, n_3156, n_3158, n_3159;
  wire n_3160, n_3161, n_3162, n_3163, n_3170, n_3171, n_3172, n_3173;
  wire n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3183, n_3186;
  wire n_3187, n_3188, n_3189, n_3190, n_3191, n_3196, n_3197, n_3198;
  wire n_3199, n_3200, n_3201, n_3202, n_3203, n_3206, n_3207, n_3208;
  wire n_3209, n_3210, n_3211, n_3216, n_3217, n_3218, n_3219, n_3220;
  wire n_3221, n_3222, n_3223, n_3226, n_3227, n_3246, n_3247, n_3248;
  wire n_3249, n_3250, n_3251, n_3252, n_3254, n_3255, n_3256, n_3257;
  wire n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265;
  wire n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273;
  wire n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281;
  wire n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289;
  wire n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297;
  wire n_3298, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305;
  wire n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313;
  wire n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321;
  wire n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329;
  wire n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337;
  wire n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345;
  wire n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353;
  wire n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361;
  wire n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369;
  wire n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377;
  wire n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385;
  wire n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393;
  wire n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401;
  wire n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409;
  wire n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417;
  wire n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425;
  wire n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433;
  wire n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441;
  wire n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449;
  wire n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457;
  wire n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465;
  wire n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473;
  wire n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481;
  wire n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489;
  wire n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497;
  wire n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505;
  wire n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513;
  wire n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521;
  wire n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529;
  wire n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537;
  wire n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545;
  wire n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553;
  wire n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561;
  wire n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569;
  wire n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577;
  wire n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585;
  wire n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593;
  wire n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601;
  wire n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609;
  wire n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617;
  wire n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625;
  wire n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633;
  wire n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641;
  wire n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g524 (n_232, A[4], A[0]);
  and g2 (n_146, A[4], A[0]);
  xor g525 (n_1212, A[1], A[5]);
  xor g526 (n_231, n_1212, A[3]);
  nand g3 (n_1213, A[1], A[5]);
  nand g527 (n_1214, A[3], A[5]);
  nand g528 (n_1215, A[1], A[3]);
  nand g529 (n_145, n_1213, n_1214, n_1215);
  xor g530 (n_323, A[6], A[4]);
  and g531 (n_324, A[6], A[4]);
  xor g532 (Z[2], A[0], A[2]);
  xor g533 (n_230, Z[2], n_323);
  nand g534 (n_1217, A[0], A[2]);
  nand g4 (n_1218, n_323, A[2]);
  nand g5 (n_1219, A[0], n_323);
  nand g535 (n_144, n_1217, n_1218, n_1219);
  xor g536 (n_1220, A[1], A[7]);
  xor g537 (n_325, n_1220, A[5]);
  nand g538 (n_1221, A[1], A[7]);
  nand g539 (n_1222, A[5], A[7]);
  nand g6 (n_327, n_1221, n_1222, n_1213);
  xor g541 (n_1224, A[3], n_324);
  xor g542 (n_229, n_1224, n_325);
  nand g543 (n_1225, A[3], n_324);
  nand g544 (n_1226, n_325, n_324);
  nand g545 (n_1227, A[3], n_325);
  nand g546 (n_143, n_1225, n_1226, n_1227);
  xor g547 (n_326, A[8], A[6]);
  and g548 (n_329, A[8], A[6]);
  xor g550 (n_328, n_232, A[2]);
  nand g552 (n_1230, A[2], A[4]);
  xor g555 (n_1232, n_326, n_327);
  xor g556 (n_228, n_1232, n_328);
  nand g557 (n_1233, n_326, n_327);
  nand g558 (n_1234, n_328, n_327);
  nand g559 (n_1235, n_326, n_328);
  nand g560 (n_142, n_1233, n_1234, n_1235);
  xor g561 (n_1236, A[1], A[9]);
  xor g562 (n_331, n_1236, A[7]);
  nand g563 (n_1237, A[1], A[9]);
  nand g564 (n_1238, A[7], A[9]);
  nand g566 (n_334, n_1237, n_1238, n_1221);
  xor g567 (n_1240, A[5], A[3]);
  xor g568 (n_332, n_1240, n_329);
  nand g570 (n_1242, n_329, A[3]);
  nand g571 (n_1243, A[5], n_329);
  nand g572 (n_336, n_1214, n_1242, n_1243);
  xor g573 (n_1244, n_330, n_331);
  xor g574 (n_227, n_1244, n_332);
  nand g575 (n_1245, n_330, n_331);
  nand g576 (n_1246, n_332, n_331);
  nand g577 (n_1247, n_330, n_332);
  nand g578 (n_141, n_1245, n_1246, n_1247);
  xor g579 (n_333, A[10], A[8]);
  and g580 (n_338, A[10], A[8]);
  xor g582 (n_335, n_323, A[0]);
  nand g584 (n_1250, A[0], A[6]);
  xor g587 (n_1252, A[2], n_333);
  xor g588 (n_337, n_1252, n_334);
  nand g589 (n_1253, A[2], n_333);
  nand g590 (n_1254, n_334, n_333);
  nand g591 (n_1255, A[2], n_334);
  nand g592 (n_342, n_1253, n_1254, n_1255);
  xor g593 (n_1256, n_335, n_336);
  xor g594 (n_226, n_1256, n_337);
  nand g595 (n_1257, n_335, n_336);
  nand g596 (n_1258, n_337, n_336);
  nand g597 (n_1259, n_335, n_337);
  nand g598 (n_140, n_1257, n_1258, n_1259);
  xor g600 (n_340, n_1236, A[5]);
  nand g602 (n_1262, A[5], A[9]);
  nand g604 (n_345, n_1237, n_1262, n_1213);
  xor g605 (n_1264, A[11], A[7]);
  xor g606 (n_341, n_1264, A[3]);
  nand g607 (n_1265, A[11], A[7]);
  nand g608 (n_1266, A[3], A[7]);
  nand g609 (n_1267, A[11], A[3]);
  nand g610 (n_346, n_1265, n_1266, n_1267);
  xor g611 (n_1268, n_338, n_339);
  xor g612 (n_343, n_1268, n_340);
  nand g613 (n_1269, n_338, n_339);
  nand g614 (n_1270, n_340, n_339);
  nand g615 (n_1271, n_338, n_340);
  nand g616 (n_349, n_1269, n_1270, n_1271);
  xor g617 (n_1272, n_341, n_342);
  xor g618 (n_225, n_1272, n_343);
  nand g619 (n_1273, n_341, n_342);
  nand g620 (n_1274, n_343, n_342);
  nand g621 (n_1275, n_341, n_343);
  nand g622 (n_139, n_1273, n_1274, n_1275);
  xor g623 (n_344, A[10], A[6]);
  and g624 (n_351, A[10], A[6]);
  xor g625 (n_1276, A[4], A[8]);
  xor g626 (n_347, n_1276, A[0]);
  nand g627 (n_1277, A[4], A[8]);
  nand g628 (n_1278, A[0], A[8]);
  xor g631 (n_1280, A[12], A[2]);
  xor g632 (n_348, n_1280, n_344);
  nand g633 (n_1281, A[12], A[2]);
  nand g634 (n_1282, n_344, A[2]);
  nand g635 (n_1283, A[12], n_344);
  nand g636 (n_355, n_1281, n_1282, n_1283);
  xor g637 (n_1284, n_345, n_346);
  xor g638 (n_350, n_1284, n_347);
  nand g639 (n_1285, n_345, n_346);
  nand g640 (n_1286, n_347, n_346);
  nand g641 (n_1287, n_345, n_347);
  nand g642 (n_357, n_1285, n_1286, n_1287);
  xor g643 (n_1288, n_348, n_349);
  xor g644 (n_224, n_1288, n_350);
  nand g645 (n_1289, n_348, n_349);
  nand g646 (n_1290, n_350, n_349);
  nand g647 (n_1291, n_348, n_350);
  nand g648 (n_138, n_1289, n_1290, n_1291);
  xor g649 (n_1292, A[1], A[11]);
  xor g650 (n_354, n_1292, A[7]);
  nand g651 (n_1293, A[1], A[11]);
  nand g654 (n_360, n_1293, n_1265, n_1221);
  xor g655 (n_1296, A[5], A[13]);
  xor g656 (n_353, n_1296, A[9]);
  nand g657 (n_1297, A[5], A[13]);
  nand g658 (n_1298, A[9], A[13]);
  nand g660 (n_361, n_1297, n_1298, n_1262);
  xor g661 (n_1300, A[3], n_351);
  xor g662 (n_356, n_1300, n_352);
  nand g663 (n_1301, A[3], n_351);
  nand g664 (n_1302, n_352, n_351);
  nand g665 (n_1303, A[3], n_352);
  nand g666 (n_364, n_1301, n_1302, n_1303);
  xor g667 (n_1304, n_353, n_354);
  xor g668 (n_358, n_1304, n_355);
  nand g669 (n_1305, n_353, n_354);
  nand g670 (n_1306, n_355, n_354);
  nand g671 (n_1307, n_353, n_355);
  nand g672 (n_366, n_1305, n_1306, n_1307);
  xor g673 (n_1308, n_356, n_357);
  xor g674 (n_223, n_1308, n_358);
  nand g675 (n_1309, n_356, n_357);
  nand g676 (n_1310, n_358, n_357);
  nand g677 (n_1311, n_356, n_358);
  nand g678 (n_137, n_1309, n_1310, n_1311);
  xor g679 (n_359, A[14], A[8]);
  and g680 (n_368, A[14], A[8]);
  xor g681 (n_1312, A[0], A[6]);
  xor g682 (n_362, n_1312, A[10]);
  nand g685 (n_1315, A[0], A[10]);
  xor g687 (n_1316, A[4], A[12]);
  xor g688 (n_363, n_1316, A[2]);
  nand g689 (n_1317, A[4], A[12]);
  nand g692 (n_372, n_1317, n_1281, n_1230);
  xor g693 (n_1320, n_359, n_360);
  xor g694 (n_365, n_1320, n_361);
  nand g695 (n_1321, n_359, n_360);
  nand g696 (n_1322, n_361, n_360);
  nand g697 (n_1323, n_359, n_361);
  nand g698 (n_374, n_1321, n_1322, n_1323);
  xor g699 (n_1324, n_362, n_363);
  xor g700 (n_367, n_1324, n_364);
  nand g701 (n_1325, n_362, n_363);
  nand g702 (n_1326, n_364, n_363);
  nand g703 (n_1327, n_362, n_364);
  nand g704 (n_377, n_1325, n_1326, n_1327);
  xor g705 (n_1328, n_365, n_366);
  xor g706 (n_222, n_1328, n_367);
  nand g707 (n_1329, n_365, n_366);
  nand g708 (n_1330, n_367, n_366);
  nand g709 (n_1331, n_365, n_367);
  nand g710 (n_136, n_1329, n_1330, n_1331);
  xor g711 (n_1332, A[1], A[15]);
  xor g712 (n_370, n_1332, A[13]);
  nand g713 (n_1333, A[1], A[15]);
  nand g714 (n_1334, A[13], A[15]);
  nand g715 (n_1335, A[1], A[13]);
  nand g716 (n_380, n_1333, n_1334, n_1335);
  xor g717 (n_1336, A[9], A[7]);
  xor g718 (n_371, n_1336, A[11]);
  nand g721 (n_1339, A[9], A[11]);
  nand g722 (n_379, n_1238, n_1265, n_1339);
  xor g724 (n_373, n_1240, n_368);
  nand g726 (n_1342, n_368, A[3]);
  nand g727 (n_1343, A[5], n_368);
  nand g728 (n_383, n_1214, n_1342, n_1343);
  xor g729 (n_1344, n_369, n_370);
  xor g730 (n_375, n_1344, n_371);
  nand g731 (n_1345, n_369, n_370);
  nand g732 (n_1346, n_371, n_370);
  nand g733 (n_1347, n_369, n_371);
  nand g734 (n_385, n_1345, n_1346, n_1347);
  xor g735 (n_1348, n_372, n_373);
  xor g736 (n_376, n_1348, n_374);
  nand g737 (n_1349, n_372, n_373);
  nand g738 (n_1350, n_374, n_373);
  nand g739 (n_1351, n_372, n_374);
  nand g740 (n_387, n_1349, n_1350, n_1351);
  xor g741 (n_1352, n_375, n_376);
  xor g742 (n_221, n_1352, n_377);
  nand g743 (n_1353, n_375, n_376);
  nand g744 (n_1354, n_377, n_376);
  nand g745 (n_1355, n_375, n_377);
  nand g746 (n_135, n_1353, n_1354, n_1355);
  xor g747 (n_378, A[16], A[14]);
  and g748 (n_389, A[16], A[14]);
  xor g749 (n_1356, A[10], A[0]);
  xor g750 (n_382, n_1356, A[8]);
  xor g756 (n_381, n_323, A[2]);
  nand g759 (n_1363, A[6], A[2]);
  xor g761 (n_1364, A[12], n_378);
  xor g762 (n_384, n_1364, n_379);
  nand g763 (n_1365, A[12], n_378);
  nand g764 (n_1366, n_379, n_378);
  nand g765 (n_1367, A[12], n_379);
  nand g766 (n_395, n_1365, n_1366, n_1367);
  xor g767 (n_1368, n_380, n_381);
  xor g768 (n_386, n_1368, n_382);
  nand g769 (n_1369, n_380, n_381);
  nand g770 (n_1370, n_382, n_381);
  nand g771 (n_1371, n_380, n_382);
  nand g772 (n_396, n_1369, n_1370, n_1371);
  xor g773 (n_1372, n_383, n_384);
  xor g774 (n_388, n_1372, n_385);
  nand g775 (n_1373, n_383, n_384);
  nand g776 (n_1374, n_385, n_384);
  nand g777 (n_1375, n_383, n_385);
  nand g778 (n_399, n_1373, n_1374, n_1375);
  xor g779 (n_1376, n_386, n_387);
  xor g780 (n_220, n_1376, n_388);
  nand g781 (n_1377, n_386, n_387);
  nand g782 (n_1378, n_388, n_387);
  nand g783 (n_1379, n_386, n_388);
  nand g784 (n_134, n_1377, n_1378, n_1379);
  xor g785 (n_1380, A[1], A[17]);
  xor g786 (n_391, n_1380, A[15]);
  nand g787 (n_1381, A[1], A[17]);
  nand g788 (n_1382, A[15], A[17]);
  nand g790 (n_402, n_1381, n_1382, n_1333);
  xor g791 (n_1384, A[11], A[9]);
  xor g792 (n_393, n_1384, A[13]);
  nand g795 (n_1387, A[11], A[13]);
  nand g796 (n_403, n_1339, n_1298, n_1387);
  xor g797 (n_1388, A[7], A[5]);
  xor g798 (n_392, n_1388, A[3]);
  nand g802 (n_405, n_1222, n_1214, n_1266);
  xor g803 (n_1392, n_389, n_390);
  xor g804 (n_397, n_1392, n_391);
  nand g805 (n_1393, n_389, n_390);
  nand g806 (n_1394, n_391, n_390);
  nand g807 (n_1395, n_389, n_391);
  nand g808 (n_408, n_1393, n_1394, n_1395);
  xor g809 (n_1396, n_392, n_393);
  xor g810 (n_398, n_1396, n_394);
  nand g811 (n_1397, n_392, n_393);
  nand g812 (n_1398, n_394, n_393);
  nand g813 (n_1399, n_392, n_394);
  nand g814 (n_409, n_1397, n_1398, n_1399);
  xor g815 (n_1400, n_395, n_396);
  xor g816 (n_400, n_1400, n_397);
  nand g817 (n_1401, n_395, n_396);
  nand g818 (n_1402, n_397, n_396);
  nand g819 (n_1403, n_395, n_397);
  nand g820 (n_412, n_1401, n_1402, n_1403);
  xor g821 (n_1404, n_398, n_399);
  xor g822 (n_219, n_1404, n_400);
  nand g823 (n_1405, n_398, n_399);
  nand g824 (n_1406, n_400, n_399);
  nand g825 (n_1407, n_398, n_400);
  nand g826 (n_133, n_1405, n_1406, n_1407);
  xor g827 (n_401, A[18], A[16]);
  and g828 (n_414, A[18], A[16]);
  xor g829 (n_1408, A[4], A[10]);
  xor g830 (n_406, n_1408, A[0]);
  nand g831 (n_1409, A[4], A[10]);
  xor g836 (n_404, n_359, A[6]);
  nand g839 (n_1415, A[14], A[6]);
  xor g842 (n_407, n_1280, n_401);
  nand g844 (n_1418, n_401, A[2]);
  nand g845 (n_1419, A[12], n_401);
  nand g846 (n_420, n_1281, n_1418, n_1419);
  xor g847 (n_1420, n_402, n_403);
  xor g848 (n_410, n_1420, n_404);
  nand g849 (n_1421, n_402, n_403);
  nand g850 (n_1422, n_404, n_403);
  nand g851 (n_1423, n_402, n_404);
  nand g852 (n_422, n_1421, n_1422, n_1423);
  xor g853 (n_1424, n_405, n_406);
  xor g854 (n_411, n_1424, n_407);
  nand g855 (n_1425, n_405, n_406);
  nand g856 (n_1426, n_407, n_406);
  nand g857 (n_1427, n_405, n_407);
  nand g858 (n_424, n_1425, n_1426, n_1427);
  xor g859 (n_1428, n_408, n_409);
  xor g860 (n_413, n_1428, n_410);
  nand g861 (n_1429, n_408, n_409);
  nand g862 (n_1430, n_410, n_409);
  nand g863 (n_1431, n_408, n_410);
  nand g864 (n_426, n_1429, n_1430, n_1431);
  xor g865 (n_1432, n_411, n_412);
  xor g866 (n_218, n_1432, n_413);
  nand g867 (n_1433, n_411, n_412);
  nand g868 (n_1434, n_413, n_412);
  nand g869 (n_1435, n_411, n_413);
  nand g870 (n_132, n_1433, n_1434, n_1435);
  xor g871 (n_1436, A[1], A[19]);
  xor g872 (n_418, n_1436, A[13]);
  nand g873 (n_1437, A[1], A[19]);
  nand g874 (n_1438, A[13], A[19]);
  nand g876 (n_428, n_1437, n_1438, n_1335);
  xor g877 (n_1440, A[5], A[17]);
  xor g878 (n_419, n_1440, A[11]);
  nand g879 (n_1441, A[5], A[17]);
  nand g880 (n_1442, A[11], A[17]);
  nand g881 (n_1443, A[5], A[11]);
  nand g882 (n_429, n_1441, n_1442, n_1443);
  xor g883 (n_1444, A[15], A[9]);
  xor g884 (n_417, n_1444, A[7]);
  nand g885 (n_1445, A[15], A[9]);
  nand g887 (n_1447, A[15], A[7]);
  nand g888 (n_430, n_1445, n_1238, n_1447);
  xor g889 (n_1448, A[3], n_414);
  xor g890 (n_421, n_1448, n_415);
  nand g891 (n_1449, A[3], n_414);
  nand g892 (n_1450, n_415, n_414);
  nand g893 (n_1451, A[3], n_415);
  nand g894 (n_434, n_1449, n_1450, n_1451);
  xor g895 (n_1452, n_416, n_417);
  xor g896 (n_423, n_1452, n_418);
  nand g897 (n_1453, n_416, n_417);
  nand g898 (n_1454, n_418, n_417);
  nand g899 (n_1455, n_416, n_418);
  nand g900 (n_436, n_1453, n_1454, n_1455);
  xor g901 (n_1456, n_419, n_420);
  xor g902 (n_425, n_1456, n_421);
  nand g903 (n_1457, n_419, n_420);
  nand g904 (n_1458, n_421, n_420);
  nand g905 (n_1459, n_419, n_421);
  nand g906 (n_438, n_1457, n_1458, n_1459);
  xor g907 (n_1460, n_422, n_423);
  xor g908 (n_427, n_1460, n_424);
  nand g909 (n_1461, n_422, n_423);
  nand g910 (n_1462, n_424, n_423);
  nand g911 (n_1463, n_422, n_424);
  nand g912 (n_440, n_1461, n_1462, n_1463);
  xor g913 (n_1464, n_425, n_426);
  xor g914 (n_217, n_1464, n_427);
  nand g915 (n_1465, n_425, n_426);
  nand g916 (n_1466, n_427, n_426);
  nand g917 (n_1467, n_425, n_427);
  nand g918 (n_131, n_1465, n_1466, n_1467);
  xor g919 (n_1468, A[20], A[18]);
  xor g920 (n_432, n_1468, A[14]);
  nand g921 (n_1469, A[20], A[18]);
  nand g922 (n_1470, A[14], A[18]);
  nand g923 (n_1471, A[20], A[14]);
  nand g924 (n_442, n_1469, n_1470, n_1471);
  xor g926 (n_433, n_323, A[16]);
  nand g928 (n_1474, A[16], A[4]);
  nand g929 (n_1475, A[6], A[16]);
  xor g932 (n_431, n_333, A[12]);
  nand g934 (n_1478, A[12], A[8]);
  nand g935 (n_1479, A[10], A[12]);
  xor g937 (n_1480, A[2], n_428);
  xor g938 (n_435, n_1480, n_429);
  nand g939 (n_1481, A[2], n_428);
  nand g940 (n_1482, n_429, n_428);
  nand g941 (n_1483, A[2], n_429);
  nand g942 (n_149, n_1481, n_1482, n_1483);
  xor g943 (n_1484, n_430, n_431);
  xor g944 (n_437, n_1484, n_432);
  nand g945 (n_1485, n_430, n_431);
  nand g946 (n_1486, n_432, n_431);
  nand g947 (n_1487, n_430, n_432);
  nand g948 (n_151, n_1485, n_1486, n_1487);
  xor g949 (n_1488, n_433, n_434);
  xor g950 (n_439, n_1488, n_435);
  nand g951 (n_1489, n_433, n_434);
  nand g952 (n_1490, n_435, n_434);
  nand g953 (n_1491, n_433, n_435);
  nand g954 (n_447, n_1489, n_1490, n_1491);
  xor g955 (n_1492, n_436, n_437);
  xor g956 (n_441, n_1492, n_438);
  nand g957 (n_1493, n_436, n_437);
  nand g958 (n_1494, n_438, n_437);
  nand g959 (n_1495, n_436, n_438);
  nand g960 (n_449, n_1493, n_1494, n_1495);
  xor g961 (n_1496, n_439, n_440);
  xor g962 (n_216, n_1496, n_441);
  nand g963 (n_1497, n_439, n_440);
  nand g964 (n_1498, n_441, n_440);
  nand g965 (n_1499, n_439, n_441);
  nand g966 (n_130, n_1497, n_1498, n_1499);
  xor g967 (n_1500, A[21], A[19]);
  xor g968 (n_445, n_1500, A[15]);
  nand g969 (n_1501, A[21], A[19]);
  nand g970 (n_1502, A[15], A[19]);
  nand g971 (n_1503, A[21], A[15]);
  nand g972 (n_451, n_1501, n_1502, n_1503);
  xor g974 (n_148, n_1388, A[13]);
  nand g977 (n_1507, A[7], A[13]);
  nand g978 (n_452, n_1222, n_1297, n_1507);
  xor g979 (n_1508, A[17], A[11]);
  xor g980 (n_444, n_1508, A[9]);
  nand g983 (n_1511, A[17], A[9]);
  nand g984 (n_453, n_1442, n_1339, n_1511);
  xor g985 (n_1512, A[3], n_442);
  xor g986 (n_150, n_1512, n_443);
  nand g987 (n_1513, A[3], n_442);
  nand g988 (n_1514, n_443, n_442);
  nand g989 (n_1515, A[3], n_443);
  nand g990 (n_457, n_1513, n_1514, n_1515);
  xor g991 (n_1516, n_444, n_445);
  xor g992 (n_446, n_1516, n_147);
  nand g993 (n_1517, n_444, n_445);
  nand g994 (n_1518, n_147, n_445);
  nand g995 (n_1519, n_444, n_147);
  nand g996 (n_459, n_1517, n_1518, n_1519);
  xor g997 (n_1520, n_148, n_149);
  xor g998 (n_448, n_1520, n_150);
  nand g999 (n_1521, n_148, n_149);
  nand g1000 (n_1522, n_150, n_149);
  nand g1001 (n_1523, n_148, n_150);
  nand g1002 (n_462, n_1521, n_1522, n_1523);
  xor g1003 (n_1524, n_151, n_446);
  xor g1004 (n_450, n_1524, n_447);
  nand g1005 (n_1525, n_151, n_446);
  nand g1006 (n_1526, n_447, n_446);
  nand g1007 (n_1527, n_151, n_447);
  nand g1008 (n_464, n_1525, n_1526, n_1527);
  xor g1009 (n_1528, n_448, n_449);
  xor g1010 (n_215, n_1528, n_450);
  nand g1011 (n_1529, n_448, n_449);
  nand g1012 (n_1530, n_450, n_449);
  nand g1013 (n_1531, n_448, n_450);
  nand g1014 (n_129, n_1529, n_1530, n_1531);
  xor g1015 (n_1532, A[22], A[20]);
  xor g1016 (n_455, n_1532, A[16]);
  nand g1017 (n_1533, A[22], A[20]);
  nand g1018 (n_1534, A[16], A[20]);
  nand g1019 (n_1535, A[22], A[16]);
  nand g1020 (n_465, n_1533, n_1534, n_1535);
  xor g1022 (n_456, n_326, A[14]);
  xor g1027 (n_1540, A[4], A[18]);
  xor g1028 (n_454, n_1540, A[10]);
  nand g1029 (n_1541, A[4], A[18]);
  nand g1030 (n_1542, A[10], A[18]);
  nand g1032 (n_467, n_1541, n_1542, n_1409);
  xor g1033 (n_1544, A[12], n_451);
  xor g1034 (n_458, n_1544, n_452);
  nand g1035 (n_1545, A[12], n_451);
  nand g1036 (n_1546, n_452, n_451);
  nand g1037 (n_1547, A[12], n_452);
  nand g1038 (n_471, n_1545, n_1546, n_1547);
  xor g1039 (n_1548, n_453, n_454);
  xor g1040 (n_460, n_1548, n_455);
  nand g1041 (n_1549, n_453, n_454);
  nand g1042 (n_1550, n_455, n_454);
  nand g1043 (n_1551, n_453, n_455);
  nand g1044 (n_473, n_1549, n_1550, n_1551);
  xor g1045 (n_1552, n_456, n_457);
  xor g1046 (n_461, n_1552, n_458);
  nand g1047 (n_1553, n_456, n_457);
  nand g1048 (n_1554, n_458, n_457);
  nand g1049 (n_1555, n_456, n_458);
  nand g1050 (n_475, n_1553, n_1554, n_1555);
  xor g1051 (n_1556, n_459, n_460);
  xor g1052 (n_463, n_1556, n_461);
  nand g1053 (n_1557, n_459, n_460);
  nand g1054 (n_1558, n_461, n_460);
  nand g1055 (n_1559, n_459, n_461);
  nand g1056 (n_478, n_1557, n_1558, n_1559);
  xor g1057 (n_1560, n_462, n_463);
  xor g1058 (n_214, n_1560, n_464);
  nand g1059 (n_1561, n_462, n_463);
  nand g1060 (n_1562, n_464, n_463);
  nand g1061 (n_1563, n_462, n_464);
  nand g1062 (n_128, n_1561, n_1562, n_1563);
  xor g1063 (n_1564, A[23], A[21]);
  xor g1064 (n_469, n_1564, A[17]);
  nand g1065 (n_1565, A[23], A[21]);
  nand g1066 (n_1566, A[17], A[21]);
  nand g1067 (n_1567, A[23], A[17]);
  nand g1068 (n_479, n_1565, n_1566, n_1567);
  xor g1070 (n_470, n_1336, A[15]);
  xor g1075 (n_1572, A[5], A[19]);
  xor g1076 (n_468, n_1572, A[13]);
  nand g1077 (n_1573, A[5], A[19]);
  nand g1080 (n_481, n_1573, n_1438, n_1297);
  xor g1081 (n_1576, A[11], n_465);
  xor g1082 (n_472, n_1576, n_415);
  nand g1083 (n_1577, A[11], n_465);
  nand g1084 (n_1578, n_415, n_465);
  nand g1085 (n_1579, A[11], n_415);
  nand g1086 (n_485, n_1577, n_1578, n_1579);
  xor g1087 (n_1580, n_467, n_468);
  xor g1088 (n_474, n_1580, n_469);
  nand g1089 (n_1581, n_467, n_468);
  nand g1090 (n_1582, n_469, n_468);
  nand g1091 (n_1583, n_467, n_469);
  nand g1092 (n_487, n_1581, n_1582, n_1583);
  xor g1093 (n_1584, n_470, n_471);
  xor g1094 (n_476, n_1584, n_472);
  nand g1095 (n_1585, n_470, n_471);
  nand g1096 (n_1586, n_472, n_471);
  nand g1097 (n_1587, n_470, n_472);
  nand g1098 (n_489, n_1585, n_1586, n_1587);
  xor g1099 (n_1588, n_473, n_474);
  xor g1100 (n_477, n_1588, n_475);
  nand g1101 (n_1589, n_473, n_474);
  nand g1102 (n_1590, n_475, n_474);
  nand g1103 (n_1591, n_473, n_475);
  nand g1104 (n_492, n_1589, n_1590, n_1591);
  xor g1105 (n_1592, n_476, n_477);
  xor g1106 (n_213, n_1592, n_478);
  nand g1107 (n_1593, n_476, n_477);
  nand g1108 (n_1594, n_478, n_477);
  nand g1109 (n_1595, n_476, n_478);
  nand g1110 (n_127, n_1593, n_1594, n_1595);
  xor g1111 (n_1596, A[24], A[22]);
  xor g1112 (n_483, n_1596, A[18]);
  nand g1113 (n_1597, A[24], A[22]);
  nand g1114 (n_1598, A[18], A[22]);
  nand g1115 (n_1599, A[24], A[18]);
  nand g1116 (n_493, n_1597, n_1598, n_1599);
  xor g1118 (n_484, n_333, A[16]);
  nand g1120 (n_1602, A[16], A[8]);
  nand g1121 (n_1603, A[10], A[16]);
  xor g1123 (n_1604, A[6], A[20]);
  xor g1124 (n_482, n_1604, A[14]);
  nand g1125 (n_1605, A[6], A[20]);
  nand g1128 (n_495, n_1605, n_1471, n_1415);
  xor g1129 (n_1608, A[12], n_479);
  xor g1130 (n_486, n_1608, n_430);
  nand g1131 (n_1609, A[12], n_479);
  nand g1132 (n_1610, n_430, n_479);
  nand g1133 (n_1611, A[12], n_430);
  nand g1134 (n_499, n_1609, n_1610, n_1611);
  xor g1135 (n_1612, n_481, n_482);
  xor g1136 (n_488, n_1612, n_483);
  nand g1137 (n_1613, n_481, n_482);
  nand g1138 (n_1614, n_483, n_482);
  nand g1139 (n_1615, n_481, n_483);
  nand g1140 (n_501, n_1613, n_1614, n_1615);
  xor g1141 (n_1616, n_484, n_485);
  xor g1142 (n_490, n_1616, n_486);
  nand g1143 (n_1617, n_484, n_485);
  nand g1144 (n_1618, n_486, n_485);
  nand g1145 (n_1619, n_484, n_486);
  nand g1146 (n_503, n_1617, n_1618, n_1619);
  xor g1147 (n_1620, n_487, n_488);
  xor g1148 (n_491, n_1620, n_489);
  nand g1149 (n_1621, n_487, n_488);
  nand g1150 (n_1622, n_489, n_488);
  nand g1151 (n_1623, n_487, n_489);
  nand g1152 (n_506, n_1621, n_1622, n_1623);
  xor g1153 (n_1624, n_490, n_491);
  xor g1154 (n_212, n_1624, n_492);
  nand g1155 (n_1625, n_490, n_491);
  nand g1156 (n_1626, n_492, n_491);
  nand g1157 (n_1627, n_490, n_492);
  nand g1158 (n_126, n_1625, n_1626, n_1627);
  xor g1159 (n_1628, A[25], A[23]);
  xor g1160 (n_497, n_1628, A[19]);
  nand g1161 (n_1629, A[25], A[23]);
  nand g1162 (n_1630, A[19], A[23]);
  nand g1163 (n_1631, A[25], A[19]);
  nand g1164 (n_507, n_1629, n_1630, n_1631);
  xor g1166 (n_498, n_1384, A[17]);
  xor g1171 (n_1636, A[7], A[21]);
  xor g1172 (n_496, n_1636, A[15]);
  nand g1173 (n_1637, A[7], A[21]);
  nand g1176 (n_508, n_1637, n_1503, n_1447);
  xor g1177 (n_1640, A[13], n_493);
  xor g1178 (n_500, n_1640, n_494);
  nand g1179 (n_1641, A[13], n_493);
  nand g1180 (n_1642, n_494, n_493);
  nand g1181 (n_1643, A[13], n_494);
  nand g1182 (n_513, n_1641, n_1642, n_1643);
  xor g1183 (n_1644, n_495, n_496);
  xor g1184 (n_502, n_1644, n_497);
  nand g1185 (n_1645, n_495, n_496);
  nand g1186 (n_1646, n_497, n_496);
  nand g1187 (n_1647, n_495, n_497);
  nand g1188 (n_515, n_1645, n_1646, n_1647);
  xor g1189 (n_1648, n_498, n_499);
  xor g1190 (n_504, n_1648, n_500);
  nand g1191 (n_1649, n_498, n_499);
  nand g1192 (n_1650, n_500, n_499);
  nand g1193 (n_1651, n_498, n_500);
  nand g1194 (n_518, n_1649, n_1650, n_1651);
  xor g1195 (n_1652, n_501, n_502);
  xor g1196 (n_505, n_1652, n_503);
  nand g1197 (n_1653, n_501, n_502);
  nand g1198 (n_1654, n_503, n_502);
  nand g1199 (n_1655, n_501, n_503);
  nand g1200 (n_520, n_1653, n_1654, n_1655);
  xor g1201 (n_1656, n_504, n_505);
  xor g1202 (n_211, n_1656, n_506);
  nand g1203 (n_1657, n_504, n_505);
  nand g1204 (n_1658, n_506, n_505);
  nand g1205 (n_1659, n_504, n_506);
  nand g1206 (n_125, n_1657, n_1658, n_1659);
  xor g1207 (n_1660, A[26], A[24]);
  xor g1208 (n_511, n_1660, A[20]);
  nand g1209 (n_1661, A[26], A[24]);
  nand g1210 (n_1662, A[20], A[24]);
  nand g1211 (n_1663, A[26], A[20]);
  nand g1212 (n_233, n_1661, n_1662, n_1663);
  xor g1213 (n_1664, A[10], A[18]);
  xor g1214 (n_512, n_1664, A[8]);
  nand g1216 (n_1666, A[8], A[18]);
  xor g1219 (n_1668, A[22], A[16]);
  xor g1220 (n_510, n_1668, A[14]);
  nand g1223 (n_1671, A[22], A[14]);
  xor g1225 (n_1672, A[12], n_507);
  xor g1226 (n_514, n_1672, n_508);
  nand g1227 (n_1673, A[12], n_507);
  nand g1228 (n_1674, n_508, n_507);
  nand g1229 (n_1675, A[12], n_508);
  nand g1230 (n_525, n_1673, n_1674, n_1675);
  xor g1231 (n_1676, n_453, n_510);
  xor g1232 (n_516, n_1676, n_511);
  nand g1233 (n_1677, n_453, n_510);
  nand g1234 (n_1678, n_511, n_510);
  nand g1235 (n_1679, n_453, n_511);
  nand g1236 (n_527, n_1677, n_1678, n_1679);
  xor g1237 (n_1680, n_512, n_513);
  xor g1238 (n_517, n_1680, n_514);
  nand g1239 (n_1681, n_512, n_513);
  nand g1240 (n_1682, n_514, n_513);
  nand g1241 (n_1683, n_512, n_514);
  nand g1242 (n_529, n_1681, n_1682, n_1683);
  xor g1243 (n_1684, n_515, n_516);
  xor g1244 (n_519, n_1684, n_517);
  nand g1245 (n_1685, n_515, n_516);
  nand g1246 (n_1686, n_517, n_516);
  nand g1247 (n_1687, n_515, n_517);
  nand g1248 (n_532, n_1685, n_1686, n_1687);
  xor g1249 (n_1688, n_518, n_519);
  xor g1250 (n_210, n_1688, n_520);
  nand g1251 (n_1689, n_518, n_519);
  nand g1252 (n_1690, n_520, n_519);
  nand g1253 (n_1691, n_518, n_520);
  nand g1254 (n_124, n_1689, n_1690, n_1691);
  xor g1255 (n_1692, A[27], A[25]);
  xor g1256 (n_523, n_1692, A[21]);
  nand g1257 (n_1693, A[27], A[25]);
  nand g1258 (n_1694, A[21], A[25]);
  nand g1259 (n_1695, A[27], A[21]);
  nand g1260 (n_533, n_1693, n_1694, n_1695);
  xor g1261 (n_1696, A[13], A[11]);
  xor g1262 (n_524, n_1696, A[19]);
  nand g1264 (n_1698, A[19], A[11]);
  nand g1266 (n_535, n_1387, n_1698, n_1438);
  xor g1267 (n_1700, A[9], A[23]);
  xor g1268 (n_522, n_1700, A[17]);
  nand g1269 (n_1701, A[9], A[23]);
  nand g1272 (n_534, n_1701, n_1567, n_1511);
  xor g1273 (n_1704, A[15], n_233);
  xor g1274 (n_526, n_1704, n_234);
  nand g1275 (n_1705, A[15], n_233);
  nand g1276 (n_1706, n_234, n_233);
  nand g1277 (n_1707, A[15], n_234);
  nand g1278 (n_539, n_1705, n_1706, n_1707);
  xor g1279 (n_1708, n_521, n_522);
  xor g1280 (n_528, n_1708, n_523);
  nand g1281 (n_1709, n_521, n_522);
  nand g1282 (n_1710, n_523, n_522);
  nand g1283 (n_1711, n_521, n_523);
  nand g1284 (n_541, n_1709, n_1710, n_1711);
  xor g1285 (n_1712, n_524, n_525);
  xor g1286 (n_530, n_1712, n_526);
  nand g1287 (n_1713, n_524, n_525);
  nand g1288 (n_1714, n_526, n_525);
  nand g1289 (n_1715, n_524, n_526);
  nand g1290 (n_544, n_1713, n_1714, n_1715);
  xor g1291 (n_1716, n_527, n_528);
  xor g1292 (n_531, n_1716, n_529);
  nand g1293 (n_1717, n_527, n_528);
  nand g1294 (n_1718, n_529, n_528);
  nand g1295 (n_1719, n_527, n_529);
  nand g1296 (n_546, n_1717, n_1718, n_1719);
  xor g1297 (n_1720, n_530, n_531);
  xor g1298 (n_209, n_1720, n_532);
  nand g1299 (n_1721, n_530, n_531);
  nand g1300 (n_1722, n_532, n_531);
  nand g1301 (n_1723, n_530, n_532);
  nand g1302 (n_123, n_1721, n_1722, n_1723);
  xor g1303 (n_1724, A[28], A[26]);
  xor g1304 (n_537, n_1724, A[22]);
  nand g1305 (n_1725, A[28], A[26]);
  nand g1306 (n_1726, A[22], A[26]);
  nand g1307 (n_1727, A[28], A[22]);
  nand g1308 (n_547, n_1725, n_1726, n_1727);
  xor g1309 (n_1728, A[14], A[20]);
  xor g1310 (n_538, n_1728, A[10]);
  nand g1312 (n_1730, A[10], A[20]);
  nand g1313 (n_1731, A[14], A[10]);
  nand g1314 (n_548, n_1471, n_1730, n_1731);
  xor g1315 (n_1732, A[24], A[18]);
  xor g1316 (n_536, n_1732, A[16]);
  nand g1319 (n_1735, A[24], A[16]);
  xor g1321 (n_1736, A[12], n_533);
  xor g1322 (n_540, n_1736, n_534);
  nand g1323 (n_1737, A[12], n_533);
  nand g1324 (n_1738, n_534, n_533);
  nand g1325 (n_1739, A[12], n_534);
  nand g1326 (n_553, n_1737, n_1738, n_1739);
  xor g1327 (n_1740, n_535, n_536);
  xor g1328 (n_542, n_1740, n_537);
  nand g1329 (n_1741, n_535, n_536);
  nand g1330 (n_1742, n_537, n_536);
  nand g1331 (n_1743, n_535, n_537);
  nand g1332 (n_555, n_1741, n_1742, n_1743);
  xor g1333 (n_1744, n_538, n_539);
  xor g1334 (n_543, n_1744, n_540);
  nand g1335 (n_1745, n_538, n_539);
  nand g1336 (n_1746, n_540, n_539);
  nand g1337 (n_1747, n_538, n_540);
  nand g1338 (n_557, n_1745, n_1746, n_1747);
  xor g1339 (n_1748, n_541, n_542);
  xor g1340 (n_545, n_1748, n_543);
  nand g1341 (n_1749, n_541, n_542);
  nand g1342 (n_1750, n_543, n_542);
  nand g1343 (n_1751, n_541, n_543);
  nand g1344 (n_560, n_1749, n_1750, n_1751);
  xor g1345 (n_1752, n_544, n_545);
  xor g1346 (n_208, n_1752, n_546);
  nand g1347 (n_1753, n_544, n_545);
  nand g1348 (n_1754, n_546, n_545);
  nand g1349 (n_1755, n_544, n_546);
  nand g1350 (n_122, n_1753, n_1754, n_1755);
  xor g1351 (n_1756, A[29], A[27]);
  xor g1352 (n_551, n_1756, A[23]);
  nand g1353 (n_1757, A[29], A[27]);
  nand g1354 (n_1758, A[23], A[27]);
  nand g1355 (n_1759, A[29], A[23]);
  nand g1356 (n_561, n_1757, n_1758, n_1759);
  xor g1357 (n_1760, A[15], A[13]);
  xor g1358 (n_552, n_1760, A[21]);
  nand g1360 (n_1762, A[21], A[13]);
  nand g1362 (n_563, n_1334, n_1762, n_1503);
  xor g1363 (n_1764, A[11], A[25]);
  xor g1364 (n_550, n_1764, A[19]);
  nand g1365 (n_1765, A[11], A[25]);
  nand g1368 (n_562, n_1765, n_1631, n_1698);
  xor g1369 (n_1768, A[17], n_547);
  xor g1370 (n_554, n_1768, n_548);
  nand g1371 (n_1769, A[17], n_547);
  nand g1372 (n_1770, n_548, n_547);
  nand g1373 (n_1771, A[17], n_548);
  nand g1374 (n_567, n_1769, n_1770, n_1771);
  xor g1375 (n_1772, n_549, n_550);
  xor g1376 (n_556, n_1772, n_551);
  nand g1377 (n_1773, n_549, n_550);
  nand g1378 (n_1774, n_551, n_550);
  nand g1379 (n_1775, n_549, n_551);
  nand g1380 (n_569, n_1773, n_1774, n_1775);
  xor g1381 (n_1776, n_552, n_553);
  xor g1382 (n_558, n_1776, n_554);
  nand g1383 (n_1777, n_552, n_553);
  nand g1384 (n_1778, n_554, n_553);
  nand g1385 (n_1779, n_552, n_554);
  nand g1386 (n_572, n_1777, n_1778, n_1779);
  xor g1387 (n_1780, n_555, n_556);
  xor g1388 (n_559, n_1780, n_557);
  nand g1389 (n_1781, n_555, n_556);
  nand g1390 (n_1782, n_557, n_556);
  nand g1391 (n_1783, n_555, n_557);
  nand g1392 (n_574, n_1781, n_1782, n_1783);
  xor g1393 (n_1784, n_558, n_559);
  xor g1394 (n_207, n_1784, n_560);
  nand g1395 (n_1785, n_558, n_559);
  nand g1396 (n_1786, n_560, n_559);
  nand g1397 (n_1787, n_558, n_560);
  nand g1398 (n_121, n_1785, n_1786, n_1787);
  xor g1399 (n_1788, A[30], A[28]);
  xor g1400 (n_565, n_1788, A[24]);
  nand g1401 (n_1789, A[30], A[28]);
  nand g1402 (n_1790, A[24], A[28]);
  nand g1403 (n_1791, A[30], A[24]);
  nand g1404 (n_575, n_1789, n_1790, n_1791);
  xor g1406 (n_566, n_378, A[22]);
  xor g1411 (n_1796, A[26], A[20]);
  xor g1412 (n_564, n_1796, A[18]);
  nand g1415 (n_1799, A[26], A[18]);
  nand g1416 (n_577, n_1663, n_1469, n_1799);
  xor g1417 (n_1800, A[12], n_561);
  xor g1418 (n_568, n_1800, n_562);
  nand g1419 (n_1801, A[12], n_561);
  nand g1420 (n_1802, n_562, n_561);
  nand g1421 (n_1803, A[12], n_562);
  nand g1422 (n_581, n_1801, n_1802, n_1803);
  xor g1423 (n_1804, n_563, n_564);
  xor g1424 (n_570, n_1804, n_565);
  nand g1425 (n_1805, n_563, n_564);
  nand g1426 (n_1806, n_565, n_564);
  nand g1427 (n_1807, n_563, n_565);
  nand g1428 (n_583, n_1805, n_1806, n_1807);
  xor g1429 (n_1808, n_566, n_567);
  xor g1430 (n_571, n_1808, n_568);
  nand g1431 (n_1809, n_566, n_567);
  nand g1432 (n_1810, n_568, n_567);
  nand g1433 (n_1811, n_566, n_568);
  nand g1434 (n_585, n_1809, n_1810, n_1811);
  xor g1435 (n_1812, n_569, n_570);
  xor g1436 (n_573, n_1812, n_571);
  nand g1437 (n_1813, n_569, n_570);
  nand g1438 (n_1814, n_571, n_570);
  nand g1439 (n_1815, n_569, n_571);
  nand g1440 (n_588, n_1813, n_1814, n_1815);
  xor g1441 (n_1816, n_572, n_573);
  xor g1442 (n_206, n_1816, n_574);
  nand g1443 (n_1817, n_572, n_573);
  nand g1444 (n_1818, n_574, n_573);
  nand g1445 (n_1819, n_572, n_574);
  nand g1446 (n_120, n_1817, n_1818, n_1819);
  xor g1447 (n_1820, A[31], A[29]);
  xor g1448 (n_579, n_1820, A[25]);
  nand g1449 (n_1821, A[31], A[29]);
  nand g1450 (n_1822, A[25], A[29]);
  nand g1451 (n_1823, A[31], A[25]);
  nand g1452 (n_589, n_1821, n_1822, n_1823);
  xor g1453 (n_1824, A[17], A[15]);
  xor g1454 (n_580, n_1824, A[23]);
  nand g1456 (n_1826, A[23], A[15]);
  nand g1458 (n_590, n_1382, n_1826, n_1567);
  xor g1459 (n_1828, A[13], A[27]);
  xor g1460 (n_578, n_1828, A[21]);
  nand g1461 (n_1829, A[13], A[27]);
  nand g1464 (n_591, n_1829, n_1695, n_1762);
  xor g1465 (n_1832, A[19], n_575);
  xor g1466 (n_582, n_1832, n_521);
  nand g1467 (n_1833, A[19], n_575);
  nand g1468 (n_1834, n_521, n_575);
  nand g1469 (n_1835, A[19], n_521);
  nand g1470 (n_595, n_1833, n_1834, n_1835);
  xor g1471 (n_1836, n_577, n_578);
  xor g1472 (n_584, n_1836, n_579);
  nand g1473 (n_1837, n_577, n_578);
  nand g1474 (n_1838, n_579, n_578);
  nand g1475 (n_1839, n_577, n_579);
  nand g1476 (n_597, n_1837, n_1838, n_1839);
  xor g1477 (n_1840, n_580, n_581);
  xor g1478 (n_586, n_1840, n_582);
  nand g1479 (n_1841, n_580, n_581);
  nand g1480 (n_1842, n_582, n_581);
  nand g1481 (n_1843, n_580, n_582);
  nand g1482 (n_599, n_1841, n_1842, n_1843);
  xor g1483 (n_1844, n_583, n_584);
  xor g1484 (n_587, n_1844, n_585);
  nand g1485 (n_1845, n_583, n_584);
  nand g1486 (n_1846, n_585, n_584);
  nand g1487 (n_1847, n_583, n_585);
  nand g1488 (n_602, n_1845, n_1846, n_1847);
  xor g1489 (n_1848, n_586, n_587);
  xor g1490 (n_205, n_1848, n_588);
  nand g1491 (n_1849, n_586, n_587);
  nand g1492 (n_1850, n_588, n_587);
  nand g1493 (n_1851, n_586, n_588);
  nand g1494 (n_119, n_1849, n_1850, n_1851);
  xor g1495 (n_1852, A[32], A[30]);
  xor g1496 (n_593, n_1852, A[26]);
  nand g1497 (n_1853, A[32], A[30]);
  nand g1498 (n_1854, A[26], A[30]);
  nand g1499 (n_1855, A[32], A[26]);
  nand g1500 (n_603, n_1853, n_1854, n_1855);
  xor g1502 (n_594, n_401, A[24]);
  xor g1507 (n_1860, A[14], A[28]);
  xor g1508 (n_592, n_1860, A[22]);
  nand g1509 (n_1861, A[14], A[28]);
  nand g1512 (n_605, n_1861, n_1727, n_1671);
  xor g1513 (n_1864, A[20], n_589);
  xor g1514 (n_596, n_1864, n_590);
  nand g1515 (n_1865, A[20], n_589);
  nand g1516 (n_1866, n_590, n_589);
  nand g1517 (n_1867, A[20], n_590);
  nand g1518 (n_609, n_1865, n_1866, n_1867);
  xor g1519 (n_1868, n_591, n_592);
  xor g1520 (n_598, n_1868, n_593);
  nand g1521 (n_1869, n_591, n_592);
  nand g1522 (n_1870, n_593, n_592);
  nand g1523 (n_1871, n_591, n_593);
  nand g1524 (n_611, n_1869, n_1870, n_1871);
  xor g1525 (n_1872, n_594, n_595);
  xor g1526 (n_600, n_1872, n_596);
  nand g1527 (n_1873, n_594, n_595);
  nand g1528 (n_1874, n_596, n_595);
  nand g1529 (n_1875, n_594, n_596);
  nand g1530 (n_613, n_1873, n_1874, n_1875);
  xor g1531 (n_1876, n_597, n_598);
  xor g1532 (n_601, n_1876, n_599);
  nand g1533 (n_1877, n_597, n_598);
  nand g1534 (n_1878, n_599, n_598);
  nand g1535 (n_1879, n_597, n_599);
  nand g1536 (n_616, n_1877, n_1878, n_1879);
  xor g1537 (n_1880, n_600, n_601);
  xor g1538 (n_204, n_1880, n_602);
  nand g1539 (n_1881, n_600, n_601);
  nand g1540 (n_1882, n_602, n_601);
  nand g1541 (n_1883, n_600, n_602);
  nand g1542 (n_118, n_1881, n_1882, n_1883);
  xor g1543 (n_1884, A[33], A[31]);
  xor g1544 (n_607, n_1884, A[27]);
  nand g1545 (n_1885, A[33], A[31]);
  nand g1546 (n_1886, A[27], A[31]);
  nand g1547 (n_1887, A[33], A[27]);
  nand g1548 (n_617, n_1885, n_1886, n_1887);
  xor g1549 (n_1888, A[19], A[17]);
  xor g1550 (n_608, n_1888, A[25]);
  nand g1551 (n_1889, A[19], A[17]);
  nand g1552 (n_1890, A[25], A[17]);
  nand g1554 (n_618, n_1889, n_1890, n_1631);
  xor g1555 (n_1892, A[15], A[29]);
  xor g1556 (n_606, n_1892, A[23]);
  nand g1557 (n_1893, A[15], A[29]);
  nand g1560 (n_619, n_1893, n_1759, n_1826);
  xor g1561 (n_1896, A[21], n_603);
  xor g1562 (n_610, n_1896, n_549);
  nand g1563 (n_1897, A[21], n_603);
  nand g1564 (n_1898, n_549, n_603);
  nand g1565 (n_1899, A[21], n_549);
  nand g1566 (n_623, n_1897, n_1898, n_1899);
  xor g1567 (n_1900, n_605, n_606);
  xor g1568 (n_612, n_1900, n_607);
  nand g1569 (n_1901, n_605, n_606);
  nand g1570 (n_1902, n_607, n_606);
  nand g1571 (n_1903, n_605, n_607);
  nand g1572 (n_625, n_1901, n_1902, n_1903);
  xor g1573 (n_1904, n_608, n_609);
  xor g1574 (n_614, n_1904, n_610);
  nand g1575 (n_1905, n_608, n_609);
  nand g1576 (n_1906, n_610, n_609);
  nand g1577 (n_1907, n_608, n_610);
  nand g1578 (n_627, n_1905, n_1906, n_1907);
  xor g1579 (n_1908, n_611, n_612);
  xor g1580 (n_615, n_1908, n_613);
  nand g1581 (n_1909, n_611, n_612);
  nand g1582 (n_1910, n_613, n_612);
  nand g1583 (n_1911, n_611, n_613);
  nand g1584 (n_630, n_1909, n_1910, n_1911);
  xor g1585 (n_1912, n_614, n_615);
  xor g1586 (n_203, n_1912, n_616);
  nand g1587 (n_1913, n_614, n_615);
  nand g1588 (n_1914, n_616, n_615);
  nand g1589 (n_1915, n_614, n_616);
  nand g1590 (n_117, n_1913, n_1914, n_1915);
  xor g1591 (n_1916, A[34], A[32]);
  xor g1592 (n_621, n_1916, A[28]);
  nand g1593 (n_1917, A[34], A[32]);
  nand g1594 (n_1918, A[28], A[32]);
  nand g1595 (n_1919, A[34], A[28]);
  nand g1596 (n_631, n_1917, n_1918, n_1919);
  xor g1598 (n_622, n_1468, A[26]);
  xor g1603 (n_1924, A[16], A[30]);
  xor g1604 (n_620, n_1924, A[24]);
  nand g1605 (n_1925, A[16], A[30]);
  nand g1608 (n_633, n_1925, n_1791, n_1735);
  xor g1609 (n_1928, A[22], n_617);
  xor g1610 (n_624, n_1928, n_618);
  nand g1611 (n_1929, A[22], n_617);
  nand g1612 (n_1930, n_618, n_617);
  nand g1613 (n_1931, A[22], n_618);
  nand g1614 (n_637, n_1929, n_1930, n_1931);
  xor g1615 (n_1932, n_619, n_620);
  xor g1616 (n_626, n_1932, n_621);
  nand g1617 (n_1933, n_619, n_620);
  nand g1618 (n_1934, n_621, n_620);
  nand g1619 (n_1935, n_619, n_621);
  nand g1620 (n_639, n_1933, n_1934, n_1935);
  xor g1621 (n_1936, n_622, n_623);
  xor g1622 (n_628, n_1936, n_624);
  nand g1623 (n_1937, n_622, n_623);
  nand g1624 (n_1938, n_624, n_623);
  nand g1625 (n_1939, n_622, n_624);
  nand g1626 (n_641, n_1937, n_1938, n_1939);
  xor g1627 (n_1940, n_625, n_626);
  xor g1628 (n_629, n_1940, n_627);
  nand g1629 (n_1941, n_625, n_626);
  nand g1630 (n_1942, n_627, n_626);
  nand g1631 (n_1943, n_625, n_627);
  nand g1632 (n_644, n_1941, n_1942, n_1943);
  xor g1633 (n_1944, n_628, n_629);
  xor g1634 (n_202, n_1944, n_630);
  nand g1635 (n_1945, n_628, n_629);
  nand g1636 (n_1946, n_630, n_629);
  nand g1637 (n_1947, n_628, n_630);
  nand g1638 (n_116, n_1945, n_1946, n_1947);
  xor g1639 (n_1948, A[35], A[33]);
  xor g1640 (n_635, n_1948, A[29]);
  nand g1641 (n_1949, A[35], A[33]);
  nand g1642 (n_1950, A[29], A[33]);
  nand g1643 (n_1951, A[35], A[29]);
  nand g1644 (n_645, n_1949, n_1950, n_1951);
  xor g1646 (n_636, n_1500, A[27]);
  nand g1648 (n_1954, A[27], A[19]);
  nand g1650 (n_646, n_1501, n_1954, n_1695);
  xor g1651 (n_1956, A[17], A[31]);
  xor g1652 (n_634, n_1956, A[25]);
  nand g1653 (n_1957, A[17], A[31]);
  nand g1656 (n_647, n_1957, n_1823, n_1890);
  xor g1657 (n_1960, A[23], n_631);
  xor g1658 (n_638, n_1960, n_577);
  nand g1659 (n_1961, A[23], n_631);
  nand g1660 (n_1962, n_577, n_631);
  nand g1661 (n_1963, A[23], n_577);
  nand g1662 (n_651, n_1961, n_1962, n_1963);
  xor g1663 (n_1964, n_633, n_634);
  xor g1664 (n_640, n_1964, n_635);
  nand g1665 (n_1965, n_633, n_634);
  nand g1666 (n_1966, n_635, n_634);
  nand g1667 (n_1967, n_633, n_635);
  nand g1668 (n_653, n_1965, n_1966, n_1967);
  xor g1669 (n_1968, n_636, n_637);
  xor g1670 (n_642, n_1968, n_638);
  nand g1671 (n_1969, n_636, n_637);
  nand g1672 (n_1970, n_638, n_637);
  nand g1673 (n_1971, n_636, n_638);
  nand g1674 (n_655, n_1969, n_1970, n_1971);
  xor g1675 (n_1972, n_639, n_640);
  xor g1676 (n_643, n_1972, n_641);
  nand g1677 (n_1973, n_639, n_640);
  nand g1678 (n_1974, n_641, n_640);
  nand g1679 (n_1975, n_639, n_641);
  nand g1680 (n_658, n_1973, n_1974, n_1975);
  xor g1681 (n_1976, n_642, n_643);
  xor g1682 (n_201, n_1976, n_644);
  nand g1683 (n_1977, n_642, n_643);
  nand g1684 (n_1978, n_644, n_643);
  nand g1685 (n_1979, n_642, n_644);
  nand g1686 (n_115, n_1977, n_1978, n_1979);
  xor g1687 (n_1980, A[36], A[34]);
  xor g1688 (n_649, n_1980, A[30]);
  nand g1689 (n_1981, A[36], A[34]);
  nand g1690 (n_1982, A[30], A[34]);
  nand g1691 (n_1983, A[36], A[30]);
  nand g1692 (n_659, n_1981, n_1982, n_1983);
  xor g1694 (n_650, n_1532, A[28]);
  nand g1696 (n_1986, A[28], A[20]);
  nand g1698 (n_660, n_1533, n_1986, n_1727);
  xor g1699 (n_1988, A[18], A[32]);
  xor g1700 (n_648, n_1988, A[26]);
  nand g1701 (n_1989, A[18], A[32]);
  nand g1704 (n_661, n_1989, n_1855, n_1799);
  xor g1705 (n_1992, A[24], n_645);
  xor g1706 (n_652, n_1992, n_646);
  nand g1707 (n_1993, A[24], n_645);
  nand g1708 (n_1994, n_646, n_645);
  nand g1709 (n_1995, A[24], n_646);
  nand g1710 (n_665, n_1993, n_1994, n_1995);
  xor g1711 (n_1996, n_647, n_648);
  xor g1712 (n_654, n_1996, n_649);
  nand g1713 (n_1997, n_647, n_648);
  nand g1714 (n_1998, n_649, n_648);
  nand g1715 (n_1999, n_647, n_649);
  nand g1716 (n_667, n_1997, n_1998, n_1999);
  xor g1717 (n_2000, n_650, n_651);
  xor g1718 (n_656, n_2000, n_652);
  nand g1719 (n_2001, n_650, n_651);
  nand g1720 (n_2002, n_652, n_651);
  nand g1721 (n_2003, n_650, n_652);
  nand g1722 (n_669, n_2001, n_2002, n_2003);
  xor g1723 (n_2004, n_653, n_654);
  xor g1724 (n_657, n_2004, n_655);
  nand g1725 (n_2005, n_653, n_654);
  nand g1726 (n_2006, n_655, n_654);
  nand g1727 (n_2007, n_653, n_655);
  nand g1728 (n_672, n_2005, n_2006, n_2007);
  xor g1729 (n_2008, n_656, n_657);
  xor g1730 (n_200, n_2008, n_658);
  nand g1731 (n_2009, n_656, n_657);
  nand g1732 (n_2010, n_658, n_657);
  nand g1733 (n_2011, n_656, n_658);
  nand g1734 (n_114, n_2009, n_2010, n_2011);
  xor g1735 (n_2012, A[37], A[35]);
  xor g1736 (n_663, n_2012, A[31]);
  nand g1737 (n_2013, A[37], A[35]);
  nand g1738 (n_2014, A[31], A[35]);
  nand g1739 (n_2015, A[37], A[31]);
  nand g1740 (n_673, n_2013, n_2014, n_2015);
  xor g1742 (n_664, n_1564, A[29]);
  nand g1744 (n_2018, A[29], A[21]);
  nand g1746 (n_674, n_1565, n_2018, n_1759);
  xor g1747 (n_2020, A[19], A[33]);
  xor g1748 (n_662, n_2020, A[27]);
  nand g1749 (n_2021, A[19], A[33]);
  nand g1752 (n_675, n_2021, n_1887, n_1954);
  xor g1753 (n_2024, A[25], n_659);
  xor g1754 (n_666, n_2024, n_660);
  nand g1755 (n_2025, A[25], n_659);
  nand g1756 (n_2026, n_660, n_659);
  nand g1757 (n_2027, A[25], n_660);
  nand g1758 (n_679, n_2025, n_2026, n_2027);
  xor g1759 (n_2028, n_661, n_662);
  xor g1760 (n_668, n_2028, n_663);
  nand g1761 (n_2029, n_661, n_662);
  nand g1762 (n_2030, n_663, n_662);
  nand g1763 (n_2031, n_661, n_663);
  nand g1764 (n_681, n_2029, n_2030, n_2031);
  xor g1765 (n_2032, n_664, n_665);
  xor g1766 (n_670, n_2032, n_666);
  nand g1767 (n_2033, n_664, n_665);
  nand g1768 (n_2034, n_666, n_665);
  nand g1769 (n_2035, n_664, n_666);
  nand g1770 (n_683, n_2033, n_2034, n_2035);
  xor g1771 (n_2036, n_667, n_668);
  xor g1772 (n_671, n_2036, n_669);
  nand g1773 (n_2037, n_667, n_668);
  nand g1774 (n_2038, n_669, n_668);
  nand g1775 (n_2039, n_667, n_669);
  nand g1776 (n_686, n_2037, n_2038, n_2039);
  xor g1777 (n_2040, n_670, n_671);
  xor g1778 (n_199, n_2040, n_672);
  nand g1779 (n_2041, n_670, n_671);
  nand g1780 (n_2042, n_672, n_671);
  nand g1781 (n_2043, n_670, n_672);
  nand g1782 (n_113, n_2041, n_2042, n_2043);
  xor g1783 (n_2044, A[38], A[36]);
  xor g1784 (n_677, n_2044, A[32]);
  nand g1785 (n_2045, A[38], A[36]);
  nand g1786 (n_2046, A[32], A[36]);
  nand g1787 (n_2047, A[38], A[32]);
  nand g1788 (n_687, n_2045, n_2046, n_2047);
  xor g1790 (n_678, n_1596, A[30]);
  nand g1792 (n_2050, A[30], A[22]);
  nand g1794 (n_688, n_1597, n_2050, n_1791);
  xor g1795 (n_2052, A[20], A[34]);
  xor g1796 (n_676, n_2052, A[28]);
  nand g1797 (n_2053, A[20], A[34]);
  nand g1800 (n_689, n_2053, n_1919, n_1986);
  xor g1801 (n_2056, A[26], n_673);
  xor g1802 (n_680, n_2056, n_674);
  nand g1803 (n_2057, A[26], n_673);
  nand g1804 (n_2058, n_674, n_673);
  nand g1805 (n_2059, A[26], n_674);
  nand g1806 (n_693, n_2057, n_2058, n_2059);
  xor g1807 (n_2060, n_675, n_676);
  xor g1808 (n_682, n_2060, n_677);
  nand g1809 (n_2061, n_675, n_676);
  nand g1810 (n_2062, n_677, n_676);
  nand g1811 (n_2063, n_675, n_677);
  nand g1812 (n_695, n_2061, n_2062, n_2063);
  xor g1813 (n_2064, n_678, n_679);
  xor g1814 (n_684, n_2064, n_680);
  nand g1815 (n_2065, n_678, n_679);
  nand g1816 (n_2066, n_680, n_679);
  nand g1817 (n_2067, n_678, n_680);
  nand g1818 (n_697, n_2065, n_2066, n_2067);
  xor g1819 (n_2068, n_681, n_682);
  xor g1820 (n_685, n_2068, n_683);
  nand g1821 (n_2069, n_681, n_682);
  nand g1822 (n_2070, n_683, n_682);
  nand g1823 (n_2071, n_681, n_683);
  nand g1824 (n_700, n_2069, n_2070, n_2071);
  xor g1825 (n_2072, n_684, n_685);
  xor g1826 (n_198, n_2072, n_686);
  nand g1827 (n_2073, n_684, n_685);
  nand g1828 (n_2074, n_686, n_685);
  nand g1829 (n_2075, n_684, n_686);
  nand g1830 (n_112, n_2073, n_2074, n_2075);
  xor g1831 (n_2076, A[39], A[37]);
  xor g1832 (n_691, n_2076, A[33]);
  nand g1833 (n_2077, A[39], A[37]);
  nand g1834 (n_2078, A[33], A[37]);
  nand g1835 (n_2079, A[39], A[33]);
  nand g1836 (n_701, n_2077, n_2078, n_2079);
  xor g1838 (n_692, n_1628, A[31]);
  nand g1840 (n_2082, A[31], A[23]);
  nand g1842 (n_702, n_1629, n_2082, n_1823);
  xor g1843 (n_2084, A[21], A[35]);
  xor g1844 (n_690, n_2084, A[29]);
  nand g1845 (n_2085, A[21], A[35]);
  nand g1848 (n_703, n_2085, n_1951, n_2018);
  xor g1849 (n_2088, A[27], n_687);
  xor g1850 (n_694, n_2088, n_688);
  nand g1851 (n_2089, A[27], n_687);
  nand g1852 (n_2090, n_688, n_687);
  nand g1853 (n_2091, A[27], n_688);
  nand g1854 (n_707, n_2089, n_2090, n_2091);
  xor g1855 (n_2092, n_689, n_690);
  xor g1856 (n_696, n_2092, n_691);
  nand g1857 (n_2093, n_689, n_690);
  nand g1858 (n_2094, n_691, n_690);
  nand g1859 (n_2095, n_689, n_691);
  nand g1860 (n_709, n_2093, n_2094, n_2095);
  xor g1861 (n_2096, n_692, n_693);
  xor g1862 (n_698, n_2096, n_694);
  nand g1863 (n_2097, n_692, n_693);
  nand g1864 (n_2098, n_694, n_693);
  nand g1865 (n_2099, n_692, n_694);
  nand g1866 (n_711, n_2097, n_2098, n_2099);
  xor g1867 (n_2100, n_695, n_696);
  xor g1868 (n_699, n_2100, n_697);
  nand g1869 (n_2101, n_695, n_696);
  nand g1870 (n_2102, n_697, n_696);
  nand g1871 (n_2103, n_695, n_697);
  nand g1872 (n_714, n_2101, n_2102, n_2103);
  xor g1873 (n_2104, n_698, n_699);
  xor g1874 (n_197, n_2104, n_700);
  nand g1875 (n_2105, n_698, n_699);
  nand g1876 (n_2106, n_700, n_699);
  nand g1877 (n_2107, n_698, n_700);
  nand g1878 (n_111, n_2105, n_2106, n_2107);
  xor g1879 (n_2108, A[40], A[38]);
  xor g1880 (n_705, n_2108, A[34]);
  nand g1881 (n_2109, A[40], A[38]);
  nand g1882 (n_2110, A[34], A[38]);
  nand g1883 (n_2111, A[40], A[34]);
  nand g1884 (n_715, n_2109, n_2110, n_2111);
  xor g1886 (n_706, n_1660, A[32]);
  nand g1888 (n_2114, A[32], A[24]);
  nand g1890 (n_716, n_1661, n_2114, n_1855);
  xor g1891 (n_2116, A[22], A[36]);
  xor g1892 (n_704, n_2116, A[30]);
  nand g1893 (n_2117, A[22], A[36]);
  nand g1896 (n_717, n_2117, n_1983, n_2050);
  xor g1897 (n_2120, A[28], n_701);
  xor g1898 (n_708, n_2120, n_702);
  nand g1899 (n_2121, A[28], n_701);
  nand g1900 (n_2122, n_702, n_701);
  nand g1901 (n_2123, A[28], n_702);
  nand g1902 (n_721, n_2121, n_2122, n_2123);
  xor g1903 (n_2124, n_703, n_704);
  xor g1904 (n_710, n_2124, n_705);
  nand g1905 (n_2125, n_703, n_704);
  nand g1906 (n_2126, n_705, n_704);
  nand g1907 (n_2127, n_703, n_705);
  nand g1908 (n_723, n_2125, n_2126, n_2127);
  xor g1909 (n_2128, n_706, n_707);
  xor g1910 (n_712, n_2128, n_708);
  nand g1911 (n_2129, n_706, n_707);
  nand g1912 (n_2130, n_708, n_707);
  nand g1913 (n_2131, n_706, n_708);
  nand g1914 (n_725, n_2129, n_2130, n_2131);
  xor g1915 (n_2132, n_709, n_710);
  xor g1916 (n_713, n_2132, n_711);
  nand g1917 (n_2133, n_709, n_710);
  nand g1918 (n_2134, n_711, n_710);
  nand g1919 (n_2135, n_709, n_711);
  nand g1920 (n_728, n_2133, n_2134, n_2135);
  xor g1921 (n_2136, n_712, n_713);
  xor g1922 (n_196, n_2136, n_714);
  nand g1923 (n_2137, n_712, n_713);
  nand g1924 (n_2138, n_714, n_713);
  nand g1925 (n_2139, n_712, n_714);
  nand g1926 (n_110, n_2137, n_2138, n_2139);
  xor g1927 (n_2140, A[41], A[39]);
  xor g1928 (n_719, n_2140, A[35]);
  nand g1929 (n_2141, A[41], A[39]);
  nand g1930 (n_2142, A[35], A[39]);
  nand g1931 (n_2143, A[41], A[35]);
  nand g1932 (n_729, n_2141, n_2142, n_2143);
  xor g1934 (n_720, n_1692, A[33]);
  nand g1936 (n_2146, A[33], A[25]);
  nand g1938 (n_731, n_1693, n_2146, n_1887);
  xor g1939 (n_2148, A[23], A[37]);
  xor g1940 (n_718, n_2148, A[31]);
  nand g1941 (n_2149, A[23], A[37]);
  nand g1944 (n_730, n_2149, n_2015, n_2082);
  xor g1945 (n_2152, A[29], n_715);
  xor g1946 (n_722, n_2152, n_716);
  nand g1947 (n_2153, A[29], n_715);
  nand g1948 (n_2154, n_716, n_715);
  nand g1949 (n_2155, A[29], n_716);
  nand g1950 (n_735, n_2153, n_2154, n_2155);
  xor g1951 (n_2156, n_717, n_718);
  xor g1952 (n_724, n_2156, n_719);
  nand g1953 (n_2157, n_717, n_718);
  nand g1954 (n_2158, n_719, n_718);
  nand g1955 (n_2159, n_717, n_719);
  nand g1956 (n_737, n_2157, n_2158, n_2159);
  xor g1957 (n_2160, n_720, n_721);
  xor g1958 (n_726, n_2160, n_722);
  nand g1959 (n_2161, n_720, n_721);
  nand g1960 (n_2162, n_722, n_721);
  nand g1961 (n_2163, n_720, n_722);
  nand g1962 (n_740, n_2161, n_2162, n_2163);
  xor g1963 (n_2164, n_723, n_724);
  xor g1964 (n_727, n_2164, n_725);
  nand g1965 (n_2165, n_723, n_724);
  nand g1966 (n_2166, n_725, n_724);
  nand g1967 (n_2167, n_723, n_725);
  nand g1968 (n_742, n_2165, n_2166, n_2167);
  xor g1969 (n_2168, n_726, n_727);
  xor g1970 (n_195, n_2168, n_728);
  nand g1971 (n_2169, n_726, n_727);
  nand g1972 (n_2170, n_728, n_727);
  nand g1973 (n_2171, n_726, n_728);
  nand g1974 (n_109, n_2169, n_2170, n_2171);
  xor g1975 (n_2172, A[40], A[36]);
  xor g1976 (n_733, n_2172, A[28]);
  nand g1977 (n_2173, A[40], A[36]);
  nand g1978 (n_2174, A[28], A[36]);
  nand g1979 (n_2175, A[40], A[28]);
  nand g1980 (n_743, n_2173, n_2174, n_2175);
  xor g1981 (n_2176, A[26], A[34]);
  xor g1982 (n_734, n_2176, A[24]);
  nand g1983 (n_2177, A[26], A[34]);
  nand g1984 (n_2178, A[24], A[34]);
  nand g1986 (n_745, n_2177, n_2178, n_1661);
  xor g1987 (n_2180, A[38], A[32]);
  xor g1988 (n_732, n_2180, A[30]);
  nand g1991 (n_2183, A[38], A[30]);
  nand g1992 (n_744, n_2047, n_1853, n_2183);
  xor g1993 (n_2184, A[42], n_729);
  xor g1994 (n_736, n_2184, n_730);
  nand g1995 (n_2185, A[42], n_729);
  nand g1996 (n_2186, n_730, n_729);
  nand g1997 (n_2187, A[42], n_730);
  nand g1998 (n_749, n_2185, n_2186, n_2187);
  xor g1999 (n_2188, n_731, n_732);
  xor g2000 (n_738, n_2188, n_733);
  nand g2001 (n_2189, n_731, n_732);
  nand g2002 (n_2190, n_733, n_732);
  nand g2003 (n_2191, n_731, n_733);
  nand g2004 (n_751, n_2189, n_2190, n_2191);
  xor g2005 (n_2192, n_734, n_735);
  xor g2006 (n_739, n_2192, n_736);
  nand g2007 (n_2193, n_734, n_735);
  nand g2008 (n_2194, n_736, n_735);
  nand g2009 (n_2195, n_734, n_736);
  nand g2010 (n_754, n_2193, n_2194, n_2195);
  xor g2011 (n_2196, n_737, n_738);
  xor g2012 (n_741, n_2196, n_739);
  nand g2013 (n_2197, n_737, n_738);
  nand g2014 (n_2198, n_739, n_738);
  nand g2015 (n_2199, n_737, n_739);
  nand g2016 (n_756, n_2197, n_2198, n_2199);
  xor g2017 (n_2200, n_740, n_741);
  xor g2018 (n_194, n_2200, n_742);
  nand g2019 (n_2201, n_740, n_741);
  nand g2020 (n_2202, n_742, n_741);
  nand g2021 (n_2203, n_740, n_742);
  nand g2022 (n_108, n_2201, n_2202, n_2203);
  xor g2023 (n_2204, A[41], A[37]);
  xor g2024 (n_747, n_2204, A[29]);
  nand g2025 (n_2205, A[41], A[37]);
  nand g2026 (n_2206, A[29], A[37]);
  nand g2027 (n_2207, A[41], A[29]);
  nand g2028 (n_757, n_2205, n_2206, n_2207);
  xor g2029 (n_2208, A[27], A[35]);
  xor g2030 (n_748, n_2208, A[25]);
  nand g2031 (n_2209, A[27], A[35]);
  nand g2032 (n_2210, A[25], A[35]);
  nand g2034 (n_759, n_2209, n_2210, n_1693);
  xor g2035 (n_2212, A[39], A[33]);
  xor g2036 (n_746, n_2212, A[31]);
  nand g2039 (n_2215, A[39], A[31]);
  nand g2040 (n_758, n_2079, n_1885, n_2215);
  xor g2041 (n_2216, A[43], n_743);
  xor g2042 (n_750, n_2216, n_744);
  nand g2043 (n_2217, A[43], n_743);
  nand g2044 (n_2218, n_744, n_743);
  nand g2045 (n_2219, A[43], n_744);
  nand g2046 (n_763, n_2217, n_2218, n_2219);
  xor g2047 (n_2220, n_745, n_746);
  xor g2048 (n_752, n_2220, n_747);
  nand g2049 (n_2221, n_745, n_746);
  nand g2050 (n_2222, n_747, n_746);
  nand g2051 (n_2223, n_745, n_747);
  nand g2052 (n_765, n_2221, n_2222, n_2223);
  xor g2053 (n_2224, n_748, n_749);
  xor g2054 (n_753, n_2224, n_750);
  nand g2055 (n_2225, n_748, n_749);
  nand g2056 (n_2226, n_750, n_749);
  nand g2057 (n_2227, n_748, n_750);
  nand g2058 (n_768, n_2225, n_2226, n_2227);
  xor g2059 (n_2228, n_751, n_752);
  xor g2060 (n_755, n_2228, n_753);
  nand g2061 (n_2229, n_751, n_752);
  nand g2062 (n_2230, n_753, n_752);
  nand g2063 (n_2231, n_751, n_753);
  nand g2064 (n_770, n_2229, n_2230, n_2231);
  xor g2065 (n_2232, n_754, n_755);
  xor g2066 (n_193, n_2232, n_756);
  nand g2067 (n_2233, n_754, n_755);
  nand g2068 (n_2234, n_756, n_755);
  nand g2069 (n_2235, n_754, n_756);
  nand g2070 (n_107, n_2233, n_2234, n_2235);
  xor g2071 (n_2236, A[44], A[38]);
  xor g2072 (n_761, n_2236, A[30]);
  nand g2073 (n_2237, A[44], A[38]);
  nand g2075 (n_2239, A[44], A[30]);
  nand g2076 (n_771, n_2237, n_2183, n_2239);
  xor g2077 (n_2240, A[28], A[36]);
  xor g2078 (n_762, n_2240, A[26]);
  nand g2080 (n_2242, A[26], A[36]);
  nand g2082 (n_773, n_2174, n_2242, n_1725);
  xor g2083 (n_2244, A[40], A[34]);
  xor g2084 (n_760, n_2244, A[32]);
  nand g2087 (n_2247, A[40], A[32]);
  nand g2088 (n_772, n_2111, n_1917, n_2247);
  xor g2089 (n_2248, A[42], n_757);
  xor g2090 (n_764, n_2248, n_758);
  nand g2091 (n_2249, A[42], n_757);
  nand g2092 (n_2250, n_758, n_757);
  nand g2093 (n_2251, A[42], n_758);
  nand g2094 (n_777, n_2249, n_2250, n_2251);
  xor g2095 (n_2252, n_759, n_760);
  xor g2096 (n_766, n_2252, n_761);
  nand g2097 (n_2253, n_759, n_760);
  nand g2098 (n_2254, n_761, n_760);
  nand g2099 (n_2255, n_759, n_761);
  nand g2100 (n_779, n_2253, n_2254, n_2255);
  xor g2101 (n_2256, n_762, n_763);
  xor g2102 (n_767, n_2256, n_764);
  nand g2103 (n_2257, n_762, n_763);
  nand g2104 (n_2258, n_764, n_763);
  nand g2105 (n_2259, n_762, n_764);
  nand g2106 (n_782, n_2257, n_2258, n_2259);
  xor g2107 (n_2260, n_765, n_766);
  xor g2108 (n_769, n_2260, n_767);
  nand g2109 (n_2261, n_765, n_766);
  nand g2110 (n_2262, n_767, n_766);
  nand g2111 (n_2263, n_765, n_767);
  nand g2112 (n_784, n_2261, n_2262, n_2263);
  xor g2113 (n_2264, n_768, n_769);
  xor g2114 (n_192, n_2264, n_770);
  nand g2115 (n_2265, n_768, n_769);
  nand g2116 (n_2266, n_770, n_769);
  nand g2117 (n_2267, n_768, n_770);
  nand g2118 (n_106, n_2265, n_2266, n_2267);
  xor g2119 (n_2268, A[45], A[39]);
  xor g2120 (n_775, n_2268, A[31]);
  nand g2121 (n_2269, A[45], A[39]);
  nand g2123 (n_2271, A[45], A[31]);
  nand g2124 (n_785, n_2269, n_2215, n_2271);
  xor g2125 (n_2272, A[29], A[37]);
  xor g2126 (n_776, n_2272, A[27]);
  nand g2128 (n_2274, A[27], A[37]);
  nand g2130 (n_786, n_2206, n_2274, n_1757);
  xor g2131 (n_2276, A[41], A[35]);
  xor g2132 (n_774, n_2276, A[33]);
  nand g2135 (n_2279, A[41], A[33]);
  nand g2136 (n_787, n_2143, n_1949, n_2279);
  xor g2137 (n_2280, A[43], n_771);
  xor g2138 (n_778, n_2280, n_772);
  nand g2139 (n_2281, A[43], n_771);
  nand g2140 (n_2282, n_772, n_771);
  nand g2141 (n_2283, A[43], n_772);
  nand g2142 (n_791, n_2281, n_2282, n_2283);
  xor g2143 (n_2284, n_773, n_774);
  xor g2144 (n_780, n_2284, n_775);
  nand g2145 (n_2285, n_773, n_774);
  nand g2146 (n_2286, n_775, n_774);
  nand g2147 (n_2287, n_773, n_775);
  nand g2148 (n_793, n_2285, n_2286, n_2287);
  xor g2149 (n_2288, n_776, n_777);
  xor g2150 (n_781, n_2288, n_778);
  nand g2151 (n_2289, n_776, n_777);
  nand g2152 (n_2290, n_778, n_777);
  nand g2153 (n_2291, n_776, n_778);
  nand g2154 (n_796, n_2289, n_2290, n_2291);
  xor g2155 (n_2292, n_779, n_780);
  xor g2156 (n_783, n_2292, n_781);
  nand g2157 (n_2293, n_779, n_780);
  nand g2158 (n_2294, n_781, n_780);
  nand g2159 (n_2295, n_779, n_781);
  nand g2160 (n_798, n_2293, n_2294, n_2295);
  xor g2161 (n_2296, n_782, n_783);
  xor g2162 (n_191, n_2296, n_784);
  nand g2163 (n_2297, n_782, n_783);
  nand g2164 (n_2298, n_784, n_783);
  nand g2165 (n_2299, n_782, n_784);
  nand g2166 (n_105, n_2297, n_2298, n_2299);
  xor g2167 (n_2300, A[46], A[44]);
  xor g2168 (n_789, n_2300, A[40]);
  nand g2169 (n_2301, A[46], A[44]);
  nand g2170 (n_2302, A[40], A[44]);
  nand g2171 (n_2303, A[46], A[40]);
  nand g2172 (n_799, n_2301, n_2302, n_2303);
  xor g2174 (n_790, n_1852, A[38]);
  xor g2180 (n_788, n_2240, A[34]);
  nand g2184 (n_801, n_2174, n_1981, n_1919);
  xor g2185 (n_2312, A[42], n_785);
  xor g2186 (n_792, n_2312, n_786);
  nand g2187 (n_2313, A[42], n_785);
  nand g2188 (n_2314, n_786, n_785);
  nand g2189 (n_2315, A[42], n_786);
  nand g2190 (n_805, n_2313, n_2314, n_2315);
  xor g2191 (n_2316, n_787, n_788);
  xor g2192 (n_794, n_2316, n_789);
  nand g2193 (n_2317, n_787, n_788);
  nand g2194 (n_2318, n_789, n_788);
  nand g2195 (n_2319, n_787, n_789);
  nand g2196 (n_807, n_2317, n_2318, n_2319);
  xor g2197 (n_2320, n_790, n_791);
  xor g2198 (n_795, n_2320, n_792);
  nand g2199 (n_2321, n_790, n_791);
  nand g2200 (n_2322, n_792, n_791);
  nand g2201 (n_2323, n_790, n_792);
  nand g2202 (n_810, n_2321, n_2322, n_2323);
  xor g2203 (n_2324, n_793, n_794);
  xor g2204 (n_797, n_2324, n_795);
  nand g2205 (n_2325, n_793, n_794);
  nand g2206 (n_2326, n_795, n_794);
  nand g2207 (n_2327, n_793, n_795);
  nand g2208 (n_812, n_2325, n_2326, n_2327);
  xor g2209 (n_2328, n_796, n_797);
  xor g2210 (n_190, n_2328, n_798);
  nand g2211 (n_2329, n_796, n_797);
  nand g2212 (n_2330, n_798, n_797);
  nand g2213 (n_2331, n_796, n_798);
  nand g2214 (n_104, n_2329, n_2330, n_2331);
  xor g2215 (n_2332, A[47], A[45]);
  xor g2216 (n_803, n_2332, A[41]);
  nand g2217 (n_2333, A[47], A[45]);
  nand g2218 (n_2334, A[41], A[45]);
  nand g2219 (n_2335, A[47], A[41]);
  nand g2220 (n_813, n_2333, n_2334, n_2335);
  xor g2222 (n_804, n_1884, A[39]);
  xor g2228 (n_802, n_2272, A[35]);
  nand g2232 (n_815, n_2206, n_2013, n_1951);
  xor g2233 (n_2344, A[43], n_799);
  xor g2234 (n_806, n_2344, n_744);
  nand g2235 (n_2345, A[43], n_799);
  nand g2236 (n_2346, n_744, n_799);
  nand g2238 (n_819, n_2345, n_2346, n_2219);
  xor g2239 (n_2348, n_801, n_802);
  xor g2240 (n_808, n_2348, n_803);
  nand g2241 (n_2349, n_801, n_802);
  nand g2242 (n_2350, n_803, n_802);
  nand g2243 (n_2351, n_801, n_803);
  nand g2244 (n_821, n_2349, n_2350, n_2351);
  xor g2245 (n_2352, n_804, n_805);
  xor g2246 (n_809, n_2352, n_806);
  nand g2247 (n_2353, n_804, n_805);
  nand g2248 (n_2354, n_806, n_805);
  nand g2249 (n_2355, n_804, n_806);
  nand g2250 (n_824, n_2353, n_2354, n_2355);
  xor g2251 (n_2356, n_807, n_808);
  xor g2252 (n_811, n_2356, n_809);
  nand g2253 (n_2357, n_807, n_808);
  nand g2254 (n_2358, n_809, n_808);
  nand g2255 (n_2359, n_807, n_809);
  nand g2256 (n_826, n_2357, n_2358, n_2359);
  xor g2257 (n_2360, n_810, n_811);
  xor g2258 (n_189, n_2360, n_812);
  nand g2259 (n_2361, n_810, n_811);
  nand g2260 (n_2362, n_812, n_811);
  nand g2261 (n_2363, n_810, n_812);
  nand g2262 (n_103, n_2361, n_2362, n_2363);
  xor g2263 (n_2364, A[46], A[40]);
  xor g2264 (n_817, n_2364, A[34]);
  nand g2267 (n_2367, A[46], A[34]);
  nand g2268 (n_827, n_2303, n_2111, n_2367);
  xor g2270 (n_818, n_1852, A[44]);
  nand g2273 (n_2371, A[32], A[44]);
  nand g2274 (n_828, n_1853, n_2239, n_2371);
  xor g2276 (n_816, n_2044, A[42]);
  nand g2278 (n_2374, A[42], A[36]);
  nand g2279 (n_2375, A[38], A[42]);
  nand g2280 (n_831, n_2045, n_2374, n_2375);
  xor g2281 (n_2376, A[48], n_813);
  xor g2282 (n_820, n_2376, n_758);
  nand g2283 (n_2377, A[48], n_813);
  nand g2284 (n_2378, n_758, n_813);
  nand g2285 (n_2379, A[48], n_758);
  nand g2286 (n_833, n_2377, n_2378, n_2379);
  xor g2287 (n_2380, n_815, n_816);
  xor g2288 (n_822, n_2380, n_817);
  nand g2289 (n_2381, n_815, n_816);
  nand g2290 (n_2382, n_817, n_816);
  nand g2291 (n_2383, n_815, n_817);
  nand g2292 (n_835, n_2381, n_2382, n_2383);
  xor g2293 (n_2384, n_818, n_819);
  xor g2294 (n_823, n_2384, n_820);
  nand g2295 (n_2385, n_818, n_819);
  nand g2296 (n_2386, n_820, n_819);
  nand g2297 (n_2387, n_818, n_820);
  nand g2298 (n_837, n_2385, n_2386, n_2387);
  xor g2299 (n_2388, n_821, n_822);
  xor g2300 (n_825, n_2388, n_823);
  nand g2301 (n_2389, n_821, n_822);
  nand g2302 (n_2390, n_823, n_822);
  nand g2303 (n_2391, n_821, n_823);
  nand g2304 (n_840, n_2389, n_2390, n_2391);
  xor g2305 (n_2392, n_824, n_825);
  xor g2306 (n_188, n_2392, n_826);
  nand g2307 (n_2393, n_824, n_825);
  nand g2308 (n_2394, n_826, n_825);
  nand g2309 (n_2395, n_824, n_826);
  nand g2310 (n_102, n_2393, n_2394, n_2395);
  xor g2311 (n_2396, A[47], A[41]);
  xor g2312 (n_830, n_2396, A[35]);
  nand g2315 (n_2399, A[47], A[35]);
  nand g2316 (n_841, n_2335, n_2143, n_2399);
  xor g2318 (n_832, n_1884, A[45]);
  nand g2321 (n_2403, A[33], A[45]);
  nand g2322 (n_842, n_1885, n_2271, n_2403);
  xor g2324 (n_829, n_2076, A[43]);
  nand g2326 (n_2406, A[43], A[37]);
  nand g2327 (n_2407, A[39], A[43]);
  nand g2328 (n_844, n_2077, n_2406, n_2407);
  xor g2329 (n_2408, A[49], n_827);
  xor g2330 (n_834, n_2408, n_828);
  nand g2331 (n_2409, A[49], n_827);
  nand g2332 (n_2410, n_828, n_827);
  nand g2333 (n_2411, A[49], n_828);
  nand g2334 (n_847, n_2409, n_2410, n_2411);
  xor g2335 (n_2412, n_829, n_830);
  xor g2336 (n_836, n_2412, n_831);
  nand g2337 (n_2413, n_829, n_830);
  nand g2338 (n_2414, n_831, n_830);
  nand g2339 (n_2415, n_829, n_831);
  nand g2340 (n_848, n_2413, n_2414, n_2415);
  xor g2341 (n_2416, n_832, n_833);
  xor g2342 (n_838, n_2416, n_834);
  nand g2343 (n_2417, n_832, n_833);
  nand g2344 (n_2418, n_834, n_833);
  nand g2345 (n_2419, n_832, n_834);
  nand g2346 (n_852, n_2417, n_2418, n_2419);
  xor g2347 (n_2420, n_835, n_836);
  xor g2348 (n_839, n_2420, n_837);
  nand g2349 (n_2421, n_835, n_836);
  nand g2350 (n_2422, n_837, n_836);
  nand g2351 (n_2423, n_835, n_837);
  nand g2352 (n_854, n_2421, n_2422, n_2423);
  xor g2353 (n_2424, n_838, n_839);
  xor g2354 (n_187, n_2424, n_840);
  nand g2355 (n_2425, n_838, n_839);
  nand g2356 (n_2426, n_840, n_839);
  nand g2357 (n_2427, n_838, n_840);
  nand g2358 (n_101, n_2425, n_2426, n_2427);
  xor g2360 (n_843, n_2300, A[36]);
  nand g2362 (n_2430, A[36], A[44]);
  nand g2363 (n_2431, A[46], A[36]);
  nand g2364 (n_855, n_2301, n_2430, n_2431);
  xor g2366 (n_845, n_1916, A[40]);
  xor g2371 (n_2436, A[38], A[48]);
  xor g2372 (n_846, n_2436, A[42]);
  nand g2373 (n_2437, A[38], A[48]);
  nand g2374 (n_2438, A[42], A[48]);
  nand g2376 (n_858, n_2437, n_2438, n_2375);
  xor g2377 (n_2440, A[50], n_841);
  xor g2378 (n_849, n_2440, n_842);
  nand g2379 (n_2441, A[50], n_841);
  nand g2380 (n_2442, n_842, n_841);
  nand g2381 (n_2443, A[50], n_842);
  nand g2382 (n_861, n_2441, n_2442, n_2443);
  xor g2383 (n_2444, n_843, n_844);
  xor g2384 (n_850, n_2444, n_845);
  nand g2385 (n_2445, n_843, n_844);
  nand g2386 (n_2446, n_845, n_844);
  nand g2387 (n_2447, n_843, n_845);
  nand g2388 (n_862, n_2445, n_2446, n_2447);
  xor g2389 (n_2448, n_846, n_847);
  xor g2390 (n_851, n_2448, n_848);
  nand g2391 (n_2449, n_846, n_847);
  nand g2392 (n_2450, n_848, n_847);
  nand g2393 (n_2451, n_846, n_848);
  nand g2394 (n_866, n_2449, n_2450, n_2451);
  xor g2395 (n_2452, n_849, n_850);
  xor g2396 (n_853, n_2452, n_851);
  nand g2397 (n_2453, n_849, n_850);
  nand g2398 (n_2454, n_851, n_850);
  nand g2399 (n_2455, n_849, n_851);
  nand g2400 (n_868, n_2453, n_2454, n_2455);
  xor g2401 (n_2456, n_852, n_853);
  xor g2402 (n_186, n_2456, n_854);
  nand g2403 (n_2457, n_852, n_853);
  nand g2404 (n_2458, n_854, n_853);
  nand g2405 (n_2459, n_852, n_854);
  nand g2406 (n_100, n_2457, n_2458, n_2459);
  xor g2408 (n_857, n_2332, A[37]);
  nand g2410 (n_2462, A[37], A[45]);
  nand g2411 (n_2463, A[47], A[37]);
  nand g2412 (n_869, n_2333, n_2462, n_2463);
  xor g2414 (n_859, n_1948, A[41]);
  xor g2419 (n_2468, A[39], A[49]);
  xor g2420 (n_860, n_2468, A[43]);
  nand g2421 (n_2469, A[39], A[49]);
  nand g2422 (n_2470, A[43], A[49]);
  nand g2424 (n_873, n_2469, n_2470, n_2407);
  xor g2425 (n_2472, A[51], n_855);
  xor g2426 (n_863, n_2472, n_772);
  nand g2427 (n_2473, A[51], n_855);
  nand g2428 (n_2474, n_772, n_855);
  nand g2429 (n_2475, A[51], n_772);
  nand g2430 (n_875, n_2473, n_2474, n_2475);
  xor g2431 (n_2476, n_857, n_858);
  xor g2432 (n_864, n_2476, n_859);
  nand g2433 (n_2477, n_857, n_858);
  nand g2434 (n_2478, n_859, n_858);
  nand g2435 (n_2479, n_857, n_859);
  nand g2436 (n_876, n_2477, n_2478, n_2479);
  xor g2437 (n_2480, n_860, n_861);
  xor g2438 (n_865, n_2480, n_862);
  nand g2439 (n_2481, n_860, n_861);
  nand g2440 (n_2482, n_862, n_861);
  nand g2441 (n_2483, n_860, n_862);
  nand g2442 (n_880, n_2481, n_2482, n_2483);
  xor g2443 (n_2484, n_863, n_864);
  xor g2444 (n_867, n_2484, n_865);
  nand g2445 (n_2485, n_863, n_864);
  nand g2446 (n_2486, n_865, n_864);
  nand g2447 (n_2487, n_863, n_865);
  nand g2448 (n_882, n_2485, n_2486, n_2487);
  xor g2449 (n_2488, n_866, n_867);
  xor g2450 (n_185, n_2488, n_868);
  nand g2451 (n_2489, n_866, n_867);
  nand g2452 (n_2490, n_868, n_867);
  nand g2453 (n_2491, n_866, n_868);
  nand g2454 (n_99, n_2489, n_2490, n_2491);
  xor g2456 (n_871, n_2300, A[38]);
  nand g2459 (n_2495, A[46], A[38]);
  nand g2460 (n_883, n_2301, n_2237, n_2495);
  xor g2462 (n_872, n_1980, A[40]);
  nand g2466 (n_884, n_1981, n_2111, n_2173);
  xor g2467 (n_2500, A[50], A[52]);
  xor g2468 (n_874, n_2500, A[42]);
  nand g2469 (n_2501, A[50], A[52]);
  nand g2470 (n_2502, A[42], A[52]);
  nand g2471 (n_2503, A[50], A[42]);
  nand g2472 (n_887, n_2501, n_2502, n_2503);
  xor g2473 (n_2504, A[48], n_869);
  xor g2474 (n_877, n_2504, n_787);
  nand g2475 (n_2505, A[48], n_869);
  nand g2476 (n_2506, n_787, n_869);
  nand g2477 (n_2507, A[48], n_787);
  nand g2478 (n_889, n_2505, n_2506, n_2507);
  xor g2479 (n_2508, n_871, n_872);
  xor g2480 (n_878, n_2508, n_873);
  nand g2481 (n_2509, n_871, n_872);
  nand g2482 (n_2510, n_873, n_872);
  nand g2483 (n_2511, n_871, n_873);
  nand g2484 (n_890, n_2509, n_2510, n_2511);
  xor g2485 (n_2512, n_874, n_875);
  xor g2486 (n_879, n_2512, n_876);
  nand g2487 (n_2513, n_874, n_875);
  nand g2488 (n_2514, n_876, n_875);
  nand g2489 (n_2515, n_874, n_876);
  nand g2490 (n_894, n_2513, n_2514, n_2515);
  xor g2491 (n_2516, n_877, n_878);
  xor g2492 (n_881, n_2516, n_879);
  nand g2493 (n_2517, n_877, n_878);
  nand g2494 (n_2518, n_879, n_878);
  nand g2495 (n_2519, n_877, n_879);
  nand g2496 (n_896, n_2517, n_2518, n_2519);
  xor g2497 (n_2520, n_880, n_881);
  xor g2498 (n_184, n_2520, n_882);
  nand g2499 (n_2521, n_880, n_881);
  nand g2500 (n_2522, n_882, n_881);
  nand g2501 (n_2523, n_880, n_882);
  nand g2502 (n_98, n_2521, n_2522, n_2523);
  xor g2504 (n_885, n_2332, A[39]);
  nand g2507 (n_2527, A[47], A[39]);
  nand g2508 (n_897, n_2333, n_2269, n_2527);
  xor g2510 (n_886, n_2012, A[41]);
  nand g2514 (n_898, n_2013, n_2143, n_2205);
  xor g2515 (n_2532, A[51], A[53]);
  xor g2516 (n_888, n_2532, A[43]);
  nand g2517 (n_2533, A[51], A[53]);
  nand g2518 (n_2534, A[43], A[53]);
  nand g2519 (n_2535, A[51], A[43]);
  nand g2520 (n_901, n_2533, n_2534, n_2535);
  xor g2521 (n_2536, A[49], n_883);
  xor g2522 (n_891, n_2536, n_884);
  nand g2523 (n_2537, A[49], n_883);
  nand g2524 (n_2538, n_884, n_883);
  nand g2525 (n_2539, A[49], n_884);
  nand g2526 (n_903, n_2537, n_2538, n_2539);
  xor g2527 (n_2540, n_885, n_886);
  xor g2528 (n_892, n_2540, n_887);
  nand g2529 (n_2541, n_885, n_886);
  nand g2530 (n_2542, n_887, n_886);
  nand g2531 (n_2543, n_885, n_887);
  nand g2532 (n_904, n_2541, n_2542, n_2543);
  xor g2533 (n_2544, n_888, n_889);
  xor g2534 (n_893, n_2544, n_890);
  nand g2535 (n_2545, n_888, n_889);
  nand g2536 (n_2546, n_890, n_889);
  nand g2537 (n_2547, n_888, n_890);
  nand g2538 (n_908, n_2545, n_2546, n_2547);
  xor g2539 (n_2548, n_891, n_892);
  xor g2540 (n_895, n_2548, n_893);
  nand g2541 (n_2549, n_891, n_892);
  nand g2542 (n_2550, n_893, n_892);
  nand g2543 (n_2551, n_891, n_893);
  nand g2544 (n_910, n_2549, n_2550, n_2551);
  xor g2545 (n_2552, n_894, n_895);
  xor g2546 (n_183, n_2552, n_896);
  nand g2547 (n_2553, n_894, n_895);
  nand g2548 (n_2554, n_896, n_895);
  nand g2549 (n_2555, n_894, n_896);
  nand g2550 (n_97, n_2553, n_2554, n_2555);
  xor g2552 (n_899, n_2364, A[38]);
  nand g2556 (n_911, n_2303, n_2109, n_2495);
  xor g2557 (n_2560, A[36], A[44]);
  xor g2558 (n_900, n_2560, A[48]);
  nand g2560 (n_2562, A[48], A[44]);
  nand g2561 (n_2563, A[36], A[48]);
  nand g2562 (n_914, n_2430, n_2562, n_2563);
  xor g2563 (n_2564, A[54], A[52]);
  xor g2564 (n_902, n_2564, A[50]);
  nand g2565 (n_2565, A[54], A[52]);
  nand g2567 (n_2567, A[54], A[50]);
  nand g2568 (n_915, n_2565, n_2501, n_2567);
  xor g2569 (n_2568, A[42], n_897);
  xor g2570 (n_905, n_2568, n_898);
  nand g2571 (n_2569, A[42], n_897);
  nand g2572 (n_2570, n_898, n_897);
  nand g2573 (n_2571, A[42], n_898);
  nand g2574 (n_917, n_2569, n_2570, n_2571);
  xor g2575 (n_2572, n_899, n_900);
  xor g2576 (n_906, n_2572, n_901);
  nand g2577 (n_2573, n_899, n_900);
  nand g2578 (n_2574, n_901, n_900);
  nand g2579 (n_2575, n_899, n_901);
  nand g2580 (n_918, n_2573, n_2574, n_2575);
  xor g2581 (n_2576, n_902, n_903);
  xor g2582 (n_907, n_2576, n_904);
  nand g2583 (n_2577, n_902, n_903);
  nand g2584 (n_2578, n_904, n_903);
  nand g2585 (n_2579, n_902, n_904);
  nand g2586 (n_922, n_2577, n_2578, n_2579);
  xor g2587 (n_2580, n_905, n_906);
  xor g2588 (n_909, n_2580, n_907);
  nand g2589 (n_2581, n_905, n_906);
  nand g2590 (n_2582, n_907, n_906);
  nand g2591 (n_2583, n_905, n_907);
  nand g2592 (n_924, n_2581, n_2582, n_2583);
  xor g2593 (n_2584, n_908, n_909);
  xor g2594 (n_182, n_2584, n_910);
  nand g2595 (n_2585, n_908, n_909);
  nand g2596 (n_2586, n_910, n_909);
  nand g2597 (n_2587, n_908, n_910);
  nand g2598 (n_96, n_2585, n_2586, n_2587);
  xor g2600 (n_912, n_2396, A[39]);
  nand g2604 (n_925, n_2335, n_2141, n_2527);
  xor g2605 (n_2592, A[37], A[45]);
  xor g2606 (n_913, n_2592, A[49]);
  nand g2608 (n_2594, A[49], A[45]);
  nand g2609 (n_2595, A[37], A[49]);
  nand g2610 (n_927, n_2462, n_2594, n_2595);
  xor g2611 (n_2596, A[55], A[53]);
  xor g2612 (n_916, n_2596, A[51]);
  nand g2613 (n_2597, A[55], A[53]);
  nand g2615 (n_2599, A[55], A[51]);
  nand g2616 (n_928, n_2597, n_2533, n_2599);
  xor g2617 (n_2600, A[43], n_911);
  xor g2618 (n_919, n_2600, n_912);
  nand g2619 (n_2601, A[43], n_911);
  nand g2620 (n_2602, n_912, n_911);
  nand g2621 (n_2603, A[43], n_912);
  nand g2622 (n_932, n_2601, n_2602, n_2603);
  xor g2623 (n_2604, n_913, n_914);
  xor g2624 (n_920, n_2604, n_915);
  nand g2625 (n_2605, n_913, n_914);
  nand g2626 (n_2606, n_915, n_914);
  nand g2627 (n_2607, n_913, n_915);
  nand g2628 (n_931, n_2605, n_2606, n_2607);
  xor g2629 (n_2608, n_916, n_917);
  xor g2630 (n_921, n_2608, n_918);
  nand g2631 (n_2609, n_916, n_917);
  nand g2632 (n_2610, n_918, n_917);
  nand g2633 (n_2611, n_916, n_918);
  nand g2634 (n_935, n_2609, n_2610, n_2611);
  xor g2635 (n_2612, n_919, n_920);
  xor g2636 (n_923, n_2612, n_921);
  nand g2637 (n_2613, n_919, n_920);
  nand g2638 (n_2614, n_921, n_920);
  nand g2639 (n_2615, n_919, n_921);
  nand g2640 (n_938, n_2613, n_2614, n_2615);
  xor g2641 (n_2616, n_922, n_923);
  xor g2642 (n_181, n_2616, n_924);
  nand g2643 (n_2617, n_922, n_923);
  nand g2644 (n_2618, n_924, n_923);
  nand g2645 (n_2619, n_922, n_924);
  nand g2646 (n_95, n_2617, n_2618, n_2619);
  xor g2653 (n_2624, A[44], A[54]);
  xor g2654 (n_929, n_2624, A[42]);
  nand g2655 (n_2625, A[44], A[54]);
  nand g2656 (n_2626, A[42], A[54]);
  nand g2657 (n_2627, A[44], A[42]);
  nand g2658 (n_941, n_2625, n_2626, n_2627);
  xor g2659 (n_2628, A[50], A[48]);
  xor g2660 (n_930, n_2628, A[52]);
  nand g2661 (n_2629, A[50], A[48]);
  nand g2662 (n_2630, A[52], A[48]);
  nand g2664 (n_942, n_2629, n_2630, n_2501);
  xor g2665 (n_2632, A[56], n_925);
  xor g2666 (n_933, n_2632, n_899);
  nand g2667 (n_2633, A[56], n_925);
  nand g2668 (n_2634, n_899, n_925);
  nand g2669 (n_2635, A[56], n_899);
  nand g2670 (n_945, n_2633, n_2634, n_2635);
  xor g2671 (n_2636, n_927, n_928);
  xor g2672 (n_934, n_2636, n_929);
  nand g2673 (n_2637, n_927, n_928);
  nand g2674 (n_2638, n_929, n_928);
  nand g2675 (n_2639, n_927, n_929);
  nand g2676 (n_948, n_2637, n_2638, n_2639);
  xor g2677 (n_2640, n_930, n_931);
  xor g2678 (n_936, n_2640, n_932);
  nand g2679 (n_2641, n_930, n_931);
  nand g2680 (n_2642, n_932, n_931);
  nand g2681 (n_2643, n_930, n_932);
  nand g2682 (n_949, n_2641, n_2642, n_2643);
  xor g2683 (n_2644, n_933, n_934);
  xor g2684 (n_937, n_2644, n_935);
  nand g2685 (n_2645, n_933, n_934);
  nand g2686 (n_2646, n_935, n_934);
  nand g2687 (n_2647, n_933, n_935);
  nand g2688 (n_952, n_2645, n_2646, n_2647);
  xor g2689 (n_2648, n_936, n_937);
  xor g2690 (n_180, n_2648, n_938);
  nand g2691 (n_2649, n_936, n_937);
  nand g2692 (n_2650, n_938, n_937);
  nand g2693 (n_2651, n_936, n_938);
  nand g2694 (n_94, n_2649, n_2650, n_2651);
  xor g2701 (n_2656, A[45], A[55]);
  xor g2702 (n_943, n_2656, A[43]);
  nand g2703 (n_2657, A[45], A[55]);
  nand g2704 (n_2658, A[43], A[55]);
  nand g2705 (n_2659, A[45], A[43]);
  nand g2706 (n_955, n_2657, n_2658, n_2659);
  xor g2707 (n_2660, A[51], A[49]);
  xor g2708 (n_944, n_2660, A[53]);
  nand g2709 (n_2661, A[51], A[49]);
  nand g2710 (n_2662, A[53], A[49]);
  nand g2712 (n_956, n_2661, n_2662, n_2533);
  xor g2713 (n_2664, A[57], n_911);
  xor g2714 (n_946, n_2664, n_912);
  nand g2715 (n_2665, A[57], n_911);
  nand g2717 (n_2667, A[57], n_912);
  nand g2718 (n_959, n_2665, n_2602, n_2667);
  xor g2719 (n_2668, n_941, n_942);
  xor g2720 (n_947, n_2668, n_943);
  nand g2721 (n_2669, n_941, n_942);
  nand g2722 (n_2670, n_943, n_942);
  nand g2723 (n_2671, n_941, n_943);
  nand g2724 (n_962, n_2669, n_2670, n_2671);
  xor g2725 (n_2672, n_944, n_945);
  xor g2726 (n_950, n_2672, n_946);
  nand g2727 (n_2673, n_944, n_945);
  nand g2728 (n_2674, n_946, n_945);
  nand g2729 (n_2675, n_944, n_946);
  nand g2730 (n_963, n_2673, n_2674, n_2675);
  xor g2731 (n_2676, n_947, n_948);
  xor g2732 (n_951, n_2676, n_949);
  nand g2733 (n_2677, n_947, n_948);
  nand g2734 (n_2678, n_949, n_948);
  nand g2735 (n_2679, n_947, n_949);
  nand g2736 (n_966, n_2677, n_2678, n_2679);
  xor g2737 (n_2680, n_950, n_951);
  xor g2738 (n_179, n_2680, n_952);
  nand g2739 (n_2681, n_950, n_951);
  nand g2740 (n_2682, n_952, n_951);
  nand g2741 (n_2683, n_950, n_952);
  nand g2742 (n_93, n_2681, n_2682, n_2683);
  xor g2749 (n_2688, A[56], A[52]);
  xor g2750 (n_958, n_2688, A[42]);
  nand g2751 (n_2689, A[56], A[52]);
  nand g2753 (n_2691, A[56], A[42]);
  nand g2754 (n_969, n_2689, n_2502, n_2691);
  xor g2755 (n_2692, A[50], A[58]);
  xor g2756 (n_957, n_2692, A[48]);
  nand g2757 (n_2693, A[50], A[58]);
  nand g2758 (n_2694, A[48], A[58]);
  nand g2760 (n_970, n_2693, n_2694, n_2629);
  xor g2761 (n_2696, A[54], n_925);
  xor g2762 (n_960, n_2696, n_789);
  nand g2763 (n_2697, A[54], n_925);
  nand g2764 (n_2698, n_789, n_925);
  nand g2765 (n_2699, A[54], n_789);
  nand g2766 (n_973, n_2697, n_2698, n_2699);
  xor g2767 (n_2700, n_955, n_956);
  xor g2768 (n_961, n_2700, n_957);
  nand g2769 (n_2701, n_955, n_956);
  nand g2770 (n_2702, n_957, n_956);
  nand g2771 (n_2703, n_955, n_957);
  nand g2772 (n_976, n_2701, n_2702, n_2703);
  xor g2773 (n_2704, n_958, n_959);
  xor g2774 (n_964, n_2704, n_960);
  nand g2775 (n_2705, n_958, n_959);
  nand g2776 (n_2706, n_960, n_959);
  nand g2777 (n_2707, n_958, n_960);
  nand g2778 (n_977, n_2705, n_2706, n_2707);
  xor g2779 (n_2708, n_961, n_962);
  xor g2780 (n_965, n_2708, n_963);
  nand g2781 (n_2709, n_961, n_962);
  nand g2782 (n_2710, n_963, n_962);
  nand g2783 (n_2711, n_961, n_963);
  nand g2784 (n_980, n_2709, n_2710, n_2711);
  xor g2785 (n_2712, n_964, n_965);
  xor g2786 (n_178, n_2712, n_966);
  nand g2787 (n_2713, n_964, n_965);
  nand g2788 (n_2714, n_966, n_965);
  nand g2789 (n_2715, n_964, n_966);
  nand g2790 (n_92, n_2713, n_2714, n_2715);
  xor g2797 (n_2720, A[57], A[53]);
  xor g2798 (n_972, n_2720, A[43]);
  nand g2799 (n_2721, A[57], A[53]);
  nand g2801 (n_2723, A[57], A[43]);
  nand g2802 (n_983, n_2721, n_2534, n_2723);
  xor g2803 (n_2724, A[51], A[59]);
  xor g2804 (n_971, n_2724, A[49]);
  nand g2805 (n_2725, A[51], A[59]);
  nand g2806 (n_2726, A[49], A[59]);
  nand g2808 (n_984, n_2725, n_2726, n_2661);
  xor g2809 (n_2728, A[55], n_799);
  xor g2810 (n_974, n_2728, n_803);
  nand g2811 (n_2729, A[55], n_799);
  nand g2812 (n_2730, n_803, n_799);
  nand g2813 (n_2731, A[55], n_803);
  nand g2814 (n_987, n_2729, n_2730, n_2731);
  xor g2815 (n_2732, n_969, n_970);
  xor g2816 (n_975, n_2732, n_971);
  nand g2817 (n_2733, n_969, n_970);
  nand g2818 (n_2734, n_971, n_970);
  nand g2819 (n_2735, n_969, n_971);
  nand g2820 (n_990, n_2733, n_2734, n_2735);
  xor g2821 (n_2736, n_972, n_973);
  xor g2822 (n_978, n_2736, n_974);
  nand g2823 (n_2737, n_972, n_973);
  nand g2824 (n_2738, n_974, n_973);
  nand g2825 (n_2739, n_972, n_974);
  nand g2826 (n_991, n_2737, n_2738, n_2739);
  xor g2827 (n_2740, n_975, n_976);
  xor g2828 (n_979, n_2740, n_977);
  nand g2829 (n_2741, n_975, n_976);
  nand g2830 (n_2742, n_977, n_976);
  nand g2831 (n_2743, n_975, n_977);
  nand g2832 (n_994, n_2741, n_2742, n_2743);
  xor g2833 (n_2744, n_978, n_979);
  xor g2834 (n_177, n_2744, n_980);
  nand g2835 (n_2745, n_978, n_979);
  nand g2836 (n_2746, n_980, n_979);
  nand g2837 (n_2747, n_978, n_980);
  nand g2838 (n_91, n_2745, n_2746, n_2747);
  xor g2840 (n_982, n_2300, A[60]);
  nand g2842 (n_2750, A[60], A[44]);
  nand g2843 (n_2751, A[46], A[60]);
  nand g2844 (n_996, n_2301, n_2750, n_2751);
  xor g2845 (n_2752, A[54], A[58]);
  xor g2846 (n_986, n_2752, A[52]);
  nand g2847 (n_2753, A[54], A[58]);
  nand g2848 (n_2754, A[52], A[58]);
  nand g2850 (n_997, n_2753, n_2754, n_2565);
  xor g2851 (n_2756, A[42], A[56]);
  xor g2852 (n_985, n_2756, A[50]);
  nand g2854 (n_2758, A[50], A[56]);
  nand g2856 (n_998, n_2691, n_2758, n_2503);
  xor g2858 (n_988, n_2376, n_982);
  nand g2860 (n_2762, n_982, n_813);
  nand g2861 (n_2763, A[48], n_982);
  nand g2862 (n_1001, n_2377, n_2762, n_2763);
  xor g2863 (n_2764, n_983, n_984);
  xor g2864 (n_989, n_2764, n_985);
  nand g2865 (n_2765, n_983, n_984);
  nand g2866 (n_2766, n_985, n_984);
  nand g2867 (n_2767, n_983, n_985);
  nand g2868 (n_1003, n_2765, n_2766, n_2767);
  xor g2869 (n_2768, n_986, n_987);
  xor g2870 (n_992, n_2768, n_988);
  nand g2871 (n_2769, n_986, n_987);
  nand g2872 (n_2770, n_988, n_987);
  nand g2873 (n_2771, n_986, n_988);
  nand g2874 (n_1005, n_2769, n_2770, n_2771);
  xor g2875 (n_2772, n_989, n_990);
  xor g2876 (n_993, n_2772, n_991);
  nand g2877 (n_2773, n_989, n_990);
  nand g2878 (n_2774, n_991, n_990);
  nand g2879 (n_2775, n_989, n_991);
  nand g2880 (n_1008, n_2773, n_2774, n_2775);
  xor g2881 (n_2776, n_992, n_993);
  xor g2882 (n_176, n_2776, n_994);
  nand g2883 (n_2777, n_992, n_993);
  nand g2884 (n_2778, n_994, n_993);
  nand g2885 (n_2779, n_992, n_994);
  nand g2886 (n_90, n_2777, n_2778, n_2779);
  xor g2888 (n_995, n_2332, A[61]);
  nand g2890 (n_2782, A[61], A[45]);
  nand g2891 (n_2783, A[47], A[61]);
  nand g2892 (n_1010, n_2333, n_2782, n_2783);
  xor g2893 (n_2784, A[55], A[59]);
  xor g2894 (n_1000, n_2784, A[53]);
  nand g2895 (n_2785, A[55], A[59]);
  nand g2896 (n_2786, A[53], A[59]);
  nand g2898 (n_1011, n_2785, n_2786, n_2597);
  xor g2899 (n_2788, A[43], A[57]);
  xor g2900 (n_999, n_2788, A[51]);
  nand g2902 (n_2790, A[51], A[57]);
  nand g2904 (n_1012, n_2723, n_2790, n_2535);
  xor g2905 (n_2792, A[49], n_995);
  xor g2906 (n_1004, n_2792, n_996);
  nand g2907 (n_2793, A[49], n_995);
  nand g2908 (n_2794, n_996, n_995);
  nand g2909 (n_2795, A[49], n_996);
  nand g2910 (n_1015, n_2793, n_2794, n_2795);
  xor g2911 (n_2796, n_997, n_998);
  xor g2912 (n_1002, n_2796, n_999);
  nand g2913 (n_2797, n_997, n_998);
  nand g2914 (n_2798, n_999, n_998);
  nand g2915 (n_2799, n_997, n_999);
  nand g2916 (n_1017, n_2797, n_2798, n_2799);
  xor g2917 (n_2800, n_1000, n_1001);
  xor g2918 (n_1006, n_2800, n_1002);
  nand g2919 (n_2801, n_1000, n_1001);
  nand g2920 (n_2802, n_1002, n_1001);
  nand g2921 (n_2803, n_1000, n_1002);
  nand g2922 (n_1019, n_2801, n_2802, n_2803);
  xor g2923 (n_2804, n_1003, n_1004);
  xor g2924 (n_1007, n_2804, n_1005);
  nand g2925 (n_2805, n_1003, n_1004);
  nand g2926 (n_2806, n_1005, n_1004);
  nand g2927 (n_2807, n_1003, n_1005);
  nand g2928 (n_1021, n_2805, n_2806, n_2807);
  xor g2929 (n_2808, n_1006, n_1007);
  xor g2930 (n_175, n_2808, n_1008);
  nand g2931 (n_2809, n_1006, n_1007);
  nand g2932 (n_2810, n_1008, n_1007);
  nand g2933 (n_2811, n_1006, n_1008);
  nand g2934 (n_89, n_2809, n_2810, n_2811);
  xor g2941 (n_2816, A[48], A[56]);
  xor g2942 (n_1014, n_2816, A[62]);
  nand g2943 (n_2817, A[48], A[56]);
  nand g2944 (n_2818, A[62], A[56]);
  nand g2945 (n_2819, A[48], A[62]);
  nand g2946 (n_1025, n_2817, n_2818, n_2819);
  xor g2953 (n_2824, A[50], n_982);
  xor g2954 (n_1018, n_2824, n_1010);
  nand g2955 (n_2825, A[50], n_982);
  nand g2956 (n_2826, n_1010, n_982);
  nand g2957 (n_2827, A[50], n_1010);
  nand g2958 (n_1029, n_2825, n_2826, n_2827);
  xor g2959 (n_2828, n_1011, n_1012);
  xor g2960 (n_1016, n_2828, n_986);
  nand g2961 (n_2829, n_1011, n_1012);
  nand g2962 (n_2830, n_986, n_1012);
  nand g2963 (n_2831, n_1011, n_986);
  nand g2964 (n_1031, n_2829, n_2830, n_2831);
  xor g2965 (n_2832, n_1014, n_1015);
  xor g2966 (n_1020, n_2832, n_1016);
  nand g2967 (n_2833, n_1014, n_1015);
  nand g2968 (n_2834, n_1016, n_1015);
  nand g2969 (n_2835, n_1014, n_1016);
  nand g2970 (n_1033, n_2833, n_2834, n_2835);
  xor g2971 (n_2836, n_1017, n_1018);
  xor g2972 (n_1022, n_2836, n_1019);
  nand g2973 (n_2837, n_1017, n_1018);
  nand g2974 (n_2838, n_1019, n_1018);
  nand g2975 (n_2839, n_1017, n_1019);
  nand g2976 (n_1036, n_2837, n_2838, n_2839);
  xor g2977 (n_2840, n_1020, n_1021);
  xor g2978 (n_174, n_2840, n_1022);
  nand g2979 (n_2841, n_1020, n_1021);
  nand g2980 (n_2842, n_1022, n_1021);
  nand g2981 (n_2843, n_1020, n_1022);
  nand g2982 (n_88, n_2841, n_2842, n_2843);
  xor g2989 (n_2848, A[49], A[57]);
  xor g2990 (n_1028, n_2848, A[63]);
  nand g2991 (n_2849, A[49], A[57]);
  nand g2992 (n_2850, A[63], A[57]);
  nand g2993 (n_2851, A[49], A[63]);
  nand g2994 (n_1038, n_2849, n_2850, n_2851);
  xor g3001 (n_2856, A[51], n_995);
  xor g3002 (n_1032, n_2856, n_996);
  nand g3003 (n_2857, A[51], n_995);
  nand g3005 (n_2859, A[51], n_996);
  nand g3006 (n_1043, n_2857, n_2794, n_2859);
  xor g3007 (n_2860, n_1025, n_997);
  xor g3008 (n_1030, n_2860, n_1000);
  nand g3009 (n_2861, n_1025, n_997);
  nand g3010 (n_2862, n_1000, n_997);
  nand g3011 (n_2863, n_1025, n_1000);
  nand g3012 (n_1045, n_2861, n_2862, n_2863);
  xor g3013 (n_2864, n_1028, n_1029);
  xor g3014 (n_1034, n_2864, n_1030);
  nand g3015 (n_2865, n_1028, n_1029);
  nand g3016 (n_2866, n_1030, n_1029);
  nand g3017 (n_2867, n_1028, n_1030);
  nand g3018 (n_1047, n_2865, n_2866, n_2867);
  xor g3019 (n_2868, n_1031, n_1032);
  xor g3020 (n_1035, n_2868, n_1033);
  nand g3021 (n_2869, n_1031, n_1032);
  nand g3022 (n_2870, n_1033, n_1032);
  nand g3023 (n_2871, n_1031, n_1033);
  nand g3024 (n_1050, n_2869, n_2870, n_2871);
  xor g3025 (n_2872, n_1034, n_1035);
  xor g3026 (n_173, n_2872, n_1036);
  nand g3027 (n_2873, n_1034, n_1035);
  nand g3028 (n_2874, n_1036, n_1035);
  nand g3029 (n_2875, n_1034, n_1036);
  nand g3030 (n_87, n_2873, n_2874, n_2875);
  xor g3031 (n_2876, A[46], A[64]);
  xor g3032 (n_1041, n_2876, A[58]);
  nand g3033 (n_2877, A[46], A[64]);
  nand g3034 (n_2878, A[58], A[64]);
  nand g3035 (n_2879, A[46], A[58]);
  nand g3036 (n_1055, n_2877, n_2878, n_2879);
  xor g3038 (n_1042, n_2628, A[62]);
  nand g3041 (n_2883, A[50], A[62]);
  nand g3042 (n_1056, n_2629, n_2819, n_2883);
  xor g3043 (n_2884, A[56], A[60]);
  xor g3044 (n_1040, n_2884, A[54]);
  nand g3045 (n_2885, A[56], A[60]);
  nand g3046 (n_2886, A[54], A[60]);
  nand g3047 (n_2887, A[56], A[54]);
  nand g3048 (n_1053, n_2885, n_2886, n_2887);
  xor g3049 (n_2888, A[52], n_1010);
  xor g3050 (n_1044, n_2888, n_1038);
  nand g3051 (n_2889, A[52], n_1010);
  nand g3052 (n_2890, n_1038, n_1010);
  nand g3053 (n_2891, A[52], n_1038);
  nand g3054 (n_1059, n_2889, n_2890, n_2891);
  xor g3055 (n_2892, n_1011, n_1040);
  xor g3056 (n_1046, n_2892, n_1041);
  nand g3057 (n_2893, n_1011, n_1040);
  nand g3058 (n_2894, n_1041, n_1040);
  nand g3059 (n_2895, n_1011, n_1041);
  nand g3060 (n_1061, n_2893, n_2894, n_2895);
  xor g3061 (n_2896, n_1042, n_1043);
  xor g3062 (n_1048, n_2896, n_1044);
  nand g3063 (n_2897, n_1042, n_1043);
  nand g3064 (n_2898, n_1044, n_1043);
  nand g3065 (n_2899, n_1042, n_1044);
  nand g3066 (n_1063, n_2897, n_2898, n_2899);
  xor g3067 (n_2900, n_1045, n_1046);
  xor g3068 (n_1049, n_2900, n_1047);
  nand g3069 (n_2901, n_1045, n_1046);
  nand g3070 (n_2902, n_1047, n_1046);
  nand g3071 (n_2903, n_1045, n_1047);
  nand g3072 (n_1066, n_2901, n_2902, n_2903);
  xor g3073 (n_2904, n_1048, n_1049);
  xor g3074 (n_172, n_2904, n_1050);
  nand g3075 (n_2905, n_1048, n_1049);
  nand g3076 (n_2906, n_1050, n_1049);
  nand g3077 (n_2907, n_1048, n_1050);
  nand g3078 (n_86, n_2905, n_2906, n_2907);
  xor g3081 (n_2908, A[65], A[47]);
  xor g3082 (n_1054, n_2908, A[49]);
  nand g3083 (n_2909, A[65], A[47]);
  nand g3084 (n_2910, A[49], A[47]);
  nand g3085 (n_2911, A[65], A[49]);
  nand g3086 (n_1071, n_2909, n_2910, n_2911);
  xor g3088 (n_1058, n_2724, A[57]);
  nand g3091 (n_2915, A[59], A[57]);
  nand g3092 (n_1072, n_2725, n_2790, n_2915);
  xor g3093 (n_2916, A[63], A[61]);
  xor g3094 (n_1057, n_2916, A[55]);
  nand g3095 (n_2917, A[63], A[61]);
  nand g3096 (n_2918, A[55], A[61]);
  nand g3097 (n_2919, A[63], A[55]);
  nand g3098 (n_1070, n_2917, n_2918, n_2919);
  xor g3099 (n_2920, A[53], n_1053);
  xor g3100 (n_1062, n_2920, n_1054);
  nand g3101 (n_2921, A[53], n_1053);
  nand g3102 (n_2922, n_1054, n_1053);
  nand g3103 (n_2923, A[53], n_1054);
  nand g3104 (n_1076, n_2921, n_2922, n_2923);
  xor g3105 (n_2924, n_1055, n_1056);
  xor g3106 (n_1060, n_2924, n_1057);
  nand g3107 (n_2925, n_1055, n_1056);
  nand g3108 (n_2926, n_1057, n_1056);
  nand g3109 (n_2927, n_1055, n_1057);
  nand g3110 (n_1078, n_2925, n_2926, n_2927);
  xor g3111 (n_2928, n_1058, n_1059);
  xor g3112 (n_1064, n_2928, n_1060);
  nand g3113 (n_2929, n_1058, n_1059);
  nand g3114 (n_2930, n_1060, n_1059);
  nand g3115 (n_2931, n_1058, n_1060);
  nand g3116 (n_1080, n_2929, n_2930, n_2931);
  xor g3117 (n_2932, n_1061, n_1062);
  xor g3118 (n_1065, n_2932, n_1063);
  nand g3119 (n_2933, n_1061, n_1062);
  nand g3120 (n_2934, n_1063, n_1062);
  nand g3121 (n_2935, n_1061, n_1063);
  nand g3122 (n_1083, n_2933, n_2934, n_2935);
  xor g3123 (n_2936, n_1064, n_1065);
  xor g3124 (n_171, n_2936, n_1066);
  nand g3125 (n_2937, n_1064, n_1065);
  nand g3126 (n_2938, n_1066, n_1065);
  nand g3127 (n_2939, n_1064, n_1066);
  nand g3128 (n_85, n_2937, n_2938, n_2939);
  nand g3139 (n_2945, A[65], A[64]);
  nand g3140 (n_2946, A[56], A[64]);
  nand g3141 (n_2947, A[65], A[56]);
  nand g3142 (n_1086, n_2945, n_2946, n_2947);
  xor g3143 (n_2948, A[62], A[60]);
  xor g3144 (n_1073, n_2948, A[54]);
  nand g3145 (n_2949, A[62], A[60]);
  nand g3147 (n_2951, A[62], A[54]);
  nand g3148 (n_1087, n_2949, n_2886, n_2951);
  xor g3149 (n_2952, A[52], n_1070);
  xor g3150 (n_1077, n_2952, n_1071);
  nand g3151 (n_2953, A[52], n_1070);
  nand g3152 (n_2954, n_1071, n_1070);
  nand g3153 (n_2955, A[52], n_1071);
  nand g3154 (n_1091, n_2953, n_2954, n_2955);
  xor g3155 (n_2956, n_1072, n_1073);
  xor g3156 (n_1079, n_2956, n_957);
  nand g3157 (n_2957, n_1072, n_1073);
  nand g3158 (n_2958, n_957, n_1073);
  nand g3159 (n_2959, n_1072, n_957);
  nand g3160 (n_1093, n_2957, n_2958, n_2959);
  xor g3161 (n_2960, n_1075, n_1076);
  xor g3162 (n_1081, n_2960, n_1077);
  nand g3163 (n_2961, n_1075, n_1076);
  nand g3164 (n_2962, n_1077, n_1076);
  nand g3165 (n_2963, n_1075, n_1077);
  nand g3166 (n_1095, n_2961, n_2962, n_2963);
  xor g3167 (n_2964, n_1078, n_1079);
  xor g3168 (n_1082, n_2964, n_1080);
  nand g3169 (n_2965, n_1078, n_1079);
  nand g3170 (n_2966, n_1080, n_1079);
  nand g3171 (n_2967, n_1078, n_1080);
  nand g3172 (n_1098, n_2965, n_2966, n_2967);
  xor g3173 (n_2968, n_1081, n_1082);
  xor g3174 (n_170, n_2968, n_1083);
  nand g3175 (n_2969, n_1081, n_1082);
  nand g3176 (n_2970, n_1083, n_1082);
  nand g3177 (n_2971, n_1081, n_1083);
  nand g3178 (n_84, n_2969, n_2970, n_2971);
  xor g3180 (n_1089, n_2972, A[59]);
  nand g3182 (n_2974, A[59], A[63]);
  nand g3184 (n_1101, n_2973, n_2974, n_2975);
  xor g3186 (n_1090, n_2660, A[57]);
  nand g3190 (n_1102, n_2661, n_2849, n_2790);
  xor g3192 (n_1088, n_2980, A[55]);
  nand g3196 (n_1103, n_2981, n_2918, n_2983);
  xor g3197 (n_2984, A[53], n_970);
  xor g3198 (n_1092, n_2984, n_1086);
  nand g3199 (n_2985, A[53], n_970);
  nand g3200 (n_2986, n_1086, n_970);
  nand g3201 (n_2987, A[53], n_1086);
  nand g3202 (n_1107, n_2985, n_2986, n_2987);
  xor g3203 (n_2988, n_1087, n_1088);
  xor g3204 (n_1094, n_2988, n_1089);
  nand g3205 (n_2989, n_1087, n_1088);
  nand g3206 (n_2990, n_1089, n_1088);
  nand g3207 (n_2991, n_1087, n_1089);
  nand g3208 (n_1109, n_2989, n_2990, n_2991);
  xor g3209 (n_2992, n_1090, n_1091);
  xor g3210 (n_1096, n_2992, n_1092);
  nand g3211 (n_2993, n_1090, n_1091);
  nand g3212 (n_2994, n_1092, n_1091);
  nand g3213 (n_2995, n_1090, n_1092);
  nand g3214 (n_1111, n_2993, n_2994, n_2995);
  xor g3215 (n_2996, n_1093, n_1094);
  xor g3216 (n_1097, n_2996, n_1095);
  nand g3217 (n_2997, n_1093, n_1094);
  nand g3218 (n_2998, n_1095, n_1094);
  nand g3219 (n_2999, n_1093, n_1095);
  nand g3220 (n_1113, n_2997, n_2998, n_2999);
  xor g3221 (n_3000, n_1096, n_1097);
  xor g3222 (n_169, n_3000, n_1098);
  nand g3223 (n_3001, n_1096, n_1097);
  nand g3224 (n_3002, n_1098, n_1097);
  nand g3225 (n_3003, n_1096, n_1098);
  nand g3226 (n_83, n_3001, n_3002, n_3003);
  xor g3229 (n_3004, A[62], A[50]);
  xor g3230 (n_1105, n_3004, A[58]);
  nand g3233 (n_3007, A[62], A[58]);
  nand g3234 (n_1116, n_2883, n_2693, n_3007);
  xor g3242 (n_1106, n_3012, n_1101);
  nand g3245 (n_3015, A[52], n_1101);
  nand g3246 (n_1120, n_3013, n_3014, n_3015);
  xor g3247 (n_3016, n_1102, n_1103);
  xor g3248 (n_1108, n_3016, n_1040);
  nand g3249 (n_3017, n_1102, n_1103);
  nand g3250 (n_3018, n_1040, n_1103);
  nand g3251 (n_3019, n_1102, n_1040);
  nand g3252 (n_1122, n_3017, n_3018, n_3019);
  xor g3253 (n_3020, n_1105, n_1106);
  xor g3254 (n_1110, n_3020, n_1107);
  nand g3255 (n_3021, n_1105, n_1106);
  nand g3256 (n_3022, n_1107, n_1106);
  nand g3257 (n_3023, n_1105, n_1107);
  nand g3258 (n_1123, n_3021, n_3022, n_3023);
  xor g3259 (n_3024, n_1108, n_1109);
  xor g3260 (n_1112, n_3024, n_1110);
  nand g3261 (n_3025, n_1108, n_1109);
  nand g3262 (n_3026, n_1110, n_1109);
  nand g3263 (n_3027, n_1108, n_1110);
  nand g3264 (n_1126, n_3025, n_3026, n_3027);
  xor g3265 (n_3028, n_1111, n_1112);
  xor g3266 (n_168, n_3028, n_1113);
  nand g3267 (n_3029, n_1111, n_1112);
  nand g3268 (n_3030, n_1113, n_1112);
  nand g3269 (n_3031, n_1111, n_1113);
  nand g3270 (n_82, n_3029, n_3030, n_3031);
  xor g3277 (n_3036, A[51], A[57]);
  xor g3278 (n_1118, n_3036, A[61]);
  nand g3280 (n_3038, A[61], A[57]);
  nand g3281 (n_3039, A[51], A[61]);
  nand g3282 (n_1130, n_2790, n_3038, n_3039);
  xor g3284 (n_1119, n_2596, A[64]);
  nand g3286 (n_3042, A[64], A[53]);
  nand g3287 (n_3043, A[55], A[64]);
  nand g3288 (n_1133, n_2597, n_3042, n_3043);
  xor g3289 (n_3044, n_1053, n_1116);
  xor g3290 (n_1121, n_3044, n_1089);
  nand g3291 (n_3045, n_1053, n_1116);
  nand g3292 (n_3046, n_1089, n_1116);
  nand g3293 (n_3047, n_1053, n_1089);
  nand g3294 (n_1135, n_3045, n_3046, n_3047);
  xor g3295 (n_3048, n_1118, n_1119);
  xor g3296 (n_1124, n_3048, n_1120);
  nand g3297 (n_3049, n_1118, n_1119);
  nand g3298 (n_3050, n_1120, n_1119);
  nand g3299 (n_3051, n_1118, n_1120);
  nand g3300 (n_1137, n_3049, n_3050, n_3051);
  xor g3301 (n_3052, n_1121, n_1122);
  xor g3302 (n_1125, n_3052, n_1123);
  nand g3303 (n_3053, n_1121, n_1122);
  nand g3304 (n_3054, n_1123, n_1122);
  nand g3305 (n_3055, n_1121, n_1123);
  nand g3306 (n_1139, n_3053, n_3054, n_3055);
  xor g3307 (n_3056, n_1124, n_1125);
  xor g3308 (n_167, n_3056, n_1126);
  nand g3309 (n_3057, n_1124, n_1125);
  nand g3310 (n_3058, n_1126, n_1125);
  nand g3311 (n_3059, n_1124, n_1126);
  nand g3312 (n_166, n_3057, n_3058, n_3059);
  xor g3315 (n_3060, A[62], A[58]);
  xor g3316 (n_1132, n_3060, A[56]);
  nand g3318 (n_3062, A[56], A[58]);
  nand g3320 (n_1141, n_3007, n_3062, n_2818);
  xor g3321 (n_3064, A[60], A[54]);
  xor g3322 (n_1131, n_3064, A[52]);
  nand g3325 (n_3067, A[60], A[52]);
  nand g3326 (n_1142, n_2886, n_2565, n_3067);
  xor g3328 (n_1134, n_3068, n_1130);
  nand g3330 (n_3070, n_1130, n_1101);
  nand g3332 (n_1146, n_3014, n_3070, n_3071);
  xor g3333 (n_3072, n_1131, n_1132);
  xor g3334 (n_1136, n_3072, n_1133);
  nand g3335 (n_3073, n_1131, n_1132);
  nand g3336 (n_3074, n_1133, n_1132);
  nand g3337 (n_3075, n_1131, n_1133);
  nand g3338 (n_1147, n_3073, n_3074, n_3075);
  xor g3339 (n_3076, n_1134, n_1135);
  xor g3340 (n_1138, n_3076, n_1136);
  nand g3341 (n_3077, n_1134, n_1135);
  nand g3342 (n_3078, n_1136, n_1135);
  nand g3343 (n_3079, n_1134, n_1136);
  nand g3344 (n_1150, n_3077, n_3078, n_3079);
  xor g3345 (n_3080, n_1137, n_1138);
  xor g3346 (n_81, n_3080, n_1139);
  nand g3347 (n_3081, n_1137, n_1138);
  nand g3348 (n_3082, n_1139, n_1138);
  nand g3349 (n_3083, n_1137, n_1139);
  nand g3350 (n_80, n_3081, n_3082, n_3083);
  xor g3357 (n_3088, A[57], A[61]);
  xor g3358 (n_1143, n_3088, A[55]);
  nand g3361 (n_3091, A[57], A[55]);
  nand g3362 (n_1153, n_3038, n_2918, n_3091);
  xor g3363 (n_3092, A[53], A[64]);
  xor g3364 (n_1145, n_3092, n_1141);
  nand g3366 (n_3094, n_1141, A[64]);
  nand g3367 (n_3095, A[53], n_1141);
  nand g3368 (n_1157, n_3042, n_3094, n_3095);
  xor g3369 (n_3096, n_1142, n_1143);
  xor g3370 (n_1148, n_3096, n_1089);
  nand g3371 (n_3097, n_1142, n_1143);
  nand g3372 (n_3098, n_1089, n_1143);
  nand g3373 (n_3099, n_1142, n_1089);
  nand g3374 (n_1158, n_3097, n_3098, n_3099);
  xor g3375 (n_3100, n_1145, n_1146);
  xor g3376 (n_1149, n_3100, n_1147);
  nand g3377 (n_3101, n_1145, n_1146);
  nand g3378 (n_3102, n_1147, n_1146);
  nand g3379 (n_3103, n_1145, n_1147);
  nand g3380 (n_1161, n_3101, n_3102, n_3103);
  xor g3381 (n_3104, n_1148, n_1149);
  xor g3382 (n_165, n_3104, n_1150);
  nand g3383 (n_3105, n_1148, n_1149);
  nand g3384 (n_3106, n_1150, n_1149);
  nand g3385 (n_3107, n_1148, n_1150);
  nand g3386 (n_79, n_3105, n_3106, n_3107);
  xor g3389 (n_3108, A[58], A[56]);
  xor g3390 (n_1155, n_3108, A[64]);
  nand g3394 (n_1163, n_3062, n_2946, n_2878);
  nand g3400 (n_1166, n_2886, n_3114, n_3115);
  xor g3401 (n_3116, n_1153, n_1101);
  xor g3402 (n_1159, n_3116, n_1155);
  nand g3403 (n_3117, n_1153, n_1101);
  nand g3404 (n_3118, n_1155, n_1101);
  nand g3405 (n_3119, n_1153, n_1155);
  nand g3406 (n_1168, n_3117, n_3118, n_3119);
  xor g3407 (n_3120, n_1156, n_1157);
  xor g3408 (n_1160, n_3120, n_1158);
  nand g3409 (n_3121, n_1156, n_1157);
  nand g3410 (n_3122, n_1158, n_1157);
  nand g3411 (n_3123, n_1156, n_1158);
  nand g3412 (n_1170, n_3121, n_3122, n_3123);
  xor g3413 (n_3124, n_1159, n_1160);
  xor g3414 (n_164, n_3124, n_1161);
  nand g3415 (n_3125, n_1159, n_1160);
  nand g3416 (n_3126, n_1161, n_1160);
  nand g3417 (n_3127, n_1159, n_1161);
  nand g3418 (n_78, n_3125, n_3126, n_3127);
  xor g3431 (n_3136, A[62], n_1163);
  xor g3432 (n_1167, n_3136, n_1143);
  nand g3433 (n_3137, A[62], n_1163);
  nand g3434 (n_3138, n_1143, n_1163);
  nand g3435 (n_3139, A[62], n_1143);
  nand g3436 (n_1177, n_3137, n_3138, n_3139);
  xor g3437 (n_3140, n_1089, n_1166);
  xor g3438 (n_1169, n_3140, n_1167);
  nand g3439 (n_3141, n_1089, n_1166);
  nand g3440 (n_3142, n_1167, n_1166);
  nand g3441 (n_3143, n_1089, n_1167);
  nand g3442 (n_1179, n_3141, n_3142, n_3143);
  xor g3443 (n_3144, n_1168, n_1169);
  xor g3444 (n_163, n_3144, n_1170);
  nand g3445 (n_3145, n_1168, n_1169);
  nand g3446 (n_3146, n_1170, n_1169);
  nand g3447 (n_3147, n_1168, n_1170);
  nand g3448 (n_77, n_3145, n_3146, n_3147);
  nand g3461 (n_3155, A[60], n_1153);
  nand g3462 (n_1184, n_3114, n_3154, n_3155);
  xor g3463 (n_3156, n_1101, n_1155);
  xor g3464 (n_1178, n_3156, n_1176);
  nand g3466 (n_3158, n_1176, n_1155);
  nand g3467 (n_3159, n_1101, n_1176);
  nand g3468 (n_1186, n_3118, n_3158, n_3159);
  xor g3469 (n_3160, n_1177, n_1178);
  xor g3470 (n_162, n_3160, n_1179);
  nand g3471 (n_3161, n_1177, n_1178);
  nand g3472 (n_3162, n_1179, n_1178);
  nand g3473 (n_3163, n_1177, n_1179);
  nand g3474 (n_161, n_3161, n_3162, n_3163);
  xor g3482 (n_1183, n_3088, A[62]);
  nand g3484 (n_3170, A[62], A[61]);
  nand g3485 (n_3171, A[57], A[62]);
  nand g3486 (n_1191, n_3038, n_3170, n_3171);
  xor g3487 (n_3172, n_1163, n_1089);
  xor g3488 (n_1185, n_3172, n_1183);
  nand g3489 (n_3173, n_1163, n_1089);
  nand g3490 (n_3174, n_1183, n_1089);
  nand g3491 (n_3175, n_1163, n_1183);
  nand g3492 (n_1193, n_3173, n_3174, n_3175);
  xor g3493 (n_3176, n_1184, n_1185);
  xor g3494 (n_76, n_3176, n_1186);
  nand g3495 (n_3177, n_1184, n_1185);
  nand g3496 (n_3178, n_1186, n_1185);
  nand g3497 (n_3179, n_1184, n_1186);
  nand g3498 (n_160, n_3177, n_3178, n_3179);
  xor g3502 (n_1190, n_3060, A[60]);
  nand g3505 (n_3183, A[58], A[60]);
  nand g3506 (n_1195, n_3007, n_2949, n_3183);
  xor g3508 (n_1192, n_3068, n_1190);
  nand g3510 (n_3186, n_1190, n_1101);
  nand g3512 (n_1198, n_3014, n_3186, n_3187);
  xor g3513 (n_3188, n_1191, n_1192);
  xor g3514 (n_75, n_3188, n_1193);
  nand g3515 (n_3189, n_1191, n_1192);
  nand g3516 (n_3190, n_1193, n_1192);
  nand g3517 (n_3191, n_1191, n_1193);
  nand g3518 (n_159, n_3189, n_3190, n_3191);
  xor g3525 (n_3196, A[61], A[64]);
  xor g3526 (n_1197, n_3196, n_1195);
  nand g3527 (n_3197, A[61], A[64]);
  nand g3528 (n_3198, n_1195, A[64]);
  nand g3529 (n_3199, A[61], n_1195);
  nand g3530 (n_1203, n_3197, n_3198, n_3199);
  xor g3531 (n_3200, n_1089, n_1197);
  xor g3532 (n_74, n_3200, n_1198);
  nand g3533 (n_3201, n_1089, n_1197);
  nand g3534 (n_3202, n_1198, n_1197);
  nand g3535 (n_3203, n_1089, n_1198);
  nand g3536 (n_158, n_3201, n_3202, n_3203);
  nand g3544 (n_1206, n_2949, n_3206, n_3207);
  xor g3545 (n_3208, n_1101, n_1202);
  xor g3546 (n_73, n_3208, n_1203);
  nand g3547 (n_3209, n_1101, n_1202);
  nand g3548 (n_3210, n_1203, n_1202);
  nand g3549 (n_3211, n_1101, n_1203);
  nand g3550 (n_157, n_3209, n_3210, n_3211);
  xor g3552 (n_1205, n_2972, A[61]);
  nand g3556 (n_1209, n_2973, n_2917, n_2981);
  xor g3557 (n_3216, A[64], n_1205);
  xor g3558 (n_72, n_3216, n_1206);
  nand g3559 (n_3217, A[64], n_1205);
  nand g3560 (n_3218, n_1206, n_1205);
  nand g3561 (n_3219, A[64], n_1206);
  nand g3562 (n_156, n_3217, n_3218, n_3219);
  xor g3566 (n_71, n_3220, n_1209);
  nand g3569 (n_3223, A[64], n_1209);
  nand g3570 (n_155, n_3221, n_3222, n_3223);
  xor g3572 (n_70, n_2972, A[62]);
  nand g3574 (n_3226, A[62], A[63]);
  nand g3576 (n_154, n_2973, n_3226, n_3227);
  nand g25 (n_3249, n_1215, n_3246, n_3247);
  xor g26 (n_3248, A[1], A[3]);
  nand g28 (n_3250, A[2], n_232);
  nand g29 (n_3251, A[2], n_3249);
  nand g30 (n_3252, n_232, n_3249);
  nand g31 (n_3254, n_3250, n_3251, n_3252);
  xor g33 (Z[4], n_3249, n_328);
  nand g34 (n_3255, n_146, n_231);
  nand g35 (n_3256, n_146, n_3254);
  nand g36 (n_3257, n_231, n_3254);
  nand g37 (n_3259, n_3255, n_3256, n_3257);
  xor g38 (n_3258, n_146, n_231);
  xor g39 (Z[5], n_3254, n_3258);
  nand g40 (n_3260, n_145, n_230);
  nand g41 (n_3261, n_145, n_3259);
  nand g42 (n_3262, n_230, n_3259);
  nand g43 (n_3264, n_3260, n_3261, n_3262);
  xor g44 (n_3263, n_145, n_230);
  xor g45 (Z[6], n_3259, n_3263);
  nand g46 (n_3265, n_144, n_229);
  nand g47 (n_3266, n_144, n_3264);
  nand g48 (n_3267, n_229, n_3264);
  nand g49 (n_3269, n_3265, n_3266, n_3267);
  xor g50 (n_3268, n_144, n_229);
  xor g51 (Z[7], n_3264, n_3268);
  nand g52 (n_3270, n_143, n_228);
  nand g53 (n_3271, n_143, n_3269);
  nand g54 (n_3272, n_228, n_3269);
  nand g55 (n_3274, n_3270, n_3271, n_3272);
  xor g56 (n_3273, n_143, n_228);
  xor g57 (Z[8], n_3269, n_3273);
  nand g58 (n_3275, n_142, n_227);
  nand g59 (n_3276, n_142, n_3274);
  nand g60 (n_3277, n_227, n_3274);
  nand g61 (n_3279, n_3275, n_3276, n_3277);
  xor g62 (n_3278, n_142, n_227);
  xor g63 (Z[9], n_3274, n_3278);
  nand g64 (n_3280, n_141, n_226);
  nand g65 (n_3281, n_141, n_3279);
  nand g66 (n_3282, n_226, n_3279);
  nand g67 (n_3284, n_3280, n_3281, n_3282);
  xor g68 (n_3283, n_141, n_226);
  xor g69 (Z[10], n_3279, n_3283);
  nand g70 (n_3285, n_140, n_225);
  nand g71 (n_3286, n_140, n_3284);
  nand g72 (n_3287, n_225, n_3284);
  nand g73 (n_3289, n_3285, n_3286, n_3287);
  xor g74 (n_3288, n_140, n_225);
  xor g75 (Z[11], n_3284, n_3288);
  nand g76 (n_3290, n_139, n_224);
  nand g77 (n_3291, n_139, n_3289);
  nand g78 (n_3292, n_224, n_3289);
  nand g79 (n_3294, n_3290, n_3291, n_3292);
  xor g80 (n_3293, n_139, n_224);
  xor g81 (Z[12], n_3289, n_3293);
  nand g82 (n_3295, n_138, n_223);
  nand g83 (n_3296, n_138, n_3294);
  nand g84 (n_3297, n_223, n_3294);
  nand g85 (n_3299, n_3295, n_3296, n_3297);
  xor g86 (n_3298, n_138, n_223);
  xor g87 (Z[13], n_3294, n_3298);
  nand g88 (n_3300, n_137, n_222);
  nand g89 (n_3301, n_137, n_3299);
  nand g90 (n_3302, n_222, n_3299);
  nand g91 (n_3304, n_3300, n_3301, n_3302);
  xor g92 (n_3303, n_137, n_222);
  xor g93 (Z[14], n_3299, n_3303);
  nand g94 (n_3305, n_136, n_221);
  nand g95 (n_3306, n_136, n_3304);
  nand g96 (n_3307, n_221, n_3304);
  nand g97 (n_3309, n_3305, n_3306, n_3307);
  xor g98 (n_3308, n_136, n_221);
  xor g99 (Z[15], n_3304, n_3308);
  nand g100 (n_3310, n_135, n_220);
  nand g101 (n_3311, n_135, n_3309);
  nand g102 (n_3312, n_220, n_3309);
  nand g103 (n_3314, n_3310, n_3311, n_3312);
  xor g104 (n_3313, n_135, n_220);
  xor g105 (Z[16], n_3309, n_3313);
  nand g106 (n_3315, n_134, n_219);
  nand g107 (n_3316, n_134, n_3314);
  nand g108 (n_3317, n_219, n_3314);
  nand g109 (n_3319, n_3315, n_3316, n_3317);
  xor g110 (n_3318, n_134, n_219);
  xor g111 (Z[17], n_3314, n_3318);
  nand g112 (n_3320, n_133, n_218);
  nand g113 (n_3321, n_133, n_3319);
  nand g114 (n_3322, n_218, n_3319);
  nand g115 (n_3324, n_3320, n_3321, n_3322);
  xor g116 (n_3323, n_133, n_218);
  xor g117 (Z[18], n_3319, n_3323);
  nand g118 (n_3325, n_132, n_217);
  nand g119 (n_3326, n_132, n_3324);
  nand g120 (n_3327, n_217, n_3324);
  nand g121 (n_3329, n_3325, n_3326, n_3327);
  xor g122 (n_3328, n_132, n_217);
  xor g123 (Z[19], n_3324, n_3328);
  nand g124 (n_3330, n_131, n_216);
  nand g125 (n_3331, n_131, n_3329);
  nand g126 (n_3332, n_216, n_3329);
  nand g127 (n_3334, n_3330, n_3331, n_3332);
  xor g128 (n_3333, n_131, n_216);
  xor g129 (Z[20], n_3329, n_3333);
  nand g130 (n_3335, n_130, n_215);
  nand g131 (n_3336, n_130, n_3334);
  nand g132 (n_3337, n_215, n_3334);
  nand g133 (n_3339, n_3335, n_3336, n_3337);
  xor g134 (n_3338, n_130, n_215);
  xor g135 (Z[21], n_3334, n_3338);
  nand g136 (n_3340, n_129, n_214);
  nand g137 (n_3341, n_129, n_3339);
  nand g138 (n_3342, n_214, n_3339);
  nand g139 (n_3344, n_3340, n_3341, n_3342);
  xor g140 (n_3343, n_129, n_214);
  xor g141 (Z[22], n_3339, n_3343);
  nand g142 (n_3345, n_128, n_213);
  nand g143 (n_3346, n_128, n_3344);
  nand g144 (n_3347, n_213, n_3344);
  nand g145 (n_3349, n_3345, n_3346, n_3347);
  xor g146 (n_3348, n_128, n_213);
  xor g147 (Z[23], n_3344, n_3348);
  nand g148 (n_3350, n_127, n_212);
  nand g149 (n_3351, n_127, n_3349);
  nand g150 (n_3352, n_212, n_3349);
  nand g151 (n_3354, n_3350, n_3351, n_3352);
  xor g152 (n_3353, n_127, n_212);
  xor g153 (Z[24], n_3349, n_3353);
  nand g154 (n_3355, n_126, n_211);
  nand g155 (n_3356, n_126, n_3354);
  nand g156 (n_3357, n_211, n_3354);
  nand g157 (n_3359, n_3355, n_3356, n_3357);
  xor g158 (n_3358, n_126, n_211);
  xor g159 (Z[25], n_3354, n_3358);
  nand g160 (n_3360, n_125, n_210);
  nand g161 (n_3361, n_125, n_3359);
  nand g162 (n_3362, n_210, n_3359);
  nand g163 (n_3364, n_3360, n_3361, n_3362);
  xor g164 (n_3363, n_125, n_210);
  xor g165 (Z[26], n_3359, n_3363);
  nand g166 (n_3365, n_124, n_209);
  nand g167 (n_3366, n_124, n_3364);
  nand g168 (n_3367, n_209, n_3364);
  nand g169 (n_3369, n_3365, n_3366, n_3367);
  xor g170 (n_3368, n_124, n_209);
  xor g171 (Z[27], n_3364, n_3368);
  nand g172 (n_3370, n_123, n_208);
  nand g173 (n_3371, n_123, n_3369);
  nand g174 (n_3372, n_208, n_3369);
  nand g175 (n_3374, n_3370, n_3371, n_3372);
  xor g176 (n_3373, n_123, n_208);
  xor g177 (Z[28], n_3369, n_3373);
  nand g178 (n_3375, n_122, n_207);
  nand g179 (n_3376, n_122, n_3374);
  nand g180 (n_3377, n_207, n_3374);
  nand g181 (n_3379, n_3375, n_3376, n_3377);
  xor g182 (n_3378, n_122, n_207);
  xor g183 (Z[29], n_3374, n_3378);
  nand g184 (n_3380, n_121, n_206);
  nand g185 (n_3381, n_121, n_3379);
  nand g186 (n_3382, n_206, n_3379);
  nand g187 (n_3384, n_3380, n_3381, n_3382);
  xor g188 (n_3383, n_121, n_206);
  xor g189 (Z[30], n_3379, n_3383);
  nand g190 (n_3385, n_120, n_205);
  nand g191 (n_3386, n_120, n_3384);
  nand g192 (n_3387, n_205, n_3384);
  nand g193 (n_3389, n_3385, n_3386, n_3387);
  xor g194 (n_3388, n_120, n_205);
  xor g195 (Z[31], n_3384, n_3388);
  nand g196 (n_3390, n_119, n_204);
  nand g197 (n_3391, n_119, n_3389);
  nand g198 (n_3392, n_204, n_3389);
  nand g199 (n_3394, n_3390, n_3391, n_3392);
  xor g200 (n_3393, n_119, n_204);
  xor g201 (Z[32], n_3389, n_3393);
  nand g202 (n_3395, n_118, n_203);
  nand g203 (n_3396, n_118, n_3394);
  nand g204 (n_3397, n_203, n_3394);
  nand g205 (n_3399, n_3395, n_3396, n_3397);
  xor g206 (n_3398, n_118, n_203);
  xor g207 (Z[33], n_3394, n_3398);
  nand g208 (n_3400, n_117, n_202);
  nand g209 (n_3401, n_117, n_3399);
  nand g210 (n_3402, n_202, n_3399);
  nand g211 (n_3404, n_3400, n_3401, n_3402);
  xor g212 (n_3403, n_117, n_202);
  xor g213 (Z[34], n_3399, n_3403);
  nand g214 (n_3405, n_116, n_201);
  nand g215 (n_3406, n_116, n_3404);
  nand g216 (n_3407, n_201, n_3404);
  nand g217 (n_3409, n_3405, n_3406, n_3407);
  xor g218 (n_3408, n_116, n_201);
  xor g219 (Z[35], n_3404, n_3408);
  nand g220 (n_3410, n_115, n_200);
  nand g221 (n_3411, n_115, n_3409);
  nand g222 (n_3412, n_200, n_3409);
  nand g223 (n_3414, n_3410, n_3411, n_3412);
  xor g224 (n_3413, n_115, n_200);
  xor g225 (Z[36], n_3409, n_3413);
  nand g226 (n_3415, n_114, n_199);
  nand g227 (n_3416, n_114, n_3414);
  nand g228 (n_3417, n_199, n_3414);
  nand g229 (n_3419, n_3415, n_3416, n_3417);
  xor g230 (n_3418, n_114, n_199);
  xor g231 (Z[37], n_3414, n_3418);
  nand g232 (n_3420, n_113, n_198);
  nand g233 (n_3421, n_113, n_3419);
  nand g234 (n_3422, n_198, n_3419);
  nand g235 (n_3424, n_3420, n_3421, n_3422);
  xor g236 (n_3423, n_113, n_198);
  xor g237 (Z[38], n_3419, n_3423);
  nand g238 (n_3425, n_112, n_197);
  nand g239 (n_3426, n_112, n_3424);
  nand g240 (n_3427, n_197, n_3424);
  nand g241 (n_3429, n_3425, n_3426, n_3427);
  xor g242 (n_3428, n_112, n_197);
  xor g243 (Z[39], n_3424, n_3428);
  nand g244 (n_3430, n_111, n_196);
  nand g245 (n_3431, n_111, n_3429);
  nand g246 (n_3432, n_196, n_3429);
  nand g247 (n_3434, n_3430, n_3431, n_3432);
  xor g248 (n_3433, n_111, n_196);
  xor g249 (Z[40], n_3429, n_3433);
  nand g250 (n_3435, n_110, n_195);
  nand g251 (n_3436, n_110, n_3434);
  nand g252 (n_3437, n_195, n_3434);
  nand g253 (n_3439, n_3435, n_3436, n_3437);
  xor g254 (n_3438, n_110, n_195);
  xor g255 (Z[41], n_3434, n_3438);
  nand g256 (n_3440, n_109, n_194);
  nand g257 (n_3441, n_109, n_3439);
  nand g258 (n_3442, n_194, n_3439);
  nand g259 (n_3444, n_3440, n_3441, n_3442);
  xor g260 (n_3443, n_109, n_194);
  xor g261 (Z[42], n_3439, n_3443);
  nand g262 (n_3445, n_108, n_193);
  nand g263 (n_3446, n_108, n_3444);
  nand g264 (n_3447, n_193, n_3444);
  nand g265 (n_3449, n_3445, n_3446, n_3447);
  xor g266 (n_3448, n_108, n_193);
  xor g267 (Z[43], n_3444, n_3448);
  nand g268 (n_3450, n_107, n_192);
  nand g269 (n_3451, n_107, n_3449);
  nand g270 (n_3452, n_192, n_3449);
  nand g271 (n_3454, n_3450, n_3451, n_3452);
  xor g272 (n_3453, n_107, n_192);
  xor g273 (Z[44], n_3449, n_3453);
  nand g274 (n_3455, n_106, n_191);
  nand g275 (n_3456, n_106, n_3454);
  nand g276 (n_3457, n_191, n_3454);
  nand g277 (n_3459, n_3455, n_3456, n_3457);
  xor g278 (n_3458, n_106, n_191);
  xor g279 (Z[45], n_3454, n_3458);
  nand g280 (n_3460, n_105, n_190);
  nand g281 (n_3461, n_105, n_3459);
  nand g282 (n_3462, n_190, n_3459);
  nand g283 (n_3464, n_3460, n_3461, n_3462);
  xor g284 (n_3463, n_105, n_190);
  xor g285 (Z[46], n_3459, n_3463);
  nand g286 (n_3465, n_104, n_189);
  nand g287 (n_3466, n_104, n_3464);
  nand g288 (n_3467, n_189, n_3464);
  nand g289 (n_3469, n_3465, n_3466, n_3467);
  xor g290 (n_3468, n_104, n_189);
  xor g291 (Z[47], n_3464, n_3468);
  nand g292 (n_3470, n_103, n_188);
  nand g293 (n_3471, n_103, n_3469);
  nand g294 (n_3472, n_188, n_3469);
  nand g295 (n_3474, n_3470, n_3471, n_3472);
  xor g296 (n_3473, n_103, n_188);
  xor g297 (Z[48], n_3469, n_3473);
  nand g298 (n_3475, n_102, n_187);
  nand g299 (n_3476, n_102, n_3474);
  nand g300 (n_3477, n_187, n_3474);
  nand g301 (n_3479, n_3475, n_3476, n_3477);
  xor g302 (n_3478, n_102, n_187);
  xor g303 (Z[49], n_3474, n_3478);
  nand g304 (n_3480, n_101, n_186);
  nand g305 (n_3481, n_101, n_3479);
  nand g306 (n_3482, n_186, n_3479);
  nand g307 (n_3484, n_3480, n_3481, n_3482);
  xor g308 (n_3483, n_101, n_186);
  xor g309 (Z[50], n_3479, n_3483);
  nand g310 (n_3485, n_100, n_185);
  nand g311 (n_3486, n_100, n_3484);
  nand g312 (n_3487, n_185, n_3484);
  nand g313 (n_3489, n_3485, n_3486, n_3487);
  xor g314 (n_3488, n_100, n_185);
  xor g315 (Z[51], n_3484, n_3488);
  nand g316 (n_3490, n_99, n_184);
  nand g317 (n_3491, n_99, n_3489);
  nand g318 (n_3492, n_184, n_3489);
  nand g319 (n_3494, n_3490, n_3491, n_3492);
  xor g320 (n_3493, n_99, n_184);
  xor g321 (Z[52], n_3489, n_3493);
  nand g322 (n_3495, n_98, n_183);
  nand g323 (n_3496, n_98, n_3494);
  nand g324 (n_3497, n_183, n_3494);
  nand g325 (n_3499, n_3495, n_3496, n_3497);
  xor g326 (n_3498, n_98, n_183);
  xor g327 (Z[53], n_3494, n_3498);
  nand g328 (n_3500, n_97, n_182);
  nand g329 (n_3501, n_97, n_3499);
  nand g330 (n_3502, n_182, n_3499);
  nand g331 (n_3504, n_3500, n_3501, n_3502);
  xor g332 (n_3503, n_97, n_182);
  xor g333 (Z[54], n_3499, n_3503);
  nand g334 (n_3505, n_96, n_181);
  nand g335 (n_3506, n_96, n_3504);
  nand g336 (n_3507, n_181, n_3504);
  nand g337 (n_3509, n_3505, n_3506, n_3507);
  xor g338 (n_3508, n_96, n_181);
  xor g339 (Z[55], n_3504, n_3508);
  nand g340 (n_3510, n_95, n_180);
  nand g341 (n_3511, n_95, n_3509);
  nand g342 (n_3512, n_180, n_3509);
  nand g343 (n_3514, n_3510, n_3511, n_3512);
  xor g344 (n_3513, n_95, n_180);
  xor g345 (Z[56], n_3509, n_3513);
  nand g346 (n_3515, n_94, n_179);
  nand g347 (n_3516, n_94, n_3514);
  nand g348 (n_3517, n_179, n_3514);
  nand g349 (n_3519, n_3515, n_3516, n_3517);
  xor g350 (n_3518, n_94, n_179);
  xor g351 (Z[57], n_3514, n_3518);
  nand g352 (n_3520, n_93, n_178);
  nand g353 (n_3521, n_93, n_3519);
  nand g354 (n_3522, n_178, n_3519);
  nand g355 (n_3524, n_3520, n_3521, n_3522);
  xor g356 (n_3523, n_93, n_178);
  xor g357 (Z[58], n_3519, n_3523);
  nand g358 (n_3525, n_92, n_177);
  nand g359 (n_3526, n_92, n_3524);
  nand g360 (n_3527, n_177, n_3524);
  nand g361 (n_3529, n_3525, n_3526, n_3527);
  xor g362 (n_3528, n_92, n_177);
  xor g363 (Z[59], n_3524, n_3528);
  nand g364 (n_3530, n_91, n_176);
  nand g365 (n_3531, n_91, n_3529);
  nand g366 (n_3532, n_176, n_3529);
  nand g367 (n_3534, n_3530, n_3531, n_3532);
  xor g368 (n_3533, n_91, n_176);
  xor g369 (Z[60], n_3529, n_3533);
  nand g370 (n_3535, n_90, n_175);
  nand g371 (n_3536, n_90, n_3534);
  nand g372 (n_3537, n_175, n_3534);
  nand g373 (n_3539, n_3535, n_3536, n_3537);
  xor g374 (n_3538, n_90, n_175);
  xor g375 (Z[61], n_3534, n_3538);
  nand g376 (n_3540, n_89, n_174);
  nand g377 (n_3541, n_89, n_3539);
  nand g378 (n_3542, n_174, n_3539);
  nand g379 (n_3544, n_3540, n_3541, n_3542);
  xor g380 (n_3543, n_89, n_174);
  xor g381 (Z[62], n_3539, n_3543);
  nand g382 (n_3545, n_88, n_173);
  nand g383 (n_3546, n_88, n_3544);
  nand g384 (n_3547, n_173, n_3544);
  nand g385 (n_3549, n_3545, n_3546, n_3547);
  xor g386 (n_3548, n_88, n_173);
  xor g387 (Z[63], n_3544, n_3548);
  nand g388 (n_3550, n_87, n_172);
  nand g389 (n_3551, n_87, n_3549);
  nand g390 (n_3552, n_172, n_3549);
  nand g391 (n_3554, n_3550, n_3551, n_3552);
  xor g392 (n_3553, n_87, n_172);
  xor g393 (Z[64], n_3549, n_3553);
  nand g394 (n_3555, n_86, n_171);
  nand g395 (n_3556, n_86, n_3554);
  nand g396 (n_3557, n_171, n_3554);
  nand g397 (n_3559, n_3555, n_3556, n_3557);
  xor g398 (n_3558, n_86, n_171);
  xor g399 (Z[65], n_3554, n_3558);
  nand g400 (n_3560, n_85, n_170);
  nand g401 (n_3561, n_85, n_3559);
  nand g402 (n_3562, n_170, n_3559);
  nand g403 (n_3564, n_3560, n_3561, n_3562);
  xor g404 (n_3563, n_85, n_170);
  xor g405 (Z[66], n_3559, n_3563);
  nand g406 (n_3565, n_84, n_169);
  nand g407 (n_3566, n_84, n_3564);
  nand g408 (n_3567, n_169, n_3564);
  nand g409 (n_3569, n_3565, n_3566, n_3567);
  xor g410 (n_3568, n_84, n_169);
  xor g411 (Z[67], n_3564, n_3568);
  nand g412 (n_3570, n_83, n_168);
  nand g413 (n_3571, n_83, n_3569);
  nand g414 (n_3572, n_168, n_3569);
  nand g415 (n_3574, n_3570, n_3571, n_3572);
  xor g416 (n_3573, n_83, n_168);
  xor g417 (Z[68], n_3569, n_3573);
  nand g418 (n_3575, n_82, n_167);
  nand g419 (n_3576, n_82, n_3574);
  nand g420 (n_3577, n_167, n_3574);
  nand g421 (n_3579, n_3575, n_3576, n_3577);
  xor g422 (n_3578, n_82, n_167);
  xor g423 (Z[69], n_3574, n_3578);
  nand g424 (n_3580, n_81, n_166);
  nand g425 (n_3581, n_81, n_3579);
  nand g426 (n_3582, n_166, n_3579);
  nand g427 (n_3584, n_3580, n_3581, n_3582);
  xor g428 (n_3583, n_81, n_166);
  xor g429 (Z[70], n_3579, n_3583);
  nand g430 (n_3585, n_80, n_165);
  nand g431 (n_3586, n_80, n_3584);
  nand g432 (n_3587, n_165, n_3584);
  nand g433 (n_3589, n_3585, n_3586, n_3587);
  xor g434 (n_3588, n_80, n_165);
  xor g435 (Z[71], n_3584, n_3588);
  nand g436 (n_3590, n_79, n_164);
  nand g437 (n_3591, n_79, n_3589);
  nand g438 (n_3592, n_164, n_3589);
  nand g439 (n_3594, n_3590, n_3591, n_3592);
  xor g440 (n_3593, n_79, n_164);
  xor g441 (Z[72], n_3589, n_3593);
  nand g442 (n_3595, n_78, n_163);
  nand g443 (n_3596, n_78, n_3594);
  nand g444 (n_3597, n_163, n_3594);
  nand g445 (n_3599, n_3595, n_3596, n_3597);
  xor g446 (n_3598, n_78, n_163);
  xor g447 (Z[73], n_3594, n_3598);
  nand g448 (n_3600, n_77, n_162);
  nand g449 (n_3601, n_77, n_3599);
  nand g450 (n_3602, n_162, n_3599);
  nand g451 (n_3604, n_3600, n_3601, n_3602);
  xor g452 (n_3603, n_77, n_162);
  xor g453 (Z[74], n_3599, n_3603);
  nand g454 (n_3605, n_76, n_161);
  nand g455 (n_3606, n_76, n_3604);
  nand g456 (n_3607, n_161, n_3604);
  nand g457 (n_3609, n_3605, n_3606, n_3607);
  xor g458 (n_3608, n_76, n_161);
  xor g459 (Z[75], n_3604, n_3608);
  nand g460 (n_3610, n_75, n_160);
  nand g461 (n_3611, n_75, n_3609);
  nand g462 (n_3612, n_160, n_3609);
  nand g463 (n_3614, n_3610, n_3611, n_3612);
  xor g464 (n_3613, n_75, n_160);
  xor g465 (Z[76], n_3609, n_3613);
  nand g466 (n_3615, n_74, n_159);
  nand g467 (n_3616, n_74, n_3614);
  nand g468 (n_3617, n_159, n_3614);
  nand g469 (n_3619, n_3615, n_3616, n_3617);
  xor g470 (n_3618, n_74, n_159);
  xor g471 (Z[77], n_3614, n_3618);
  nand g472 (n_3620, n_73, n_158);
  nand g473 (n_3621, n_73, n_3619);
  nand g474 (n_3622, n_158, n_3619);
  nand g475 (n_3624, n_3620, n_3621, n_3622);
  xor g476 (n_3623, n_73, n_158);
  xor g477 (Z[78], n_3619, n_3623);
  nand g478 (n_3625, n_72, n_157);
  nand g479 (n_3626, n_72, n_3624);
  nand g480 (n_3627, n_157, n_3624);
  nand g481 (n_3629, n_3625, n_3626, n_3627);
  xor g482 (n_3628, n_72, n_157);
  xor g483 (Z[79], n_3624, n_3628);
  nand g484 (n_3630, n_71, n_156);
  nand g485 (n_3631, n_71, n_3629);
  nand g486 (n_3632, n_156, n_3629);
  nand g487 (n_3634, n_3630, n_3631, n_3632);
  xor g488 (n_3633, n_71, n_156);
  xor g489 (Z[80], n_3629, n_3633);
  nand g490 (n_3635, n_70, n_155);
  nand g491 (n_3636, n_70, n_3634);
  nand g492 (n_3637, n_155, n_3634);
  nand g493 (n_3639, n_3635, n_3636, n_3637);
  xor g494 (n_3638, n_70, n_155);
  xor g495 (Z[81], n_3634, n_3638);
  nand g498 (n_3642, n_154, n_3639);
  nand g499 (n_3644, n_3640, n_3641, n_3642);
  xor g501 (Z[82], n_3639, n_3643);
  nand g504 (n_3647, A[64], n_3644);
  nand g505 (n_3649, n_3645, n_3646, n_3647);
  xor g507 (Z[83], n_3644, n_3648);
  or g3594 (n_330, wc, wc0, n_146);
  not gc0 (wc0, n_1217);
  not gc (wc, n_1230);
  or g3595 (n_339, wc1, n_324, n_146);
  not gc1 (wc1, n_1250);
  or g3596 (n_352, wc2, wc3, n_146);
  not gc3 (wc3, n_1277);
  not gc2 (wc2, n_1278);
  or g3597 (n_369, wc4, n_351, wc5);
  not gc5 (wc5, n_1250);
  not gc4 (wc4, n_1315);
  or g3598 (n_390, wc6, wc7, n_338);
  not gc7 (wc7, n_1278);
  not gc6 (wc6, n_1315);
  or g3599 (n_394, wc8, wc9, n_324);
  not gc9 (wc9, n_1230);
  not gc8 (wc8, n_1363);
  or g3600 (n_416, wc10, wc11, n_146);
  not gc11 (wc11, n_1315);
  not gc10 (wc10, n_1409);
  or g3601 (n_415, wc12, n_368, n_329);
  not gc12 (wc12, n_1415);
  or g3602 (n_443, wc13, wc14, n_324);
  not gc14 (wc14, n_1474);
  not gc13 (wc13, n_1475);
  or g3603 (n_147, wc15, wc16, n_338);
  not gc16 (wc16, n_1478);
  not gc15 (wc15, n_1479);
  or g3604 (n_494, wc17, wc18, n_338);
  not gc18 (wc18, n_1602);
  not gc17 (wc17, n_1603);
  or g3605 (n_234, wc19, wc20, n_338);
  not gc20 (wc20, n_1542);
  not gc19 (wc19, n_1666);
  or g3606 (n_521, wc21, wc22, n_389);
  not gc22 (wc22, n_1535);
  not gc21 (wc21, n_1671);
  or g3607 (n_549, wc23, wc24, n_414);
  not gc24 (wc24, n_1599);
  not gc23 (wc23, n_1735);
  xnor g3608 (n_2972, A[65], A[63]);
  or g3609 (n_2973, wc25, A[65]);
  not gc25 (wc25, A[63]);
  or g3610 (n_2975, wc26, A[65]);
  not gc26 (wc26, A[59]);
  xnor g3611 (n_3012, A[64], A[52]);
  or g3612 (n_3013, wc27, A[64]);
  not gc27 (wc27, A[52]);
  xnor g3613 (n_1156, n_3064, A[62]);
  or g3614 (n_3114, wc28, A[62]);
  not gc28 (wc28, A[60]);
  or g3615 (n_3115, wc29, A[62]);
  not gc29 (wc29, A[54]);
  xnor g3617 (n_1202, n_2948, A[64]);
  or g3618 (n_3206, wc30, A[64]);
  not gc30 (wc30, A[60]);
  or g3619 (n_3207, wc31, A[64]);
  not gc31 (wc31, A[62]);
  or g3620 (n_2981, wc32, A[65]);
  not gc32 (wc32, A[61]);
  xnor g3621 (n_3220, A[64], A[62]);
  or g3622 (n_3221, A[62], wc33);
  not gc33 (wc33, A[64]);
  or g3623 (n_3227, wc34, A[65]);
  not gc34 (wc34, A[62]);
  or g3624 (n_3645, wc35, A[65]);
  not gc35 (wc35, A[64]);
  xnor g3625 (n_3648, A[65], A[64]);
  or g3626 (n_3071, A[64], wc36);
  not gc36 (wc36, n_1130);
  xnor g3627 (n_1176, n_2948, n_1153);
  or g3628 (n_3154, A[62], wc37);
  not gc37 (wc37, n_1153);
  or g3629 (n_3187, A[64], wc38);
  not gc38 (wc38, n_1190);
  xnor g3631 (n_2980, A[65], A[61]);
  or g3632 (n_2983, wc39, A[65]);
  not gc39 (wc39, A[55]);
  or g3633 (n_3014, A[64], wc40);
  not gc40 (wc40, n_1101);
  xnor g3634 (n_3068, n_1101, A[64]);
  or g3635 (n_3222, A[62], wc41);
  not gc41 (wc41, n_1209);
  or g3636 (n_3640, A[64], wc42);
  not gc42 (wc42, n_154);
  xnor g3637 (n_3643, n_154, A[64]);
  xnor g3638 (n_1075, n_3648, A[56]);
  or g3640 (n_3246, wc43, n_1217);
  not gc43 (wc43, A[1]);
  or g3641 (n_3247, wc44, n_1217);
  not gc44 (wc44, A[3]);
  xnor g3642 (Z[3], n_1217, n_3248);
  or g3643 (n_3641, A[64], wc45);
  not gc45 (wc45, n_3639);
  or g3644 (n_3646, A[65], wc46);
  not gc46 (wc46, n_3644);
  not g3645 (Z[84], n_3649);
endmodule

module mult_signed_const_15762_GENERIC(A, Z);
  input [65:0] A;
  output [84:0] Z;
  wire [65:0] A;
  wire [84:0] Z;
  mult_signed_const_15762_GENERIC_REAL g1(.A ({A[65:2], A[0], A[0]}),
       .Z (Z));
endmodule

module mult_signed_const_16293_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [66:0] A;
  output [85:0] Z;
  wire [66:0] A;
  wire [85:0] Z;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78;
  wire n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_454, n_455, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538;
  wire n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562;
  wire n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578;
  wire n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586;
  wire n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594;
  wire n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602;
  wire n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610;
  wire n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618;
  wire n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626;
  wire n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634;
  wire n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642;
  wire n_643, n_644, n_645, n_646, n_647, n_648, n_649, n_650;
  wire n_651, n_652, n_653, n_654, n_655, n_656, n_657, n_658;
  wire n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666;
  wire n_667, n_668, n_669, n_670, n_671, n_672, n_673, n_674;
  wire n_675, n_676, n_677, n_678, n_679, n_680, n_681, n_682;
  wire n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690;
  wire n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698;
  wire n_699, n_700, n_701, n_702, n_703, n_704, n_705, n_706;
  wire n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714;
  wire n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722;
  wire n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730;
  wire n_731, n_732, n_733, n_734, n_735, n_736, n_737, n_738;
  wire n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746;
  wire n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754;
  wire n_755, n_756, n_757, n_758, n_759, n_760, n_761, n_762;
  wire n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770;
  wire n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778;
  wire n_779, n_780, n_781, n_782, n_783, n_784, n_785, n_786;
  wire n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794;
  wire n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802;
  wire n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810;
  wire n_811, n_812, n_813, n_814, n_815, n_816, n_817, n_818;
  wire n_819, n_820, n_821, n_822, n_823, n_824, n_825, n_826;
  wire n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834;
  wire n_835, n_836, n_837, n_838, n_839, n_840, n_841, n_842;
  wire n_843, n_844, n_845, n_846, n_847, n_848, n_849, n_850;
  wire n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858;
  wire n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866;
  wire n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874;
  wire n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882;
  wire n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890;
  wire n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898;
  wire n_899, n_900, n_901, n_902, n_903, n_904, n_905, n_906;
  wire n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914;
  wire n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922;
  wire n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_930;
  wire n_931, n_932, n_933, n_934, n_935, n_936, n_937, n_938;
  wire n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946;
  wire n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954;
  wire n_955, n_956, n_957, n_958, n_959, n_960, n_961, n_962;
  wire n_963, n_964, n_965, n_966, n_967, n_968, n_969, n_970;
  wire n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978;
  wire n_979, n_980, n_981, n_982, n_983, n_984, n_985, n_986;
  wire n_987, n_988, n_989, n_990, n_991, n_992, n_993, n_994;
  wire n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002;
  wire n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010;
  wire n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018;
  wire n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026;
  wire n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034;
  wire n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042;
  wire n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050;
  wire n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058;
  wire n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066;
  wire n_1067, n_1068, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
  wire n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084;
  wire n_1088, n_1089, n_1090, n_1092, n_1093, n_1094, n_1095, n_1096;
  wire n_1097, n_1098, n_1099, n_1100, n_1101, n_1103, n_1105, n_1107;
  wire n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115;
  wire n_1116, n_1119, n_1120, n_1123, n_1124, n_1125, n_1126, n_1127;
  wire n_1128, n_1129, n_1130, n_1131, n_1134, n_1136, n_1137, n_1138;
  wire n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1148, n_1149;
  wire n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157;
  wire n_1159, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167;
  wire n_1168, n_1171, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178;
  wire n_1179, n_1181, n_1182, n_1184, n_1185, n_1186, n_1187, n_1188;
  wire n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1201, n_1202;
  wire n_1203, n_1204, n_1208, n_1209, n_1210, n_1211, n_1213, n_1214;
  wire n_1215, n_1216, n_1219, n_1220, n_1221, n_1223, n_1224, n_1227;
  wire n_1230, n_1231, n_1232, n_1233, n_1235, n_1236, n_1237, n_1238;
  wire n_1239, n_1241, n_1242, n_1243, n_1244, n_1245, n_1249, n_1250;
  wire n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258;
  wire n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1268;
  wire n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
  wire n_1278, n_1279, n_1280, n_1281, n_1282, n_1286, n_1287, n_1288;
  wire n_1289, n_1290, n_1291, n_1292, n_1293, n_1296, n_1300, n_1301;
  wire n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309;
  wire n_1310, n_1311, n_1312, n_1313, n_1314, n_1318, n_1319, n_1320;
  wire n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328;
  wire n_1329, n_1330, n_1331, n_1332, n_1334, n_1335, n_1337, n_1338;
  wire n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346;
  wire n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354;
  wire n_1357, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366;
  wire n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374;
  wire n_1377, n_1378, n_1379, n_1380, n_1382, n_1383, n_1384, n_1385;
  wire n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393;
  wire n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401;
  wire n_1402, n_1404, n_1406, n_1409, n_1410, n_1411, n_1412, n_1413;
  wire n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421;
  wire n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1429, n_1430;
  wire n_1432, n_1433, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441;
  wire n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449;
  wire n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457;
  wire n_1460, n_1462, n_1463, n_1466, n_1467, n_1468, n_1469, n_1470;
  wire n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478;
  wire n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486;
  wire n_1487, n_1488, n_1489, n_1494, n_1495, n_1496, n_1498, n_1499;
  wire n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507;
  wire n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515;
  wire n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1526, n_1527;
  wire n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537;
  wire n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545;
  wire n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553;
  wire n_1556, n_1557, n_1558, n_1559, n_1560, n_1562, n_1563, n_1564;
  wire n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572;
  wire n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580;
  wire n_1581, n_1582, n_1583, n_1584, n_1585, n_1588, n_1590, n_1591;
  wire n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601;
  wire n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609;
  wire n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617;
  wire n_1620, n_1622, n_1623, n_1626, n_1627, n_1628, n_1629, n_1630;
  wire n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638;
  wire n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646;
  wire n_1647, n_1648, n_1649, n_1652, n_1654, n_1655, n_1658, n_1659;
  wire n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667;
  wire n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675;
  wire n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1684, n_1686;
  wire n_1687, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696;
  wire n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704;
  wire n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712;
  wire n_1713, n_1716, n_1718, n_1719, n_1722, n_1723, n_1724, n_1725;
  wire n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733;
  wire n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741;
  wire n_1742, n_1743, n_1744, n_1745, n_1748, n_1750, n_1751, n_1754;
  wire n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762;
  wire n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770;
  wire n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1780;
  wire n_1782, n_1783, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
  wire n_1808, n_1809, n_1812, n_1814, n_1815, n_1818, n_1819, n_1820;
  wire n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
  wire n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836;
  wire n_1837, n_1838, n_1839, n_1840, n_1841, n_1844, n_1846, n_1847;
  wire n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857;
  wire n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865;
  wire n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873;
  wire n_1876, n_1878, n_1879, n_1882, n_1883, n_1884, n_1885, n_1886;
  wire n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894;
  wire n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902;
  wire n_1903, n_1904, n_1905, n_1908, n_1910, n_1911, n_1914, n_1915;
  wire n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923;
  wire n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931;
  wire n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1940, n_1942;
  wire n_1943, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952;
  wire n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960;
  wire n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968;
  wire n_1969, n_1972, n_1974, n_1975, n_1978, n_1979, n_1980, n_1981;
  wire n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989;
  wire n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997;
  wire n_1998, n_1999, n_2000, n_2001, n_2004, n_2006, n_2007, n_2010;
  wire n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018;
  wire n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026;
  wire n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2036;
  wire n_2038, n_2039, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047;
  wire n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055;
  wire n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063;
  wire n_2064, n_2065, n_2068, n_2070, n_2071, n_2074, n_2075, n_2076;
  wire n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084;
  wire n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092;
  wire n_2093, n_2094, n_2095, n_2096, n_2097, n_2100, n_2102, n_2103;
  wire n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113;
  wire n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121;
  wire n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129;
  wire n_2132, n_2134, n_2135, n_2138, n_2139, n_2140, n_2141, n_2142;
  wire n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150;
  wire n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158;
  wire n_2159, n_2160, n_2161, n_2164, n_2166, n_2167, n_2170, n_2171;
  wire n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179;
  wire n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187;
  wire n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2196, n_2198;
  wire n_2199, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208;
  wire n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216;
  wire n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224;
  wire n_2225, n_2228, n_2230, n_2231, n_2234, n_2235, n_2236, n_2237;
  wire n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245;
  wire n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253;
  wire n_2254, n_2255, n_2256, n_2257, n_2260, n_2262, n_2263, n_2266;
  wire n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274;
  wire n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282;
  wire n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2292;
  wire n_2294, n_2295, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303;
  wire n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311;
  wire n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319;
  wire n_2320, n_2321, n_2324, n_2326, n_2327, n_2330, n_2331, n_2332;
  wire n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340;
  wire n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348;
  wire n_2349, n_2350, n_2351, n_2352, n_2353, n_2356, n_2358, n_2359;
  wire n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369;
  wire n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377;
  wire n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385;
  wire n_2388, n_2390, n_2391, n_2394, n_2395, n_2396, n_2397, n_2398;
  wire n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406;
  wire n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414;
  wire n_2415, n_2416, n_2417, n_2420, n_2422, n_2423, n_2426, n_2427;
  wire n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435;
  wire n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443;
  wire n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2452, n_2454;
  wire n_2455, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464;
  wire n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472;
  wire n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480;
  wire n_2481, n_2484, n_2486, n_2487, n_2490, n_2491, n_2492, n_2493;
  wire n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501;
  wire n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509;
  wire n_2510, n_2511, n_2512, n_2513, n_2516, n_2518, n_2519, n_2522;
  wire n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530;
  wire n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538;
  wire n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2548;
  wire n_2550, n_2551, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559;
  wire n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567;
  wire n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575;
  wire n_2576, n_2577, n_2580, n_2582, n_2583, n_2586, n_2587, n_2588;
  wire n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596;
  wire n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604;
  wire n_2605, n_2606, n_2607, n_2608, n_2609, n_2612, n_2614, n_2615;
  wire n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625;
  wire n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, n_2633;
  wire n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641;
  wire n_2644, n_2646, n_2647, n_2650, n_2651, n_2652, n_2653, n_2654;
  wire n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662;
  wire n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670;
  wire n_2671, n_2672, n_2673, n_2676, n_2678, n_2679, n_2682, n_2683;
  wire n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691;
  wire n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699;
  wire n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2708, n_2710;
  wire n_2711, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720;
  wire n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728;
  wire n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736;
  wire n_2737, n_2740, n_2742, n_2743, n_2746, n_2747, n_2748, n_2749;
  wire n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757;
  wire n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765;
  wire n_2766, n_2767, n_2768, n_2769, n_2772, n_2774, n_2775, n_2778;
  wire n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2786;
  wire n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794;
  wire n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2804;
  wire n_2806, n_2807, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815;
  wire n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823;
  wire n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831;
  wire n_2832, n_2833, n_2836, n_2838, n_2839, n_2842, n_2843, n_2844;
  wire n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852;
  wire n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860;
  wire n_2861, n_2862, n_2863, n_2864, n_2865, n_2868, n_2870, n_2871;
  wire n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881;
  wire n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889;
  wire n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897;
  wire n_2898, n_2899, n_2900, n_2902, n_2905, n_2906, n_2907, n_2908;
  wire n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916;
  wire n_2917, n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924;
  wire n_2925, n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932;
  wire n_2934, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943;
  wire n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951;
  wire n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959;
  wire n_2961, n_2962, n_2963, n_2964, n_2966, n_2969, n_2970, n_2971;
  wire n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979;
  wire n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987;
  wire n_2988, n_2989, n_2992, n_2993, n_2994, n_3002, n_3003, n_3004;
  wire n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012;
  wire n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020;
  wire n_3021, n_3022, n_3023, n_3025, n_3026, n_3028, n_3029, n_3034;
  wire n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042;
  wire n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050;
  wire n_3051, n_3052, n_3053, n_3054, n_3062, n_3063, n_3064, n_3065;
  wire n_3066, n_3067, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074;
  wire n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3090;
  wire n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098;
  wire n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106;
  wire n_3107, n_3108, n_3109, n_3116, n_3117, n_3118, n_3120, n_3121;
  wire n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129;
  wire n_3130, n_3131, n_3132, n_3133, n_3142, n_3144, n_3145, n_3146;
  wire n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154;
  wire n_3155, n_3156, n_3157, n_3160, n_3162, n_3163, n_3164, n_3165;
  wire n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173;
  wire n_3174, n_3175, n_3176, n_3177, n_3184, n_3185, n_3186, n_3187;
  wire n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195;
  wire n_3196, n_3197, n_3202, n_3204, n_3205, n_3206, n_3207, n_3208;
  wire n_3209, n_3210, n_3211, n_3212, n_3213, n_3218, n_3220, n_3221;
  wire n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229;
  wire n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, n_3240;
  wire n_3241, n_3245, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253;
  wire n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, n_3265, n_3266;
  wire n_3267, n_3268, n_3269, n_3272, n_3273, n_3274, n_3277, n_3296;
  wire n_3297, n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305;
  wire n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313;
  wire n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321;
  wire n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329;
  wire n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337;
  wire n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345;
  wire n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353;
  wire n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361;
  wire n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369;
  wire n_3370, n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377;
  wire n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385;
  wire n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393;
  wire n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401;
  wire n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409;
  wire n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417;
  wire n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425;
  wire n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433;
  wire n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441;
  wire n_3442, n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449;
  wire n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, n_3456, n_3457;
  wire n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, n_3465;
  wire n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473;
  wire n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481;
  wire n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489;
  wire n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497;
  wire n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505;
  wire n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513;
  wire n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521;
  wire n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529;
  wire n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537;
  wire n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545;
  wire n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553;
  wire n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561;
  wire n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569;
  wire n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577;
  wire n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585;
  wire n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593;
  wire n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601;
  wire n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609;
  wire n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617;
  wire n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625;
  wire n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633;
  wire n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641;
  wire n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649;
  wire n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657;
  wire n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665;
  wire n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673;
  wire n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681;
  wire n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689;
  wire n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697;
  wire n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g532 (n_235, A[4], A[0]);
  and g2 (n_148, A[4], A[0]);
  xor g533 (n_1230, A[5], A[3]);
  xor g534 (n_234, n_1230, A[1]);
  nand g3 (n_1231, A[5], A[3]);
  nand g535 (n_1232, A[1], A[3]);
  nand g536 (n_1233, A[5], A[1]);
  nand g537 (n_147, n_1231, n_1232, n_1233);
  xor g538 (n_327, A[6], A[4]);
  and g539 (n_328, A[6], A[4]);
  xor g540 (Z[2], A[0], A[2]);
  xor g541 (n_233, Z[2], n_327);
  nand g542 (n_1235, A[0], A[2]);
  nand g4 (n_1236, n_327, A[2]);
  nand g5 (n_1237, A[0], n_327);
  nand g543 (n_146, n_1235, n_1236, n_1237);
  xor g544 (n_1238, A[7], A[5]);
  xor g545 (n_329, n_1238, A[1]);
  nand g546 (n_1239, A[7], A[5]);
  nand g548 (n_1241, A[7], A[1]);
  nand g6 (n_331, n_1239, n_1233, n_1241);
  xor g549 (n_1242, A[3], n_328);
  xor g550 (n_232, n_1242, n_329);
  nand g551 (n_1243, A[3], n_328);
  nand g552 (n_1244, n_329, n_328);
  nand g553 (n_1245, A[3], n_329);
  nand g554 (n_145, n_1243, n_1244, n_1245);
  xor g555 (n_330, A[8], A[6]);
  and g556 (n_333, A[8], A[6]);
  xor g558 (n_332, Z[2], A[4]);
  nand g561 (n_1249, A[2], A[4]);
  xor g563 (n_1250, n_330, n_331);
  xor g564 (n_231, n_1250, n_332);
  nand g565 (n_1251, n_330, n_331);
  nand g566 (n_1252, n_332, n_331);
  nand g567 (n_1253, n_330, n_332);
  nand g568 (n_144, n_1251, n_1252, n_1253);
  xor g569 (n_1254, A[9], A[7]);
  xor g570 (n_335, n_1254, A[3]);
  nand g571 (n_1255, A[9], A[7]);
  nand g572 (n_1256, A[3], A[7]);
  nand g573 (n_1257, A[9], A[3]);
  nand g574 (n_338, n_1255, n_1256, n_1257);
  xor g575 (n_1258, A[1], A[5]);
  xor g576 (n_336, n_1258, n_333);
  nand g578 (n_1260, n_333, A[5]);
  nand g579 (n_1261, A[1], n_333);
  nand g580 (n_340, n_1233, n_1260, n_1261);
  xor g581 (n_1262, n_334, n_335);
  xor g582 (n_230, n_1262, n_336);
  nand g583 (n_1263, n_334, n_335);
  nand g584 (n_1264, n_336, n_335);
  nand g585 (n_1265, n_334, n_336);
  nand g586 (n_143, n_1263, n_1264, n_1265);
  xor g587 (n_337, A[10], A[8]);
  and g588 (n_342, A[10], A[8]);
  xor g589 (n_1266, A[4], A[2]);
  xor g590 (n_339, n_1266, A[6]);
  nand g592 (n_1268, A[6], A[2]);
  xor g595 (n_1270, A[0], n_337);
  xor g596 (n_341, n_1270, n_338);
  nand g597 (n_1271, A[0], n_337);
  nand g598 (n_1272, n_338, n_337);
  nand g599 (n_1273, A[0], n_338);
  nand g600 (n_346, n_1271, n_1272, n_1273);
  xor g601 (n_1274, n_339, n_340);
  xor g602 (n_229, n_1274, n_341);
  nand g603 (n_1275, n_339, n_340);
  nand g604 (n_1276, n_341, n_340);
  nand g605 (n_1277, n_339, n_341);
  nand g606 (n_142, n_1275, n_1276, n_1277);
  xor g607 (n_1278, A[11], A[9]);
  xor g608 (n_344, n_1278, A[5]);
  nand g609 (n_1279, A[11], A[9]);
  nand g610 (n_1280, A[5], A[9]);
  nand g611 (n_1281, A[11], A[5]);
  nand g612 (n_349, n_1279, n_1280, n_1281);
  xor g613 (n_1282, A[3], A[7]);
  xor g614 (n_345, n_1282, A[1]);
  nand g618 (n_350, n_1256, n_1241, n_1232);
  xor g619 (n_1286, n_342, n_343);
  xor g620 (n_347, n_1286, n_344);
  nand g621 (n_1287, n_342, n_343);
  nand g622 (n_1288, n_344, n_343);
  nand g623 (n_1289, n_342, n_344);
  nand g624 (n_354, n_1287, n_1288, n_1289);
  xor g625 (n_1290, n_345, n_346);
  xor g626 (n_228, n_1290, n_347);
  nand g627 (n_1291, n_345, n_346);
  nand g628 (n_1292, n_347, n_346);
  nand g629 (n_1293, n_345, n_347);
  nand g630 (n_141, n_1291, n_1292, n_1293);
  xor g631 (n_348, A[12], A[10]);
  and g632 (n_355, A[12], A[10]);
  xor g634 (n_351, n_327, A[8]);
  nand g636 (n_1296, A[8], A[4]);
  xor g640 (n_352, Z[2], n_348);
  nand g642 (n_1300, n_348, A[0]);
  nand g643 (n_1301, A[2], n_348);
  nand g644 (n_359, n_1235, n_1300, n_1301);
  xor g645 (n_1302, n_349, n_350);
  xor g646 (n_353, n_1302, n_351);
  nand g647 (n_1303, n_349, n_350);
  nand g648 (n_1304, n_351, n_350);
  nand g649 (n_1305, n_349, n_351);
  nand g650 (n_361, n_1303, n_1304, n_1305);
  xor g651 (n_1306, n_352, n_353);
  xor g652 (n_227, n_1306, n_354);
  nand g653 (n_1307, n_352, n_353);
  nand g654 (n_1308, n_354, n_353);
  nand g655 (n_1309, n_352, n_354);
  nand g656 (n_140, n_1307, n_1308, n_1309);
  xor g657 (n_1310, A[13], A[11]);
  xor g658 (n_358, n_1310, A[7]);
  nand g659 (n_1311, A[13], A[11]);
  nand g660 (n_1312, A[7], A[11]);
  nand g661 (n_1313, A[13], A[7]);
  nand g662 (n_364, n_1311, n_1312, n_1313);
  xor g663 (n_1314, A[5], A[9]);
  xor g664 (n_357, n_1314, A[3]);
  nand g668 (n_365, n_1280, n_1257, n_1231);
  xor g669 (n_1318, A[1], n_355);
  xor g670 (n_360, n_1318, n_356);
  nand g671 (n_1319, A[1], n_355);
  nand g672 (n_1320, n_356, n_355);
  nand g673 (n_1321, A[1], n_356);
  nand g674 (n_368, n_1319, n_1320, n_1321);
  xor g675 (n_1322, n_357, n_358);
  xor g676 (n_362, n_1322, n_359);
  nand g677 (n_1323, n_357, n_358);
  nand g678 (n_1324, n_359, n_358);
  nand g679 (n_1325, n_357, n_359);
  nand g680 (n_370, n_1323, n_1324, n_1325);
  xor g681 (n_1326, n_360, n_361);
  xor g682 (n_226, n_1326, n_362);
  nand g683 (n_1327, n_360, n_361);
  nand g684 (n_1328, n_362, n_361);
  nand g685 (n_1329, n_360, n_362);
  nand g686 (n_139, n_1327, n_1328, n_1329);
  xor g687 (n_363, A[14], A[12]);
  and g688 (n_372, A[14], A[12]);
  xor g689 (n_1330, A[8], A[0]);
  xor g690 (n_367, n_1330, A[6]);
  nand g691 (n_1331, A[8], A[0]);
  nand g692 (n_1332, A[6], A[0]);
  xor g695 (n_1334, A[10], A[4]);
  xor g696 (n_366, n_1334, A[2]);
  nand g697 (n_1335, A[10], A[4]);
  nand g699 (n_1337, A[10], A[2]);
  nand g700 (n_374, n_1335, n_1249, n_1337);
  xor g701 (n_1338, n_363, n_364);
  xor g702 (n_369, n_1338, n_365);
  nand g703 (n_1339, n_363, n_364);
  nand g704 (n_1340, n_365, n_364);
  nand g705 (n_1341, n_363, n_365);
  nand g706 (n_378, n_1339, n_1340, n_1341);
  xor g707 (n_1342, n_366, n_367);
  xor g708 (n_371, n_1342, n_368);
  nand g709 (n_1343, n_366, n_367);
  nand g710 (n_1344, n_368, n_367);
  nand g711 (n_1345, n_366, n_368);
  nand g712 (n_381, n_1343, n_1344, n_1345);
  xor g713 (n_1346, n_369, n_370);
  xor g714 (n_225, n_1346, n_371);
  nand g715 (n_1347, n_369, n_370);
  nand g716 (n_1348, n_371, n_370);
  nand g717 (n_1349, n_369, n_371);
  nand g718 (n_138, n_1347, n_1348, n_1349);
  xor g719 (n_1350, A[15], A[13]);
  xor g720 (n_375, n_1350, A[9]);
  nand g721 (n_1351, A[15], A[13]);
  nand g722 (n_1352, A[9], A[13]);
  nand g723 (n_1353, A[15], A[9]);
  nand g724 (n_383, n_1351, n_1352, n_1353);
  xor g725 (n_1354, A[1], A[7]);
  xor g726 (n_376, n_1354, A[11]);
  nand g729 (n_1357, A[1], A[11]);
  nand g730 (n_384, n_1241, n_1312, n_1357);
  xor g732 (n_377, n_1230, n_372);
  nand g734 (n_1360, n_372, A[3]);
  nand g735 (n_1361, A[5], n_372);
  nand g736 (n_387, n_1231, n_1360, n_1361);
  xor g737 (n_1362, n_373, n_374);
  xor g738 (n_379, n_1362, n_375);
  nand g739 (n_1363, n_373, n_374);
  nand g740 (n_1364, n_375, n_374);
  nand g741 (n_1365, n_373, n_375);
  nand g742 (n_389, n_1363, n_1364, n_1365);
  xor g743 (n_1366, n_376, n_377);
  xor g744 (n_380, n_1366, n_378);
  nand g745 (n_1367, n_376, n_377);
  nand g746 (n_1368, n_378, n_377);
  nand g747 (n_1369, n_376, n_378);
  nand g748 (n_391, n_1367, n_1368, n_1369);
  xor g749 (n_1370, n_379, n_380);
  xor g750 (n_224, n_1370, n_381);
  nand g751 (n_1371, n_379, n_380);
  nand g752 (n_1372, n_381, n_380);
  nand g753 (n_1373, n_379, n_381);
  nand g754 (n_137, n_1371, n_1372, n_1373);
  xor g755 (n_382, A[16], A[14]);
  and g756 (n_393, A[16], A[14]);
  xor g757 (n_1374, A[10], A[2]);
  xor g758 (n_386, n_1374, A[0]);
  nand g761 (n_1377, A[10], A[0]);
  nand g762 (n_394, n_1337, n_1235, n_1377);
  xor g763 (n_1378, A[8], A[12]);
  xor g764 (n_385, n_1378, A[6]);
  nand g765 (n_1379, A[8], A[12]);
  nand g766 (n_1380, A[6], A[12]);
  xor g769 (n_1382, A[4], n_382);
  xor g770 (n_388, n_1382, n_383);
  nand g771 (n_1383, A[4], n_382);
  nand g772 (n_1384, n_383, n_382);
  nand g773 (n_1385, A[4], n_383);
  nand g774 (n_399, n_1383, n_1384, n_1385);
  xor g775 (n_1386, n_384, n_385);
  xor g776 (n_390, n_1386, n_386);
  nand g777 (n_1387, n_384, n_385);
  nand g778 (n_1388, n_386, n_385);
  nand g779 (n_1389, n_384, n_386);
  nand g780 (n_401, n_1387, n_1388, n_1389);
  xor g781 (n_1390, n_387, n_388);
  xor g782 (n_392, n_1390, n_389);
  nand g783 (n_1391, n_387, n_388);
  nand g784 (n_1392, n_389, n_388);
  nand g785 (n_1393, n_387, n_389);
  nand g786 (n_403, n_1391, n_1392, n_1393);
  xor g787 (n_1394, n_390, n_391);
  xor g788 (n_223, n_1394, n_392);
  nand g789 (n_1395, n_390, n_391);
  nand g790 (n_1396, n_392, n_391);
  nand g791 (n_1397, n_390, n_392);
  nand g792 (n_136, n_1395, n_1396, n_1397);
  xor g793 (n_1398, A[17], A[15]);
  xor g794 (n_397, n_1398, A[11]);
  nand g795 (n_1399, A[17], A[15]);
  nand g796 (n_1400, A[11], A[15]);
  nand g797 (n_1401, A[17], A[11]);
  nand g798 (n_406, n_1399, n_1400, n_1401);
  xor g799 (n_1402, A[3], A[1]);
  xor g800 (n_398, n_1402, A[9]);
  nand g802 (n_1404, A[9], A[1]);
  nand g804 (n_408, n_1232, n_1404, n_1257);
  xor g805 (n_1406, A[13], A[7]);
  xor g806 (n_396, n_1406, A[5]);
  nand g809 (n_1409, A[13], A[5]);
  nand g810 (n_407, n_1313, n_1239, n_1409);
  xor g811 (n_1410, n_393, n_394);
  xor g812 (n_400, n_1410, n_395);
  nand g813 (n_1411, n_393, n_394);
  nand g814 (n_1412, n_395, n_394);
  nand g815 (n_1413, n_393, n_395);
  nand g816 (n_412, n_1411, n_1412, n_1413);
  xor g817 (n_1414, n_396, n_397);
  xor g818 (n_402, n_1414, n_398);
  nand g819 (n_1415, n_396, n_397);
  nand g820 (n_1416, n_398, n_397);
  nand g821 (n_1417, n_396, n_398);
  nand g822 (n_414, n_1415, n_1416, n_1417);
  xor g823 (n_1418, n_399, n_400);
  xor g824 (n_404, n_1418, n_401);
  nand g825 (n_1419, n_399, n_400);
  nand g826 (n_1420, n_401, n_400);
  nand g827 (n_1421, n_399, n_401);
  nand g828 (n_416, n_1419, n_1420, n_1421);
  xor g829 (n_1422, n_402, n_403);
  xor g830 (n_222, n_1422, n_404);
  nand g831 (n_1423, n_402, n_403);
  nand g832 (n_1424, n_404, n_403);
  nand g833 (n_1425, n_402, n_404);
  nand g834 (n_135, n_1423, n_1424, n_1425);
  xor g835 (n_405, A[18], A[16]);
  and g836 (n_418, A[18], A[16]);
  xor g837 (n_1426, A[12], A[4]);
  xor g838 (n_409, n_1426, A[2]);
  nand g839 (n_1427, A[12], A[4]);
  nand g841 (n_1429, A[12], A[2]);
  nand g842 (n_419, n_1427, n_1249, n_1429);
  xor g843 (n_1430, A[10], A[0]);
  xor g844 (n_410, n_1430, A[14]);
  nand g846 (n_1432, A[14], A[0]);
  nand g847 (n_1433, A[10], A[14]);
  nand g848 (n_420, n_1377, n_1432, n_1433);
  xor g850 (n_411, n_330, n_405);
  nand g852 (n_1436, n_405, A[6]);
  nand g853 (n_1437, A[8], n_405);
  xor g855 (n_1438, n_406, n_407);
  xor g856 (n_413, n_1438, n_408);
  nand g857 (n_1439, n_406, n_407);
  nand g858 (n_1440, n_408, n_407);
  nand g859 (n_1441, n_406, n_408);
  nand g860 (n_426, n_1439, n_1440, n_1441);
  xor g861 (n_1442, n_409, n_410);
  xor g862 (n_415, n_1442, n_411);
  nand g863 (n_1443, n_409, n_410);
  nand g864 (n_1444, n_411, n_410);
  nand g865 (n_1445, n_409, n_411);
  nand g866 (n_427, n_1443, n_1444, n_1445);
  xor g867 (n_1446, n_412, n_413);
  xor g868 (n_417, n_1446, n_414);
  nand g869 (n_1447, n_412, n_413);
  nand g870 (n_1448, n_414, n_413);
  nand g871 (n_1449, n_412, n_414);
  nand g872 (n_430, n_1447, n_1448, n_1449);
  xor g873 (n_1450, n_415, n_416);
  xor g874 (n_221, n_1450, n_417);
  nand g875 (n_1451, n_415, n_416);
  nand g876 (n_1452, n_417, n_416);
  nand g877 (n_1453, n_415, n_417);
  nand g878 (n_134, n_1451, n_1452, n_1453);
  xor g879 (n_1454, A[19], A[17]);
  xor g880 (n_422, n_1454, A[13]);
  nand g881 (n_1455, A[19], A[17]);
  nand g882 (n_1456, A[13], A[17]);
  nand g883 (n_1457, A[19], A[13]);
  nand g884 (n_432, n_1455, n_1456, n_1457);
  xor g886 (n_423, n_1230, A[11]);
  nand g888 (n_1460, A[11], A[3]);
  nand g890 (n_433, n_1231, n_1460, n_1281);
  xor g891 (n_1462, A[1], A[15]);
  xor g892 (n_421, n_1462, A[9]);
  nand g893 (n_1463, A[1], A[15]);
  nand g896 (n_434, n_1463, n_1353, n_1404);
  xor g897 (n_1466, A[7], n_418);
  xor g898 (n_425, n_1466, n_419);
  nand g899 (n_1467, A[7], n_418);
  nand g900 (n_1468, n_419, n_418);
  nand g901 (n_1469, A[7], n_419);
  nand g902 (n_438, n_1467, n_1468, n_1469);
  xor g903 (n_1470, n_420, n_421);
  xor g904 (n_428, n_1470, n_422);
  nand g905 (n_1471, n_420, n_421);
  nand g906 (n_1472, n_422, n_421);
  nand g907 (n_1473, n_420, n_422);
  nand g908 (n_440, n_1471, n_1472, n_1473);
  xor g909 (n_1474, n_423, n_424);
  xor g910 (n_429, n_1474, n_425);
  nand g911 (n_1475, n_423, n_424);
  nand g912 (n_1476, n_425, n_424);
  nand g913 (n_1477, n_423, n_425);
  nand g914 (n_442, n_1475, n_1476, n_1477);
  xor g915 (n_1478, n_426, n_427);
  xor g916 (n_431, n_1478, n_428);
  nand g917 (n_1479, n_426, n_427);
  nand g918 (n_1480, n_428, n_427);
  nand g919 (n_1481, n_426, n_428);
  nand g920 (n_444, n_1479, n_1480, n_1481);
  xor g921 (n_1482, n_429, n_430);
  xor g922 (n_220, n_1482, n_431);
  nand g923 (n_1483, n_429, n_430);
  nand g924 (n_1484, n_431, n_430);
  nand g925 (n_1485, n_429, n_431);
  nand g926 (n_133, n_1483, n_1484, n_1485);
  xor g927 (n_1486, A[20], A[18]);
  xor g928 (n_436, n_1486, A[14]);
  nand g929 (n_1487, A[20], A[18]);
  nand g930 (n_1488, A[14], A[18]);
  nand g931 (n_1489, A[20], A[14]);
  nand g932 (n_446, n_1487, n_1488, n_1489);
  xor g934 (n_437, n_327, A[12]);
  xor g939 (n_1494, A[2], A[16]);
  xor g940 (n_435, n_1494, A[10]);
  nand g941 (n_1495, A[2], A[16]);
  nand g942 (n_1496, A[10], A[16]);
  nand g944 (n_448, n_1495, n_1496, n_1337);
  xor g945 (n_1498, A[8], n_432);
  xor g946 (n_439, n_1498, n_433);
  nand g947 (n_1499, A[8], n_432);
  nand g948 (n_1500, n_433, n_432);
  nand g949 (n_1501, A[8], n_433);
  nand g950 (n_149, n_1499, n_1500, n_1501);
  xor g951 (n_1502, n_434, n_435);
  xor g952 (n_441, n_1502, n_436);
  nand g953 (n_1503, n_434, n_435);
  nand g954 (n_1504, n_436, n_435);
  nand g955 (n_1505, n_434, n_436);
  nand g956 (n_151, n_1503, n_1504, n_1505);
  xor g957 (n_1506, n_437, n_438);
  xor g958 (n_443, n_1506, n_439);
  nand g959 (n_1507, n_437, n_438);
  nand g960 (n_1508, n_439, n_438);
  nand g961 (n_1509, n_437, n_439);
  nand g962 (n_153, n_1507, n_1508, n_1509);
  xor g963 (n_1510, n_440, n_441);
  xor g964 (n_445, n_1510, n_442);
  nand g965 (n_1511, n_440, n_441);
  nand g966 (n_1512, n_442, n_441);
  nand g967 (n_1513, n_440, n_442);
  nand g968 (n_453, n_1511, n_1512, n_1513);
  xor g969 (n_1514, n_443, n_444);
  xor g970 (n_219, n_1514, n_445);
  nand g971 (n_1515, n_443, n_444);
  nand g972 (n_1516, n_445, n_444);
  nand g973 (n_1517, n_443, n_445);
  nand g974 (n_132, n_1515, n_1516, n_1517);
  xor g975 (n_1518, A[21], A[19]);
  xor g976 (n_450, n_1518, A[15]);
  nand g977 (n_1519, A[21], A[19]);
  nand g978 (n_1520, A[15], A[19]);
  nand g979 (n_1521, A[21], A[15]);
  nand g980 (n_455, n_1519, n_1520, n_1521);
  xor g982 (n_451, n_1238, A[13]);
  xor g987 (n_1526, A[3], A[17]);
  xor g988 (n_449, n_1526, A[11]);
  nand g989 (n_1527, A[3], A[17]);
  nand g992 (n_457, n_1527, n_1401, n_1460);
  xor g993 (n_1530, A[9], n_446);
  xor g994 (n_150, n_1530, n_447);
  nand g995 (n_1531, A[9], n_446);
  nand g996 (n_1532, n_447, n_446);
  nand g997 (n_1533, A[9], n_447);
  nand g998 (n_461, n_1531, n_1532, n_1533);
  xor g999 (n_1534, n_448, n_449);
  xor g1000 (n_152, n_1534, n_450);
  nand g1001 (n_1535, n_448, n_449);
  nand g1002 (n_1536, n_450, n_449);
  nand g1003 (n_1537, n_448, n_450);
  nand g1004 (n_463, n_1535, n_1536, n_1537);
  xor g1005 (n_1538, n_451, n_149);
  xor g1006 (n_452, n_1538, n_150);
  nand g1007 (n_1539, n_451, n_149);
  nand g1008 (n_1540, n_150, n_149);
  nand g1009 (n_1541, n_451, n_150);
  nand g1010 (n_465, n_1539, n_1540, n_1541);
  xor g1011 (n_1542, n_151, n_152);
  xor g1012 (n_454, n_1542, n_153);
  nand g1013 (n_1543, n_151, n_152);
  nand g1014 (n_1544, n_153, n_152);
  nand g1015 (n_1545, n_151, n_153);
  nand g1016 (n_468, n_1543, n_1544, n_1545);
  xor g1017 (n_1546, n_452, n_453);
  xor g1018 (n_218, n_1546, n_454);
  nand g1019 (n_1547, n_452, n_453);
  nand g1020 (n_1548, n_454, n_453);
  nand g1021 (n_1549, n_452, n_454);
  nand g1022 (n_131, n_1547, n_1548, n_1549);
  xor g1023 (n_1550, A[22], A[20]);
  xor g1024 (n_459, n_1550, A[16]);
  nand g1025 (n_1551, A[22], A[20]);
  nand g1026 (n_1552, A[16], A[20]);
  nand g1027 (n_1553, A[22], A[16]);
  nand g1028 (n_469, n_1551, n_1552, n_1553);
  xor g1030 (n_460, n_330, A[14]);
  nand g1032 (n_1556, A[14], A[6]);
  nand g1033 (n_1557, A[8], A[14]);
  xor g1035 (n_1558, A[4], A[18]);
  xor g1036 (n_458, n_1558, A[12]);
  nand g1037 (n_1559, A[4], A[18]);
  nand g1038 (n_1560, A[12], A[18]);
  nand g1040 (n_471, n_1559, n_1560, n_1427);
  xor g1041 (n_1562, A[10], n_455);
  xor g1042 (n_462, n_1562, n_407);
  nand g1043 (n_1563, A[10], n_455);
  nand g1044 (n_1564, n_407, n_455);
  nand g1045 (n_1565, A[10], n_407);
  nand g1046 (n_475, n_1563, n_1564, n_1565);
  xor g1047 (n_1566, n_457, n_458);
  xor g1048 (n_464, n_1566, n_459);
  nand g1049 (n_1567, n_457, n_458);
  nand g1050 (n_1568, n_459, n_458);
  nand g1051 (n_1569, n_457, n_459);
  nand g1052 (n_477, n_1567, n_1568, n_1569);
  xor g1053 (n_1570, n_460, n_461);
  xor g1054 (n_466, n_1570, n_462);
  nand g1055 (n_1571, n_460, n_461);
  nand g1056 (n_1572, n_462, n_461);
  nand g1057 (n_1573, n_460, n_462);
  nand g1058 (n_479, n_1571, n_1572, n_1573);
  xor g1059 (n_1574, n_463, n_464);
  xor g1060 (n_467, n_1574, n_465);
  nand g1061 (n_1575, n_463, n_464);
  nand g1062 (n_1576, n_465, n_464);
  nand g1063 (n_1577, n_463, n_465);
  nand g1064 (n_482, n_1575, n_1576, n_1577);
  xor g1065 (n_1578, n_466, n_467);
  xor g1066 (n_217, n_1578, n_468);
  nand g1067 (n_1579, n_466, n_467);
  nand g1068 (n_1580, n_468, n_467);
  nand g1069 (n_1581, n_466, n_468);
  nand g1070 (n_130, n_1579, n_1580, n_1581);
  xor g1071 (n_1582, A[23], A[21]);
  xor g1072 (n_473, n_1582, A[17]);
  nand g1073 (n_1583, A[23], A[21]);
  nand g1074 (n_1584, A[17], A[21]);
  nand g1075 (n_1585, A[23], A[17]);
  nand g1076 (n_483, n_1583, n_1584, n_1585);
  xor g1078 (n_474, n_1254, A[15]);
  nand g1080 (n_1588, A[15], A[7]);
  nand g1082 (n_484, n_1255, n_1588, n_1353);
  xor g1083 (n_1590, A[5], A[19]);
  xor g1084 (n_472, n_1590, A[13]);
  nand g1085 (n_1591, A[5], A[19]);
  nand g1088 (n_485, n_1591, n_1457, n_1409);
  xor g1089 (n_1594, A[11], n_469);
  xor g1090 (n_476, n_1594, n_470);
  nand g1091 (n_1595, A[11], n_469);
  nand g1092 (n_1596, n_470, n_469);
  nand g1093 (n_1597, A[11], n_470);
  nand g1094 (n_489, n_1595, n_1596, n_1597);
  xor g1095 (n_1598, n_471, n_472);
  xor g1096 (n_478, n_1598, n_473);
  nand g1097 (n_1599, n_471, n_472);
  nand g1098 (n_1600, n_473, n_472);
  nand g1099 (n_1601, n_471, n_473);
  nand g1100 (n_491, n_1599, n_1600, n_1601);
  xor g1101 (n_1602, n_474, n_475);
  xor g1102 (n_480, n_1602, n_476);
  nand g1103 (n_1603, n_474, n_475);
  nand g1104 (n_1604, n_476, n_475);
  nand g1105 (n_1605, n_474, n_476);
  nand g1106 (n_493, n_1603, n_1604, n_1605);
  xor g1107 (n_1606, n_477, n_478);
  xor g1108 (n_481, n_1606, n_479);
  nand g1109 (n_1607, n_477, n_478);
  nand g1110 (n_1608, n_479, n_478);
  nand g1111 (n_1609, n_477, n_479);
  nand g1112 (n_496, n_1607, n_1608, n_1609);
  xor g1113 (n_1610, n_480, n_481);
  xor g1114 (n_216, n_1610, n_482);
  nand g1115 (n_1611, n_480, n_481);
  nand g1116 (n_1612, n_482, n_481);
  nand g1117 (n_1613, n_480, n_482);
  nand g1118 (n_129, n_1611, n_1612, n_1613);
  xor g1119 (n_1614, A[24], A[22]);
  xor g1120 (n_487, n_1614, A[18]);
  nand g1121 (n_1615, A[24], A[22]);
  nand g1122 (n_1616, A[18], A[22]);
  nand g1123 (n_1617, A[24], A[18]);
  nand g1124 (n_497, n_1615, n_1616, n_1617);
  xor g1126 (n_488, n_337, A[16]);
  nand g1128 (n_1620, A[16], A[8]);
  xor g1131 (n_1622, A[6], A[20]);
  xor g1132 (n_486, n_1622, A[14]);
  nand g1133 (n_1623, A[6], A[20]);
  nand g1136 (n_499, n_1623, n_1489, n_1556);
  xor g1137 (n_1626, A[12], n_483);
  xor g1138 (n_490, n_1626, n_484);
  nand g1139 (n_1627, A[12], n_483);
  nand g1140 (n_1628, n_484, n_483);
  nand g1141 (n_1629, A[12], n_484);
  nand g1142 (n_503, n_1627, n_1628, n_1629);
  xor g1143 (n_1630, n_485, n_486);
  xor g1144 (n_492, n_1630, n_487);
  nand g1145 (n_1631, n_485, n_486);
  nand g1146 (n_1632, n_487, n_486);
  nand g1147 (n_1633, n_485, n_487);
  nand g1148 (n_505, n_1631, n_1632, n_1633);
  xor g1149 (n_1634, n_488, n_489);
  xor g1150 (n_494, n_1634, n_490);
  nand g1151 (n_1635, n_488, n_489);
  nand g1152 (n_1636, n_490, n_489);
  nand g1153 (n_1637, n_488, n_490);
  nand g1154 (n_507, n_1635, n_1636, n_1637);
  xor g1155 (n_1638, n_491, n_492);
  xor g1156 (n_495, n_1638, n_493);
  nand g1157 (n_1639, n_491, n_492);
  nand g1158 (n_1640, n_493, n_492);
  nand g1159 (n_1641, n_491, n_493);
  nand g1160 (n_510, n_1639, n_1640, n_1641);
  xor g1161 (n_1642, n_494, n_495);
  xor g1162 (n_215, n_1642, n_496);
  nand g1163 (n_1643, n_494, n_495);
  nand g1164 (n_1644, n_496, n_495);
  nand g1165 (n_1645, n_494, n_496);
  nand g1166 (n_128, n_1643, n_1644, n_1645);
  xor g1167 (n_1646, A[25], A[23]);
  xor g1168 (n_501, n_1646, A[19]);
  nand g1169 (n_1647, A[25], A[23]);
  nand g1170 (n_1648, A[19], A[23]);
  nand g1171 (n_1649, A[25], A[19]);
  nand g1172 (n_511, n_1647, n_1648, n_1649);
  xor g1174 (n_502, n_1278, A[17]);
  nand g1176 (n_1652, A[17], A[9]);
  nand g1178 (n_512, n_1279, n_1652, n_1401);
  xor g1179 (n_1654, A[7], A[21]);
  xor g1180 (n_500, n_1654, A[15]);
  nand g1181 (n_1655, A[7], A[21]);
  nand g1184 (n_513, n_1655, n_1521, n_1588);
  xor g1185 (n_1658, A[13], n_497);
  xor g1186 (n_504, n_1658, n_498);
  nand g1187 (n_1659, A[13], n_497);
  nand g1188 (n_1660, n_498, n_497);
  nand g1189 (n_1661, A[13], n_498);
  nand g1190 (n_517, n_1659, n_1660, n_1661);
  xor g1191 (n_1662, n_499, n_500);
  xor g1192 (n_506, n_1662, n_501);
  nand g1193 (n_1663, n_499, n_500);
  nand g1194 (n_1664, n_501, n_500);
  nand g1195 (n_1665, n_499, n_501);
  nand g1196 (n_519, n_1663, n_1664, n_1665);
  xor g1197 (n_1666, n_502, n_503);
  xor g1198 (n_508, n_1666, n_504);
  nand g1199 (n_1667, n_502, n_503);
  nand g1200 (n_1668, n_504, n_503);
  nand g1201 (n_1669, n_502, n_504);
  nand g1202 (n_521, n_1667, n_1668, n_1669);
  xor g1203 (n_1670, n_505, n_506);
  xor g1204 (n_509, n_1670, n_507);
  nand g1205 (n_1671, n_505, n_506);
  nand g1206 (n_1672, n_507, n_506);
  nand g1207 (n_1673, n_505, n_507);
  nand g1208 (n_524, n_1671, n_1672, n_1673);
  xor g1209 (n_1674, n_508, n_509);
  xor g1210 (n_214, n_1674, n_510);
  nand g1211 (n_1675, n_508, n_509);
  nand g1212 (n_1676, n_510, n_509);
  nand g1213 (n_1677, n_508, n_510);
  nand g1214 (n_127, n_1675, n_1676, n_1677);
  xor g1215 (n_1678, A[26], A[24]);
  xor g1216 (n_515, n_1678, A[20]);
  nand g1217 (n_1679, A[26], A[24]);
  nand g1218 (n_1680, A[20], A[24]);
  nand g1219 (n_1681, A[26], A[20]);
  nand g1220 (n_525, n_1679, n_1680, n_1681);
  xor g1222 (n_516, n_348, A[18]);
  nand g1224 (n_1684, A[18], A[10]);
  xor g1227 (n_1686, A[8], A[22]);
  xor g1228 (n_514, n_1686, A[16]);
  nand g1229 (n_1687, A[8], A[22]);
  nand g1232 (n_527, n_1687, n_1553, n_1620);
  xor g1233 (n_1690, A[14], n_511);
  xor g1234 (n_518, n_1690, n_512);
  nand g1235 (n_1691, A[14], n_511);
  nand g1236 (n_1692, n_512, n_511);
  nand g1237 (n_1693, A[14], n_512);
  nand g1238 (n_529, n_1691, n_1692, n_1693);
  xor g1239 (n_1694, n_513, n_514);
  xor g1240 (n_520, n_1694, n_515);
  nand g1241 (n_1695, n_513, n_514);
  nand g1242 (n_1696, n_515, n_514);
  nand g1243 (n_1697, n_513, n_515);
  nand g1244 (n_531, n_1695, n_1696, n_1697);
  xor g1245 (n_1698, n_516, n_517);
  xor g1246 (n_522, n_1698, n_518);
  nand g1247 (n_1699, n_516, n_517);
  nand g1248 (n_1700, n_518, n_517);
  nand g1249 (n_1701, n_516, n_518);
  nand g1250 (n_533, n_1699, n_1700, n_1701);
  xor g1251 (n_1702, n_519, n_520);
  xor g1252 (n_523, n_1702, n_521);
  nand g1253 (n_1703, n_519, n_520);
  nand g1254 (n_1704, n_521, n_520);
  nand g1255 (n_1705, n_519, n_521);
  nand g1256 (n_536, n_1703, n_1704, n_1705);
  xor g1257 (n_1706, n_522, n_523);
  xor g1258 (n_213, n_1706, n_524);
  nand g1259 (n_1707, n_522, n_523);
  nand g1260 (n_1708, n_524, n_523);
  nand g1261 (n_1709, n_522, n_524);
  nand g1262 (n_126, n_1707, n_1708, n_1709);
  xor g1263 (n_1710, A[27], A[25]);
  xor g1264 (n_237, n_1710, A[21]);
  nand g1265 (n_1711, A[27], A[25]);
  nand g1266 (n_1712, A[21], A[25]);
  nand g1267 (n_1713, A[27], A[21]);
  nand g1268 (n_537, n_1711, n_1712, n_1713);
  xor g1270 (n_528, n_1310, A[19]);
  nand g1272 (n_1716, A[19], A[11]);
  nand g1274 (n_538, n_1311, n_1716, n_1457);
  xor g1275 (n_1718, A[9], A[23]);
  xor g1276 (n_236, n_1718, A[17]);
  nand g1277 (n_1719, A[9], A[23]);
  nand g1280 (n_539, n_1719, n_1585, n_1652);
  xor g1281 (n_1722, A[15], n_525);
  xor g1282 (n_530, n_1722, n_526);
  nand g1283 (n_1723, A[15], n_525);
  nand g1284 (n_1724, n_526, n_525);
  nand g1285 (n_1725, A[15], n_526);
  nand g1286 (n_543, n_1723, n_1724, n_1725);
  xor g1287 (n_1726, n_527, n_236);
  xor g1288 (n_532, n_1726, n_237);
  nand g1289 (n_1727, n_527, n_236);
  nand g1290 (n_1728, n_237, n_236);
  nand g1291 (n_1729, n_527, n_237);
  nand g1292 (n_545, n_1727, n_1728, n_1729);
  xor g1293 (n_1730, n_528, n_529);
  xor g1294 (n_534, n_1730, n_530);
  nand g1295 (n_1731, n_528, n_529);
  nand g1296 (n_1732, n_530, n_529);
  nand g1297 (n_1733, n_528, n_530);
  nand g1298 (n_547, n_1731, n_1732, n_1733);
  xor g1299 (n_1734, n_531, n_532);
  xor g1300 (n_535, n_1734, n_533);
  nand g1301 (n_1735, n_531, n_532);
  nand g1302 (n_1736, n_533, n_532);
  nand g1303 (n_1737, n_531, n_533);
  nand g1304 (n_550, n_1735, n_1736, n_1737);
  xor g1305 (n_1738, n_534, n_535);
  xor g1306 (n_212, n_1738, n_536);
  nand g1307 (n_1739, n_534, n_535);
  nand g1308 (n_1740, n_536, n_535);
  nand g1309 (n_1741, n_534, n_536);
  nand g1310 (n_125, n_1739, n_1740, n_1741);
  xor g1311 (n_1742, A[28], A[26]);
  xor g1312 (n_541, n_1742, A[22]);
  nand g1313 (n_1743, A[28], A[26]);
  nand g1314 (n_1744, A[22], A[26]);
  nand g1315 (n_1745, A[28], A[22]);
  nand g1316 (n_551, n_1743, n_1744, n_1745);
  xor g1318 (n_542, n_363, A[20]);
  nand g1320 (n_1748, A[20], A[12]);
  xor g1323 (n_1750, A[10], A[24]);
  xor g1324 (n_540, n_1750, A[18]);
  nand g1325 (n_1751, A[10], A[24]);
  nand g1328 (n_553, n_1751, n_1617, n_1684);
  xor g1329 (n_1754, A[16], n_537);
  xor g1330 (n_544, n_1754, n_538);
  nand g1331 (n_1755, A[16], n_537);
  nand g1332 (n_1756, n_538, n_537);
  nand g1333 (n_1757, A[16], n_538);
  nand g1334 (n_557, n_1755, n_1756, n_1757);
  xor g1335 (n_1758, n_539, n_540);
  xor g1336 (n_546, n_1758, n_541);
  nand g1337 (n_1759, n_539, n_540);
  nand g1338 (n_1760, n_541, n_540);
  nand g1339 (n_1761, n_539, n_541);
  nand g1340 (n_559, n_1759, n_1760, n_1761);
  xor g1341 (n_1762, n_542, n_543);
  xor g1342 (n_548, n_1762, n_544);
  nand g1343 (n_1763, n_542, n_543);
  nand g1344 (n_1764, n_544, n_543);
  nand g1345 (n_1765, n_542, n_544);
  nand g1346 (n_561, n_1763, n_1764, n_1765);
  xor g1347 (n_1766, n_545, n_546);
  xor g1348 (n_549, n_1766, n_547);
  nand g1349 (n_1767, n_545, n_546);
  nand g1350 (n_1768, n_547, n_546);
  nand g1351 (n_1769, n_545, n_547);
  nand g1352 (n_564, n_1767, n_1768, n_1769);
  xor g1353 (n_1770, n_548, n_549);
  xor g1354 (n_211, n_1770, n_550);
  nand g1355 (n_1771, n_548, n_549);
  nand g1356 (n_1772, n_550, n_549);
  nand g1357 (n_1773, n_548, n_550);
  nand g1358 (n_124, n_1771, n_1772, n_1773);
  xor g1359 (n_1774, A[29], A[27]);
  xor g1360 (n_555, n_1774, A[23]);
  nand g1361 (n_1775, A[29], A[27]);
  nand g1362 (n_1776, A[23], A[27]);
  nand g1363 (n_1777, A[29], A[23]);
  nand g1364 (n_565, n_1775, n_1776, n_1777);
  xor g1366 (n_556, n_1350, A[21]);
  nand g1368 (n_1780, A[21], A[13]);
  nand g1370 (n_566, n_1351, n_1780, n_1521);
  xor g1371 (n_1782, A[11], A[25]);
  xor g1372 (n_554, n_1782, A[19]);
  nand g1373 (n_1783, A[11], A[25]);
  nand g1376 (n_567, n_1783, n_1649, n_1716);
  xor g1377 (n_1786, A[17], n_551);
  xor g1378 (n_558, n_1786, n_552);
  nand g1379 (n_1787, A[17], n_551);
  nand g1380 (n_1788, n_552, n_551);
  nand g1381 (n_1789, A[17], n_552);
  nand g1382 (n_571, n_1787, n_1788, n_1789);
  xor g1383 (n_1790, n_553, n_554);
  xor g1384 (n_560, n_1790, n_555);
  nand g1385 (n_1791, n_553, n_554);
  nand g1386 (n_1792, n_555, n_554);
  nand g1387 (n_1793, n_553, n_555);
  nand g1388 (n_573, n_1791, n_1792, n_1793);
  xor g1389 (n_1794, n_556, n_557);
  xor g1390 (n_562, n_1794, n_558);
  nand g1391 (n_1795, n_556, n_557);
  nand g1392 (n_1796, n_558, n_557);
  nand g1393 (n_1797, n_556, n_558);
  nand g1394 (n_575, n_1795, n_1796, n_1797);
  xor g1395 (n_1798, n_559, n_560);
  xor g1396 (n_563, n_1798, n_561);
  nand g1397 (n_1799, n_559, n_560);
  nand g1398 (n_1800, n_561, n_560);
  nand g1399 (n_1801, n_559, n_561);
  nand g1400 (n_578, n_1799, n_1800, n_1801);
  xor g1401 (n_1802, n_562, n_563);
  xor g1402 (n_210, n_1802, n_564);
  nand g1403 (n_1803, n_562, n_563);
  nand g1404 (n_1804, n_564, n_563);
  nand g1405 (n_1805, n_562, n_564);
  nand g1406 (n_123, n_1803, n_1804, n_1805);
  xor g1407 (n_1806, A[30], A[28]);
  xor g1408 (n_569, n_1806, A[24]);
  nand g1409 (n_1807, A[30], A[28]);
  nand g1410 (n_1808, A[24], A[28]);
  nand g1411 (n_1809, A[30], A[24]);
  nand g1412 (n_579, n_1807, n_1808, n_1809);
  xor g1414 (n_570, n_382, A[22]);
  nand g1416 (n_1812, A[22], A[14]);
  xor g1419 (n_1814, A[12], A[26]);
  xor g1420 (n_568, n_1814, A[20]);
  nand g1421 (n_1815, A[12], A[26]);
  nand g1424 (n_581, n_1815, n_1681, n_1748);
  xor g1425 (n_1818, A[18], n_565);
  xor g1426 (n_572, n_1818, n_566);
  nand g1427 (n_1819, A[18], n_565);
  nand g1428 (n_1820, n_566, n_565);
  nand g1429 (n_1821, A[18], n_566);
  nand g1430 (n_585, n_1819, n_1820, n_1821);
  xor g1431 (n_1822, n_567, n_568);
  xor g1432 (n_574, n_1822, n_569);
  nand g1433 (n_1823, n_567, n_568);
  nand g1434 (n_1824, n_569, n_568);
  nand g1435 (n_1825, n_567, n_569);
  nand g1436 (n_587, n_1823, n_1824, n_1825);
  xor g1437 (n_1826, n_570, n_571);
  xor g1438 (n_576, n_1826, n_572);
  nand g1439 (n_1827, n_570, n_571);
  nand g1440 (n_1828, n_572, n_571);
  nand g1441 (n_1829, n_570, n_572);
  nand g1442 (n_589, n_1827, n_1828, n_1829);
  xor g1443 (n_1830, n_573, n_574);
  xor g1444 (n_577, n_1830, n_575);
  nand g1445 (n_1831, n_573, n_574);
  nand g1446 (n_1832, n_575, n_574);
  nand g1447 (n_1833, n_573, n_575);
  nand g1448 (n_592, n_1831, n_1832, n_1833);
  xor g1449 (n_1834, n_576, n_577);
  xor g1450 (n_209, n_1834, n_578);
  nand g1451 (n_1835, n_576, n_577);
  nand g1452 (n_1836, n_578, n_577);
  nand g1453 (n_1837, n_576, n_578);
  nand g1454 (n_122, n_1835, n_1836, n_1837);
  xor g1455 (n_1838, A[31], A[29]);
  xor g1456 (n_583, n_1838, A[25]);
  nand g1457 (n_1839, A[31], A[29]);
  nand g1458 (n_1840, A[25], A[29]);
  nand g1459 (n_1841, A[31], A[25]);
  nand g1460 (n_593, n_1839, n_1840, n_1841);
  xor g1462 (n_584, n_1398, A[23]);
  nand g1464 (n_1844, A[23], A[15]);
  nand g1466 (n_594, n_1399, n_1844, n_1585);
  xor g1467 (n_1846, A[13], A[27]);
  xor g1468 (n_582, n_1846, A[21]);
  nand g1469 (n_1847, A[13], A[27]);
  nand g1472 (n_595, n_1847, n_1713, n_1780);
  xor g1473 (n_1850, A[19], n_579);
  xor g1474 (n_586, n_1850, n_580);
  nand g1475 (n_1851, A[19], n_579);
  nand g1476 (n_1852, n_580, n_579);
  nand g1477 (n_1853, A[19], n_580);
  nand g1478 (n_599, n_1851, n_1852, n_1853);
  xor g1479 (n_1854, n_581, n_582);
  xor g1480 (n_588, n_1854, n_583);
  nand g1481 (n_1855, n_581, n_582);
  nand g1482 (n_1856, n_583, n_582);
  nand g1483 (n_1857, n_581, n_583);
  nand g1484 (n_601, n_1855, n_1856, n_1857);
  xor g1485 (n_1858, n_584, n_585);
  xor g1486 (n_590, n_1858, n_586);
  nand g1487 (n_1859, n_584, n_585);
  nand g1488 (n_1860, n_586, n_585);
  nand g1489 (n_1861, n_584, n_586);
  nand g1490 (n_603, n_1859, n_1860, n_1861);
  xor g1491 (n_1862, n_587, n_588);
  xor g1492 (n_591, n_1862, n_589);
  nand g1493 (n_1863, n_587, n_588);
  nand g1494 (n_1864, n_589, n_588);
  nand g1495 (n_1865, n_587, n_589);
  nand g1496 (n_606, n_1863, n_1864, n_1865);
  xor g1497 (n_1866, n_590, n_591);
  xor g1498 (n_208, n_1866, n_592);
  nand g1499 (n_1867, n_590, n_591);
  nand g1500 (n_1868, n_592, n_591);
  nand g1501 (n_1869, n_590, n_592);
  nand g1502 (n_121, n_1867, n_1868, n_1869);
  xor g1503 (n_1870, A[32], A[30]);
  xor g1504 (n_597, n_1870, A[26]);
  nand g1505 (n_1871, A[32], A[30]);
  nand g1506 (n_1872, A[26], A[30]);
  nand g1507 (n_1873, A[32], A[26]);
  nand g1508 (n_607, n_1871, n_1872, n_1873);
  xor g1510 (n_598, n_405, A[24]);
  nand g1512 (n_1876, A[24], A[16]);
  xor g1515 (n_1878, A[14], A[28]);
  xor g1516 (n_596, n_1878, A[22]);
  nand g1517 (n_1879, A[14], A[28]);
  nand g1520 (n_609, n_1879, n_1745, n_1812);
  xor g1521 (n_1882, A[20], n_593);
  xor g1522 (n_600, n_1882, n_594);
  nand g1523 (n_1883, A[20], n_593);
  nand g1524 (n_1884, n_594, n_593);
  nand g1525 (n_1885, A[20], n_594);
  nand g1526 (n_613, n_1883, n_1884, n_1885);
  xor g1527 (n_1886, n_595, n_596);
  xor g1528 (n_602, n_1886, n_597);
  nand g1529 (n_1887, n_595, n_596);
  nand g1530 (n_1888, n_597, n_596);
  nand g1531 (n_1889, n_595, n_597);
  nand g1532 (n_615, n_1887, n_1888, n_1889);
  xor g1533 (n_1890, n_598, n_599);
  xor g1534 (n_604, n_1890, n_600);
  nand g1535 (n_1891, n_598, n_599);
  nand g1536 (n_1892, n_600, n_599);
  nand g1537 (n_1893, n_598, n_600);
  nand g1538 (n_617, n_1891, n_1892, n_1893);
  xor g1539 (n_1894, n_601, n_602);
  xor g1540 (n_605, n_1894, n_603);
  nand g1541 (n_1895, n_601, n_602);
  nand g1542 (n_1896, n_603, n_602);
  nand g1543 (n_1897, n_601, n_603);
  nand g1544 (n_620, n_1895, n_1896, n_1897);
  xor g1545 (n_1898, n_604, n_605);
  xor g1546 (n_207, n_1898, n_606);
  nand g1547 (n_1899, n_604, n_605);
  nand g1548 (n_1900, n_606, n_605);
  nand g1549 (n_1901, n_604, n_606);
  nand g1550 (n_120, n_1899, n_1900, n_1901);
  xor g1551 (n_1902, A[33], A[31]);
  xor g1552 (n_611, n_1902, A[27]);
  nand g1553 (n_1903, A[33], A[31]);
  nand g1554 (n_1904, A[27], A[31]);
  nand g1555 (n_1905, A[33], A[27]);
  nand g1556 (n_621, n_1903, n_1904, n_1905);
  xor g1558 (n_612, n_1454, A[25]);
  nand g1560 (n_1908, A[25], A[17]);
  nand g1562 (n_622, n_1455, n_1908, n_1649);
  xor g1563 (n_1910, A[15], A[29]);
  xor g1564 (n_610, n_1910, A[23]);
  nand g1565 (n_1911, A[15], A[29]);
  nand g1568 (n_623, n_1911, n_1777, n_1844);
  xor g1569 (n_1914, A[21], n_607);
  xor g1570 (n_614, n_1914, n_608);
  nand g1571 (n_1915, A[21], n_607);
  nand g1572 (n_1916, n_608, n_607);
  nand g1573 (n_1917, A[21], n_608);
  nand g1574 (n_627, n_1915, n_1916, n_1917);
  xor g1575 (n_1918, n_609, n_610);
  xor g1576 (n_616, n_1918, n_611);
  nand g1577 (n_1919, n_609, n_610);
  nand g1578 (n_1920, n_611, n_610);
  nand g1579 (n_1921, n_609, n_611);
  nand g1580 (n_629, n_1919, n_1920, n_1921);
  xor g1581 (n_1922, n_612, n_613);
  xor g1582 (n_618, n_1922, n_614);
  nand g1583 (n_1923, n_612, n_613);
  nand g1584 (n_1924, n_614, n_613);
  nand g1585 (n_1925, n_612, n_614);
  nand g1586 (n_631, n_1923, n_1924, n_1925);
  xor g1587 (n_1926, n_615, n_616);
  xor g1588 (n_619, n_1926, n_617);
  nand g1589 (n_1927, n_615, n_616);
  nand g1590 (n_1928, n_617, n_616);
  nand g1591 (n_1929, n_615, n_617);
  nand g1592 (n_634, n_1927, n_1928, n_1929);
  xor g1593 (n_1930, n_618, n_619);
  xor g1594 (n_206, n_1930, n_620);
  nand g1595 (n_1931, n_618, n_619);
  nand g1596 (n_1932, n_620, n_619);
  nand g1597 (n_1933, n_618, n_620);
  nand g1598 (n_119, n_1931, n_1932, n_1933);
  xor g1599 (n_1934, A[34], A[32]);
  xor g1600 (n_625, n_1934, A[28]);
  nand g1601 (n_1935, A[34], A[32]);
  nand g1602 (n_1936, A[28], A[32]);
  nand g1603 (n_1937, A[34], A[28]);
  nand g1604 (n_635, n_1935, n_1936, n_1937);
  xor g1606 (n_626, n_1486, A[26]);
  nand g1608 (n_1940, A[26], A[18]);
  nand g1610 (n_636, n_1487, n_1940, n_1681);
  xor g1611 (n_1942, A[16], A[30]);
  xor g1612 (n_624, n_1942, A[24]);
  nand g1613 (n_1943, A[16], A[30]);
  nand g1616 (n_637, n_1943, n_1809, n_1876);
  xor g1617 (n_1946, A[22], n_621);
  xor g1618 (n_628, n_1946, n_622);
  nand g1619 (n_1947, A[22], n_621);
  nand g1620 (n_1948, n_622, n_621);
  nand g1621 (n_1949, A[22], n_622);
  nand g1622 (n_641, n_1947, n_1948, n_1949);
  xor g1623 (n_1950, n_623, n_624);
  xor g1624 (n_630, n_1950, n_625);
  nand g1625 (n_1951, n_623, n_624);
  nand g1626 (n_1952, n_625, n_624);
  nand g1627 (n_1953, n_623, n_625);
  nand g1628 (n_643, n_1951, n_1952, n_1953);
  xor g1629 (n_1954, n_626, n_627);
  xor g1630 (n_632, n_1954, n_628);
  nand g1631 (n_1955, n_626, n_627);
  nand g1632 (n_1956, n_628, n_627);
  nand g1633 (n_1957, n_626, n_628);
  nand g1634 (n_645, n_1955, n_1956, n_1957);
  xor g1635 (n_1958, n_629, n_630);
  xor g1636 (n_633, n_1958, n_631);
  nand g1637 (n_1959, n_629, n_630);
  nand g1638 (n_1960, n_631, n_630);
  nand g1639 (n_1961, n_629, n_631);
  nand g1640 (n_648, n_1959, n_1960, n_1961);
  xor g1641 (n_1962, n_632, n_633);
  xor g1642 (n_205, n_1962, n_634);
  nand g1643 (n_1963, n_632, n_633);
  nand g1644 (n_1964, n_634, n_633);
  nand g1645 (n_1965, n_632, n_634);
  nand g1646 (n_118, n_1963, n_1964, n_1965);
  xor g1647 (n_1966, A[35], A[33]);
  xor g1648 (n_639, n_1966, A[29]);
  nand g1649 (n_1967, A[35], A[33]);
  nand g1650 (n_1968, A[29], A[33]);
  nand g1651 (n_1969, A[35], A[29]);
  nand g1652 (n_649, n_1967, n_1968, n_1969);
  xor g1654 (n_640, n_1518, A[27]);
  nand g1656 (n_1972, A[27], A[19]);
  nand g1658 (n_650, n_1519, n_1972, n_1713);
  xor g1659 (n_1974, A[17], A[31]);
  xor g1660 (n_638, n_1974, A[25]);
  nand g1661 (n_1975, A[17], A[31]);
  nand g1664 (n_651, n_1975, n_1841, n_1908);
  xor g1665 (n_1978, A[23], n_635);
  xor g1666 (n_642, n_1978, n_636);
  nand g1667 (n_1979, A[23], n_635);
  nand g1668 (n_1980, n_636, n_635);
  nand g1669 (n_1981, A[23], n_636);
  nand g1670 (n_655, n_1979, n_1980, n_1981);
  xor g1671 (n_1982, n_637, n_638);
  xor g1672 (n_644, n_1982, n_639);
  nand g1673 (n_1983, n_637, n_638);
  nand g1674 (n_1984, n_639, n_638);
  nand g1675 (n_1985, n_637, n_639);
  nand g1676 (n_657, n_1983, n_1984, n_1985);
  xor g1677 (n_1986, n_640, n_641);
  xor g1678 (n_646, n_1986, n_642);
  nand g1679 (n_1987, n_640, n_641);
  nand g1680 (n_1988, n_642, n_641);
  nand g1681 (n_1989, n_640, n_642);
  nand g1682 (n_659, n_1987, n_1988, n_1989);
  xor g1683 (n_1990, n_643, n_644);
  xor g1684 (n_647, n_1990, n_645);
  nand g1685 (n_1991, n_643, n_644);
  nand g1686 (n_1992, n_645, n_644);
  nand g1687 (n_1993, n_643, n_645);
  nand g1688 (n_662, n_1991, n_1992, n_1993);
  xor g1689 (n_1994, n_646, n_647);
  xor g1690 (n_204, n_1994, n_648);
  nand g1691 (n_1995, n_646, n_647);
  nand g1692 (n_1996, n_648, n_647);
  nand g1693 (n_1997, n_646, n_648);
  nand g1694 (n_117, n_1995, n_1996, n_1997);
  xor g1695 (n_1998, A[36], A[34]);
  xor g1696 (n_653, n_1998, A[30]);
  nand g1697 (n_1999, A[36], A[34]);
  nand g1698 (n_2000, A[30], A[34]);
  nand g1699 (n_2001, A[36], A[30]);
  nand g1700 (n_663, n_1999, n_2000, n_2001);
  xor g1702 (n_654, n_1550, A[28]);
  nand g1704 (n_2004, A[28], A[20]);
  nand g1706 (n_664, n_1551, n_2004, n_1745);
  xor g1707 (n_2006, A[18], A[32]);
  xor g1708 (n_652, n_2006, A[26]);
  nand g1709 (n_2007, A[18], A[32]);
  nand g1712 (n_665, n_2007, n_1873, n_1940);
  xor g1713 (n_2010, A[24], n_649);
  xor g1714 (n_656, n_2010, n_650);
  nand g1715 (n_2011, A[24], n_649);
  nand g1716 (n_2012, n_650, n_649);
  nand g1717 (n_2013, A[24], n_650);
  nand g1718 (n_669, n_2011, n_2012, n_2013);
  xor g1719 (n_2014, n_651, n_652);
  xor g1720 (n_658, n_2014, n_653);
  nand g1721 (n_2015, n_651, n_652);
  nand g1722 (n_2016, n_653, n_652);
  nand g1723 (n_2017, n_651, n_653);
  nand g1724 (n_671, n_2015, n_2016, n_2017);
  xor g1725 (n_2018, n_654, n_655);
  xor g1726 (n_660, n_2018, n_656);
  nand g1727 (n_2019, n_654, n_655);
  nand g1728 (n_2020, n_656, n_655);
  nand g1729 (n_2021, n_654, n_656);
  nand g1730 (n_673, n_2019, n_2020, n_2021);
  xor g1731 (n_2022, n_657, n_658);
  xor g1732 (n_661, n_2022, n_659);
  nand g1733 (n_2023, n_657, n_658);
  nand g1734 (n_2024, n_659, n_658);
  nand g1735 (n_2025, n_657, n_659);
  nand g1736 (n_676, n_2023, n_2024, n_2025);
  xor g1737 (n_2026, n_660, n_661);
  xor g1738 (n_203, n_2026, n_662);
  nand g1739 (n_2027, n_660, n_661);
  nand g1740 (n_2028, n_662, n_661);
  nand g1741 (n_2029, n_660, n_662);
  nand g1742 (n_116, n_2027, n_2028, n_2029);
  xor g1743 (n_2030, A[37], A[35]);
  xor g1744 (n_667, n_2030, A[31]);
  nand g1745 (n_2031, A[37], A[35]);
  nand g1746 (n_2032, A[31], A[35]);
  nand g1747 (n_2033, A[37], A[31]);
  nand g1748 (n_677, n_2031, n_2032, n_2033);
  xor g1750 (n_668, n_1582, A[29]);
  nand g1752 (n_2036, A[29], A[21]);
  nand g1754 (n_678, n_1583, n_2036, n_1777);
  xor g1755 (n_2038, A[19], A[33]);
  xor g1756 (n_666, n_2038, A[27]);
  nand g1757 (n_2039, A[19], A[33]);
  nand g1760 (n_679, n_2039, n_1905, n_1972);
  xor g1761 (n_2042, A[25], n_663);
  xor g1762 (n_670, n_2042, n_664);
  nand g1763 (n_2043, A[25], n_663);
  nand g1764 (n_2044, n_664, n_663);
  nand g1765 (n_2045, A[25], n_664);
  nand g1766 (n_683, n_2043, n_2044, n_2045);
  xor g1767 (n_2046, n_665, n_666);
  xor g1768 (n_672, n_2046, n_667);
  nand g1769 (n_2047, n_665, n_666);
  nand g1770 (n_2048, n_667, n_666);
  nand g1771 (n_2049, n_665, n_667);
  nand g1772 (n_685, n_2047, n_2048, n_2049);
  xor g1773 (n_2050, n_668, n_669);
  xor g1774 (n_674, n_2050, n_670);
  nand g1775 (n_2051, n_668, n_669);
  nand g1776 (n_2052, n_670, n_669);
  nand g1777 (n_2053, n_668, n_670);
  nand g1778 (n_687, n_2051, n_2052, n_2053);
  xor g1779 (n_2054, n_671, n_672);
  xor g1780 (n_675, n_2054, n_673);
  nand g1781 (n_2055, n_671, n_672);
  nand g1782 (n_2056, n_673, n_672);
  nand g1783 (n_2057, n_671, n_673);
  nand g1784 (n_690, n_2055, n_2056, n_2057);
  xor g1785 (n_2058, n_674, n_675);
  xor g1786 (n_202, n_2058, n_676);
  nand g1787 (n_2059, n_674, n_675);
  nand g1788 (n_2060, n_676, n_675);
  nand g1789 (n_2061, n_674, n_676);
  nand g1790 (n_115, n_2059, n_2060, n_2061);
  xor g1791 (n_2062, A[38], A[36]);
  xor g1792 (n_681, n_2062, A[32]);
  nand g1793 (n_2063, A[38], A[36]);
  nand g1794 (n_2064, A[32], A[36]);
  nand g1795 (n_2065, A[38], A[32]);
  nand g1796 (n_691, n_2063, n_2064, n_2065);
  xor g1798 (n_682, n_1614, A[30]);
  nand g1800 (n_2068, A[30], A[22]);
  nand g1802 (n_692, n_1615, n_2068, n_1809);
  xor g1803 (n_2070, A[20], A[34]);
  xor g1804 (n_680, n_2070, A[28]);
  nand g1805 (n_2071, A[20], A[34]);
  nand g1808 (n_693, n_2071, n_1937, n_2004);
  xor g1809 (n_2074, A[26], n_677);
  xor g1810 (n_684, n_2074, n_678);
  nand g1811 (n_2075, A[26], n_677);
  nand g1812 (n_2076, n_678, n_677);
  nand g1813 (n_2077, A[26], n_678);
  nand g1814 (n_697, n_2075, n_2076, n_2077);
  xor g1815 (n_2078, n_679, n_680);
  xor g1816 (n_686, n_2078, n_681);
  nand g1817 (n_2079, n_679, n_680);
  nand g1818 (n_2080, n_681, n_680);
  nand g1819 (n_2081, n_679, n_681);
  nand g1820 (n_699, n_2079, n_2080, n_2081);
  xor g1821 (n_2082, n_682, n_683);
  xor g1822 (n_688, n_2082, n_684);
  nand g1823 (n_2083, n_682, n_683);
  nand g1824 (n_2084, n_684, n_683);
  nand g1825 (n_2085, n_682, n_684);
  nand g1826 (n_701, n_2083, n_2084, n_2085);
  xor g1827 (n_2086, n_685, n_686);
  xor g1828 (n_689, n_2086, n_687);
  nand g1829 (n_2087, n_685, n_686);
  nand g1830 (n_2088, n_687, n_686);
  nand g1831 (n_2089, n_685, n_687);
  nand g1832 (n_704, n_2087, n_2088, n_2089);
  xor g1833 (n_2090, n_688, n_689);
  xor g1834 (n_201, n_2090, n_690);
  nand g1835 (n_2091, n_688, n_689);
  nand g1836 (n_2092, n_690, n_689);
  nand g1837 (n_2093, n_688, n_690);
  nand g1838 (n_114, n_2091, n_2092, n_2093);
  xor g1839 (n_2094, A[39], A[37]);
  xor g1840 (n_695, n_2094, A[33]);
  nand g1841 (n_2095, A[39], A[37]);
  nand g1842 (n_2096, A[33], A[37]);
  nand g1843 (n_2097, A[39], A[33]);
  nand g1844 (n_705, n_2095, n_2096, n_2097);
  xor g1846 (n_696, n_1646, A[31]);
  nand g1848 (n_2100, A[31], A[23]);
  nand g1850 (n_706, n_1647, n_2100, n_1841);
  xor g1851 (n_2102, A[21], A[35]);
  xor g1852 (n_694, n_2102, A[29]);
  nand g1853 (n_2103, A[21], A[35]);
  nand g1856 (n_707, n_2103, n_1969, n_2036);
  xor g1857 (n_2106, A[27], n_691);
  xor g1858 (n_698, n_2106, n_692);
  nand g1859 (n_2107, A[27], n_691);
  nand g1860 (n_2108, n_692, n_691);
  nand g1861 (n_2109, A[27], n_692);
  nand g1862 (n_711, n_2107, n_2108, n_2109);
  xor g1863 (n_2110, n_693, n_694);
  xor g1864 (n_700, n_2110, n_695);
  nand g1865 (n_2111, n_693, n_694);
  nand g1866 (n_2112, n_695, n_694);
  nand g1867 (n_2113, n_693, n_695);
  nand g1868 (n_713, n_2111, n_2112, n_2113);
  xor g1869 (n_2114, n_696, n_697);
  xor g1870 (n_702, n_2114, n_698);
  nand g1871 (n_2115, n_696, n_697);
  nand g1872 (n_2116, n_698, n_697);
  nand g1873 (n_2117, n_696, n_698);
  nand g1874 (n_715, n_2115, n_2116, n_2117);
  xor g1875 (n_2118, n_699, n_700);
  xor g1876 (n_703, n_2118, n_701);
  nand g1877 (n_2119, n_699, n_700);
  nand g1878 (n_2120, n_701, n_700);
  nand g1879 (n_2121, n_699, n_701);
  nand g1880 (n_718, n_2119, n_2120, n_2121);
  xor g1881 (n_2122, n_702, n_703);
  xor g1882 (n_200, n_2122, n_704);
  nand g1883 (n_2123, n_702, n_703);
  nand g1884 (n_2124, n_704, n_703);
  nand g1885 (n_2125, n_702, n_704);
  nand g1886 (n_113, n_2123, n_2124, n_2125);
  xor g1887 (n_2126, A[40], A[38]);
  xor g1888 (n_709, n_2126, A[34]);
  nand g1889 (n_2127, A[40], A[38]);
  nand g1890 (n_2128, A[34], A[38]);
  nand g1891 (n_2129, A[40], A[34]);
  nand g1892 (n_719, n_2127, n_2128, n_2129);
  xor g1894 (n_710, n_1678, A[32]);
  nand g1896 (n_2132, A[32], A[24]);
  nand g1898 (n_720, n_1679, n_2132, n_1873);
  xor g1899 (n_2134, A[22], A[36]);
  xor g1900 (n_708, n_2134, A[30]);
  nand g1901 (n_2135, A[22], A[36]);
  nand g1904 (n_721, n_2135, n_2001, n_2068);
  xor g1905 (n_2138, A[28], n_705);
  xor g1906 (n_712, n_2138, n_706);
  nand g1907 (n_2139, A[28], n_705);
  nand g1908 (n_2140, n_706, n_705);
  nand g1909 (n_2141, A[28], n_706);
  nand g1910 (n_725, n_2139, n_2140, n_2141);
  xor g1911 (n_2142, n_707, n_708);
  xor g1912 (n_714, n_2142, n_709);
  nand g1913 (n_2143, n_707, n_708);
  nand g1914 (n_2144, n_709, n_708);
  nand g1915 (n_2145, n_707, n_709);
  nand g1916 (n_727, n_2143, n_2144, n_2145);
  xor g1917 (n_2146, n_710, n_711);
  xor g1918 (n_716, n_2146, n_712);
  nand g1919 (n_2147, n_710, n_711);
  nand g1920 (n_2148, n_712, n_711);
  nand g1921 (n_2149, n_710, n_712);
  nand g1922 (n_729, n_2147, n_2148, n_2149);
  xor g1923 (n_2150, n_713, n_714);
  xor g1924 (n_717, n_2150, n_715);
  nand g1925 (n_2151, n_713, n_714);
  nand g1926 (n_2152, n_715, n_714);
  nand g1927 (n_2153, n_713, n_715);
  nand g1928 (n_732, n_2151, n_2152, n_2153);
  xor g1929 (n_2154, n_716, n_717);
  xor g1930 (n_199, n_2154, n_718);
  nand g1931 (n_2155, n_716, n_717);
  nand g1932 (n_2156, n_718, n_717);
  nand g1933 (n_2157, n_716, n_718);
  nand g1934 (n_112, n_2155, n_2156, n_2157);
  xor g1935 (n_2158, A[41], A[39]);
  xor g1936 (n_723, n_2158, A[35]);
  nand g1937 (n_2159, A[41], A[39]);
  nand g1938 (n_2160, A[35], A[39]);
  nand g1939 (n_2161, A[41], A[35]);
  nand g1940 (n_733, n_2159, n_2160, n_2161);
  xor g1942 (n_724, n_1710, A[33]);
  nand g1944 (n_2164, A[33], A[25]);
  nand g1946 (n_734, n_1711, n_2164, n_1905);
  xor g1947 (n_2166, A[23], A[37]);
  xor g1948 (n_722, n_2166, A[31]);
  nand g1949 (n_2167, A[23], A[37]);
  nand g1952 (n_735, n_2167, n_2033, n_2100);
  xor g1953 (n_2170, A[29], n_719);
  xor g1954 (n_726, n_2170, n_720);
  nand g1955 (n_2171, A[29], n_719);
  nand g1956 (n_2172, n_720, n_719);
  nand g1957 (n_2173, A[29], n_720);
  nand g1958 (n_739, n_2171, n_2172, n_2173);
  xor g1959 (n_2174, n_721, n_722);
  xor g1960 (n_728, n_2174, n_723);
  nand g1961 (n_2175, n_721, n_722);
  nand g1962 (n_2176, n_723, n_722);
  nand g1963 (n_2177, n_721, n_723);
  nand g1964 (n_741, n_2175, n_2176, n_2177);
  xor g1965 (n_2178, n_724, n_725);
  xor g1966 (n_730, n_2178, n_726);
  nand g1967 (n_2179, n_724, n_725);
  nand g1968 (n_2180, n_726, n_725);
  nand g1969 (n_2181, n_724, n_726);
  nand g1970 (n_743, n_2179, n_2180, n_2181);
  xor g1971 (n_2182, n_727, n_728);
  xor g1972 (n_731, n_2182, n_729);
  nand g1973 (n_2183, n_727, n_728);
  nand g1974 (n_2184, n_729, n_728);
  nand g1975 (n_2185, n_727, n_729);
  nand g1976 (n_746, n_2183, n_2184, n_2185);
  xor g1977 (n_2186, n_730, n_731);
  xor g1978 (n_198, n_2186, n_732);
  nand g1979 (n_2187, n_730, n_731);
  nand g1980 (n_2188, n_732, n_731);
  nand g1981 (n_2189, n_730, n_732);
  nand g1982 (n_111, n_2187, n_2188, n_2189);
  xor g1983 (n_2190, A[42], A[40]);
  xor g1984 (n_737, n_2190, A[36]);
  nand g1985 (n_2191, A[42], A[40]);
  nand g1986 (n_2192, A[36], A[40]);
  nand g1987 (n_2193, A[42], A[36]);
  nand g1988 (n_747, n_2191, n_2192, n_2193);
  xor g1990 (n_738, n_1742, A[34]);
  nand g1992 (n_2196, A[34], A[26]);
  nand g1994 (n_748, n_1743, n_2196, n_1937);
  xor g1995 (n_2198, A[24], A[38]);
  xor g1996 (n_736, n_2198, A[32]);
  nand g1997 (n_2199, A[24], A[38]);
  nand g2000 (n_749, n_2199, n_2065, n_2132);
  xor g2001 (n_2202, A[30], n_733);
  xor g2002 (n_740, n_2202, n_734);
  nand g2003 (n_2203, A[30], n_733);
  nand g2004 (n_2204, n_734, n_733);
  nand g2005 (n_2205, A[30], n_734);
  nand g2006 (n_753, n_2203, n_2204, n_2205);
  xor g2007 (n_2206, n_735, n_736);
  xor g2008 (n_742, n_2206, n_737);
  nand g2009 (n_2207, n_735, n_736);
  nand g2010 (n_2208, n_737, n_736);
  nand g2011 (n_2209, n_735, n_737);
  nand g2012 (n_755, n_2207, n_2208, n_2209);
  xor g2013 (n_2210, n_738, n_739);
  xor g2014 (n_744, n_2210, n_740);
  nand g2015 (n_2211, n_738, n_739);
  nand g2016 (n_2212, n_740, n_739);
  nand g2017 (n_2213, n_738, n_740);
  nand g2018 (n_757, n_2211, n_2212, n_2213);
  xor g2019 (n_2214, n_741, n_742);
  xor g2020 (n_745, n_2214, n_743);
  nand g2021 (n_2215, n_741, n_742);
  nand g2022 (n_2216, n_743, n_742);
  nand g2023 (n_2217, n_741, n_743);
  nand g2024 (n_760, n_2215, n_2216, n_2217);
  xor g2025 (n_2218, n_744, n_745);
  xor g2026 (n_197, n_2218, n_746);
  nand g2027 (n_2219, n_744, n_745);
  nand g2028 (n_2220, n_746, n_745);
  nand g2029 (n_2221, n_744, n_746);
  nand g2030 (n_110, n_2219, n_2220, n_2221);
  xor g2031 (n_2222, A[43], A[41]);
  xor g2032 (n_751, n_2222, A[37]);
  nand g2033 (n_2223, A[43], A[41]);
  nand g2034 (n_2224, A[37], A[41]);
  nand g2035 (n_2225, A[43], A[37]);
  nand g2036 (n_761, n_2223, n_2224, n_2225);
  xor g2038 (n_752, n_1774, A[35]);
  nand g2040 (n_2228, A[35], A[27]);
  nand g2042 (n_762, n_1775, n_2228, n_1969);
  xor g2043 (n_2230, A[25], A[39]);
  xor g2044 (n_750, n_2230, A[33]);
  nand g2045 (n_2231, A[25], A[39]);
  nand g2048 (n_763, n_2231, n_2097, n_2164);
  xor g2049 (n_2234, A[31], n_747);
  xor g2050 (n_754, n_2234, n_748);
  nand g2051 (n_2235, A[31], n_747);
  nand g2052 (n_2236, n_748, n_747);
  nand g2053 (n_2237, A[31], n_748);
  nand g2054 (n_767, n_2235, n_2236, n_2237);
  xor g2055 (n_2238, n_749, n_750);
  xor g2056 (n_756, n_2238, n_751);
  nand g2057 (n_2239, n_749, n_750);
  nand g2058 (n_2240, n_751, n_750);
  nand g2059 (n_2241, n_749, n_751);
  nand g2060 (n_769, n_2239, n_2240, n_2241);
  xor g2061 (n_2242, n_752, n_753);
  xor g2062 (n_758, n_2242, n_754);
  nand g2063 (n_2243, n_752, n_753);
  nand g2064 (n_2244, n_754, n_753);
  nand g2065 (n_2245, n_752, n_754);
  nand g2066 (n_771, n_2243, n_2244, n_2245);
  xor g2067 (n_2246, n_755, n_756);
  xor g2068 (n_759, n_2246, n_757);
  nand g2069 (n_2247, n_755, n_756);
  nand g2070 (n_2248, n_757, n_756);
  nand g2071 (n_2249, n_755, n_757);
  nand g2072 (n_774, n_2247, n_2248, n_2249);
  xor g2073 (n_2250, n_758, n_759);
  xor g2074 (n_196, n_2250, n_760);
  nand g2075 (n_2251, n_758, n_759);
  nand g2076 (n_2252, n_760, n_759);
  nand g2077 (n_2253, n_758, n_760);
  nand g2078 (n_109, n_2251, n_2252, n_2253);
  xor g2079 (n_2254, A[44], A[42]);
  xor g2080 (n_765, n_2254, A[38]);
  nand g2081 (n_2255, A[44], A[42]);
  nand g2082 (n_2256, A[38], A[42]);
  nand g2083 (n_2257, A[44], A[38]);
  nand g2084 (n_775, n_2255, n_2256, n_2257);
  xor g2086 (n_766, n_1806, A[36]);
  nand g2088 (n_2260, A[36], A[28]);
  nand g2090 (n_776, n_1807, n_2260, n_2001);
  xor g2091 (n_2262, A[26], A[40]);
  xor g2092 (n_764, n_2262, A[34]);
  nand g2093 (n_2263, A[26], A[40]);
  nand g2096 (n_777, n_2263, n_2129, n_2196);
  xor g2097 (n_2266, A[32], n_761);
  xor g2098 (n_768, n_2266, n_762);
  nand g2099 (n_2267, A[32], n_761);
  nand g2100 (n_2268, n_762, n_761);
  nand g2101 (n_2269, A[32], n_762);
  nand g2102 (n_781, n_2267, n_2268, n_2269);
  xor g2103 (n_2270, n_763, n_764);
  xor g2104 (n_770, n_2270, n_765);
  nand g2105 (n_2271, n_763, n_764);
  nand g2106 (n_2272, n_765, n_764);
  nand g2107 (n_2273, n_763, n_765);
  nand g2108 (n_783, n_2271, n_2272, n_2273);
  xor g2109 (n_2274, n_766, n_767);
  xor g2110 (n_772, n_2274, n_768);
  nand g2111 (n_2275, n_766, n_767);
  nand g2112 (n_2276, n_768, n_767);
  nand g2113 (n_2277, n_766, n_768);
  nand g2114 (n_785, n_2275, n_2276, n_2277);
  xor g2115 (n_2278, n_769, n_770);
  xor g2116 (n_773, n_2278, n_771);
  nand g2117 (n_2279, n_769, n_770);
  nand g2118 (n_2280, n_771, n_770);
  nand g2119 (n_2281, n_769, n_771);
  nand g2120 (n_788, n_2279, n_2280, n_2281);
  xor g2121 (n_2282, n_772, n_773);
  xor g2122 (n_195, n_2282, n_774);
  nand g2123 (n_2283, n_772, n_773);
  nand g2124 (n_2284, n_774, n_773);
  nand g2125 (n_2285, n_772, n_774);
  nand g2126 (n_108, n_2283, n_2284, n_2285);
  xor g2127 (n_2286, A[45], A[43]);
  xor g2128 (n_779, n_2286, A[39]);
  nand g2129 (n_2287, A[45], A[43]);
  nand g2130 (n_2288, A[39], A[43]);
  nand g2131 (n_2289, A[45], A[39]);
  nand g2132 (n_789, n_2287, n_2288, n_2289);
  xor g2134 (n_780, n_1838, A[37]);
  nand g2136 (n_2292, A[37], A[29]);
  nand g2138 (n_790, n_1839, n_2292, n_2033);
  xor g2139 (n_2294, A[27], A[41]);
  xor g2140 (n_778, n_2294, A[35]);
  nand g2141 (n_2295, A[27], A[41]);
  nand g2144 (n_791, n_2295, n_2161, n_2228);
  xor g2145 (n_2298, A[33], n_775);
  xor g2146 (n_782, n_2298, n_776);
  nand g2147 (n_2299, A[33], n_775);
  nand g2148 (n_2300, n_776, n_775);
  nand g2149 (n_2301, A[33], n_776);
  nand g2150 (n_795, n_2299, n_2300, n_2301);
  xor g2151 (n_2302, n_777, n_778);
  xor g2152 (n_784, n_2302, n_779);
  nand g2153 (n_2303, n_777, n_778);
  nand g2154 (n_2304, n_779, n_778);
  nand g2155 (n_2305, n_777, n_779);
  nand g2156 (n_797, n_2303, n_2304, n_2305);
  xor g2157 (n_2306, n_780, n_781);
  xor g2158 (n_786, n_2306, n_782);
  nand g2159 (n_2307, n_780, n_781);
  nand g2160 (n_2308, n_782, n_781);
  nand g2161 (n_2309, n_780, n_782);
  nand g2162 (n_799, n_2307, n_2308, n_2309);
  xor g2163 (n_2310, n_783, n_784);
  xor g2164 (n_787, n_2310, n_785);
  nand g2165 (n_2311, n_783, n_784);
  nand g2166 (n_2312, n_785, n_784);
  nand g2167 (n_2313, n_783, n_785);
  nand g2168 (n_802, n_2311, n_2312, n_2313);
  xor g2169 (n_2314, n_786, n_787);
  xor g2170 (n_194, n_2314, n_788);
  nand g2171 (n_2315, n_786, n_787);
  nand g2172 (n_2316, n_788, n_787);
  nand g2173 (n_2317, n_786, n_788);
  nand g2174 (n_107, n_2315, n_2316, n_2317);
  xor g2175 (n_2318, A[46], A[44]);
  xor g2176 (n_793, n_2318, A[40]);
  nand g2177 (n_2319, A[46], A[44]);
  nand g2178 (n_2320, A[40], A[44]);
  nand g2179 (n_2321, A[46], A[40]);
  nand g2180 (n_803, n_2319, n_2320, n_2321);
  xor g2182 (n_794, n_1870, A[38]);
  nand g2184 (n_2324, A[38], A[30]);
  nand g2186 (n_804, n_1871, n_2324, n_2065);
  xor g2187 (n_2326, A[28], A[42]);
  xor g2188 (n_792, n_2326, A[36]);
  nand g2189 (n_2327, A[28], A[42]);
  nand g2192 (n_805, n_2327, n_2193, n_2260);
  xor g2193 (n_2330, A[34], n_789);
  xor g2194 (n_796, n_2330, n_790);
  nand g2195 (n_2331, A[34], n_789);
  nand g2196 (n_2332, n_790, n_789);
  nand g2197 (n_2333, A[34], n_790);
  nand g2198 (n_809, n_2331, n_2332, n_2333);
  xor g2199 (n_2334, n_791, n_792);
  xor g2200 (n_798, n_2334, n_793);
  nand g2201 (n_2335, n_791, n_792);
  nand g2202 (n_2336, n_793, n_792);
  nand g2203 (n_2337, n_791, n_793);
  nand g2204 (n_811, n_2335, n_2336, n_2337);
  xor g2205 (n_2338, n_794, n_795);
  xor g2206 (n_800, n_2338, n_796);
  nand g2207 (n_2339, n_794, n_795);
  nand g2208 (n_2340, n_796, n_795);
  nand g2209 (n_2341, n_794, n_796);
  nand g2210 (n_813, n_2339, n_2340, n_2341);
  xor g2211 (n_2342, n_797, n_798);
  xor g2212 (n_801, n_2342, n_799);
  nand g2213 (n_2343, n_797, n_798);
  nand g2214 (n_2344, n_799, n_798);
  nand g2215 (n_2345, n_797, n_799);
  nand g2216 (n_816, n_2343, n_2344, n_2345);
  xor g2217 (n_2346, n_800, n_801);
  xor g2218 (n_193, n_2346, n_802);
  nand g2219 (n_2347, n_800, n_801);
  nand g2220 (n_2348, n_802, n_801);
  nand g2221 (n_2349, n_800, n_802);
  nand g2222 (n_106, n_2347, n_2348, n_2349);
  xor g2223 (n_2350, A[47], A[45]);
  xor g2224 (n_807, n_2350, A[41]);
  nand g2225 (n_2351, A[47], A[45]);
  nand g2226 (n_2352, A[41], A[45]);
  nand g2227 (n_2353, A[47], A[41]);
  nand g2228 (n_817, n_2351, n_2352, n_2353);
  xor g2230 (n_808, n_1902, A[39]);
  nand g2232 (n_2356, A[39], A[31]);
  nand g2234 (n_818, n_1903, n_2356, n_2097);
  xor g2235 (n_2358, A[29], A[43]);
  xor g2236 (n_806, n_2358, A[37]);
  nand g2237 (n_2359, A[29], A[43]);
  nand g2240 (n_819, n_2359, n_2225, n_2292);
  xor g2241 (n_2362, A[35], n_803);
  xor g2242 (n_810, n_2362, n_804);
  nand g2243 (n_2363, A[35], n_803);
  nand g2244 (n_2364, n_804, n_803);
  nand g2245 (n_2365, A[35], n_804);
  nand g2246 (n_823, n_2363, n_2364, n_2365);
  xor g2247 (n_2366, n_805, n_806);
  xor g2248 (n_812, n_2366, n_807);
  nand g2249 (n_2367, n_805, n_806);
  nand g2250 (n_2368, n_807, n_806);
  nand g2251 (n_2369, n_805, n_807);
  nand g2252 (n_825, n_2367, n_2368, n_2369);
  xor g2253 (n_2370, n_808, n_809);
  xor g2254 (n_814, n_2370, n_810);
  nand g2255 (n_2371, n_808, n_809);
  nand g2256 (n_2372, n_810, n_809);
  nand g2257 (n_2373, n_808, n_810);
  nand g2258 (n_827, n_2371, n_2372, n_2373);
  xor g2259 (n_2374, n_811, n_812);
  xor g2260 (n_815, n_2374, n_813);
  nand g2261 (n_2375, n_811, n_812);
  nand g2262 (n_2376, n_813, n_812);
  nand g2263 (n_2377, n_811, n_813);
  nand g2264 (n_830, n_2375, n_2376, n_2377);
  xor g2265 (n_2378, n_814, n_815);
  xor g2266 (n_192, n_2378, n_816);
  nand g2267 (n_2379, n_814, n_815);
  nand g2268 (n_2380, n_816, n_815);
  nand g2269 (n_2381, n_814, n_816);
  nand g2270 (n_105, n_2379, n_2380, n_2381);
  xor g2271 (n_2382, A[48], A[46]);
  xor g2272 (n_821, n_2382, A[42]);
  nand g2273 (n_2383, A[48], A[46]);
  nand g2274 (n_2384, A[42], A[46]);
  nand g2275 (n_2385, A[48], A[42]);
  nand g2276 (n_831, n_2383, n_2384, n_2385);
  xor g2278 (n_822, n_1934, A[40]);
  nand g2280 (n_2388, A[40], A[32]);
  nand g2282 (n_832, n_1935, n_2388, n_2129);
  xor g2283 (n_2390, A[30], A[44]);
  xor g2284 (n_820, n_2390, A[38]);
  nand g2285 (n_2391, A[30], A[44]);
  nand g2288 (n_833, n_2391, n_2257, n_2324);
  xor g2289 (n_2394, A[36], n_817);
  xor g2290 (n_824, n_2394, n_818);
  nand g2291 (n_2395, A[36], n_817);
  nand g2292 (n_2396, n_818, n_817);
  nand g2293 (n_2397, A[36], n_818);
  nand g2294 (n_837, n_2395, n_2396, n_2397);
  xor g2295 (n_2398, n_819, n_820);
  xor g2296 (n_826, n_2398, n_821);
  nand g2297 (n_2399, n_819, n_820);
  nand g2298 (n_2400, n_821, n_820);
  nand g2299 (n_2401, n_819, n_821);
  nand g2300 (n_839, n_2399, n_2400, n_2401);
  xor g2301 (n_2402, n_822, n_823);
  xor g2302 (n_828, n_2402, n_824);
  nand g2303 (n_2403, n_822, n_823);
  nand g2304 (n_2404, n_824, n_823);
  nand g2305 (n_2405, n_822, n_824);
  nand g2306 (n_841, n_2403, n_2404, n_2405);
  xor g2307 (n_2406, n_825, n_826);
  xor g2308 (n_829, n_2406, n_827);
  nand g2309 (n_2407, n_825, n_826);
  nand g2310 (n_2408, n_827, n_826);
  nand g2311 (n_2409, n_825, n_827);
  nand g2312 (n_844, n_2407, n_2408, n_2409);
  xor g2313 (n_2410, n_828, n_829);
  xor g2314 (n_191, n_2410, n_830);
  nand g2315 (n_2411, n_828, n_829);
  nand g2316 (n_2412, n_830, n_829);
  nand g2317 (n_2413, n_828, n_830);
  nand g2318 (n_104, n_2411, n_2412, n_2413);
  xor g2319 (n_2414, A[49], A[47]);
  xor g2320 (n_835, n_2414, A[43]);
  nand g2321 (n_2415, A[49], A[47]);
  nand g2322 (n_2416, A[43], A[47]);
  nand g2323 (n_2417, A[49], A[43]);
  nand g2324 (n_845, n_2415, n_2416, n_2417);
  xor g2326 (n_836, n_1966, A[41]);
  nand g2328 (n_2420, A[41], A[33]);
  nand g2330 (n_846, n_1967, n_2420, n_2161);
  xor g2331 (n_2422, A[31], A[45]);
  xor g2332 (n_834, n_2422, A[39]);
  nand g2333 (n_2423, A[31], A[45]);
  nand g2336 (n_847, n_2423, n_2289, n_2356);
  xor g2337 (n_2426, A[37], n_831);
  xor g2338 (n_838, n_2426, n_832);
  nand g2339 (n_2427, A[37], n_831);
  nand g2340 (n_2428, n_832, n_831);
  nand g2341 (n_2429, A[37], n_832);
  nand g2342 (n_851, n_2427, n_2428, n_2429);
  xor g2343 (n_2430, n_833, n_834);
  xor g2344 (n_840, n_2430, n_835);
  nand g2345 (n_2431, n_833, n_834);
  nand g2346 (n_2432, n_835, n_834);
  nand g2347 (n_2433, n_833, n_835);
  nand g2348 (n_853, n_2431, n_2432, n_2433);
  xor g2349 (n_2434, n_836, n_837);
  xor g2350 (n_842, n_2434, n_838);
  nand g2351 (n_2435, n_836, n_837);
  nand g2352 (n_2436, n_838, n_837);
  nand g2353 (n_2437, n_836, n_838);
  nand g2354 (n_855, n_2435, n_2436, n_2437);
  xor g2355 (n_2438, n_839, n_840);
  xor g2356 (n_843, n_2438, n_841);
  nand g2357 (n_2439, n_839, n_840);
  nand g2358 (n_2440, n_841, n_840);
  nand g2359 (n_2441, n_839, n_841);
  nand g2360 (n_858, n_2439, n_2440, n_2441);
  xor g2361 (n_2442, n_842, n_843);
  xor g2362 (n_190, n_2442, n_844);
  nand g2363 (n_2443, n_842, n_843);
  nand g2364 (n_2444, n_844, n_843);
  nand g2365 (n_2445, n_842, n_844);
  nand g2366 (n_103, n_2443, n_2444, n_2445);
  xor g2367 (n_2446, A[50], A[48]);
  xor g2368 (n_849, n_2446, A[44]);
  nand g2369 (n_2447, A[50], A[48]);
  nand g2370 (n_2448, A[44], A[48]);
  nand g2371 (n_2449, A[50], A[44]);
  nand g2372 (n_859, n_2447, n_2448, n_2449);
  xor g2374 (n_850, n_1998, A[42]);
  nand g2376 (n_2452, A[42], A[34]);
  nand g2378 (n_860, n_1999, n_2452, n_2193);
  xor g2379 (n_2454, A[32], A[46]);
  xor g2380 (n_848, n_2454, A[40]);
  nand g2381 (n_2455, A[32], A[46]);
  nand g2384 (n_861, n_2455, n_2321, n_2388);
  xor g2385 (n_2458, A[38], n_845);
  xor g2386 (n_852, n_2458, n_846);
  nand g2387 (n_2459, A[38], n_845);
  nand g2388 (n_2460, n_846, n_845);
  nand g2389 (n_2461, A[38], n_846);
  nand g2390 (n_865, n_2459, n_2460, n_2461);
  xor g2391 (n_2462, n_847, n_848);
  xor g2392 (n_854, n_2462, n_849);
  nand g2393 (n_2463, n_847, n_848);
  nand g2394 (n_2464, n_849, n_848);
  nand g2395 (n_2465, n_847, n_849);
  nand g2396 (n_867, n_2463, n_2464, n_2465);
  xor g2397 (n_2466, n_850, n_851);
  xor g2398 (n_856, n_2466, n_852);
  nand g2399 (n_2467, n_850, n_851);
  nand g2400 (n_2468, n_852, n_851);
  nand g2401 (n_2469, n_850, n_852);
  nand g2402 (n_869, n_2467, n_2468, n_2469);
  xor g2403 (n_2470, n_853, n_854);
  xor g2404 (n_857, n_2470, n_855);
  nand g2405 (n_2471, n_853, n_854);
  nand g2406 (n_2472, n_855, n_854);
  nand g2407 (n_2473, n_853, n_855);
  nand g2408 (n_872, n_2471, n_2472, n_2473);
  xor g2409 (n_2474, n_856, n_857);
  xor g2410 (n_189, n_2474, n_858);
  nand g2411 (n_2475, n_856, n_857);
  nand g2412 (n_2476, n_858, n_857);
  nand g2413 (n_2477, n_856, n_858);
  nand g2414 (n_102, n_2475, n_2476, n_2477);
  xor g2415 (n_2478, A[51], A[49]);
  xor g2416 (n_863, n_2478, A[45]);
  nand g2417 (n_2479, A[51], A[49]);
  nand g2418 (n_2480, A[45], A[49]);
  nand g2419 (n_2481, A[51], A[45]);
  nand g2420 (n_873, n_2479, n_2480, n_2481);
  xor g2422 (n_864, n_2030, A[43]);
  nand g2424 (n_2484, A[43], A[35]);
  nand g2426 (n_874, n_2031, n_2484, n_2225);
  xor g2427 (n_2486, A[33], A[47]);
  xor g2428 (n_862, n_2486, A[41]);
  nand g2429 (n_2487, A[33], A[47]);
  nand g2432 (n_875, n_2487, n_2353, n_2420);
  xor g2433 (n_2490, A[39], n_859);
  xor g2434 (n_866, n_2490, n_860);
  nand g2435 (n_2491, A[39], n_859);
  nand g2436 (n_2492, n_860, n_859);
  nand g2437 (n_2493, A[39], n_860);
  nand g2438 (n_879, n_2491, n_2492, n_2493);
  xor g2439 (n_2494, n_861, n_862);
  xor g2440 (n_868, n_2494, n_863);
  nand g2441 (n_2495, n_861, n_862);
  nand g2442 (n_2496, n_863, n_862);
  nand g2443 (n_2497, n_861, n_863);
  nand g2444 (n_881, n_2495, n_2496, n_2497);
  xor g2445 (n_2498, n_864, n_865);
  xor g2446 (n_870, n_2498, n_866);
  nand g2447 (n_2499, n_864, n_865);
  nand g2448 (n_2500, n_866, n_865);
  nand g2449 (n_2501, n_864, n_866);
  nand g2450 (n_883, n_2499, n_2500, n_2501);
  xor g2451 (n_2502, n_867, n_868);
  xor g2452 (n_871, n_2502, n_869);
  nand g2453 (n_2503, n_867, n_868);
  nand g2454 (n_2504, n_869, n_868);
  nand g2455 (n_2505, n_867, n_869);
  nand g2456 (n_886, n_2503, n_2504, n_2505);
  xor g2457 (n_2506, n_870, n_871);
  xor g2458 (n_188, n_2506, n_872);
  nand g2459 (n_2507, n_870, n_871);
  nand g2460 (n_2508, n_872, n_871);
  nand g2461 (n_2509, n_870, n_872);
  nand g2462 (n_101, n_2507, n_2508, n_2509);
  xor g2463 (n_2510, A[52], A[50]);
  xor g2464 (n_877, n_2510, A[46]);
  nand g2465 (n_2511, A[52], A[50]);
  nand g2466 (n_2512, A[46], A[50]);
  nand g2467 (n_2513, A[52], A[46]);
  nand g2468 (n_887, n_2511, n_2512, n_2513);
  xor g2470 (n_878, n_2062, A[44]);
  nand g2472 (n_2516, A[44], A[36]);
  nand g2474 (n_888, n_2063, n_2516, n_2257);
  xor g2475 (n_2518, A[34], A[48]);
  xor g2476 (n_876, n_2518, A[42]);
  nand g2477 (n_2519, A[34], A[48]);
  nand g2480 (n_889, n_2519, n_2385, n_2452);
  xor g2481 (n_2522, A[40], n_873);
  xor g2482 (n_880, n_2522, n_874);
  nand g2483 (n_2523, A[40], n_873);
  nand g2484 (n_2524, n_874, n_873);
  nand g2485 (n_2525, A[40], n_874);
  nand g2486 (n_893, n_2523, n_2524, n_2525);
  xor g2487 (n_2526, n_875, n_876);
  xor g2488 (n_882, n_2526, n_877);
  nand g2489 (n_2527, n_875, n_876);
  nand g2490 (n_2528, n_877, n_876);
  nand g2491 (n_2529, n_875, n_877);
  nand g2492 (n_895, n_2527, n_2528, n_2529);
  xor g2493 (n_2530, n_878, n_879);
  xor g2494 (n_884, n_2530, n_880);
  nand g2495 (n_2531, n_878, n_879);
  nand g2496 (n_2532, n_880, n_879);
  nand g2497 (n_2533, n_878, n_880);
  nand g2498 (n_897, n_2531, n_2532, n_2533);
  xor g2499 (n_2534, n_881, n_882);
  xor g2500 (n_885, n_2534, n_883);
  nand g2501 (n_2535, n_881, n_882);
  nand g2502 (n_2536, n_883, n_882);
  nand g2503 (n_2537, n_881, n_883);
  nand g2504 (n_900, n_2535, n_2536, n_2537);
  xor g2505 (n_2538, n_884, n_885);
  xor g2506 (n_187, n_2538, n_886);
  nand g2507 (n_2539, n_884, n_885);
  nand g2508 (n_2540, n_886, n_885);
  nand g2509 (n_2541, n_884, n_886);
  nand g2510 (n_100, n_2539, n_2540, n_2541);
  xor g2511 (n_2542, A[53], A[51]);
  xor g2512 (n_891, n_2542, A[47]);
  nand g2513 (n_2543, A[53], A[51]);
  nand g2514 (n_2544, A[47], A[51]);
  nand g2515 (n_2545, A[53], A[47]);
  nand g2516 (n_901, n_2543, n_2544, n_2545);
  xor g2518 (n_892, n_2094, A[45]);
  nand g2520 (n_2548, A[45], A[37]);
  nand g2522 (n_902, n_2095, n_2548, n_2289);
  xor g2523 (n_2550, A[35], A[49]);
  xor g2524 (n_890, n_2550, A[43]);
  nand g2525 (n_2551, A[35], A[49]);
  nand g2528 (n_903, n_2551, n_2417, n_2484);
  xor g2529 (n_2554, A[41], n_887);
  xor g2530 (n_894, n_2554, n_888);
  nand g2531 (n_2555, A[41], n_887);
  nand g2532 (n_2556, n_888, n_887);
  nand g2533 (n_2557, A[41], n_888);
  nand g2534 (n_907, n_2555, n_2556, n_2557);
  xor g2535 (n_2558, n_889, n_890);
  xor g2536 (n_896, n_2558, n_891);
  nand g2537 (n_2559, n_889, n_890);
  nand g2538 (n_2560, n_891, n_890);
  nand g2539 (n_2561, n_889, n_891);
  nand g2540 (n_909, n_2559, n_2560, n_2561);
  xor g2541 (n_2562, n_892, n_893);
  xor g2542 (n_898, n_2562, n_894);
  nand g2543 (n_2563, n_892, n_893);
  nand g2544 (n_2564, n_894, n_893);
  nand g2545 (n_2565, n_892, n_894);
  nand g2546 (n_911, n_2563, n_2564, n_2565);
  xor g2547 (n_2566, n_895, n_896);
  xor g2548 (n_899, n_2566, n_897);
  nand g2549 (n_2567, n_895, n_896);
  nand g2550 (n_2568, n_897, n_896);
  nand g2551 (n_2569, n_895, n_897);
  nand g2552 (n_914, n_2567, n_2568, n_2569);
  xor g2553 (n_2570, n_898, n_899);
  xor g2554 (n_186, n_2570, n_900);
  nand g2555 (n_2571, n_898, n_899);
  nand g2556 (n_2572, n_900, n_899);
  nand g2557 (n_2573, n_898, n_900);
  nand g2558 (n_99, n_2571, n_2572, n_2573);
  xor g2559 (n_2574, A[54], A[52]);
  xor g2560 (n_905, n_2574, A[48]);
  nand g2561 (n_2575, A[54], A[52]);
  nand g2562 (n_2576, A[48], A[52]);
  nand g2563 (n_2577, A[54], A[48]);
  nand g2564 (n_915, n_2575, n_2576, n_2577);
  xor g2566 (n_906, n_2126, A[46]);
  nand g2568 (n_2580, A[46], A[38]);
  nand g2570 (n_916, n_2127, n_2580, n_2321);
  xor g2571 (n_2582, A[36], A[50]);
  xor g2572 (n_904, n_2582, A[44]);
  nand g2573 (n_2583, A[36], A[50]);
  nand g2576 (n_917, n_2583, n_2449, n_2516);
  xor g2577 (n_2586, A[42], n_901);
  xor g2578 (n_908, n_2586, n_902);
  nand g2579 (n_2587, A[42], n_901);
  nand g2580 (n_2588, n_902, n_901);
  nand g2581 (n_2589, A[42], n_902);
  nand g2582 (n_921, n_2587, n_2588, n_2589);
  xor g2583 (n_2590, n_903, n_904);
  xor g2584 (n_910, n_2590, n_905);
  nand g2585 (n_2591, n_903, n_904);
  nand g2586 (n_2592, n_905, n_904);
  nand g2587 (n_2593, n_903, n_905);
  nand g2588 (n_923, n_2591, n_2592, n_2593);
  xor g2589 (n_2594, n_906, n_907);
  xor g2590 (n_912, n_2594, n_908);
  nand g2591 (n_2595, n_906, n_907);
  nand g2592 (n_2596, n_908, n_907);
  nand g2593 (n_2597, n_906, n_908);
  nand g2594 (n_925, n_2595, n_2596, n_2597);
  xor g2595 (n_2598, n_909, n_910);
  xor g2596 (n_913, n_2598, n_911);
  nand g2597 (n_2599, n_909, n_910);
  nand g2598 (n_2600, n_911, n_910);
  nand g2599 (n_2601, n_909, n_911);
  nand g2600 (n_928, n_2599, n_2600, n_2601);
  xor g2601 (n_2602, n_912, n_913);
  xor g2602 (n_185, n_2602, n_914);
  nand g2603 (n_2603, n_912, n_913);
  nand g2604 (n_2604, n_914, n_913);
  nand g2605 (n_2605, n_912, n_914);
  nand g2606 (n_98, n_2603, n_2604, n_2605);
  xor g2607 (n_2606, A[55], A[53]);
  xor g2608 (n_919, n_2606, A[49]);
  nand g2609 (n_2607, A[55], A[53]);
  nand g2610 (n_2608, A[49], A[53]);
  nand g2611 (n_2609, A[55], A[49]);
  nand g2612 (n_929, n_2607, n_2608, n_2609);
  xor g2614 (n_920, n_2158, A[47]);
  nand g2616 (n_2612, A[47], A[39]);
  nand g2618 (n_930, n_2159, n_2612, n_2353);
  xor g2619 (n_2614, A[37], A[51]);
  xor g2620 (n_918, n_2614, A[45]);
  nand g2621 (n_2615, A[37], A[51]);
  nand g2624 (n_931, n_2615, n_2481, n_2548);
  xor g2625 (n_2618, A[43], n_915);
  xor g2626 (n_922, n_2618, n_916);
  nand g2627 (n_2619, A[43], n_915);
  nand g2628 (n_2620, n_916, n_915);
  nand g2629 (n_2621, A[43], n_916);
  nand g2630 (n_935, n_2619, n_2620, n_2621);
  xor g2631 (n_2622, n_917, n_918);
  xor g2632 (n_924, n_2622, n_919);
  nand g2633 (n_2623, n_917, n_918);
  nand g2634 (n_2624, n_919, n_918);
  nand g2635 (n_2625, n_917, n_919);
  nand g2636 (n_937, n_2623, n_2624, n_2625);
  xor g2637 (n_2626, n_920, n_921);
  xor g2638 (n_926, n_2626, n_922);
  nand g2639 (n_2627, n_920, n_921);
  nand g2640 (n_2628, n_922, n_921);
  nand g2641 (n_2629, n_920, n_922);
  nand g2642 (n_939, n_2627, n_2628, n_2629);
  xor g2643 (n_2630, n_923, n_924);
  xor g2644 (n_927, n_2630, n_925);
  nand g2645 (n_2631, n_923, n_924);
  nand g2646 (n_2632, n_925, n_924);
  nand g2647 (n_2633, n_923, n_925);
  nand g2648 (n_942, n_2631, n_2632, n_2633);
  xor g2649 (n_2634, n_926, n_927);
  xor g2650 (n_184, n_2634, n_928);
  nand g2651 (n_2635, n_926, n_927);
  nand g2652 (n_2636, n_928, n_927);
  nand g2653 (n_2637, n_926, n_928);
  nand g2654 (n_97, n_2635, n_2636, n_2637);
  xor g2655 (n_2638, A[56], A[54]);
  xor g2656 (n_933, n_2638, A[50]);
  nand g2657 (n_2639, A[56], A[54]);
  nand g2658 (n_2640, A[50], A[54]);
  nand g2659 (n_2641, A[56], A[50]);
  nand g2660 (n_943, n_2639, n_2640, n_2641);
  xor g2662 (n_934, n_2190, A[48]);
  nand g2664 (n_2644, A[48], A[40]);
  nand g2666 (n_944, n_2191, n_2644, n_2385);
  xor g2667 (n_2646, A[38], A[52]);
  xor g2668 (n_932, n_2646, A[46]);
  nand g2669 (n_2647, A[38], A[52]);
  nand g2672 (n_945, n_2647, n_2513, n_2580);
  xor g2673 (n_2650, A[44], n_929);
  xor g2674 (n_936, n_2650, n_930);
  nand g2675 (n_2651, A[44], n_929);
  nand g2676 (n_2652, n_930, n_929);
  nand g2677 (n_2653, A[44], n_930);
  nand g2678 (n_949, n_2651, n_2652, n_2653);
  xor g2679 (n_2654, n_931, n_932);
  xor g2680 (n_938, n_2654, n_933);
  nand g2681 (n_2655, n_931, n_932);
  nand g2682 (n_2656, n_933, n_932);
  nand g2683 (n_2657, n_931, n_933);
  nand g2684 (n_951, n_2655, n_2656, n_2657);
  xor g2685 (n_2658, n_934, n_935);
  xor g2686 (n_940, n_2658, n_936);
  nand g2687 (n_2659, n_934, n_935);
  nand g2688 (n_2660, n_936, n_935);
  nand g2689 (n_2661, n_934, n_936);
  nand g2690 (n_953, n_2659, n_2660, n_2661);
  xor g2691 (n_2662, n_937, n_938);
  xor g2692 (n_941, n_2662, n_939);
  nand g2693 (n_2663, n_937, n_938);
  nand g2694 (n_2664, n_939, n_938);
  nand g2695 (n_2665, n_937, n_939);
  nand g2696 (n_956, n_2663, n_2664, n_2665);
  xor g2697 (n_2666, n_940, n_941);
  xor g2698 (n_183, n_2666, n_942);
  nand g2699 (n_2667, n_940, n_941);
  nand g2700 (n_2668, n_942, n_941);
  nand g2701 (n_2669, n_940, n_942);
  nand g2702 (n_96, n_2667, n_2668, n_2669);
  xor g2703 (n_2670, A[57], A[55]);
  xor g2704 (n_947, n_2670, A[51]);
  nand g2705 (n_2671, A[57], A[55]);
  nand g2706 (n_2672, A[51], A[55]);
  nand g2707 (n_2673, A[57], A[51]);
  nand g2708 (n_957, n_2671, n_2672, n_2673);
  xor g2710 (n_948, n_2222, A[49]);
  nand g2712 (n_2676, A[49], A[41]);
  nand g2714 (n_958, n_2223, n_2676, n_2417);
  xor g2715 (n_2678, A[39], A[53]);
  xor g2716 (n_946, n_2678, A[47]);
  nand g2717 (n_2679, A[39], A[53]);
  nand g2720 (n_959, n_2679, n_2545, n_2612);
  xor g2721 (n_2682, A[45], n_943);
  xor g2722 (n_950, n_2682, n_944);
  nand g2723 (n_2683, A[45], n_943);
  nand g2724 (n_2684, n_944, n_943);
  nand g2725 (n_2685, A[45], n_944);
  nand g2726 (n_963, n_2683, n_2684, n_2685);
  xor g2727 (n_2686, n_945, n_946);
  xor g2728 (n_952, n_2686, n_947);
  nand g2729 (n_2687, n_945, n_946);
  nand g2730 (n_2688, n_947, n_946);
  nand g2731 (n_2689, n_945, n_947);
  nand g2732 (n_965, n_2687, n_2688, n_2689);
  xor g2733 (n_2690, n_948, n_949);
  xor g2734 (n_954, n_2690, n_950);
  nand g2735 (n_2691, n_948, n_949);
  nand g2736 (n_2692, n_950, n_949);
  nand g2737 (n_2693, n_948, n_950);
  nand g2738 (n_967, n_2691, n_2692, n_2693);
  xor g2739 (n_2694, n_951, n_952);
  xor g2740 (n_955, n_2694, n_953);
  nand g2741 (n_2695, n_951, n_952);
  nand g2742 (n_2696, n_953, n_952);
  nand g2743 (n_2697, n_951, n_953);
  nand g2744 (n_970, n_2695, n_2696, n_2697);
  xor g2745 (n_2698, n_954, n_955);
  xor g2746 (n_182, n_2698, n_956);
  nand g2747 (n_2699, n_954, n_955);
  nand g2748 (n_2700, n_956, n_955);
  nand g2749 (n_2701, n_954, n_956);
  nand g2750 (n_95, n_2699, n_2700, n_2701);
  xor g2751 (n_2702, A[58], A[56]);
  xor g2752 (n_961, n_2702, A[52]);
  nand g2753 (n_2703, A[58], A[56]);
  nand g2754 (n_2704, A[52], A[56]);
  nand g2755 (n_2705, A[58], A[52]);
  nand g2756 (n_971, n_2703, n_2704, n_2705);
  xor g2758 (n_962, n_2254, A[50]);
  nand g2760 (n_2708, A[50], A[42]);
  nand g2762 (n_972, n_2255, n_2708, n_2449);
  xor g2763 (n_2710, A[40], A[54]);
  xor g2764 (n_960, n_2710, A[48]);
  nand g2765 (n_2711, A[40], A[54]);
  nand g2768 (n_973, n_2711, n_2577, n_2644);
  xor g2769 (n_2714, A[46], n_957);
  xor g2770 (n_964, n_2714, n_958);
  nand g2771 (n_2715, A[46], n_957);
  nand g2772 (n_2716, n_958, n_957);
  nand g2773 (n_2717, A[46], n_958);
  nand g2774 (n_977, n_2715, n_2716, n_2717);
  xor g2775 (n_2718, n_959, n_960);
  xor g2776 (n_966, n_2718, n_961);
  nand g2777 (n_2719, n_959, n_960);
  nand g2778 (n_2720, n_961, n_960);
  nand g2779 (n_2721, n_959, n_961);
  nand g2780 (n_979, n_2719, n_2720, n_2721);
  xor g2781 (n_2722, n_962, n_963);
  xor g2782 (n_968, n_2722, n_964);
  nand g2783 (n_2723, n_962, n_963);
  nand g2784 (n_2724, n_964, n_963);
  nand g2785 (n_2725, n_962, n_964);
  nand g2786 (n_981, n_2723, n_2724, n_2725);
  xor g2787 (n_2726, n_965, n_966);
  xor g2788 (n_969, n_2726, n_967);
  nand g2789 (n_2727, n_965, n_966);
  nand g2790 (n_2728, n_967, n_966);
  nand g2791 (n_2729, n_965, n_967);
  nand g2792 (n_984, n_2727, n_2728, n_2729);
  xor g2793 (n_2730, n_968, n_969);
  xor g2794 (n_181, n_2730, n_970);
  nand g2795 (n_2731, n_968, n_969);
  nand g2796 (n_2732, n_970, n_969);
  nand g2797 (n_2733, n_968, n_970);
  nand g2798 (n_94, n_2731, n_2732, n_2733);
  xor g2799 (n_2734, A[59], A[57]);
  xor g2800 (n_975, n_2734, A[53]);
  nand g2801 (n_2735, A[59], A[57]);
  nand g2802 (n_2736, A[53], A[57]);
  nand g2803 (n_2737, A[59], A[53]);
  nand g2804 (n_985, n_2735, n_2736, n_2737);
  xor g2806 (n_976, n_2286, A[51]);
  nand g2808 (n_2740, A[51], A[43]);
  nand g2810 (n_986, n_2287, n_2740, n_2481);
  xor g2811 (n_2742, A[41], A[55]);
  xor g2812 (n_974, n_2742, A[49]);
  nand g2813 (n_2743, A[41], A[55]);
  nand g2816 (n_987, n_2743, n_2609, n_2676);
  xor g2817 (n_2746, A[47], n_971);
  xor g2818 (n_978, n_2746, n_972);
  nand g2819 (n_2747, A[47], n_971);
  nand g2820 (n_2748, n_972, n_971);
  nand g2821 (n_2749, A[47], n_972);
  nand g2822 (n_991, n_2747, n_2748, n_2749);
  xor g2823 (n_2750, n_973, n_974);
  xor g2824 (n_980, n_2750, n_975);
  nand g2825 (n_2751, n_973, n_974);
  nand g2826 (n_2752, n_975, n_974);
  nand g2827 (n_2753, n_973, n_975);
  nand g2828 (n_993, n_2751, n_2752, n_2753);
  xor g2829 (n_2754, n_976, n_977);
  xor g2830 (n_982, n_2754, n_978);
  nand g2831 (n_2755, n_976, n_977);
  nand g2832 (n_2756, n_978, n_977);
  nand g2833 (n_2757, n_976, n_978);
  nand g2834 (n_995, n_2755, n_2756, n_2757);
  xor g2835 (n_2758, n_979, n_980);
  xor g2836 (n_983, n_2758, n_981);
  nand g2837 (n_2759, n_979, n_980);
  nand g2838 (n_2760, n_981, n_980);
  nand g2839 (n_2761, n_979, n_981);
  nand g2840 (n_998, n_2759, n_2760, n_2761);
  xor g2841 (n_2762, n_982, n_983);
  xor g2842 (n_180, n_2762, n_984);
  nand g2843 (n_2763, n_982, n_983);
  nand g2844 (n_2764, n_984, n_983);
  nand g2845 (n_2765, n_982, n_984);
  nand g2846 (n_93, n_2763, n_2764, n_2765);
  xor g2847 (n_2766, A[60], A[58]);
  xor g2848 (n_989, n_2766, A[54]);
  nand g2849 (n_2767, A[60], A[58]);
  nand g2850 (n_2768, A[54], A[58]);
  nand g2851 (n_2769, A[60], A[54]);
  nand g2852 (n_999, n_2767, n_2768, n_2769);
  xor g2854 (n_990, n_2318, A[52]);
  nand g2856 (n_2772, A[52], A[44]);
  nand g2858 (n_1000, n_2319, n_2772, n_2513);
  xor g2859 (n_2774, A[42], A[56]);
  xor g2860 (n_988, n_2774, A[50]);
  nand g2861 (n_2775, A[42], A[56]);
  nand g2864 (n_1001, n_2775, n_2641, n_2708);
  xor g2865 (n_2778, A[48], n_985);
  xor g2866 (n_992, n_2778, n_986);
  nand g2867 (n_2779, A[48], n_985);
  nand g2868 (n_2780, n_986, n_985);
  nand g2869 (n_2781, A[48], n_986);
  nand g2870 (n_1005, n_2779, n_2780, n_2781);
  xor g2871 (n_2782, n_987, n_988);
  xor g2872 (n_994, n_2782, n_989);
  nand g2873 (n_2783, n_987, n_988);
  nand g2874 (n_2784, n_989, n_988);
  nand g2875 (n_2785, n_987, n_989);
  nand g2876 (n_1007, n_2783, n_2784, n_2785);
  xor g2877 (n_2786, n_990, n_991);
  xor g2878 (n_996, n_2786, n_992);
  nand g2879 (n_2787, n_990, n_991);
  nand g2880 (n_2788, n_992, n_991);
  nand g2881 (n_2789, n_990, n_992);
  nand g2882 (n_1009, n_2787, n_2788, n_2789);
  xor g2883 (n_2790, n_993, n_994);
  xor g2884 (n_997, n_2790, n_995);
  nand g2885 (n_2791, n_993, n_994);
  nand g2886 (n_2792, n_995, n_994);
  nand g2887 (n_2793, n_993, n_995);
  nand g2888 (n_1012, n_2791, n_2792, n_2793);
  xor g2889 (n_2794, n_996, n_997);
  xor g2890 (n_179, n_2794, n_998);
  nand g2891 (n_2795, n_996, n_997);
  nand g2892 (n_2796, n_998, n_997);
  nand g2893 (n_2797, n_996, n_998);
  nand g2894 (n_92, n_2795, n_2796, n_2797);
  xor g2895 (n_2798, A[61], A[59]);
  xor g2896 (n_1003, n_2798, A[55]);
  nand g2897 (n_2799, A[61], A[59]);
  nand g2898 (n_2800, A[55], A[59]);
  nand g2899 (n_2801, A[61], A[55]);
  nand g2900 (n_1013, n_2799, n_2800, n_2801);
  xor g2902 (n_1004, n_2350, A[53]);
  nand g2904 (n_2804, A[53], A[45]);
  nand g2906 (n_1014, n_2351, n_2804, n_2545);
  xor g2907 (n_2806, A[43], A[57]);
  xor g2908 (n_1002, n_2806, A[51]);
  nand g2909 (n_2807, A[43], A[57]);
  nand g2912 (n_1015, n_2807, n_2673, n_2740);
  xor g2913 (n_2810, A[49], n_999);
  xor g2914 (n_1006, n_2810, n_1000);
  nand g2915 (n_2811, A[49], n_999);
  nand g2916 (n_2812, n_1000, n_999);
  nand g2917 (n_2813, A[49], n_1000);
  nand g2918 (n_1019, n_2811, n_2812, n_2813);
  xor g2919 (n_2814, n_1001, n_1002);
  xor g2920 (n_1008, n_2814, n_1003);
  nand g2921 (n_2815, n_1001, n_1002);
  nand g2922 (n_2816, n_1003, n_1002);
  nand g2923 (n_2817, n_1001, n_1003);
  nand g2924 (n_1021, n_2815, n_2816, n_2817);
  xor g2925 (n_2818, n_1004, n_1005);
  xor g2926 (n_1010, n_2818, n_1006);
  nand g2927 (n_2819, n_1004, n_1005);
  nand g2928 (n_2820, n_1006, n_1005);
  nand g2929 (n_2821, n_1004, n_1006);
  nand g2930 (n_1023, n_2819, n_2820, n_2821);
  xor g2931 (n_2822, n_1007, n_1008);
  xor g2932 (n_1011, n_2822, n_1009);
  nand g2933 (n_2823, n_1007, n_1008);
  nand g2934 (n_2824, n_1009, n_1008);
  nand g2935 (n_2825, n_1007, n_1009);
  nand g2936 (n_1026, n_2823, n_2824, n_2825);
  xor g2937 (n_2826, n_1010, n_1011);
  xor g2938 (n_178, n_2826, n_1012);
  nand g2939 (n_2827, n_1010, n_1011);
  nand g2940 (n_2828, n_1012, n_1011);
  nand g2941 (n_2829, n_1010, n_1012);
  nand g2942 (n_91, n_2827, n_2828, n_2829);
  xor g2943 (n_2830, A[62], A[60]);
  xor g2944 (n_1017, n_2830, A[56]);
  nand g2945 (n_2831, A[62], A[60]);
  nand g2946 (n_2832, A[56], A[60]);
  nand g2947 (n_2833, A[62], A[56]);
  nand g2948 (n_1027, n_2831, n_2832, n_2833);
  xor g2950 (n_1018, n_2382, A[54]);
  nand g2952 (n_2836, A[54], A[46]);
  nand g2954 (n_1028, n_2383, n_2836, n_2577);
  xor g2955 (n_2838, A[44], A[58]);
  xor g2956 (n_1016, n_2838, A[52]);
  nand g2957 (n_2839, A[44], A[58]);
  nand g2960 (n_1029, n_2839, n_2705, n_2772);
  xor g2961 (n_2842, A[50], n_1013);
  xor g2962 (n_1020, n_2842, n_1014);
  nand g2963 (n_2843, A[50], n_1013);
  nand g2964 (n_2844, n_1014, n_1013);
  nand g2965 (n_2845, A[50], n_1014);
  nand g2966 (n_1033, n_2843, n_2844, n_2845);
  xor g2967 (n_2846, n_1015, n_1016);
  xor g2968 (n_1022, n_2846, n_1017);
  nand g2969 (n_2847, n_1015, n_1016);
  nand g2970 (n_2848, n_1017, n_1016);
  nand g2971 (n_2849, n_1015, n_1017);
  nand g2972 (n_1035, n_2847, n_2848, n_2849);
  xor g2973 (n_2850, n_1018, n_1019);
  xor g2974 (n_1024, n_2850, n_1020);
  nand g2975 (n_2851, n_1018, n_1019);
  nand g2976 (n_2852, n_1020, n_1019);
  nand g2977 (n_2853, n_1018, n_1020);
  nand g2978 (n_1037, n_2851, n_2852, n_2853);
  xor g2979 (n_2854, n_1021, n_1022);
  xor g2980 (n_1025, n_2854, n_1023);
  nand g2981 (n_2855, n_1021, n_1022);
  nand g2982 (n_2856, n_1023, n_1022);
  nand g2983 (n_2857, n_1021, n_1023);
  nand g2984 (n_1040, n_2855, n_2856, n_2857);
  xor g2985 (n_2858, n_1024, n_1025);
  xor g2986 (n_177, n_2858, n_1026);
  nand g2987 (n_2859, n_1024, n_1025);
  nand g2988 (n_2860, n_1026, n_1025);
  nand g2989 (n_2861, n_1024, n_1026);
  nand g2990 (n_90, n_2859, n_2860, n_2861);
  xor g2991 (n_2862, A[63], A[61]);
  xor g2992 (n_1031, n_2862, A[57]);
  nand g2993 (n_2863, A[63], A[61]);
  nand g2994 (n_2864, A[57], A[61]);
  nand g2995 (n_2865, A[63], A[57]);
  nand g2996 (n_1041, n_2863, n_2864, n_2865);
  xor g2998 (n_1032, n_2414, A[55]);
  nand g3000 (n_2868, A[55], A[47]);
  nand g3002 (n_1043, n_2415, n_2868, n_2609);
  xor g3003 (n_2870, A[45], A[59]);
  xor g3004 (n_1030, n_2870, A[53]);
  nand g3005 (n_2871, A[45], A[59]);
  nand g3008 (n_1042, n_2871, n_2737, n_2804);
  xor g3009 (n_2874, A[51], n_1027);
  xor g3010 (n_1034, n_2874, n_1028);
  nand g3011 (n_2875, A[51], n_1027);
  nand g3012 (n_2876, n_1028, n_1027);
  nand g3013 (n_2877, A[51], n_1028);
  nand g3014 (n_1047, n_2875, n_2876, n_2877);
  xor g3015 (n_2878, n_1029, n_1030);
  xor g3016 (n_1036, n_2878, n_1031);
  nand g3017 (n_2879, n_1029, n_1030);
  nand g3018 (n_2880, n_1031, n_1030);
  nand g3019 (n_2881, n_1029, n_1031);
  nand g3020 (n_1049, n_2879, n_2880, n_2881);
  xor g3021 (n_2882, n_1032, n_1033);
  xor g3022 (n_1038, n_2882, n_1034);
  nand g3023 (n_2883, n_1032, n_1033);
  nand g3024 (n_2884, n_1034, n_1033);
  nand g3025 (n_2885, n_1032, n_1034);
  nand g3026 (n_1052, n_2883, n_2884, n_2885);
  xor g3027 (n_2886, n_1035, n_1036);
  xor g3028 (n_1039, n_2886, n_1037);
  nand g3029 (n_2887, n_1035, n_1036);
  nand g3030 (n_2888, n_1037, n_1036);
  nand g3031 (n_2889, n_1035, n_1037);
  nand g3032 (n_1054, n_2887, n_2888, n_2889);
  xor g3033 (n_2890, n_1038, n_1039);
  xor g3034 (n_176, n_2890, n_1040);
  nand g3035 (n_2891, n_1038, n_1039);
  nand g3036 (n_2892, n_1040, n_1039);
  nand g3037 (n_2893, n_1038, n_1040);
  nand g3038 (n_89, n_2891, n_2892, n_2893);
  xor g3039 (n_2894, A[62], A[58]);
  xor g3040 (n_1045, n_2894, A[50]);
  nand g3041 (n_2895, A[62], A[58]);
  nand g3042 (n_2896, A[50], A[58]);
  nand g3043 (n_2897, A[62], A[50]);
  nand g3044 (n_1055, n_2895, n_2896, n_2897);
  xor g3045 (n_2898, A[48], A[56]);
  xor g3046 (n_1046, n_2898, A[46]);
  nand g3047 (n_2899, A[48], A[56]);
  nand g3048 (n_2900, A[46], A[56]);
  nand g3050 (n_1057, n_2899, n_2900, n_2383);
  xor g3051 (n_2902, A[60], A[54]);
  xor g3052 (n_1044, n_2902, A[52]);
  nand g3055 (n_2905, A[60], A[52]);
  nand g3056 (n_1056, n_2769, n_2575, n_2905);
  xor g3057 (n_2906, A[64], n_1041);
  xor g3058 (n_1048, n_2906, n_1042);
  nand g3059 (n_2907, A[64], n_1041);
  nand g3060 (n_2908, n_1042, n_1041);
  nand g3061 (n_2909, A[64], n_1042);
  nand g3062 (n_1061, n_2907, n_2908, n_2909);
  xor g3063 (n_2910, n_1043, n_1044);
  xor g3064 (n_1050, n_2910, n_1045);
  nand g3065 (n_2911, n_1043, n_1044);
  nand g3066 (n_2912, n_1045, n_1044);
  nand g3067 (n_2913, n_1043, n_1045);
  nand g3068 (n_1063, n_2911, n_2912, n_2913);
  xor g3069 (n_2914, n_1046, n_1047);
  xor g3070 (n_1051, n_2914, n_1048);
  nand g3071 (n_2915, n_1046, n_1047);
  nand g3072 (n_2916, n_1048, n_1047);
  nand g3073 (n_2917, n_1046, n_1048);
  nand g3074 (n_1066, n_2915, n_2916, n_2917);
  xor g3075 (n_2918, n_1049, n_1050);
  xor g3076 (n_1053, n_2918, n_1051);
  nand g3077 (n_2919, n_1049, n_1050);
  nand g3078 (n_2920, n_1051, n_1050);
  nand g3079 (n_2921, n_1049, n_1051);
  nand g3080 (n_1068, n_2919, n_2920, n_2921);
  xor g3081 (n_2922, n_1052, n_1053);
  xor g3082 (n_175, n_2922, n_1054);
  nand g3083 (n_2923, n_1052, n_1053);
  nand g3084 (n_2924, n_1054, n_1053);
  nand g3085 (n_2925, n_1052, n_1054);
  nand g3086 (n_88, n_2923, n_2924, n_2925);
  xor g3087 (n_2926, A[63], A[59]);
  xor g3088 (n_1059, n_2926, A[51]);
  nand g3089 (n_2927, A[63], A[59]);
  nand g3090 (n_2928, A[51], A[59]);
  nand g3091 (n_2929, A[63], A[51]);
  nand g3092 (n_1071, n_2927, n_2928, n_2929);
  xor g3093 (n_2930, A[49], A[57]);
  xor g3094 (n_1060, n_2930, A[47]);
  nand g3095 (n_2931, A[49], A[57]);
  nand g3096 (n_2932, A[47], A[57]);
  nand g3098 (n_1072, n_2931, n_2932, n_2415);
  xor g3099 (n_2934, A[61], A[55]);
  xor g3100 (n_1058, n_2934, A[53]);
  nand g3103 (n_2937, A[61], A[53]);
  nand g3104 (n_1073, n_2801, n_2607, n_2937);
  xor g3105 (n_2938, A[65], n_1055);
  xor g3106 (n_1062, n_2938, n_1056);
  nand g3107 (n_2939, A[65], n_1055);
  nand g3108 (n_2940, n_1056, n_1055);
  nand g3109 (n_2941, A[65], n_1056);
  nand g3110 (n_1077, n_2939, n_2940, n_2941);
  xor g3111 (n_2942, n_1057, n_1058);
  xor g3112 (n_1064, n_2942, n_1059);
  nand g3113 (n_2943, n_1057, n_1058);
  nand g3114 (n_2944, n_1059, n_1058);
  nand g3115 (n_2945, n_1057, n_1059);
  nand g3116 (n_1079, n_2943, n_2944, n_2945);
  xor g3117 (n_2946, n_1060, n_1061);
  xor g3118 (n_1065, n_2946, n_1062);
  nand g3119 (n_2947, n_1060, n_1061);
  nand g3120 (n_2948, n_1062, n_1061);
  nand g3121 (n_2949, n_1060, n_1062);
  nand g3122 (n_1082, n_2947, n_2948, n_2949);
  xor g3123 (n_2950, n_1063, n_1064);
  xor g3124 (n_1067, n_2950, n_1065);
  nand g3125 (n_2951, n_1063, n_1064);
  nand g3126 (n_2952, n_1065, n_1064);
  nand g3127 (n_2953, n_1063, n_1065);
  nand g3128 (n_1084, n_2951, n_2952, n_2953);
  xor g3129 (n_2954, n_1066, n_1067);
  xor g3130 (n_174, n_2954, n_1068);
  nand g3131 (n_2955, n_1066, n_1067);
  nand g3132 (n_2956, n_1068, n_1067);
  nand g3133 (n_2957, n_1066, n_1068);
  nand g3134 (n_87, n_2955, n_2956, n_2957);
  xor g3137 (n_2958, A[66], A[52]);
  xor g3138 (n_1075, n_2958, A[50]);
  nand g3139 (n_2959, A[66], A[52]);
  nand g3141 (n_2961, A[66], A[50]);
  nand g3142 (n_1088, n_2959, n_2511, n_2961);
  xor g3143 (n_2962, A[60], A[48]);
  xor g3144 (n_1076, n_2962, A[58]);
  nand g3145 (n_2963, A[60], A[48]);
  nand g3146 (n_2964, A[58], A[48]);
  nand g3148 (n_1089, n_2963, n_2964, n_2767);
  xor g3149 (n_2966, A[62], A[56]);
  xor g3150 (n_1074, n_2966, A[54]);
  nand g3153 (n_2969, A[62], A[54]);
  nand g3154 (n_1090, n_2833, n_2639, n_2969);
  xor g3155 (n_2970, A[64], n_1071);
  xor g3156 (n_1078, n_2970, n_1072);
  nand g3157 (n_2971, A[64], n_1071);
  nand g3158 (n_2972, n_1072, n_1071);
  nand g3159 (n_2973, A[64], n_1072);
  nand g3160 (n_1094, n_2971, n_2972, n_2973);
  xor g3161 (n_2974, n_1073, n_1074);
  xor g3162 (n_1080, n_2974, n_1075);
  nand g3163 (n_2975, n_1073, n_1074);
  nand g3164 (n_2976, n_1075, n_1074);
  nand g3165 (n_2977, n_1073, n_1075);
  nand g3166 (n_1096, n_2975, n_2976, n_2977);
  xor g3167 (n_2978, n_1076, n_1077);
  xor g3168 (n_1081, n_2978, n_1078);
  nand g3169 (n_2979, n_1076, n_1077);
  nand g3170 (n_2980, n_1078, n_1077);
  nand g3171 (n_2981, n_1076, n_1078);
  nand g3172 (n_1099, n_2979, n_2980, n_2981);
  xor g3173 (n_2982, n_1079, n_1080);
  xor g3174 (n_1083, n_2982, n_1081);
  nand g3175 (n_2983, n_1079, n_1080);
  nand g3176 (n_2984, n_1081, n_1080);
  nand g3177 (n_2985, n_1079, n_1081);
  nand g3178 (n_1101, n_2983, n_2984, n_2985);
  xor g3179 (n_2986, n_1082, n_1083);
  xor g3180 (n_173, n_2986, n_1084);
  nand g3181 (n_2987, n_1082, n_1083);
  nand g3182 (n_2988, n_1084, n_1083);
  nand g3183 (n_2989, n_1082, n_1084);
  nand g3184 (n_86, n_2987, n_2988, n_2989);
  xor g3188 (n_1092, n_2478, A[66]);
  nand g3190 (n_2992, A[66], A[49]);
  nand g3191 (n_2993, A[51], A[66]);
  nand g3192 (n_1103, n_2479, n_2992, n_2993);
  xor g3193 (n_2994, A[63], A[57]);
  xor g3194 (n_1093, n_2994, A[59]);
  nand g3198 (n_1105, n_2865, n_2735, n_2927);
  xor g3205 (n_3002, A[65], n_1088);
  xor g3206 (n_1095, n_3002, n_1089);
  nand g3207 (n_3003, A[65], n_1088);
  nand g3208 (n_3004, n_1089, n_1088);
  nand g3209 (n_3005, A[65], n_1089);
  nand g3210 (n_1109, n_3003, n_3004, n_3005);
  xor g3211 (n_3006, n_1090, n_1058);
  xor g3212 (n_1097, n_3006, n_1092);
  nand g3213 (n_3007, n_1090, n_1058);
  nand g3214 (n_3008, n_1092, n_1058);
  nand g3215 (n_3009, n_1090, n_1092);
  nand g3216 (n_1111, n_3007, n_3008, n_3009);
  xor g3217 (n_3010, n_1093, n_1094);
  xor g3218 (n_1098, n_3010, n_1095);
  nand g3219 (n_3011, n_1093, n_1094);
  nand g3220 (n_3012, n_1095, n_1094);
  nand g3221 (n_3013, n_1093, n_1095);
  nand g3222 (n_1114, n_3011, n_3012, n_3013);
  xor g3223 (n_3014, n_1096, n_1097);
  xor g3224 (n_1100, n_3014, n_1098);
  nand g3225 (n_3015, n_1096, n_1097);
  nand g3226 (n_3016, n_1098, n_1097);
  nand g3227 (n_3017, n_1096, n_1098);
  nand g3228 (n_1116, n_3015, n_3016, n_3017);
  xor g3229 (n_3018, n_1099, n_1100);
  xor g3230 (n_172, n_3018, n_1101);
  nand g3231 (n_3019, n_1099, n_1100);
  nand g3232 (n_3020, n_1101, n_1100);
  nand g3233 (n_3021, n_1099, n_1101);
  nand g3234 (n_85, n_3019, n_3020, n_3021);
  xor g3236 (n_1107, n_3022, A[52]);
  nand g3240 (n_1119, n_3023, n_2905, n_3025);
  xor g3241 (n_3026, A[50], A[58]);
  nand g3246 (n_1120, n_2896, n_3028, n_3029);
  xor g3253 (n_3034, A[64], n_1103);
  xor g3254 (n_1110, n_3034, n_1073);
  nand g3255 (n_3035, A[64], n_1103);
  nand g3256 (n_3036, n_1073, n_1103);
  nand g3257 (n_3037, A[64], n_1073);
  nand g3258 (n_1124, n_3035, n_3036, n_3037);
  xor g3259 (n_3038, n_1105, n_1074);
  xor g3260 (n_1112, n_3038, n_1107);
  nand g3261 (n_3039, n_1105, n_1074);
  nand g3262 (n_3040, n_1107, n_1074);
  nand g3263 (n_3041, n_1105, n_1107);
  nand g3264 (n_1126, n_3039, n_3040, n_3041);
  xor g3265 (n_3042, n_1108, n_1109);
  xor g3266 (n_1113, n_3042, n_1110);
  nand g3267 (n_3043, n_1108, n_1109);
  nand g3268 (n_3044, n_1110, n_1109);
  nand g3269 (n_3045, n_1108, n_1110);
  nand g3270 (n_1129, n_3043, n_3044, n_3045);
  xor g3271 (n_3046, n_1111, n_1112);
  xor g3272 (n_1115, n_3046, n_1113);
  nand g3273 (n_3047, n_1111, n_1112);
  nand g3274 (n_3048, n_1113, n_1112);
  nand g3275 (n_3049, n_1111, n_1113);
  nand g3276 (n_1131, n_3047, n_3048, n_3049);
  xor g3277 (n_3050, n_1114, n_1115);
  xor g3278 (n_171, n_3050, n_1116);
  nand g3279 (n_3051, n_1114, n_1115);
  nand g3280 (n_3052, n_1116, n_1115);
  nand g3281 (n_3053, n_1114, n_1116);
  nand g3282 (n_84, n_3051, n_3052, n_3053);
  xor g3285 (n_3054, A[59], A[51]);
  xor g3286 (n_1123, n_3054, A[57]);
  nand g3290 (n_1134, n_2928, n_2673, n_2735);
  xor g3298 (n_1125, n_3062, n_1119);
  nand g3301 (n_3065, A[65], n_1119);
  nand g3302 (n_1138, n_3063, n_3064, n_3065);
  xor g3303 (n_3066, n_1120, n_1090);
  xor g3304 (n_1127, n_3066, n_1058);
  nand g3305 (n_3067, n_1120, n_1090);
  nand g3307 (n_3069, n_1120, n_1058);
  nand g3308 (n_1140, n_3067, n_3007, n_3069);
  xor g3309 (n_3070, n_1123, n_1124);
  xor g3310 (n_1128, n_3070, n_1125);
  nand g3311 (n_3071, n_1123, n_1124);
  nand g3312 (n_3072, n_1125, n_1124);
  nand g3313 (n_3073, n_1123, n_1125);
  nand g3314 (n_1141, n_3071, n_3072, n_3073);
  xor g3315 (n_3074, n_1126, n_1127);
  xor g3316 (n_1130, n_3074, n_1128);
  nand g3317 (n_3075, n_1126, n_1127);
  nand g3318 (n_3076, n_1128, n_1127);
  nand g3319 (n_3077, n_1126, n_1128);
  nand g3320 (n_1144, n_3075, n_3076, n_3077);
  xor g3321 (n_3078, n_1129, n_1130);
  xor g3322 (n_170, n_3078, n_1131);
  nand g3323 (n_3079, n_1129, n_1130);
  nand g3324 (n_3080, n_1131, n_1130);
  nand g3325 (n_3081, n_1129, n_1131);
  nand g3326 (n_83, n_3079, n_3080, n_3081);
  xor g3334 (n_1136, n_2894, A[56]);
  nand g3338 (n_1148, n_2895, n_2833, n_2703);
  xor g3339 (n_3090, A[54], A[64]);
  xor g3340 (n_1137, n_3090, A[63]);
  nand g3341 (n_3091, A[54], A[64]);
  nand g3342 (n_3092, A[63], A[64]);
  nand g3343 (n_3093, A[54], A[63]);
  nand g3344 (n_1151, n_3091, n_3092, n_3093);
  xor g3345 (n_3094, n_1073, n_1134);
  xor g3346 (n_1139, n_3094, n_1107);
  nand g3347 (n_3095, n_1073, n_1134);
  nand g3348 (n_3096, n_1107, n_1134);
  nand g3349 (n_3097, n_1073, n_1107);
  nand g3350 (n_1153, n_3095, n_3096, n_3097);
  xor g3351 (n_3098, n_1136, n_1137);
  xor g3352 (n_1142, n_3098, n_1138);
  nand g3353 (n_3099, n_1136, n_1137);
  nand g3354 (n_3100, n_1138, n_1137);
  nand g3355 (n_3101, n_1136, n_1138);
  nand g3356 (n_1155, n_3099, n_3100, n_3101);
  xor g3357 (n_3102, n_1139, n_1140);
  xor g3358 (n_1143, n_3102, n_1141);
  nand g3359 (n_3103, n_1139, n_1140);
  nand g3360 (n_3104, n_1141, n_1140);
  nand g3361 (n_3105, n_1139, n_1141);
  nand g3362 (n_1157, n_3103, n_3104, n_3105);
  xor g3363 (n_3106, n_1142, n_1143);
  xor g3364 (n_169, n_3106, n_1144);
  nand g3365 (n_3107, n_1142, n_1143);
  nand g3366 (n_3108, n_1144, n_1143);
  nand g3367 (n_3109, n_1142, n_1144);
  nand g3368 (n_168, n_3107, n_3108, n_3109);
  xor g3372 (n_1150, n_2734, A[61]);
  nand g3376 (n_1159, n_2735, n_2864, n_2799);
  xor g3378 (n_1149, n_2606, A[65]);
  nand g3380 (n_3116, A[65], A[53]);
  nand g3381 (n_3117, A[55], A[65]);
  nand g3382 (n_1161, n_2607, n_3116, n_3117);
  xor g3384 (n_1152, n_3118, n_1148);
  nand g3386 (n_3120, n_1148, n_1119);
  nand g3388 (n_1164, n_3064, n_3120, n_3121);
  xor g3389 (n_3122, n_1149, n_1150);
  xor g3390 (n_1154, n_3122, n_1151);
  nand g3391 (n_3123, n_1149, n_1150);
  nand g3392 (n_3124, n_1151, n_1150);
  nand g3393 (n_3125, n_1149, n_1151);
  nand g3394 (n_1165, n_3123, n_3124, n_3125);
  xor g3395 (n_3126, n_1152, n_1153);
  xor g3396 (n_1156, n_3126, n_1154);
  nand g3397 (n_3127, n_1152, n_1153);
  nand g3398 (n_3128, n_1154, n_1153);
  nand g3399 (n_3129, n_1152, n_1154);
  nand g3400 (n_1168, n_3127, n_3128, n_3129);
  xor g3401 (n_3130, n_1155, n_1156);
  xor g3402 (n_82, n_3130, n_1157);
  nand g3403 (n_3131, n_1155, n_1156);
  nand g3404 (n_3132, n_1157, n_1156);
  nand g3405 (n_3133, n_1155, n_1157);
  nand g3406 (n_81, n_3131, n_3132, n_3133);
  xor g3408 (n_1162, n_3022, A[58]);
  nand g3412 (n_1171, n_3023, n_2767, n_3028);
  xor g3419 (n_3142, A[64], A[63]);
  xor g3420 (n_1163, n_3142, n_1159);
  nand g3422 (n_3144, n_1159, A[63]);
  nand g3423 (n_3145, A[64], n_1159);
  nand g3424 (n_1175, n_3092, n_3144, n_3145);
  xor g3425 (n_3146, n_1074, n_1161);
  xor g3426 (n_1166, n_3146, n_1162);
  nand g3427 (n_3147, n_1074, n_1161);
  nand g3428 (n_3148, n_1162, n_1161);
  nand g3429 (n_3149, n_1074, n_1162);
  nand g3430 (n_1176, n_3147, n_3148, n_3149);
  xor g3431 (n_3150, n_1163, n_1164);
  xor g3432 (n_1167, n_3150, n_1165);
  nand g3433 (n_3151, n_1163, n_1164);
  nand g3434 (n_3152, n_1165, n_1164);
  nand g3435 (n_3153, n_1163, n_1165);
  nand g3436 (n_1179, n_3151, n_3152, n_3153);
  xor g3437 (n_3154, n_1166, n_1167);
  xor g3438 (n_167, n_3154, n_1168);
  nand g3439 (n_3155, n_1166, n_1167);
  nand g3440 (n_3156, n_1168, n_1167);
  nand g3441 (n_3157, n_1166, n_1168);
  nand g3442 (n_80, n_3155, n_3156, n_3157);
  xor g3446 (n_1173, n_2994, A[55]);
  nand g3448 (n_3160, A[55], A[63]);
  nand g3450 (n_1181, n_2865, n_3160, n_2671);
  xor g3451 (n_3162, A[61], A[65]);
  nand g3453 (n_3163, A[61], A[65]);
  nand g3456 (n_1184, n_3163, n_3164, n_3165);
  xor g3457 (n_3166, n_1171, n_1090);
  xor g3458 (n_1177, n_3166, n_1173);
  nand g3459 (n_3167, n_1171, n_1090);
  nand g3460 (n_3168, n_1173, n_1090);
  nand g3461 (n_3169, n_1171, n_1173);
  nand g3462 (n_1186, n_3167, n_3168, n_3169);
  xor g3463 (n_3170, n_1174, n_1175);
  xor g3464 (n_1178, n_3170, n_1176);
  nand g3465 (n_3171, n_1174, n_1175);
  nand g3466 (n_3172, n_1176, n_1175);
  nand g3467 (n_3173, n_1174, n_1176);
  nand g3468 (n_1188, n_3171, n_3172, n_3173);
  xor g3469 (n_3174, n_1177, n_1178);
  xor g3470 (n_166, n_3174, n_1179);
  nand g3471 (n_3175, n_1177, n_1178);
  nand g3472 (n_3176, n_1179, n_1178);
  nand g3473 (n_3177, n_1177, n_1179);
  nand g3474 (n_79, n_3175, n_3176, n_3177);
  xor g3482 (n_1182, n_2966, A[64]);
  nand g3484 (n_3184, A[64], A[56]);
  nand g3485 (n_3185, A[62], A[64]);
  nand g3486 (n_1193, n_2833, n_3184, n_3185);
  xor g3487 (n_3186, A[59], n_1181);
  xor g3488 (n_1185, n_3186, n_1182);
  nand g3489 (n_3187, A[59], n_1181);
  nand g3490 (n_3188, n_1182, n_1181);
  nand g3491 (n_3189, A[59], n_1182);
  nand g3492 (n_1195, n_3187, n_3188, n_3189);
  xor g3493 (n_3190, n_1162, n_1184);
  xor g3494 (n_1187, n_3190, n_1185);
  nand g3495 (n_3191, n_1162, n_1184);
  nand g3496 (n_3192, n_1185, n_1184);
  nand g3497 (n_3193, n_1162, n_1185);
  nand g3498 (n_1197, n_3191, n_3192, n_3193);
  xor g3499 (n_3194, n_1186, n_1187);
  xor g3500 (n_165, n_3194, n_1188);
  nand g3501 (n_3195, n_1186, n_1187);
  nand g3502 (n_3196, n_1188, n_1187);
  nand g3503 (n_3197, n_1186, n_1188);
  nand g3504 (n_78, n_3195, n_3196, n_3197);
  xor g3508 (n_1192, n_2994, A[61]);
  xor g3514 (n_1194, n_3202, n_1171);
  nand g3517 (n_3205, A[65], n_1171);
  nand g3518 (n_1202, n_3164, n_3204, n_3205);
  xor g3519 (n_3206, n_1192, n_1193);
  xor g3520 (n_1196, n_3206, n_1194);
  nand g3521 (n_3207, n_1192, n_1193);
  nand g3522 (n_3208, n_1194, n_1193);
  nand g3523 (n_3209, n_1192, n_1194);
  nand g3524 (n_1204, n_3207, n_3208, n_3209);
  xor g3525 (n_3210, n_1195, n_1196);
  xor g3526 (n_164, n_3210, n_1197);
  nand g3527 (n_3211, n_1195, n_1196);
  nand g3528 (n_3212, n_1197, n_1196);
  nand g3529 (n_3213, n_1195, n_1197);
  nand g3530 (n_163, n_3211, n_3212, n_3213);
  xor g3537 (n_3218, A[62], A[64]);
  xor g3538 (n_1201, n_3218, A[59]);
  nand g3540 (n_3220, A[59], A[64]);
  nand g3541 (n_3221, A[62], A[59]);
  nand g3542 (n_1209, n_3185, n_3220, n_3221);
  xor g3543 (n_3222, n_1041, n_1162);
  xor g3544 (n_1203, n_3222, n_1201);
  nand g3545 (n_3223, n_1041, n_1162);
  nand g3546 (n_3224, n_1201, n_1162);
  nand g3547 (n_3225, n_1041, n_1201);
  nand g3548 (n_1211, n_3223, n_3224, n_3225);
  xor g3549 (n_3226, n_1202, n_1203);
  xor g3550 (n_77, n_3226, n_1204);
  nand g3551 (n_3227, n_1202, n_1203);
  nand g3552 (n_3228, n_1204, n_1203);
  nand g3553 (n_3229, n_1202, n_1204);
  nand g3554 (n_162, n_3227, n_3228, n_3229);
  xor g3558 (n_1208, n_2798, A[65]);
  nand g3561 (n_3233, A[59], A[65]);
  nand g3562 (n_1214, n_2799, n_3163, n_3233);
  xor g3564 (n_1210, n_3234, n_1208);
  nand g3566 (n_3236, n_1208, n_1171);
  nand g3568 (n_1216, n_3235, n_3236, n_3237);
  xor g3569 (n_3238, n_1209, n_1210);
  xor g3570 (n_76, n_3238, n_1211);
  nand g3571 (n_3239, n_1209, n_1210);
  nand g3572 (n_3240, n_1211, n_1210);
  nand g3573 (n_3241, n_1209, n_1211);
  nand g3574 (n_75, n_3239, n_3240, n_3241);
  xor g3576 (n_1213, n_3022, A[62]);
  nand g3580 (n_1219, n_3023, n_2831, n_3245);
  xor g3582 (n_1215, n_3142, n_1213);
  nand g3584 (n_3248, n_1213, A[63]);
  nand g3585 (n_3249, A[64], n_1213);
  nand g3586 (n_1221, n_3092, n_3248, n_3249);
  xor g3587 (n_3250, n_1214, n_1215);
  xor g3588 (n_161, n_3250, n_1216);
  nand g3589 (n_3251, n_1214, n_1215);
  nand g3590 (n_3252, n_1216, n_1215);
  nand g3591 (n_3253, n_1214, n_1216);
  nand g3592 (n_74, n_3251, n_3252, n_3253);
  nand g3600 (n_1224, n_3163, n_3063, n_3257);
  xor g3601 (n_3258, n_1219, n_1220);
  xor g3602 (n_160, n_3258, n_1221);
  nand g3603 (n_3259, n_1219, n_1220);
  nand g3604 (n_3260, n_1221, n_1220);
  nand g3605 (n_3261, n_1219, n_1221);
  nand g3606 (n_159, n_3259, n_3260, n_3261);
  xor g3608 (n_1223, n_3262, A[64]);
  nand g3612 (n_1227, n_3245, n_3185, n_3265);
  xor g3613 (n_3266, A[63], n_1223);
  xor g3614 (n_73, n_3266, n_1224);
  nand g3615 (n_3267, A[63], n_1223);
  nand g3616 (n_3268, n_1224, n_1223);
  nand g3617 (n_3269, A[63], n_1224);
  nand g3618 (n_158, n_3267, n_3268, n_3269);
  xor g3622 (n_72, n_3062, n_1227);
  nand g3625 (n_3273, A[65], n_1227);
  nand g3626 (n_157, n_3063, n_3272, n_3273);
  xor g3628 (n_71, n_3274, A[63]);
  nand g3632 (n_156, n_3265, n_3092, n_3277);
  nand g25 (n_3299, n_1232, n_3296, n_3297);
  nand g28 (n_3300, A[2], n_235);
  nand g29 (n_3301, A[2], n_3299);
  nand g30 (n_3302, n_235, n_3299);
  nand g31 (n_3304, n_3300, n_3301, n_3302);
  xor g32 (n_3303, A[2], n_235);
  xor g33 (Z[4], n_3299, n_3303);
  nand g34 (n_3305, n_148, n_234);
  nand g35 (n_3306, n_148, n_3304);
  nand g36 (n_3307, n_234, n_3304);
  nand g37 (n_3309, n_3305, n_3306, n_3307);
  xor g38 (n_3308, n_148, n_234);
  xor g39 (Z[5], n_3304, n_3308);
  nand g40 (n_3310, n_147, n_233);
  nand g41 (n_3311, n_147, n_3309);
  nand g42 (n_3312, n_233, n_3309);
  nand g43 (n_3314, n_3310, n_3311, n_3312);
  xor g44 (n_3313, n_147, n_233);
  xor g45 (Z[6], n_3309, n_3313);
  nand g46 (n_3315, n_146, n_232);
  nand g47 (n_3316, n_146, n_3314);
  nand g48 (n_3317, n_232, n_3314);
  nand g49 (n_3319, n_3315, n_3316, n_3317);
  xor g50 (n_3318, n_146, n_232);
  xor g51 (Z[7], n_3314, n_3318);
  nand g52 (n_3320, n_145, n_231);
  nand g53 (n_3321, n_145, n_3319);
  nand g54 (n_3322, n_231, n_3319);
  nand g55 (n_3324, n_3320, n_3321, n_3322);
  xor g56 (n_3323, n_145, n_231);
  xor g57 (Z[8], n_3319, n_3323);
  nand g58 (n_3325, n_144, n_230);
  nand g59 (n_3326, n_144, n_3324);
  nand g60 (n_3327, n_230, n_3324);
  nand g61 (n_3329, n_3325, n_3326, n_3327);
  xor g62 (n_3328, n_144, n_230);
  xor g63 (Z[9], n_3324, n_3328);
  nand g64 (n_3330, n_143, n_229);
  nand g65 (n_3331, n_143, n_3329);
  nand g66 (n_3332, n_229, n_3329);
  nand g67 (n_3334, n_3330, n_3331, n_3332);
  xor g68 (n_3333, n_143, n_229);
  xor g69 (Z[10], n_3329, n_3333);
  nand g70 (n_3335, n_142, n_228);
  nand g71 (n_3336, n_142, n_3334);
  nand g72 (n_3337, n_228, n_3334);
  nand g73 (n_3339, n_3335, n_3336, n_3337);
  xor g74 (n_3338, n_142, n_228);
  xor g75 (Z[11], n_3334, n_3338);
  nand g76 (n_3340, n_141, n_227);
  nand g77 (n_3341, n_141, n_3339);
  nand g78 (n_3342, n_227, n_3339);
  nand g79 (n_3344, n_3340, n_3341, n_3342);
  xor g80 (n_3343, n_141, n_227);
  xor g81 (Z[12], n_3339, n_3343);
  nand g82 (n_3345, n_140, n_226);
  nand g83 (n_3346, n_140, n_3344);
  nand g84 (n_3347, n_226, n_3344);
  nand g85 (n_3349, n_3345, n_3346, n_3347);
  xor g86 (n_3348, n_140, n_226);
  xor g87 (Z[13], n_3344, n_3348);
  nand g88 (n_3350, n_139, n_225);
  nand g89 (n_3351, n_139, n_3349);
  nand g90 (n_3352, n_225, n_3349);
  nand g91 (n_3354, n_3350, n_3351, n_3352);
  xor g92 (n_3353, n_139, n_225);
  xor g93 (Z[14], n_3349, n_3353);
  nand g94 (n_3355, n_138, n_224);
  nand g95 (n_3356, n_138, n_3354);
  nand g96 (n_3357, n_224, n_3354);
  nand g97 (n_3359, n_3355, n_3356, n_3357);
  xor g98 (n_3358, n_138, n_224);
  xor g99 (Z[15], n_3354, n_3358);
  nand g100 (n_3360, n_137, n_223);
  nand g101 (n_3361, n_137, n_3359);
  nand g102 (n_3362, n_223, n_3359);
  nand g103 (n_3364, n_3360, n_3361, n_3362);
  xor g104 (n_3363, n_137, n_223);
  xor g105 (Z[16], n_3359, n_3363);
  nand g106 (n_3365, n_136, n_222);
  nand g107 (n_3366, n_136, n_3364);
  nand g108 (n_3367, n_222, n_3364);
  nand g109 (n_3369, n_3365, n_3366, n_3367);
  xor g110 (n_3368, n_136, n_222);
  xor g111 (Z[17], n_3364, n_3368);
  nand g112 (n_3370, n_135, n_221);
  nand g113 (n_3371, n_135, n_3369);
  nand g114 (n_3372, n_221, n_3369);
  nand g115 (n_3374, n_3370, n_3371, n_3372);
  xor g116 (n_3373, n_135, n_221);
  xor g117 (Z[18], n_3369, n_3373);
  nand g118 (n_3375, n_134, n_220);
  nand g119 (n_3376, n_134, n_3374);
  nand g120 (n_3377, n_220, n_3374);
  nand g121 (n_3379, n_3375, n_3376, n_3377);
  xor g122 (n_3378, n_134, n_220);
  xor g123 (Z[19], n_3374, n_3378);
  nand g124 (n_3380, n_133, n_219);
  nand g125 (n_3381, n_133, n_3379);
  nand g126 (n_3382, n_219, n_3379);
  nand g127 (n_3384, n_3380, n_3381, n_3382);
  xor g128 (n_3383, n_133, n_219);
  xor g129 (Z[20], n_3379, n_3383);
  nand g130 (n_3385, n_132, n_218);
  nand g131 (n_3386, n_132, n_3384);
  nand g132 (n_3387, n_218, n_3384);
  nand g133 (n_3389, n_3385, n_3386, n_3387);
  xor g134 (n_3388, n_132, n_218);
  xor g135 (Z[21], n_3384, n_3388);
  nand g136 (n_3390, n_131, n_217);
  nand g137 (n_3391, n_131, n_3389);
  nand g138 (n_3392, n_217, n_3389);
  nand g139 (n_3394, n_3390, n_3391, n_3392);
  xor g140 (n_3393, n_131, n_217);
  xor g141 (Z[22], n_3389, n_3393);
  nand g142 (n_3395, n_130, n_216);
  nand g143 (n_3396, n_130, n_3394);
  nand g144 (n_3397, n_216, n_3394);
  nand g145 (n_3399, n_3395, n_3396, n_3397);
  xor g146 (n_3398, n_130, n_216);
  xor g147 (Z[23], n_3394, n_3398);
  nand g148 (n_3400, n_129, n_215);
  nand g149 (n_3401, n_129, n_3399);
  nand g150 (n_3402, n_215, n_3399);
  nand g151 (n_3404, n_3400, n_3401, n_3402);
  xor g152 (n_3403, n_129, n_215);
  xor g153 (Z[24], n_3399, n_3403);
  nand g154 (n_3405, n_128, n_214);
  nand g155 (n_3406, n_128, n_3404);
  nand g156 (n_3407, n_214, n_3404);
  nand g157 (n_3409, n_3405, n_3406, n_3407);
  xor g158 (n_3408, n_128, n_214);
  xor g159 (Z[25], n_3404, n_3408);
  nand g160 (n_3410, n_127, n_213);
  nand g161 (n_3411, n_127, n_3409);
  nand g162 (n_3412, n_213, n_3409);
  nand g163 (n_3414, n_3410, n_3411, n_3412);
  xor g164 (n_3413, n_127, n_213);
  xor g165 (Z[26], n_3409, n_3413);
  nand g166 (n_3415, n_126, n_212);
  nand g167 (n_3416, n_126, n_3414);
  nand g168 (n_3417, n_212, n_3414);
  nand g169 (n_3419, n_3415, n_3416, n_3417);
  xor g170 (n_3418, n_126, n_212);
  xor g171 (Z[27], n_3414, n_3418);
  nand g172 (n_3420, n_125, n_211);
  nand g173 (n_3421, n_125, n_3419);
  nand g174 (n_3422, n_211, n_3419);
  nand g175 (n_3424, n_3420, n_3421, n_3422);
  xor g176 (n_3423, n_125, n_211);
  xor g177 (Z[28], n_3419, n_3423);
  nand g178 (n_3425, n_124, n_210);
  nand g179 (n_3426, n_124, n_3424);
  nand g180 (n_3427, n_210, n_3424);
  nand g181 (n_3429, n_3425, n_3426, n_3427);
  xor g182 (n_3428, n_124, n_210);
  xor g183 (Z[29], n_3424, n_3428);
  nand g184 (n_3430, n_123, n_209);
  nand g185 (n_3431, n_123, n_3429);
  nand g186 (n_3432, n_209, n_3429);
  nand g187 (n_3434, n_3430, n_3431, n_3432);
  xor g188 (n_3433, n_123, n_209);
  xor g189 (Z[30], n_3429, n_3433);
  nand g190 (n_3435, n_122, n_208);
  nand g191 (n_3436, n_122, n_3434);
  nand g192 (n_3437, n_208, n_3434);
  nand g193 (n_3439, n_3435, n_3436, n_3437);
  xor g194 (n_3438, n_122, n_208);
  xor g195 (Z[31], n_3434, n_3438);
  nand g196 (n_3440, n_121, n_207);
  nand g197 (n_3441, n_121, n_3439);
  nand g198 (n_3442, n_207, n_3439);
  nand g199 (n_3444, n_3440, n_3441, n_3442);
  xor g200 (n_3443, n_121, n_207);
  xor g201 (Z[32], n_3439, n_3443);
  nand g202 (n_3445, n_120, n_206);
  nand g203 (n_3446, n_120, n_3444);
  nand g204 (n_3447, n_206, n_3444);
  nand g205 (n_3449, n_3445, n_3446, n_3447);
  xor g206 (n_3448, n_120, n_206);
  xor g207 (Z[33], n_3444, n_3448);
  nand g208 (n_3450, n_119, n_205);
  nand g209 (n_3451, n_119, n_3449);
  nand g210 (n_3452, n_205, n_3449);
  nand g211 (n_3454, n_3450, n_3451, n_3452);
  xor g212 (n_3453, n_119, n_205);
  xor g213 (Z[34], n_3449, n_3453);
  nand g214 (n_3455, n_118, n_204);
  nand g215 (n_3456, n_118, n_3454);
  nand g216 (n_3457, n_204, n_3454);
  nand g217 (n_3459, n_3455, n_3456, n_3457);
  xor g218 (n_3458, n_118, n_204);
  xor g219 (Z[35], n_3454, n_3458);
  nand g220 (n_3460, n_117, n_203);
  nand g221 (n_3461, n_117, n_3459);
  nand g222 (n_3462, n_203, n_3459);
  nand g223 (n_3464, n_3460, n_3461, n_3462);
  xor g224 (n_3463, n_117, n_203);
  xor g225 (Z[36], n_3459, n_3463);
  nand g226 (n_3465, n_116, n_202);
  nand g227 (n_3466, n_116, n_3464);
  nand g228 (n_3467, n_202, n_3464);
  nand g229 (n_3469, n_3465, n_3466, n_3467);
  xor g230 (n_3468, n_116, n_202);
  xor g231 (Z[37], n_3464, n_3468);
  nand g232 (n_3470, n_115, n_201);
  nand g233 (n_3471, n_115, n_3469);
  nand g234 (n_3472, n_201, n_3469);
  nand g235 (n_3474, n_3470, n_3471, n_3472);
  xor g236 (n_3473, n_115, n_201);
  xor g237 (Z[38], n_3469, n_3473);
  nand g238 (n_3475, n_114, n_200);
  nand g239 (n_3476, n_114, n_3474);
  nand g240 (n_3477, n_200, n_3474);
  nand g241 (n_3479, n_3475, n_3476, n_3477);
  xor g242 (n_3478, n_114, n_200);
  xor g243 (Z[39], n_3474, n_3478);
  nand g244 (n_3480, n_113, n_199);
  nand g245 (n_3481, n_113, n_3479);
  nand g246 (n_3482, n_199, n_3479);
  nand g247 (n_3484, n_3480, n_3481, n_3482);
  xor g248 (n_3483, n_113, n_199);
  xor g249 (Z[40], n_3479, n_3483);
  nand g250 (n_3485, n_112, n_198);
  nand g251 (n_3486, n_112, n_3484);
  nand g252 (n_3487, n_198, n_3484);
  nand g253 (n_3489, n_3485, n_3486, n_3487);
  xor g254 (n_3488, n_112, n_198);
  xor g255 (Z[41], n_3484, n_3488);
  nand g256 (n_3490, n_111, n_197);
  nand g257 (n_3491, n_111, n_3489);
  nand g258 (n_3492, n_197, n_3489);
  nand g259 (n_3494, n_3490, n_3491, n_3492);
  xor g260 (n_3493, n_111, n_197);
  xor g261 (Z[42], n_3489, n_3493);
  nand g262 (n_3495, n_110, n_196);
  nand g263 (n_3496, n_110, n_3494);
  nand g264 (n_3497, n_196, n_3494);
  nand g265 (n_3499, n_3495, n_3496, n_3497);
  xor g266 (n_3498, n_110, n_196);
  xor g267 (Z[43], n_3494, n_3498);
  nand g268 (n_3500, n_109, n_195);
  nand g269 (n_3501, n_109, n_3499);
  nand g270 (n_3502, n_195, n_3499);
  nand g271 (n_3504, n_3500, n_3501, n_3502);
  xor g272 (n_3503, n_109, n_195);
  xor g273 (Z[44], n_3499, n_3503);
  nand g274 (n_3505, n_108, n_194);
  nand g275 (n_3506, n_108, n_3504);
  nand g276 (n_3507, n_194, n_3504);
  nand g277 (n_3509, n_3505, n_3506, n_3507);
  xor g278 (n_3508, n_108, n_194);
  xor g279 (Z[45], n_3504, n_3508);
  nand g280 (n_3510, n_107, n_193);
  nand g281 (n_3511, n_107, n_3509);
  nand g282 (n_3512, n_193, n_3509);
  nand g283 (n_3514, n_3510, n_3511, n_3512);
  xor g284 (n_3513, n_107, n_193);
  xor g285 (Z[46], n_3509, n_3513);
  nand g286 (n_3515, n_106, n_192);
  nand g287 (n_3516, n_106, n_3514);
  nand g288 (n_3517, n_192, n_3514);
  nand g289 (n_3519, n_3515, n_3516, n_3517);
  xor g290 (n_3518, n_106, n_192);
  xor g291 (Z[47], n_3514, n_3518);
  nand g292 (n_3520, n_105, n_191);
  nand g293 (n_3521, n_105, n_3519);
  nand g294 (n_3522, n_191, n_3519);
  nand g295 (n_3524, n_3520, n_3521, n_3522);
  xor g296 (n_3523, n_105, n_191);
  xor g297 (Z[48], n_3519, n_3523);
  nand g298 (n_3525, n_104, n_190);
  nand g299 (n_3526, n_104, n_3524);
  nand g300 (n_3527, n_190, n_3524);
  nand g301 (n_3529, n_3525, n_3526, n_3527);
  xor g302 (n_3528, n_104, n_190);
  xor g303 (Z[49], n_3524, n_3528);
  nand g304 (n_3530, n_103, n_189);
  nand g305 (n_3531, n_103, n_3529);
  nand g306 (n_3532, n_189, n_3529);
  nand g307 (n_3534, n_3530, n_3531, n_3532);
  xor g308 (n_3533, n_103, n_189);
  xor g309 (Z[50], n_3529, n_3533);
  nand g310 (n_3535, n_102, n_188);
  nand g311 (n_3536, n_102, n_3534);
  nand g312 (n_3537, n_188, n_3534);
  nand g313 (n_3539, n_3535, n_3536, n_3537);
  xor g314 (n_3538, n_102, n_188);
  xor g315 (Z[51], n_3534, n_3538);
  nand g316 (n_3540, n_101, n_187);
  nand g317 (n_3541, n_101, n_3539);
  nand g318 (n_3542, n_187, n_3539);
  nand g319 (n_3544, n_3540, n_3541, n_3542);
  xor g320 (n_3543, n_101, n_187);
  xor g321 (Z[52], n_3539, n_3543);
  nand g322 (n_3545, n_100, n_186);
  nand g323 (n_3546, n_100, n_3544);
  nand g324 (n_3547, n_186, n_3544);
  nand g325 (n_3549, n_3545, n_3546, n_3547);
  xor g326 (n_3548, n_100, n_186);
  xor g327 (Z[53], n_3544, n_3548);
  nand g328 (n_3550, n_99, n_185);
  nand g329 (n_3551, n_99, n_3549);
  nand g330 (n_3552, n_185, n_3549);
  nand g331 (n_3554, n_3550, n_3551, n_3552);
  xor g332 (n_3553, n_99, n_185);
  xor g333 (Z[54], n_3549, n_3553);
  nand g334 (n_3555, n_98, n_184);
  nand g335 (n_3556, n_98, n_3554);
  nand g336 (n_3557, n_184, n_3554);
  nand g337 (n_3559, n_3555, n_3556, n_3557);
  xor g338 (n_3558, n_98, n_184);
  xor g339 (Z[55], n_3554, n_3558);
  nand g340 (n_3560, n_97, n_183);
  nand g341 (n_3561, n_97, n_3559);
  nand g342 (n_3562, n_183, n_3559);
  nand g343 (n_3564, n_3560, n_3561, n_3562);
  xor g344 (n_3563, n_97, n_183);
  xor g345 (Z[56], n_3559, n_3563);
  nand g346 (n_3565, n_96, n_182);
  nand g347 (n_3566, n_96, n_3564);
  nand g348 (n_3567, n_182, n_3564);
  nand g349 (n_3569, n_3565, n_3566, n_3567);
  xor g350 (n_3568, n_96, n_182);
  xor g351 (Z[57], n_3564, n_3568);
  nand g352 (n_3570, n_95, n_181);
  nand g353 (n_3571, n_95, n_3569);
  nand g354 (n_3572, n_181, n_3569);
  nand g355 (n_3574, n_3570, n_3571, n_3572);
  xor g356 (n_3573, n_95, n_181);
  xor g357 (Z[58], n_3569, n_3573);
  nand g358 (n_3575, n_94, n_180);
  nand g359 (n_3576, n_94, n_3574);
  nand g360 (n_3577, n_180, n_3574);
  nand g361 (n_3579, n_3575, n_3576, n_3577);
  xor g362 (n_3578, n_94, n_180);
  xor g363 (Z[59], n_3574, n_3578);
  nand g364 (n_3580, n_93, n_179);
  nand g365 (n_3581, n_93, n_3579);
  nand g366 (n_3582, n_179, n_3579);
  nand g367 (n_3584, n_3580, n_3581, n_3582);
  xor g368 (n_3583, n_93, n_179);
  xor g369 (Z[60], n_3579, n_3583);
  nand g370 (n_3585, n_92, n_178);
  nand g371 (n_3586, n_92, n_3584);
  nand g372 (n_3587, n_178, n_3584);
  nand g373 (n_3589, n_3585, n_3586, n_3587);
  xor g374 (n_3588, n_92, n_178);
  xor g375 (Z[61], n_3584, n_3588);
  nand g376 (n_3590, n_91, n_177);
  nand g377 (n_3591, n_91, n_3589);
  nand g378 (n_3592, n_177, n_3589);
  nand g379 (n_3594, n_3590, n_3591, n_3592);
  xor g380 (n_3593, n_91, n_177);
  xor g381 (Z[62], n_3589, n_3593);
  nand g382 (n_3595, n_90, n_176);
  nand g383 (n_3596, n_90, n_3594);
  nand g384 (n_3597, n_176, n_3594);
  nand g385 (n_3599, n_3595, n_3596, n_3597);
  xor g386 (n_3598, n_90, n_176);
  xor g387 (Z[63], n_3594, n_3598);
  nand g388 (n_3600, n_89, n_175);
  nand g389 (n_3601, n_89, n_3599);
  nand g390 (n_3602, n_175, n_3599);
  nand g391 (n_3604, n_3600, n_3601, n_3602);
  xor g392 (n_3603, n_89, n_175);
  xor g393 (Z[64], n_3599, n_3603);
  nand g394 (n_3605, n_88, n_174);
  nand g395 (n_3606, n_88, n_3604);
  nand g396 (n_3607, n_174, n_3604);
  nand g397 (n_3609, n_3605, n_3606, n_3607);
  xor g398 (n_3608, n_88, n_174);
  xor g399 (Z[65], n_3604, n_3608);
  nand g400 (n_3610, n_87, n_173);
  nand g401 (n_3611, n_87, n_3609);
  nand g402 (n_3612, n_173, n_3609);
  nand g403 (n_3614, n_3610, n_3611, n_3612);
  xor g404 (n_3613, n_87, n_173);
  xor g405 (Z[66], n_3609, n_3613);
  nand g406 (n_3615, n_86, n_172);
  nand g407 (n_3616, n_86, n_3614);
  nand g408 (n_3617, n_172, n_3614);
  nand g409 (n_3619, n_3615, n_3616, n_3617);
  xor g410 (n_3618, n_86, n_172);
  xor g411 (Z[67], n_3614, n_3618);
  nand g412 (n_3620, n_85, n_171);
  nand g413 (n_3621, n_85, n_3619);
  nand g414 (n_3622, n_171, n_3619);
  nand g415 (n_3624, n_3620, n_3621, n_3622);
  xor g416 (n_3623, n_85, n_171);
  xor g417 (Z[68], n_3619, n_3623);
  nand g418 (n_3625, n_84, n_170);
  nand g419 (n_3626, n_84, n_3624);
  nand g420 (n_3627, n_170, n_3624);
  nand g421 (n_3629, n_3625, n_3626, n_3627);
  xor g422 (n_3628, n_84, n_170);
  xor g423 (Z[69], n_3624, n_3628);
  nand g424 (n_3630, n_83, n_169);
  nand g425 (n_3631, n_83, n_3629);
  nand g426 (n_3632, n_169, n_3629);
  nand g427 (n_3634, n_3630, n_3631, n_3632);
  xor g428 (n_3633, n_83, n_169);
  xor g429 (Z[70], n_3629, n_3633);
  nand g430 (n_3635, n_82, n_168);
  nand g431 (n_3636, n_82, n_3634);
  nand g432 (n_3637, n_168, n_3634);
  nand g433 (n_3639, n_3635, n_3636, n_3637);
  xor g434 (n_3638, n_82, n_168);
  xor g435 (Z[71], n_3634, n_3638);
  nand g436 (n_3640, n_81, n_167);
  nand g437 (n_3641, n_81, n_3639);
  nand g438 (n_3642, n_167, n_3639);
  nand g439 (n_3644, n_3640, n_3641, n_3642);
  xor g440 (n_3643, n_81, n_167);
  xor g441 (Z[72], n_3639, n_3643);
  nand g442 (n_3645, n_80, n_166);
  nand g443 (n_3646, n_80, n_3644);
  nand g444 (n_3647, n_166, n_3644);
  nand g445 (n_3649, n_3645, n_3646, n_3647);
  xor g446 (n_3648, n_80, n_166);
  xor g447 (Z[73], n_3644, n_3648);
  nand g448 (n_3650, n_79, n_165);
  nand g449 (n_3651, n_79, n_3649);
  nand g450 (n_3652, n_165, n_3649);
  nand g451 (n_3654, n_3650, n_3651, n_3652);
  xor g452 (n_3653, n_79, n_165);
  xor g453 (Z[74], n_3649, n_3653);
  nand g454 (n_3655, n_78, n_164);
  nand g455 (n_3656, n_78, n_3654);
  nand g456 (n_3657, n_164, n_3654);
  nand g457 (n_3659, n_3655, n_3656, n_3657);
  xor g458 (n_3658, n_78, n_164);
  xor g459 (Z[75], n_3654, n_3658);
  nand g460 (n_3660, n_77, n_163);
  nand g461 (n_3661, n_77, n_3659);
  nand g462 (n_3662, n_163, n_3659);
  nand g463 (n_3664, n_3660, n_3661, n_3662);
  xor g464 (n_3663, n_77, n_163);
  xor g465 (Z[76], n_3659, n_3663);
  nand g466 (n_3665, n_76, n_162);
  nand g467 (n_3666, n_76, n_3664);
  nand g468 (n_3667, n_162, n_3664);
  nand g469 (n_3669, n_3665, n_3666, n_3667);
  xor g470 (n_3668, n_76, n_162);
  xor g471 (Z[77], n_3664, n_3668);
  nand g472 (n_3670, n_75, n_161);
  nand g473 (n_3671, n_75, n_3669);
  nand g474 (n_3672, n_161, n_3669);
  nand g475 (n_3674, n_3670, n_3671, n_3672);
  xor g476 (n_3673, n_75, n_161);
  xor g477 (Z[78], n_3669, n_3673);
  nand g478 (n_3675, n_74, n_160);
  nand g479 (n_3676, n_74, n_3674);
  nand g480 (n_3677, n_160, n_3674);
  nand g481 (n_3679, n_3675, n_3676, n_3677);
  xor g482 (n_3678, n_74, n_160);
  xor g483 (Z[79], n_3674, n_3678);
  nand g484 (n_3680, n_73, n_159);
  nand g485 (n_3681, n_73, n_3679);
  nand g486 (n_3682, n_159, n_3679);
  nand g487 (n_3684, n_3680, n_3681, n_3682);
  xor g488 (n_3683, n_73, n_159);
  xor g489 (Z[80], n_3679, n_3683);
  nand g490 (n_3685, n_72, n_158);
  nand g491 (n_3686, n_72, n_3684);
  nand g492 (n_3687, n_158, n_3684);
  nand g493 (n_3689, n_3685, n_3686, n_3687);
  xor g494 (n_3688, n_72, n_158);
  xor g495 (Z[81], n_3684, n_3688);
  nand g496 (n_3690, n_71, n_157);
  nand g497 (n_3691, n_71, n_3689);
  nand g498 (n_3692, n_157, n_3689);
  nand g499 (n_3694, n_3690, n_3691, n_3692);
  xor g500 (n_3693, n_71, n_157);
  xor g501 (Z[82], n_3689, n_3693);
  nand g504 (n_3697, n_156, n_3694);
  nand g505 (n_3699, n_3695, n_3696, n_3697);
  xor g507 (Z[83], n_3694, n_3698);
  nand g510 (n_3702, A[65], n_3699);
  nand g511 (n_3704, n_3700, n_3701, n_3702);
  xor g513 (Z[84], n_3699, n_3703);
  or g3651 (n_334, wc, wc0, n_148);
  not gc0 (wc0, n_1235);
  not gc (wc, n_1249);
  or g3652 (n_343, wc1, wc2, n_328);
  not gc2 (wc2, n_1249);
  not gc1 (wc1, n_1268);
  or g3653 (n_356, wc3, n_333, n_328);
  not gc3 (wc3, n_1296);
  or g3654 (n_373, wc4, wc5, n_333);
  not gc5 (wc5, n_1331);
  not gc4 (wc4, n_1332);
  or g3655 (n_395, wc6, wc7, n_333);
  not gc7 (wc7, n_1379);
  not gc6 (wc6, n_1380);
  or g3656 (n_447, wc8, wc9, n_328);
  not gc9 (wc9, n_1380);
  not gc8 (wc8, n_1427);
  or g3657 (n_470, wc10, wc11, n_333);
  not gc11 (wc11, n_1556);
  not gc10 (wc10, n_1557);
  or g3658 (n_498, wc12, wc13, n_342);
  not gc13 (wc13, n_1496);
  not gc12 (wc12, n_1620);
  or g3659 (n_526, wc14, wc15, n_355);
  not gc15 (wc15, n_1560);
  not gc14 (wc14, n_1684);
  or g3660 (n_552, wc16, wc17, n_372);
  not gc17 (wc17, n_1489);
  not gc16 (wc16, n_1748);
  or g3661 (n_580, wc18, wc19, n_393);
  not gc19 (wc19, n_1553);
  not gc18 (wc18, n_1812);
  or g3662 (n_608, wc20, wc21, n_418);
  not gc21 (wc21, n_1617);
  not gc20 (wc20, n_1876);
  xnor g3663 (n_3022, A[66], A[60]);
  or g3664 (n_3023, wc22, A[66]);
  not gc22 (wc22, A[60]);
  or g3665 (n_3025, wc23, A[66]);
  not gc23 (wc23, A[52]);
  xnor g3666 (n_3062, A[65], A[63]);
  or g3667 (n_3063, A[63], wc24);
  not gc24 (wc24, A[65]);
  or g3668 (n_3028, wc25, A[66]);
  not gc25 (wc25, A[58]);
  xnor g3669 (n_1174, n_3162, A[59]);
  or g3670 (n_3164, A[59], wc26);
  not gc26 (wc26, A[65]);
  or g3671 (n_3165, A[59], wc27);
  not gc27 (wc27, A[61]);
  xnor g3672 (n_3202, A[65], A[59]);
  or g3673 (n_3245, wc28, A[66]);
  not gc28 (wc28, A[62]);
  xnor g3674 (n_1220, n_3162, A[63]);
  or g3675 (n_3257, wc29, A[63]);
  not gc29 (wc29, A[61]);
  xnor g3676 (n_3262, A[66], A[62]);
  or g3677 (n_3265, wc30, A[66]);
  not gc30 (wc30, A[64]);
  xnor g3678 (n_3274, A[66], A[64]);
  or g3679 (n_3277, wc31, A[66]);
  not gc31 (wc31, A[63]);
  or g3680 (n_3700, wc32, A[66]);
  not gc32 (wc32, A[65]);
  xnor g3681 (n_3703, A[66], A[65]);
  or g3682 (n_424, wc33, wc34, n_333);
  not gc34 (wc34, n_1436);
  not gc33 (wc33, n_1437);
  or g3683 (n_3121, A[63], wc35);
  not gc35 (wc35, n_1148);
  or g3684 (n_3237, A[63], wc36);
  not gc36 (wc36, n_1208);
  xnor g3685 (n_1108, n_3026, A[66]);
  or g3686 (n_3029, wc37, A[66]);
  not gc37 (wc37, A[50]);
  or g3687 (n_3064, A[63], wc38);
  not gc38 (wc38, n_1119);
  xnor g3688 (n_3118, n_1119, A[63]);
  or g3689 (n_3204, A[59], wc39);
  not gc39 (wc39, n_1171);
  xnor g3690 (n_3234, n_1171, A[63]);
  or g3691 (n_3235, A[63], wc40);
  not gc40 (wc40, n_1171);
  or g3692 (n_3272, A[63], wc41);
  not gc41 (wc41, n_1227);
  or g3693 (n_3695, A[65], wc42);
  not gc42 (wc42, n_156);
  xnor g3694 (n_3698, n_156, A[65]);
  or g3696 (n_3296, wc43, n_1235);
  not gc43 (wc43, A[3]);
  or g3697 (n_3297, wc44, n_1235);
  not gc44 (wc44, A[1]);
  xnor g3698 (Z[3], n_1235, n_1402);
  or g3699 (n_3696, A[65], wc45);
  not gc45 (wc45, n_3694);
  or g3700 (n_3701, A[66], wc46);
  not gc46 (wc46, n_3699);
  not g3701 (Z[85], n_3704);
endmodule

module mult_signed_const_16293_GENERIC(A, Z);
  input [66:0] A;
  output [85:0] Z;
  wire [66:0] A;
  wire [85:0] Z;
  mult_signed_const_16293_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_16824_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [66:0] A;
  output [85:0] Z;
  wire [66:0] A;
  wire [85:0] Z;
  wire n_71, n_72, n_73, n_74, n_75, n_76, n_77, n_78;
  wire n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176;
  wire n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184;
  wire n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192;
  wire n_193, n_194, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_327, n_328, n_329;
  wire n_330, n_331, n_332, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353;
  wire n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361;
  wire n_362, n_363, n_364, n_365, n_366, n_367, n_368, n_369;
  wire n_370, n_371, n_372, n_373, n_374, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_386, n_387;
  wire n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395;
  wire n_397, n_399, n_400, n_401, n_402, n_403, n_404, n_405;
  wire n_406, n_407, n_408, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_513;
  wire n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593;
  wire n_594, n_595, n_596, n_597, n_598, n_599, n_600, n_601;
  wire n_602, n_603, n_604, n_605, n_606, n_607, n_608, n_609;
  wire n_610, n_611, n_612, n_613, n_614, n_615, n_616, n_617;
  wire n_618, n_619, n_620, n_621, n_622, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_642, n_643, n_644, n_645, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_655, n_656, n_657;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_666, n_667, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681;
  wire n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_694, n_695, n_696, n_697;
  wire n_698, n_699, n_700, n_701, n_702, n_703, n_704, n_705;
  wire n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_714, n_715, n_716, n_717, n_718, n_719, n_720, n_721;
  wire n_722, n_723, n_724, n_725, n_726, n_727, n_728, n_729;
  wire n_730, n_731, n_732, n_733, n_734, n_735, n_736, n_737;
  wire n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745;
  wire n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753;
  wire n_754, n_755, n_756, n_757, n_758, n_759, n_760, n_761;
  wire n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769;
  wire n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777;
  wire n_778, n_779, n_780, n_781, n_782, n_783, n_784, n_785;
  wire n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793;
  wire n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801;
  wire n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809;
  wire n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817;
  wire n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825;
  wire n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833;
  wire n_834, n_835, n_836, n_837, n_838, n_839, n_840, n_841;
  wire n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865;
  wire n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873;
  wire n_874, n_875, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_895, n_896, n_897;
  wire n_898, n_899, n_900, n_901, n_902, n_903, n_904, n_905;
  wire n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913;
  wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
  wire n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929;
  wire n_930, n_931, n_932, n_933, n_934, n_935, n_936, n_937;
  wire n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945;
  wire n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953;
  wire n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961;
  wire n_962, n_963, n_964, n_965, n_966, n_967, n_968, n_969;
  wire n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977;
  wire n_978, n_979, n_980, n_981, n_982, n_983, n_984, n_985;
  wire n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993;
  wire n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001;
  wire n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009;
  wire n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017;
  wire n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025;
  wire n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033;
  wire n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041;
  wire n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049;
  wire n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057;
  wire n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065;
  wire n_1066, n_1067, n_1068, n_1071, n_1072, n_1073, n_1074, n_1075;
  wire n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083;
  wire n_1084, n_1089, n_1090, n_1091, n_1092, n_1094, n_1095, n_1096;
  wire n_1097, n_1098, n_1099, n_1100, n_1101, n_1103, n_1104, n_1105;
  wire n_1107, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115;
  wire n_1116, n_1119, n_1120, n_1122, n_1124, n_1125, n_1126, n_1127;
  wire n_1128, n_1129, n_1130, n_1131, n_1135, n_1137, n_1138, n_1139;
  wire n_1140, n_1141, n_1142, n_1143, n_1144, n_1148, n_1149, n_1150;
  wire n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1159;
  wire n_1160, n_1161, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168;
  wire n_1171, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179;
  wire n_1181, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1192;
  wire n_1193, n_1194, n_1195, n_1196, n_1197, n_1199, n_1200, n_1201;
  wire n_1202, n_1203, n_1204, n_1207, n_1208, n_1210, n_1211, n_1214;
  wire n_1215, n_1216, n_1219, n_1220, n_1221, n_1223, n_1224, n_1227;
  wire n_1230, n_1231, n_1232, n_1233, n_1235, n_1236, n_1237, n_1238;
  wire n_1239, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247;
  wire n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1257, n_1258;
  wire n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1268, n_1270;
  wire n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278;
  wire n_1279, n_1281, n_1282, n_1283, n_1286, n_1287, n_1288, n_1289;
  wire n_1290, n_1291, n_1292, n_1293, n_1296, n_1300, n_1301, n_1302;
  wire n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310;
  wire n_1311, n_1312, n_1313, n_1314, n_1316, n_1318, n_1319, n_1320;
  wire n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328;
  wire n_1329, n_1332, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343;
  wire n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351;
  wire n_1352, n_1353, n_1354, n_1360, n_1361, n_1362, n_1363, n_1364;
  wire n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372;
  wire n_1373, n_1376, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387;
  wire n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395;
  wire n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1410;
  wire n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418;
  wire n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426;
  wire n_1427, n_1428, n_1430, n_1431, n_1433, n_1436, n_1437, n_1438;
  wire n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446;
  wire n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454;
  wire n_1455, n_1456, n_1457, n_1458, n_1461, n_1466, n_1467, n_1468;
  wire n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476;
  wire n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484;
  wire n_1485, n_1486, n_1487, n_1488, n_1489, n_1493, n_1494, n_1495;
  wire n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504;
  wire n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512;
  wire n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520;
  wire n_1521, n_1524, n_1526, n_1529, n_1530, n_1531, n_1532, n_1533;
  wire n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541;
  wire n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1551, n_1552, n_1553, n_1558, n_1559, n_1560, n_1562;
  wire n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570;
  wire n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578;
  wire n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1588;
  wire n_1590, n_1591, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599;
  wire n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607;
  wire n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615;
  wire n_1616, n_1617, n_1622, n_1623, n_1626, n_1627, n_1628, n_1629;
  wire n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637;
  wire n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645;
  wire n_1646, n_1647, n_1648, n_1649, n_1654, n_1655, n_1658, n_1659;
  wire n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667;
  wire n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675;
  wire n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1684, n_1686;
  wire n_1687, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696;
  wire n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704;
  wire n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712;
  wire n_1713, n_1716, n_1718, n_1719, n_1722, n_1723, n_1724, n_1725;
  wire n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733;
  wire n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741;
  wire n_1742, n_1743, n_1744, n_1745, n_1748, n_1750, n_1751, n_1754;
  wire n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762;
  wire n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770;
  wire n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1780;
  wire n_1782, n_1783, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
  wire n_1808, n_1809, n_1812, n_1814, n_1815, n_1818, n_1819, n_1820;
  wire n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
  wire n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836;
  wire n_1837, n_1838, n_1839, n_1840, n_1841, n_1844, n_1846, n_1847;
  wire n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857;
  wire n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865;
  wire n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873;
  wire n_1876, n_1878, n_1879, n_1882, n_1883, n_1884, n_1885, n_1886;
  wire n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894;
  wire n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902;
  wire n_1903, n_1904, n_1905, n_1908, n_1910, n_1911, n_1914, n_1915;
  wire n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923;
  wire n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931;
  wire n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1940, n_1942;
  wire n_1943, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952;
  wire n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960;
  wire n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968;
  wire n_1969, n_1972, n_1974, n_1975, n_1978, n_1979, n_1980, n_1981;
  wire n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989;
  wire n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997;
  wire n_1998, n_1999, n_2000, n_2001, n_2004, n_2006, n_2007, n_2010;
  wire n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018;
  wire n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026;
  wire n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2036;
  wire n_2038, n_2039, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047;
  wire n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055;
  wire n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063;
  wire n_2064, n_2065, n_2068, n_2070, n_2071, n_2074, n_2075, n_2076;
  wire n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084;
  wire n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092;
  wire n_2093, n_2094, n_2095, n_2096, n_2097, n_2100, n_2102, n_2103;
  wire n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113;
  wire n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121;
  wire n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129;
  wire n_2132, n_2134, n_2135, n_2138, n_2139, n_2140, n_2141, n_2142;
  wire n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150;
  wire n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158;
  wire n_2159, n_2160, n_2161, n_2164, n_2166, n_2167, n_2170, n_2171;
  wire n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179;
  wire n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187;
  wire n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2196, n_2198;
  wire n_2199, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208;
  wire n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216;
  wire n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224;
  wire n_2225, n_2228, n_2230, n_2231, n_2234, n_2235, n_2236, n_2237;
  wire n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245;
  wire n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253;
  wire n_2254, n_2255, n_2256, n_2257, n_2260, n_2262, n_2263, n_2266;
  wire n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274;
  wire n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282;
  wire n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2292;
  wire n_2294, n_2295, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303;
  wire n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311;
  wire n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319;
  wire n_2320, n_2321, n_2324, n_2326, n_2327, n_2330, n_2331, n_2332;
  wire n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340;
  wire n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348;
  wire n_2349, n_2350, n_2351, n_2352, n_2353, n_2356, n_2358, n_2359;
  wire n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369;
  wire n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377;
  wire n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385;
  wire n_2388, n_2390, n_2391, n_2394, n_2395, n_2396, n_2397, n_2398;
  wire n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406;
  wire n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414;
  wire n_2415, n_2416, n_2417, n_2420, n_2422, n_2423, n_2426, n_2427;
  wire n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435;
  wire n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443;
  wire n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2452, n_2454;
  wire n_2455, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464;
  wire n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472;
  wire n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480;
  wire n_2481, n_2484, n_2486, n_2487, n_2490, n_2491, n_2492, n_2493;
  wire n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501;
  wire n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509;
  wire n_2510, n_2511, n_2512, n_2513, n_2516, n_2518, n_2519, n_2522;
  wire n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530;
  wire n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538;
  wire n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2548;
  wire n_2550, n_2551, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559;
  wire n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567;
  wire n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575;
  wire n_2576, n_2577, n_2580, n_2582, n_2583, n_2586, n_2587, n_2588;
  wire n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596;
  wire n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604;
  wire n_2605, n_2606, n_2607, n_2608, n_2609, n_2612, n_2614, n_2615;
  wire n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625;
  wire n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, n_2633;
  wire n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641;
  wire n_2644, n_2646, n_2647, n_2650, n_2651, n_2652, n_2653, n_2654;
  wire n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662;
  wire n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670;
  wire n_2671, n_2672, n_2673, n_2676, n_2678, n_2679, n_2682, n_2683;
  wire n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691;
  wire n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699;
  wire n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2708, n_2710;
  wire n_2711, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720;
  wire n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728;
  wire n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736;
  wire n_2737, n_2740, n_2742, n_2743, n_2746, n_2747, n_2748, n_2749;
  wire n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757;
  wire n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765;
  wire n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2774;
  wire n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784;
  wire n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792;
  wire n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800;
  wire n_2801, n_2802, n_2803, n_2804, n_2806, n_2809, n_2810, n_2811;
  wire n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819;
  wire n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827;
  wire n_2828, n_2829, n_2833, n_2834, n_2836, n_2840, n_2841, n_2842;
  wire n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850;
  wire n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, n_2858;
  wire n_2859, n_2860, n_2861, n_2865, n_2866, n_2868, n_2872, n_2873;
  wire n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881;
  wire n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889;
  wire n_2890, n_2891, n_2892, n_2893, n_2897, n_2902, n_2903, n_2904;
  wire n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912;
  wire n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920;
  wire n_2921, n_2922, n_2923, n_2924, n_2925, n_2929, n_2934, n_2935;
  wire n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943;
  wire n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951;
  wire n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959;
  wire n_2961, n_2962, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971;
  wire n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979;
  wire n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987;
  wire n_2988, n_2989, n_2992, n_2993, n_3002, n_3003, n_3004, n_3005;
  wire n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013;
  wire n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021;
  wire n_3022, n_3023, n_3025, n_3026, n_3027, n_3028, n_3034, n_3035;
  wire n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043;
  wire n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, n_3051;
  wire n_3052, n_3053, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067;
  wire n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075;
  wire n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3089, n_3090;
  wire n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099;
  wire n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107;
  wire n_3108, n_3109, n_3114, n_3116, n_3117, n_3118, n_3120, n_3121;
  wire n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129;
  wire n_3130, n_3131, n_3132, n_3133, n_3142, n_3144, n_3145, n_3146;
  wire n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154;
  wire n_3155, n_3156, n_3157, n_3160, n_3161, n_3162, n_3164, n_3165;
  wire n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, n_3173;
  wire n_3174, n_3175, n_3176, n_3177, n_3182, n_3185, n_3186, n_3187;
  wire n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195;
  wire n_3196, n_3197, n_3198, n_3201, n_3202, n_3204, n_3205, n_3206;
  wire n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3216;
  wire n_3217, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226;
  wire n_3227, n_3228, n_3229, n_3234, n_3235, n_3236, n_3237, n_3238;
  wire n_3239, n_3240, n_3241, n_3242, n_3243, n_3248, n_3249, n_3250;
  wire n_3251, n_3252, n_3253, n_3254, n_3256, n_3257, n_3258, n_3259;
  wire n_3260, n_3261, n_3265, n_3266, n_3267, n_3268, n_3269, n_3271;
  wire n_3272, n_3273, n_3276, n_3277, n_3296, n_3297, n_3299, n_3300;
  wire n_3301, n_3302, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309;
  wire n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317;
  wire n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325;
  wire n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333;
  wire n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341;
  wire n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, n_3348, n_3349;
  wire n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, n_3357;
  wire n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365;
  wire n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373;
  wire n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381;
  wire n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, n_3389;
  wire n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397;
  wire n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405;
  wire n_3406, n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413;
  wire n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, n_3420, n_3421;
  wire n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, n_3429;
  wire n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437;
  wire n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445;
  wire n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453;
  wire n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, n_3461;
  wire n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469;
  wire n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477;
  wire n_3478, n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485;
  wire n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, n_3492, n_3493;
  wire n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, n_3501;
  wire n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509;
  wire n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517;
  wire n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525;
  wire n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, n_3533;
  wire n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541;
  wire n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549;
  wire n_3550, n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557;
  wire n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, n_3564, n_3565;
  wire n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572, n_3573;
  wire n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581;
  wire n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, n_3589;
  wire n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, n_3596, n_3597;
  wire n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, n_3605;
  wire n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613;
  wire n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621;
  wire n_3622, n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629;
  wire n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, n_3636, n_3637;
  wire n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644, n_3645;
  wire n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653;
  wire n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661;
  wire n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3668, n_3669;
  wire n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, n_3677;
  wire n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685;
  wire n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693;
  wire n_3694, n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701;
  wire n_3702, n_3703, n_3704;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g532 (n_235, A[4], A[0]);
  and g2 (n_148, A[4], A[0]);
  xor g533 (n_1230, A[5], A[3]);
  xor g534 (n_234, n_1230, A[1]);
  nand g3 (n_1231, A[5], A[3]);
  nand g535 (n_1232, A[1], A[3]);
  nand g536 (n_1233, A[5], A[1]);
  nand g537 (n_147, n_1231, n_1232, n_1233);
  xor g538 (n_327, A[6], A[4]);
  and g539 (n_328, A[6], A[4]);
  xor g540 (Z[2], A[0], A[2]);
  xor g541 (n_233, Z[2], n_327);
  nand g542 (n_1235, A[0], A[2]);
  nand g4 (n_1236, n_327, A[2]);
  nand g5 (n_1237, A[0], n_327);
  nand g543 (n_146, n_1235, n_1236, n_1237);
  xor g544 (n_1238, A[7], A[5]);
  xor g545 (n_329, n_1238, A[1]);
  nand g546 (n_1239, A[7], A[5]);
  nand g548 (n_1241, A[7], A[1]);
  nand g6 (n_331, n_1239, n_1233, n_1241);
  xor g549 (n_1242, A[3], n_328);
  xor g550 (n_232, n_1242, n_329);
  nand g551 (n_1243, A[3], n_328);
  nand g552 (n_1244, n_329, n_328);
  nand g553 (n_1245, A[3], n_329);
  nand g554 (n_145, n_1243, n_1244, n_1245);
  xor g555 (n_330, A[8], A[6]);
  and g556 (n_333, A[8], A[6]);
  xor g557 (n_1246, A[4], A[2]);
  xor g558 (n_332, n_1246, A[0]);
  nand g559 (n_1247, A[4], A[2]);
  xor g563 (n_1250, n_330, n_331);
  xor g564 (n_231, n_1250, n_332);
  nand g565 (n_1251, n_330, n_331);
  nand g566 (n_1252, n_332, n_331);
  nand g567 (n_1253, n_330, n_332);
  nand g568 (n_144, n_1251, n_1252, n_1253);
  xor g569 (n_1254, A[9], A[7]);
  xor g570 (n_334, n_1254, A[5]);
  nand g571 (n_1255, A[9], A[7]);
  nand g573 (n_1257, A[9], A[5]);
  nand g574 (n_338, n_1255, n_1239, n_1257);
  xor g575 (n_1258, A[3], A[1]);
  xor g576 (n_336, n_1258, n_333);
  nand g578 (n_1260, n_333, A[1]);
  nand g579 (n_1261, A[3], n_333);
  nand g580 (n_340, n_1232, n_1260, n_1261);
  xor g581 (n_1262, n_334, n_335);
  xor g582 (n_230, n_1262, n_336);
  nand g583 (n_1263, n_334, n_335);
  nand g584 (n_1264, n_336, n_335);
  nand g585 (n_1265, n_334, n_336);
  nand g586 (n_143, n_1263, n_1264, n_1265);
  xor g587 (n_337, A[10], A[8]);
  and g588 (n_342, A[10], A[8]);
  xor g590 (n_339, n_327, A[2]);
  nand g592 (n_1268, A[2], A[6]);
  xor g595 (n_1270, A[0], n_337);
  xor g596 (n_341, n_1270, n_338);
  nand g597 (n_1271, A[0], n_337);
  nand g598 (n_1272, n_338, n_337);
  nand g599 (n_1273, A[0], n_338);
  nand g600 (n_346, n_1271, n_1272, n_1273);
  xor g601 (n_1274, n_339, n_340);
  xor g602 (n_229, n_1274, n_341);
  nand g603 (n_1275, n_339, n_340);
  nand g604 (n_1276, n_341, n_340);
  nand g605 (n_1277, n_339, n_341);
  nand g606 (n_142, n_1275, n_1276, n_1277);
  xor g607 (n_1278, A[11], A[9]);
  xor g608 (n_343, n_1278, A[5]);
  nand g609 (n_1279, A[11], A[9]);
  nand g611 (n_1281, A[11], A[5]);
  nand g612 (n_349, n_1279, n_1257, n_1281);
  xor g613 (n_1282, A[7], A[3]);
  xor g614 (n_345, n_1282, A[1]);
  nand g615 (n_1283, A[7], A[3]);
  nand g618 (n_350, n_1283, n_1232, n_1241);
  xor g619 (n_1286, n_342, n_343);
  xor g620 (n_347, n_1286, n_344);
  nand g621 (n_1287, n_342, n_343);
  nand g622 (n_1288, n_344, n_343);
  nand g623 (n_1289, n_342, n_344);
  nand g624 (n_353, n_1287, n_1288, n_1289);
  xor g625 (n_1290, n_345, n_346);
  xor g626 (n_228, n_1290, n_347);
  nand g627 (n_1291, n_345, n_346);
  nand g628 (n_1292, n_347, n_346);
  nand g629 (n_1293, n_345, n_347);
  nand g630 (n_141, n_1291, n_1292, n_1293);
  xor g631 (n_348, A[12], A[10]);
  and g632 (n_355, A[12], A[10]);
  xor g634 (n_351, n_327, A[8]);
  nand g636 (n_1296, A[8], A[4]);
  xor g640 (n_352, Z[2], n_348);
  nand g642 (n_1300, n_348, A[0]);
  nand g643 (n_1301, A[2], n_348);
  nand g644 (n_359, n_1235, n_1300, n_1301);
  xor g645 (n_1302, n_349, n_350);
  xor g646 (n_354, n_1302, n_351);
  nand g647 (n_1303, n_349, n_350);
  nand g648 (n_1304, n_351, n_350);
  nand g649 (n_1305, n_349, n_351);
  nand g650 (n_361, n_1303, n_1304, n_1305);
  xor g651 (n_1306, n_352, n_353);
  xor g652 (n_227, n_1306, n_354);
  nand g653 (n_1307, n_352, n_353);
  nand g654 (n_1308, n_354, n_353);
  nand g655 (n_1309, n_352, n_354);
  nand g656 (n_140, n_1307, n_1308, n_1309);
  xor g657 (n_1310, A[13], A[11]);
  xor g658 (n_358, n_1310, A[7]);
  nand g659 (n_1311, A[13], A[11]);
  nand g660 (n_1312, A[7], A[11]);
  nand g661 (n_1313, A[13], A[7]);
  nand g662 (n_364, n_1311, n_1312, n_1313);
  xor g663 (n_1314, A[5], A[9]);
  xor g664 (n_357, n_1314, A[3]);
  nand g666 (n_1316, A[3], A[9]);
  nand g668 (n_365, n_1257, n_1316, n_1231);
  xor g669 (n_1318, A[1], n_355);
  xor g670 (n_360, n_1318, n_356);
  nand g671 (n_1319, A[1], n_355);
  nand g672 (n_1320, n_356, n_355);
  nand g673 (n_1321, A[1], n_356);
  nand g674 (n_368, n_1319, n_1320, n_1321);
  xor g675 (n_1322, n_357, n_358);
  xor g676 (n_362, n_1322, n_359);
  nand g677 (n_1323, n_357, n_358);
  nand g678 (n_1324, n_359, n_358);
  nand g679 (n_1325, n_357, n_359);
  nand g680 (n_370, n_1323, n_1324, n_1325);
  xor g681 (n_1326, n_360, n_361);
  xor g682 (n_226, n_1326, n_362);
  nand g683 (n_1327, n_360, n_361);
  nand g684 (n_1328, n_362, n_361);
  nand g685 (n_1329, n_360, n_362);
  nand g686 (n_139, n_1327, n_1328, n_1329);
  xor g687 (n_363, A[14], A[12]);
  and g688 (n_372, A[14], A[12]);
  xor g690 (n_366, n_330, A[10]);
  nand g692 (n_1332, A[10], A[6]);
  xor g696 (n_367, n_235, A[2]);
  xor g701 (n_1338, n_363, n_364);
  xor g702 (n_369, n_1338, n_365);
  nand g703 (n_1339, n_363, n_364);
  nand g704 (n_1340, n_365, n_364);
  nand g705 (n_1341, n_363, n_365);
  nand g706 (n_378, n_1339, n_1340, n_1341);
  xor g707 (n_1342, n_366, n_367);
  xor g708 (n_371, n_1342, n_368);
  nand g709 (n_1343, n_366, n_367);
  nand g710 (n_1344, n_368, n_367);
  nand g711 (n_1345, n_366, n_368);
  nand g712 (n_380, n_1343, n_1344, n_1345);
  xor g713 (n_1346, n_369, n_370);
  xor g714 (n_225, n_1346, n_371);
  nand g715 (n_1347, n_369, n_370);
  nand g716 (n_1348, n_371, n_370);
  nand g717 (n_1349, n_369, n_371);
  nand g718 (n_138, n_1347, n_1348, n_1349);
  xor g719 (n_1350, A[15], A[13]);
  xor g720 (n_376, n_1350, A[9]);
  nand g721 (n_1351, A[15], A[13]);
  nand g722 (n_1352, A[9], A[13]);
  nand g723 (n_1353, A[15], A[9]);
  nand g724 (n_384, n_1351, n_1352, n_1353);
  xor g725 (n_1354, A[7], A[11]);
  xor g726 (n_374, n_1354, A[5]);
  nand g730 (n_383, n_1312, n_1281, n_1239);
  xor g732 (n_377, n_1258, n_372);
  nand g734 (n_1360, n_372, A[3]);
  nand g735 (n_1361, A[1], n_372);
  nand g736 (n_387, n_1232, n_1360, n_1361);
  xor g737 (n_1362, n_373, n_374);
  xor g738 (n_379, n_1362, n_335);
  nand g739 (n_1363, n_373, n_374);
  nand g740 (n_1364, n_335, n_374);
  nand g741 (n_1365, n_373, n_335);
  nand g742 (n_389, n_1363, n_1364, n_1365);
  xor g743 (n_1366, n_376, n_377);
  xor g744 (n_381, n_1366, n_378);
  nand g745 (n_1367, n_376, n_377);
  nand g746 (n_1368, n_378, n_377);
  nand g747 (n_1369, n_376, n_378);
  nand g748 (n_392, n_1367, n_1368, n_1369);
  xor g749 (n_1370, n_379, n_380);
  xor g750 (n_224, n_1370, n_381);
  nand g751 (n_1371, n_379, n_380);
  nand g752 (n_1372, n_381, n_380);
  nand g753 (n_1373, n_379, n_381);
  nand g754 (n_137, n_1371, n_1372, n_1373);
  xor g755 (n_382, A[16], A[14]);
  and g756 (n_393, A[16], A[14]);
  xor g758 (n_386, n_337, A[12]);
  nand g760 (n_1376, A[12], A[8]);
  xor g769 (n_1382, A[0], n_382);
  xor g770 (n_388, n_1382, n_383);
  nand g771 (n_1383, A[0], n_382);
  nand g772 (n_1384, n_383, n_382);
  nand g773 (n_1385, A[0], n_383);
  nand g774 (n_399, n_1383, n_1384, n_1385);
  xor g775 (n_1386, n_384, n_339);
  xor g776 (n_390, n_1386, n_386);
  nand g777 (n_1387, n_384, n_339);
  nand g778 (n_1388, n_386, n_339);
  nand g779 (n_1389, n_384, n_386);
  nand g780 (n_401, n_1387, n_1388, n_1389);
  xor g781 (n_1390, n_387, n_388);
  xor g782 (n_391, n_1390, n_389);
  nand g783 (n_1391, n_387, n_388);
  nand g784 (n_1392, n_389, n_388);
  nand g785 (n_1393, n_387, n_389);
  nand g786 (n_403, n_1391, n_1392, n_1393);
  xor g787 (n_1394, n_390, n_391);
  xor g788 (n_223, n_1394, n_392);
  nand g789 (n_1395, n_390, n_391);
  nand g790 (n_1396, n_392, n_391);
  nand g791 (n_1397, n_390, n_392);
  nand g792 (n_136, n_1395, n_1396, n_1397);
  xor g793 (n_1398, A[17], A[15]);
  xor g794 (n_397, n_1398, A[11]);
  nand g795 (n_1399, A[17], A[15]);
  nand g796 (n_1400, A[11], A[15]);
  nand g797 (n_1401, A[17], A[11]);
  nand g798 (n_406, n_1399, n_1400, n_1401);
  xor g799 (n_1402, A[9], A[13]);
  xor g800 (n_395, n_1402, A[7]);
  nand g804 (n_407, n_1352, n_1313, n_1255);
  xor g811 (n_1410, n_393, n_394);
  xor g812 (n_400, n_1410, n_395);
  nand g813 (n_1411, n_393, n_394);
  nand g814 (n_1412, n_395, n_394);
  nand g815 (n_1413, n_393, n_395);
  nand g816 (n_413, n_1411, n_1412, n_1413);
  xor g817 (n_1414, n_344, n_397);
  xor g818 (n_402, n_1414, n_234);
  nand g819 (n_1415, n_344, n_397);
  nand g820 (n_1416, n_234, n_397);
  nand g821 (n_1417, n_344, n_234);
  nand g822 (n_414, n_1415, n_1416, n_1417);
  xor g823 (n_1418, n_399, n_400);
  xor g824 (n_404, n_1418, n_401);
  nand g825 (n_1419, n_399, n_400);
  nand g826 (n_1420, n_401, n_400);
  nand g827 (n_1421, n_399, n_401);
  nand g828 (n_416, n_1419, n_1420, n_1421);
  xor g829 (n_1422, n_402, n_403);
  xor g830 (n_222, n_1422, n_404);
  nand g831 (n_1423, n_402, n_403);
  nand g832 (n_1424, n_404, n_403);
  nand g833 (n_1425, n_402, n_404);
  nand g834 (n_135, n_1423, n_1424, n_1425);
  xor g835 (n_405, A[18], A[16]);
  and g836 (n_418, A[18], A[16]);
  xor g837 (n_1426, A[12], A[4]);
  xor g838 (n_410, n_1426, A[10]);
  nand g839 (n_1427, A[12], A[4]);
  nand g840 (n_1428, A[10], A[4]);
  xor g843 (n_1430, A[14], A[8]);
  xor g844 (n_408, n_1430, A[6]);
  nand g845 (n_1431, A[14], A[8]);
  nand g847 (n_1433, A[14], A[6]);
  xor g850 (n_411, Z[2], n_405);
  nand g852 (n_1436, n_405, A[0]);
  nand g853 (n_1437, A[2], n_405);
  nand g854 (n_424, n_1235, n_1436, n_1437);
  xor g855 (n_1438, n_406, n_407);
  xor g856 (n_412, n_1438, n_408);
  nand g857 (n_1439, n_406, n_407);
  nand g858 (n_1440, n_408, n_407);
  nand g859 (n_1441, n_406, n_408);
  nand g860 (n_426, n_1439, n_1440, n_1441);
  xor g861 (n_1442, n_147, n_410);
  xor g862 (n_415, n_1442, n_411);
  nand g863 (n_1443, n_147, n_410);
  nand g864 (n_1444, n_411, n_410);
  nand g865 (n_1445, n_147, n_411);
  nand g866 (n_428, n_1443, n_1444, n_1445);
  xor g867 (n_1446, n_412, n_413);
  xor g868 (n_417, n_1446, n_414);
  nand g869 (n_1447, n_412, n_413);
  nand g870 (n_1448, n_414, n_413);
  nand g871 (n_1449, n_412, n_414);
  nand g872 (n_430, n_1447, n_1448, n_1449);
  xor g873 (n_1450, n_415, n_416);
  xor g874 (n_221, n_1450, n_417);
  nand g875 (n_1451, n_415, n_416);
  nand g876 (n_1452, n_417, n_416);
  nand g877 (n_1453, n_415, n_417);
  nand g878 (n_134, n_1451, n_1452, n_1453);
  xor g879 (n_1454, A[19], A[17]);
  xor g880 (n_422, n_1454, A[13]);
  nand g881 (n_1455, A[19], A[17]);
  nand g882 (n_1456, A[13], A[17]);
  nand g883 (n_1457, A[19], A[13]);
  nand g884 (n_432, n_1455, n_1456, n_1457);
  xor g885 (n_1458, A[5], A[11]);
  xor g886 (n_423, n_1458, A[15]);
  nand g889 (n_1461, A[5], A[15]);
  nand g890 (n_433, n_1281, n_1400, n_1461);
  xor g892 (n_421, n_1254, A[3]);
  nand g896 (n_436, n_1255, n_1283, n_1316);
  xor g897 (n_1466, A[1], n_418);
  xor g898 (n_425, n_1466, n_419);
  nand g899 (n_1467, A[1], n_418);
  nand g900 (n_1468, n_419, n_418);
  nand g901 (n_1469, A[1], n_419);
  nand g902 (n_438, n_1467, n_1468, n_1469);
  xor g903 (n_1470, n_420, n_421);
  xor g904 (n_427, n_1470, n_422);
  nand g905 (n_1471, n_420, n_421);
  nand g906 (n_1472, n_422, n_421);
  nand g907 (n_1473, n_420, n_422);
  nand g908 (n_440, n_1471, n_1472, n_1473);
  xor g909 (n_1474, n_423, n_424);
  xor g910 (n_429, n_1474, n_425);
  nand g911 (n_1475, n_423, n_424);
  nand g912 (n_1476, n_425, n_424);
  nand g913 (n_1477, n_423, n_425);
  nand g914 (n_442, n_1475, n_1476, n_1477);
  xor g915 (n_1478, n_426, n_427);
  xor g916 (n_431, n_1478, n_428);
  nand g917 (n_1479, n_426, n_427);
  nand g918 (n_1480, n_428, n_427);
  nand g919 (n_1481, n_426, n_428);
  nand g920 (n_444, n_1479, n_1480, n_1481);
  xor g921 (n_1482, n_429, n_430);
  xor g922 (n_220, n_1482, n_431);
  nand g923 (n_1483, n_429, n_430);
  nand g924 (n_1484, n_431, n_430);
  nand g925 (n_1485, n_429, n_431);
  nand g926 (n_133, n_1483, n_1484, n_1485);
  xor g927 (n_1486, A[20], A[18]);
  xor g928 (n_435, n_1486, A[14]);
  nand g929 (n_1487, A[20], A[18]);
  nand g930 (n_1488, A[14], A[18]);
  nand g931 (n_1489, A[20], A[14]);
  nand g932 (n_446, n_1487, n_1488, n_1489);
  xor g934 (n_437, n_327, A[12]);
  nand g937 (n_1493, A[6], A[12]);
  xor g939 (n_1494, A[16], A[10]);
  xor g940 (n_434, n_1494, A[8]);
  nand g941 (n_1495, A[16], A[10]);
  nand g943 (n_1497, A[16], A[8]);
  xor g945 (n_1498, A[2], n_432);
  xor g946 (n_439, n_1498, n_433);
  nand g947 (n_1499, A[2], n_432);
  nand g948 (n_1500, n_433, n_432);
  nand g949 (n_1501, A[2], n_433);
  nand g950 (n_149, n_1499, n_1500, n_1501);
  xor g951 (n_1502, n_434, n_435);
  xor g952 (n_441, n_1502, n_436);
  nand g953 (n_1503, n_434, n_435);
  nand g954 (n_1504, n_436, n_435);
  nand g955 (n_1505, n_434, n_436);
  nand g956 (n_151, n_1503, n_1504, n_1505);
  xor g957 (n_1506, n_437, n_438);
  xor g958 (n_443, n_1506, n_439);
  nand g959 (n_1507, n_437, n_438);
  nand g960 (n_1508, n_439, n_438);
  nand g961 (n_1509, n_437, n_439);
  nand g962 (n_452, n_1507, n_1508, n_1509);
  xor g963 (n_1510, n_440, n_441);
  xor g964 (n_445, n_1510, n_442);
  nand g965 (n_1511, n_440, n_441);
  nand g966 (n_1512, n_442, n_441);
  nand g967 (n_1513, n_440, n_442);
  nand g968 (n_453, n_1511, n_1512, n_1513);
  xor g969 (n_1514, n_443, n_444);
  xor g970 (n_219, n_1514, n_445);
  nand g971 (n_1515, n_443, n_444);
  nand g972 (n_1516, n_445, n_444);
  nand g973 (n_1517, n_443, n_445);
  nand g974 (n_132, n_1515, n_1516, n_1517);
  xor g975 (n_1518, A[21], A[19]);
  xor g976 (n_450, n_1518, A[15]);
  nand g977 (n_1519, A[21], A[19]);
  nand g978 (n_1520, A[15], A[19]);
  nand g979 (n_1521, A[21], A[15]);
  nand g980 (n_455, n_1519, n_1520, n_1521);
  xor g982 (n_451, n_1238, A[13]);
  nand g984 (n_1524, A[13], A[5]);
  nand g986 (n_456, n_1239, n_1524, n_1313);
  xor g987 (n_1526, A[17], A[11]);
  xor g988 (n_449, n_1526, A[9]);
  nand g991 (n_1529, A[17], A[9]);
  nand g992 (n_457, n_1401, n_1279, n_1529);
  xor g993 (n_1530, A[3], n_446);
  xor g994 (n_150, n_1530, n_447);
  nand g995 (n_1531, A[3], n_446);
  nand g996 (n_1532, n_447, n_446);
  nand g997 (n_1533, A[3], n_447);
  nand g998 (n_461, n_1531, n_1532, n_1533);
  xor g999 (n_1534, n_448, n_449);
  xor g1000 (n_152, n_1534, n_450);
  nand g1001 (n_1535, n_448, n_449);
  nand g1002 (n_1536, n_450, n_449);
  nand g1003 (n_1537, n_448, n_450);
  nand g1004 (n_463, n_1535, n_1536, n_1537);
  xor g1005 (n_1538, n_451, n_149);
  xor g1006 (n_153, n_1538, n_150);
  nand g1007 (n_1539, n_451, n_149);
  nand g1008 (n_1540, n_150, n_149);
  nand g1009 (n_1541, n_451, n_150);
  nand g1010 (n_465, n_1539, n_1540, n_1541);
  xor g1011 (n_1542, n_151, n_152);
  xor g1012 (n_454, n_1542, n_153);
  nand g1013 (n_1543, n_151, n_152);
  nand g1014 (n_1544, n_153, n_152);
  nand g1015 (n_1545, n_151, n_153);
  nand g1016 (n_468, n_1543, n_1544, n_1545);
  xor g1017 (n_1546, n_452, n_453);
  xor g1018 (n_218, n_1546, n_454);
  nand g1019 (n_1547, n_452, n_453);
  nand g1020 (n_1548, n_454, n_453);
  nand g1021 (n_1549, n_452, n_454);
  nand g1022 (n_131, n_1547, n_1548, n_1549);
  xor g1023 (n_1550, A[22], A[20]);
  xor g1024 (n_459, n_1550, A[16]);
  nand g1025 (n_1551, A[22], A[20]);
  nand g1026 (n_1552, A[16], A[20]);
  nand g1027 (n_1553, A[22], A[16]);
  nand g1028 (n_469, n_1551, n_1552, n_1553);
  xor g1030 (n_460, n_330, A[14]);
  xor g1035 (n_1558, A[4], A[18]);
  xor g1036 (n_458, n_1558, A[12]);
  nand g1037 (n_1559, A[4], A[18]);
  nand g1038 (n_1560, A[12], A[18]);
  nand g1040 (n_471, n_1559, n_1560, n_1427);
  xor g1041 (n_1562, A[10], n_455);
  xor g1042 (n_462, n_1562, n_456);
  nand g1043 (n_1563, A[10], n_455);
  nand g1044 (n_1564, n_456, n_455);
  nand g1045 (n_1565, A[10], n_456);
  nand g1046 (n_475, n_1563, n_1564, n_1565);
  xor g1047 (n_1566, n_457, n_458);
  xor g1048 (n_464, n_1566, n_459);
  nand g1049 (n_1567, n_457, n_458);
  nand g1050 (n_1568, n_459, n_458);
  nand g1051 (n_1569, n_457, n_459);
  nand g1052 (n_477, n_1567, n_1568, n_1569);
  xor g1053 (n_1570, n_460, n_461);
  xor g1054 (n_466, n_1570, n_462);
  nand g1055 (n_1571, n_460, n_461);
  nand g1056 (n_1572, n_462, n_461);
  nand g1057 (n_1573, n_460, n_462);
  nand g1058 (n_479, n_1571, n_1572, n_1573);
  xor g1059 (n_1574, n_463, n_464);
  xor g1060 (n_467, n_1574, n_465);
  nand g1061 (n_1575, n_463, n_464);
  nand g1062 (n_1576, n_465, n_464);
  nand g1063 (n_1577, n_463, n_465);
  nand g1064 (n_482, n_1575, n_1576, n_1577);
  xor g1065 (n_1578, n_466, n_467);
  xor g1066 (n_217, n_1578, n_468);
  nand g1067 (n_1579, n_466, n_467);
  nand g1068 (n_1580, n_468, n_467);
  nand g1069 (n_1581, n_466, n_468);
  nand g1070 (n_130, n_1579, n_1580, n_1581);
  xor g1071 (n_1582, A[23], A[21]);
  xor g1072 (n_473, n_1582, A[17]);
  nand g1073 (n_1583, A[23], A[21]);
  nand g1074 (n_1584, A[17], A[21]);
  nand g1075 (n_1585, A[23], A[17]);
  nand g1076 (n_483, n_1583, n_1584, n_1585);
  xor g1078 (n_474, n_1254, A[15]);
  nand g1080 (n_1588, A[15], A[7]);
  nand g1082 (n_484, n_1255, n_1588, n_1353);
  xor g1083 (n_1590, A[5], A[19]);
  xor g1084 (n_472, n_1590, A[13]);
  nand g1085 (n_1591, A[5], A[19]);
  nand g1088 (n_485, n_1591, n_1457, n_1524);
  xor g1089 (n_1594, A[11], n_469);
  xor g1090 (n_476, n_1594, n_420);
  nand g1091 (n_1595, A[11], n_469);
  nand g1092 (n_1596, n_420, n_469);
  nand g1093 (n_1597, A[11], n_420);
  nand g1094 (n_489, n_1595, n_1596, n_1597);
  xor g1095 (n_1598, n_471, n_472);
  xor g1096 (n_478, n_1598, n_473);
  nand g1097 (n_1599, n_471, n_472);
  nand g1098 (n_1600, n_473, n_472);
  nand g1099 (n_1601, n_471, n_473);
  nand g1100 (n_491, n_1599, n_1600, n_1601);
  xor g1101 (n_1602, n_474, n_475);
  xor g1102 (n_480, n_1602, n_476);
  nand g1103 (n_1603, n_474, n_475);
  nand g1104 (n_1604, n_476, n_475);
  nand g1105 (n_1605, n_474, n_476);
  nand g1106 (n_493, n_1603, n_1604, n_1605);
  xor g1107 (n_1606, n_477, n_478);
  xor g1108 (n_481, n_1606, n_479);
  nand g1109 (n_1607, n_477, n_478);
  nand g1110 (n_1608, n_479, n_478);
  nand g1111 (n_1609, n_477, n_479);
  nand g1112 (n_496, n_1607, n_1608, n_1609);
  xor g1113 (n_1610, n_480, n_481);
  xor g1114 (n_216, n_1610, n_482);
  nand g1115 (n_1611, n_480, n_481);
  nand g1116 (n_1612, n_482, n_481);
  nand g1117 (n_1613, n_480, n_482);
  nand g1118 (n_129, n_1611, n_1612, n_1613);
  xor g1119 (n_1614, A[24], A[22]);
  xor g1120 (n_487, n_1614, A[18]);
  nand g1121 (n_1615, A[24], A[22]);
  nand g1122 (n_1616, A[18], A[22]);
  nand g1123 (n_1617, A[24], A[18]);
  nand g1124 (n_497, n_1615, n_1616, n_1617);
  xor g1126 (n_488, n_337, A[16]);
  xor g1131 (n_1622, A[6], A[20]);
  xor g1132 (n_486, n_1622, A[14]);
  nand g1133 (n_1623, A[6], A[20]);
  nand g1136 (n_499, n_1623, n_1489, n_1433);
  xor g1137 (n_1626, A[12], n_483);
  xor g1138 (n_490, n_1626, n_484);
  nand g1139 (n_1627, A[12], n_483);
  nand g1140 (n_1628, n_484, n_483);
  nand g1141 (n_1629, A[12], n_484);
  nand g1142 (n_503, n_1627, n_1628, n_1629);
  xor g1143 (n_1630, n_485, n_486);
  xor g1144 (n_492, n_1630, n_487);
  nand g1145 (n_1631, n_485, n_486);
  nand g1146 (n_1632, n_487, n_486);
  nand g1147 (n_1633, n_485, n_487);
  nand g1148 (n_505, n_1631, n_1632, n_1633);
  xor g1149 (n_1634, n_488, n_489);
  xor g1150 (n_494, n_1634, n_490);
  nand g1151 (n_1635, n_488, n_489);
  nand g1152 (n_1636, n_490, n_489);
  nand g1153 (n_1637, n_488, n_490);
  nand g1154 (n_507, n_1635, n_1636, n_1637);
  xor g1155 (n_1638, n_491, n_492);
  xor g1156 (n_495, n_1638, n_493);
  nand g1157 (n_1639, n_491, n_492);
  nand g1158 (n_1640, n_493, n_492);
  nand g1159 (n_1641, n_491, n_493);
  nand g1160 (n_510, n_1639, n_1640, n_1641);
  xor g1161 (n_1642, n_494, n_495);
  xor g1162 (n_215, n_1642, n_496);
  nand g1163 (n_1643, n_494, n_495);
  nand g1164 (n_1644, n_496, n_495);
  nand g1165 (n_1645, n_494, n_496);
  nand g1166 (n_128, n_1643, n_1644, n_1645);
  xor g1167 (n_1646, A[25], A[23]);
  xor g1168 (n_501, n_1646, A[19]);
  nand g1169 (n_1647, A[25], A[23]);
  nand g1170 (n_1648, A[19], A[23]);
  nand g1171 (n_1649, A[25], A[19]);
  nand g1172 (n_511, n_1647, n_1648, n_1649);
  xor g1174 (n_502, n_1278, A[17]);
  xor g1179 (n_1654, A[7], A[21]);
  xor g1180 (n_500, n_1654, A[15]);
  nand g1181 (n_1655, A[7], A[21]);
  nand g1184 (n_513, n_1655, n_1521, n_1588);
  xor g1185 (n_1658, A[13], n_497);
  xor g1186 (n_504, n_1658, n_447);
  nand g1187 (n_1659, A[13], n_497);
  nand g1188 (n_1660, n_447, n_497);
  nand g1189 (n_1661, A[13], n_447);
  nand g1190 (n_517, n_1659, n_1660, n_1661);
  xor g1191 (n_1662, n_499, n_500);
  xor g1192 (n_506, n_1662, n_501);
  nand g1193 (n_1663, n_499, n_500);
  nand g1194 (n_1664, n_501, n_500);
  nand g1195 (n_1665, n_499, n_501);
  nand g1196 (n_519, n_1663, n_1664, n_1665);
  xor g1197 (n_1666, n_502, n_503);
  xor g1198 (n_508, n_1666, n_504);
  nand g1199 (n_1667, n_502, n_503);
  nand g1200 (n_1668, n_504, n_503);
  nand g1201 (n_1669, n_502, n_504);
  nand g1202 (n_521, n_1667, n_1668, n_1669);
  xor g1203 (n_1670, n_505, n_506);
  xor g1204 (n_509, n_1670, n_507);
  nand g1205 (n_1671, n_505, n_506);
  nand g1206 (n_1672, n_507, n_506);
  nand g1207 (n_1673, n_505, n_507);
  nand g1208 (n_524, n_1671, n_1672, n_1673);
  xor g1209 (n_1674, n_508, n_509);
  xor g1210 (n_214, n_1674, n_510);
  nand g1211 (n_1675, n_508, n_509);
  nand g1212 (n_1676, n_510, n_509);
  nand g1213 (n_1677, n_508, n_510);
  nand g1214 (n_127, n_1675, n_1676, n_1677);
  xor g1215 (n_1678, A[26], A[24]);
  xor g1216 (n_515, n_1678, A[20]);
  nand g1217 (n_1679, A[26], A[24]);
  nand g1218 (n_1680, A[20], A[24]);
  nand g1219 (n_1681, A[26], A[20]);
  nand g1220 (n_525, n_1679, n_1680, n_1681);
  xor g1222 (n_516, n_348, A[18]);
  nand g1224 (n_1684, A[18], A[10]);
  xor g1227 (n_1686, A[8], A[22]);
  xor g1228 (n_514, n_1686, A[16]);
  nand g1229 (n_1687, A[8], A[22]);
  nand g1232 (n_527, n_1687, n_1553, n_1497);
  xor g1233 (n_1690, A[14], n_511);
  xor g1234 (n_518, n_1690, n_457);
  nand g1235 (n_1691, A[14], n_511);
  nand g1236 (n_1692, n_457, n_511);
  nand g1237 (n_1693, A[14], n_457);
  nand g1238 (n_529, n_1691, n_1692, n_1693);
  xor g1239 (n_1694, n_513, n_514);
  xor g1240 (n_520, n_1694, n_515);
  nand g1241 (n_1695, n_513, n_514);
  nand g1242 (n_1696, n_515, n_514);
  nand g1243 (n_1697, n_513, n_515);
  nand g1244 (n_531, n_1695, n_1696, n_1697);
  xor g1245 (n_1698, n_516, n_517);
  xor g1246 (n_522, n_1698, n_518);
  nand g1247 (n_1699, n_516, n_517);
  nand g1248 (n_1700, n_518, n_517);
  nand g1249 (n_1701, n_516, n_518);
  nand g1250 (n_533, n_1699, n_1700, n_1701);
  xor g1251 (n_1702, n_519, n_520);
  xor g1252 (n_523, n_1702, n_521);
  nand g1253 (n_1703, n_519, n_520);
  nand g1254 (n_1704, n_521, n_520);
  nand g1255 (n_1705, n_519, n_521);
  nand g1256 (n_536, n_1703, n_1704, n_1705);
  xor g1257 (n_1706, n_522, n_523);
  xor g1258 (n_213, n_1706, n_524);
  nand g1259 (n_1707, n_522, n_523);
  nand g1260 (n_1708, n_524, n_523);
  nand g1261 (n_1709, n_522, n_524);
  nand g1262 (n_126, n_1707, n_1708, n_1709);
  xor g1263 (n_1710, A[27], A[25]);
  xor g1264 (n_237, n_1710, A[21]);
  nand g1265 (n_1711, A[27], A[25]);
  nand g1266 (n_1712, A[21], A[25]);
  nand g1267 (n_1713, A[27], A[21]);
  nand g1268 (n_537, n_1711, n_1712, n_1713);
  xor g1270 (n_528, n_1310, A[19]);
  nand g1272 (n_1716, A[19], A[11]);
  nand g1274 (n_538, n_1311, n_1716, n_1457);
  xor g1275 (n_1718, A[9], A[23]);
  xor g1276 (n_236, n_1718, A[17]);
  nand g1277 (n_1719, A[9], A[23]);
  nand g1280 (n_539, n_1719, n_1585, n_1529);
  xor g1281 (n_1722, A[15], n_525);
  xor g1282 (n_530, n_1722, n_526);
  nand g1283 (n_1723, A[15], n_525);
  nand g1284 (n_1724, n_526, n_525);
  nand g1285 (n_1725, A[15], n_526);
  nand g1286 (n_543, n_1723, n_1724, n_1725);
  xor g1287 (n_1726, n_527, n_236);
  xor g1288 (n_532, n_1726, n_237);
  nand g1289 (n_1727, n_527, n_236);
  nand g1290 (n_1728, n_237, n_236);
  nand g1291 (n_1729, n_527, n_237);
  nand g1292 (n_545, n_1727, n_1728, n_1729);
  xor g1293 (n_1730, n_528, n_529);
  xor g1294 (n_534, n_1730, n_530);
  nand g1295 (n_1731, n_528, n_529);
  nand g1296 (n_1732, n_530, n_529);
  nand g1297 (n_1733, n_528, n_530);
  nand g1298 (n_547, n_1731, n_1732, n_1733);
  xor g1299 (n_1734, n_531, n_532);
  xor g1300 (n_535, n_1734, n_533);
  nand g1301 (n_1735, n_531, n_532);
  nand g1302 (n_1736, n_533, n_532);
  nand g1303 (n_1737, n_531, n_533);
  nand g1304 (n_550, n_1735, n_1736, n_1737);
  xor g1305 (n_1738, n_534, n_535);
  xor g1306 (n_212, n_1738, n_536);
  nand g1307 (n_1739, n_534, n_535);
  nand g1308 (n_1740, n_536, n_535);
  nand g1309 (n_1741, n_534, n_536);
  nand g1310 (n_125, n_1739, n_1740, n_1741);
  xor g1311 (n_1742, A[28], A[26]);
  xor g1312 (n_541, n_1742, A[22]);
  nand g1313 (n_1743, A[28], A[26]);
  nand g1314 (n_1744, A[22], A[26]);
  nand g1315 (n_1745, A[28], A[22]);
  nand g1316 (n_551, n_1743, n_1744, n_1745);
  xor g1318 (n_542, n_363, A[20]);
  nand g1320 (n_1748, A[20], A[12]);
  xor g1323 (n_1750, A[10], A[24]);
  xor g1324 (n_540, n_1750, A[18]);
  nand g1325 (n_1751, A[10], A[24]);
  nand g1328 (n_553, n_1751, n_1617, n_1684);
  xor g1329 (n_1754, A[16], n_537);
  xor g1330 (n_544, n_1754, n_538);
  nand g1331 (n_1755, A[16], n_537);
  nand g1332 (n_1756, n_538, n_537);
  nand g1333 (n_1757, A[16], n_538);
  nand g1334 (n_557, n_1755, n_1756, n_1757);
  xor g1335 (n_1758, n_539, n_540);
  xor g1336 (n_546, n_1758, n_541);
  nand g1337 (n_1759, n_539, n_540);
  nand g1338 (n_1760, n_541, n_540);
  nand g1339 (n_1761, n_539, n_541);
  nand g1340 (n_559, n_1759, n_1760, n_1761);
  xor g1341 (n_1762, n_542, n_543);
  xor g1342 (n_548, n_1762, n_544);
  nand g1343 (n_1763, n_542, n_543);
  nand g1344 (n_1764, n_544, n_543);
  nand g1345 (n_1765, n_542, n_544);
  nand g1346 (n_561, n_1763, n_1764, n_1765);
  xor g1347 (n_1766, n_545, n_546);
  xor g1348 (n_549, n_1766, n_547);
  nand g1349 (n_1767, n_545, n_546);
  nand g1350 (n_1768, n_547, n_546);
  nand g1351 (n_1769, n_545, n_547);
  nand g1352 (n_564, n_1767, n_1768, n_1769);
  xor g1353 (n_1770, n_548, n_549);
  xor g1354 (n_211, n_1770, n_550);
  nand g1355 (n_1771, n_548, n_549);
  nand g1356 (n_1772, n_550, n_549);
  nand g1357 (n_1773, n_548, n_550);
  nand g1358 (n_124, n_1771, n_1772, n_1773);
  xor g1359 (n_1774, A[29], A[27]);
  xor g1360 (n_555, n_1774, A[23]);
  nand g1361 (n_1775, A[29], A[27]);
  nand g1362 (n_1776, A[23], A[27]);
  nand g1363 (n_1777, A[29], A[23]);
  nand g1364 (n_565, n_1775, n_1776, n_1777);
  xor g1366 (n_556, n_1350, A[21]);
  nand g1368 (n_1780, A[21], A[13]);
  nand g1370 (n_566, n_1351, n_1780, n_1521);
  xor g1371 (n_1782, A[11], A[25]);
  xor g1372 (n_554, n_1782, A[19]);
  nand g1373 (n_1783, A[11], A[25]);
  nand g1376 (n_567, n_1783, n_1649, n_1716);
  xor g1377 (n_1786, A[17], n_551);
  xor g1378 (n_558, n_1786, n_552);
  nand g1379 (n_1787, A[17], n_551);
  nand g1380 (n_1788, n_552, n_551);
  nand g1381 (n_1789, A[17], n_552);
  nand g1382 (n_571, n_1787, n_1788, n_1789);
  xor g1383 (n_1790, n_553, n_554);
  xor g1384 (n_560, n_1790, n_555);
  nand g1385 (n_1791, n_553, n_554);
  nand g1386 (n_1792, n_555, n_554);
  nand g1387 (n_1793, n_553, n_555);
  nand g1388 (n_573, n_1791, n_1792, n_1793);
  xor g1389 (n_1794, n_556, n_557);
  xor g1390 (n_562, n_1794, n_558);
  nand g1391 (n_1795, n_556, n_557);
  nand g1392 (n_1796, n_558, n_557);
  nand g1393 (n_1797, n_556, n_558);
  nand g1394 (n_575, n_1795, n_1796, n_1797);
  xor g1395 (n_1798, n_559, n_560);
  xor g1396 (n_563, n_1798, n_561);
  nand g1397 (n_1799, n_559, n_560);
  nand g1398 (n_1800, n_561, n_560);
  nand g1399 (n_1801, n_559, n_561);
  nand g1400 (n_578, n_1799, n_1800, n_1801);
  xor g1401 (n_1802, n_562, n_563);
  xor g1402 (n_210, n_1802, n_564);
  nand g1403 (n_1803, n_562, n_563);
  nand g1404 (n_1804, n_564, n_563);
  nand g1405 (n_1805, n_562, n_564);
  nand g1406 (n_123, n_1803, n_1804, n_1805);
  xor g1407 (n_1806, A[30], A[28]);
  xor g1408 (n_569, n_1806, A[24]);
  nand g1409 (n_1807, A[30], A[28]);
  nand g1410 (n_1808, A[24], A[28]);
  nand g1411 (n_1809, A[30], A[24]);
  nand g1412 (n_579, n_1807, n_1808, n_1809);
  xor g1414 (n_570, n_382, A[22]);
  nand g1416 (n_1812, A[22], A[14]);
  xor g1419 (n_1814, A[12], A[26]);
  xor g1420 (n_568, n_1814, A[20]);
  nand g1421 (n_1815, A[12], A[26]);
  nand g1424 (n_581, n_1815, n_1681, n_1748);
  xor g1425 (n_1818, A[18], n_565);
  xor g1426 (n_572, n_1818, n_566);
  nand g1427 (n_1819, A[18], n_565);
  nand g1428 (n_1820, n_566, n_565);
  nand g1429 (n_1821, A[18], n_566);
  nand g1430 (n_585, n_1819, n_1820, n_1821);
  xor g1431 (n_1822, n_567, n_568);
  xor g1432 (n_574, n_1822, n_569);
  nand g1433 (n_1823, n_567, n_568);
  nand g1434 (n_1824, n_569, n_568);
  nand g1435 (n_1825, n_567, n_569);
  nand g1436 (n_587, n_1823, n_1824, n_1825);
  xor g1437 (n_1826, n_570, n_571);
  xor g1438 (n_576, n_1826, n_572);
  nand g1439 (n_1827, n_570, n_571);
  nand g1440 (n_1828, n_572, n_571);
  nand g1441 (n_1829, n_570, n_572);
  nand g1442 (n_589, n_1827, n_1828, n_1829);
  xor g1443 (n_1830, n_573, n_574);
  xor g1444 (n_577, n_1830, n_575);
  nand g1445 (n_1831, n_573, n_574);
  nand g1446 (n_1832, n_575, n_574);
  nand g1447 (n_1833, n_573, n_575);
  nand g1448 (n_592, n_1831, n_1832, n_1833);
  xor g1449 (n_1834, n_576, n_577);
  xor g1450 (n_209, n_1834, n_578);
  nand g1451 (n_1835, n_576, n_577);
  nand g1452 (n_1836, n_578, n_577);
  nand g1453 (n_1837, n_576, n_578);
  nand g1454 (n_122, n_1835, n_1836, n_1837);
  xor g1455 (n_1838, A[31], A[29]);
  xor g1456 (n_583, n_1838, A[25]);
  nand g1457 (n_1839, A[31], A[29]);
  nand g1458 (n_1840, A[25], A[29]);
  nand g1459 (n_1841, A[31], A[25]);
  nand g1460 (n_593, n_1839, n_1840, n_1841);
  xor g1462 (n_584, n_1398, A[23]);
  nand g1464 (n_1844, A[23], A[15]);
  nand g1466 (n_594, n_1399, n_1844, n_1585);
  xor g1467 (n_1846, A[13], A[27]);
  xor g1468 (n_582, n_1846, A[21]);
  nand g1469 (n_1847, A[13], A[27]);
  nand g1472 (n_595, n_1847, n_1713, n_1780);
  xor g1473 (n_1850, A[19], n_579);
  xor g1474 (n_586, n_1850, n_580);
  nand g1475 (n_1851, A[19], n_579);
  nand g1476 (n_1852, n_580, n_579);
  nand g1477 (n_1853, A[19], n_580);
  nand g1478 (n_599, n_1851, n_1852, n_1853);
  xor g1479 (n_1854, n_581, n_582);
  xor g1480 (n_588, n_1854, n_583);
  nand g1481 (n_1855, n_581, n_582);
  nand g1482 (n_1856, n_583, n_582);
  nand g1483 (n_1857, n_581, n_583);
  nand g1484 (n_601, n_1855, n_1856, n_1857);
  xor g1485 (n_1858, n_584, n_585);
  xor g1486 (n_590, n_1858, n_586);
  nand g1487 (n_1859, n_584, n_585);
  nand g1488 (n_1860, n_586, n_585);
  nand g1489 (n_1861, n_584, n_586);
  nand g1490 (n_603, n_1859, n_1860, n_1861);
  xor g1491 (n_1862, n_587, n_588);
  xor g1492 (n_591, n_1862, n_589);
  nand g1493 (n_1863, n_587, n_588);
  nand g1494 (n_1864, n_589, n_588);
  nand g1495 (n_1865, n_587, n_589);
  nand g1496 (n_606, n_1863, n_1864, n_1865);
  xor g1497 (n_1866, n_590, n_591);
  xor g1498 (n_208, n_1866, n_592);
  nand g1499 (n_1867, n_590, n_591);
  nand g1500 (n_1868, n_592, n_591);
  nand g1501 (n_1869, n_590, n_592);
  nand g1502 (n_121, n_1867, n_1868, n_1869);
  xor g1503 (n_1870, A[32], A[30]);
  xor g1504 (n_597, n_1870, A[26]);
  nand g1505 (n_1871, A[32], A[30]);
  nand g1506 (n_1872, A[26], A[30]);
  nand g1507 (n_1873, A[32], A[26]);
  nand g1508 (n_607, n_1871, n_1872, n_1873);
  xor g1510 (n_598, n_405, A[24]);
  nand g1512 (n_1876, A[24], A[16]);
  xor g1515 (n_1878, A[14], A[28]);
  xor g1516 (n_596, n_1878, A[22]);
  nand g1517 (n_1879, A[14], A[28]);
  nand g1520 (n_609, n_1879, n_1745, n_1812);
  xor g1521 (n_1882, A[20], n_593);
  xor g1522 (n_600, n_1882, n_594);
  nand g1523 (n_1883, A[20], n_593);
  nand g1524 (n_1884, n_594, n_593);
  nand g1525 (n_1885, A[20], n_594);
  nand g1526 (n_613, n_1883, n_1884, n_1885);
  xor g1527 (n_1886, n_595, n_596);
  xor g1528 (n_602, n_1886, n_597);
  nand g1529 (n_1887, n_595, n_596);
  nand g1530 (n_1888, n_597, n_596);
  nand g1531 (n_1889, n_595, n_597);
  nand g1532 (n_615, n_1887, n_1888, n_1889);
  xor g1533 (n_1890, n_598, n_599);
  xor g1534 (n_604, n_1890, n_600);
  nand g1535 (n_1891, n_598, n_599);
  nand g1536 (n_1892, n_600, n_599);
  nand g1537 (n_1893, n_598, n_600);
  nand g1538 (n_617, n_1891, n_1892, n_1893);
  xor g1539 (n_1894, n_601, n_602);
  xor g1540 (n_605, n_1894, n_603);
  nand g1541 (n_1895, n_601, n_602);
  nand g1542 (n_1896, n_603, n_602);
  nand g1543 (n_1897, n_601, n_603);
  nand g1544 (n_620, n_1895, n_1896, n_1897);
  xor g1545 (n_1898, n_604, n_605);
  xor g1546 (n_207, n_1898, n_606);
  nand g1547 (n_1899, n_604, n_605);
  nand g1548 (n_1900, n_606, n_605);
  nand g1549 (n_1901, n_604, n_606);
  nand g1550 (n_120, n_1899, n_1900, n_1901);
  xor g1551 (n_1902, A[33], A[31]);
  xor g1552 (n_611, n_1902, A[27]);
  nand g1553 (n_1903, A[33], A[31]);
  nand g1554 (n_1904, A[27], A[31]);
  nand g1555 (n_1905, A[33], A[27]);
  nand g1556 (n_621, n_1903, n_1904, n_1905);
  xor g1558 (n_612, n_1454, A[25]);
  nand g1560 (n_1908, A[25], A[17]);
  nand g1562 (n_622, n_1455, n_1908, n_1649);
  xor g1563 (n_1910, A[15], A[29]);
  xor g1564 (n_610, n_1910, A[23]);
  nand g1565 (n_1911, A[15], A[29]);
  nand g1568 (n_623, n_1911, n_1777, n_1844);
  xor g1569 (n_1914, A[21], n_607);
  xor g1570 (n_614, n_1914, n_608);
  nand g1571 (n_1915, A[21], n_607);
  nand g1572 (n_1916, n_608, n_607);
  nand g1573 (n_1917, A[21], n_608);
  nand g1574 (n_627, n_1915, n_1916, n_1917);
  xor g1575 (n_1918, n_609, n_610);
  xor g1576 (n_616, n_1918, n_611);
  nand g1577 (n_1919, n_609, n_610);
  nand g1578 (n_1920, n_611, n_610);
  nand g1579 (n_1921, n_609, n_611);
  nand g1580 (n_629, n_1919, n_1920, n_1921);
  xor g1581 (n_1922, n_612, n_613);
  xor g1582 (n_618, n_1922, n_614);
  nand g1583 (n_1923, n_612, n_613);
  nand g1584 (n_1924, n_614, n_613);
  nand g1585 (n_1925, n_612, n_614);
  nand g1586 (n_631, n_1923, n_1924, n_1925);
  xor g1587 (n_1926, n_615, n_616);
  xor g1588 (n_619, n_1926, n_617);
  nand g1589 (n_1927, n_615, n_616);
  nand g1590 (n_1928, n_617, n_616);
  nand g1591 (n_1929, n_615, n_617);
  nand g1592 (n_634, n_1927, n_1928, n_1929);
  xor g1593 (n_1930, n_618, n_619);
  xor g1594 (n_206, n_1930, n_620);
  nand g1595 (n_1931, n_618, n_619);
  nand g1596 (n_1932, n_620, n_619);
  nand g1597 (n_1933, n_618, n_620);
  nand g1598 (n_119, n_1931, n_1932, n_1933);
  xor g1599 (n_1934, A[34], A[32]);
  xor g1600 (n_625, n_1934, A[28]);
  nand g1601 (n_1935, A[34], A[32]);
  nand g1602 (n_1936, A[28], A[32]);
  nand g1603 (n_1937, A[34], A[28]);
  nand g1604 (n_635, n_1935, n_1936, n_1937);
  xor g1606 (n_626, n_1486, A[26]);
  nand g1608 (n_1940, A[26], A[18]);
  nand g1610 (n_636, n_1487, n_1940, n_1681);
  xor g1611 (n_1942, A[16], A[30]);
  xor g1612 (n_624, n_1942, A[24]);
  nand g1613 (n_1943, A[16], A[30]);
  nand g1616 (n_637, n_1943, n_1809, n_1876);
  xor g1617 (n_1946, A[22], n_621);
  xor g1618 (n_628, n_1946, n_622);
  nand g1619 (n_1947, A[22], n_621);
  nand g1620 (n_1948, n_622, n_621);
  nand g1621 (n_1949, A[22], n_622);
  nand g1622 (n_641, n_1947, n_1948, n_1949);
  xor g1623 (n_1950, n_623, n_624);
  xor g1624 (n_630, n_1950, n_625);
  nand g1625 (n_1951, n_623, n_624);
  nand g1626 (n_1952, n_625, n_624);
  nand g1627 (n_1953, n_623, n_625);
  nand g1628 (n_643, n_1951, n_1952, n_1953);
  xor g1629 (n_1954, n_626, n_627);
  xor g1630 (n_632, n_1954, n_628);
  nand g1631 (n_1955, n_626, n_627);
  nand g1632 (n_1956, n_628, n_627);
  nand g1633 (n_1957, n_626, n_628);
  nand g1634 (n_645, n_1955, n_1956, n_1957);
  xor g1635 (n_1958, n_629, n_630);
  xor g1636 (n_633, n_1958, n_631);
  nand g1637 (n_1959, n_629, n_630);
  nand g1638 (n_1960, n_631, n_630);
  nand g1639 (n_1961, n_629, n_631);
  nand g1640 (n_648, n_1959, n_1960, n_1961);
  xor g1641 (n_1962, n_632, n_633);
  xor g1642 (n_205, n_1962, n_634);
  nand g1643 (n_1963, n_632, n_633);
  nand g1644 (n_1964, n_634, n_633);
  nand g1645 (n_1965, n_632, n_634);
  nand g1646 (n_118, n_1963, n_1964, n_1965);
  xor g1647 (n_1966, A[35], A[33]);
  xor g1648 (n_639, n_1966, A[29]);
  nand g1649 (n_1967, A[35], A[33]);
  nand g1650 (n_1968, A[29], A[33]);
  nand g1651 (n_1969, A[35], A[29]);
  nand g1652 (n_649, n_1967, n_1968, n_1969);
  xor g1654 (n_640, n_1518, A[27]);
  nand g1656 (n_1972, A[27], A[19]);
  nand g1658 (n_650, n_1519, n_1972, n_1713);
  xor g1659 (n_1974, A[17], A[31]);
  xor g1660 (n_638, n_1974, A[25]);
  nand g1661 (n_1975, A[17], A[31]);
  nand g1664 (n_651, n_1975, n_1841, n_1908);
  xor g1665 (n_1978, A[23], n_635);
  xor g1666 (n_642, n_1978, n_636);
  nand g1667 (n_1979, A[23], n_635);
  nand g1668 (n_1980, n_636, n_635);
  nand g1669 (n_1981, A[23], n_636);
  nand g1670 (n_655, n_1979, n_1980, n_1981);
  xor g1671 (n_1982, n_637, n_638);
  xor g1672 (n_644, n_1982, n_639);
  nand g1673 (n_1983, n_637, n_638);
  nand g1674 (n_1984, n_639, n_638);
  nand g1675 (n_1985, n_637, n_639);
  nand g1676 (n_657, n_1983, n_1984, n_1985);
  xor g1677 (n_1986, n_640, n_641);
  xor g1678 (n_646, n_1986, n_642);
  nand g1679 (n_1987, n_640, n_641);
  nand g1680 (n_1988, n_642, n_641);
  nand g1681 (n_1989, n_640, n_642);
  nand g1682 (n_659, n_1987, n_1988, n_1989);
  xor g1683 (n_1990, n_643, n_644);
  xor g1684 (n_647, n_1990, n_645);
  nand g1685 (n_1991, n_643, n_644);
  nand g1686 (n_1992, n_645, n_644);
  nand g1687 (n_1993, n_643, n_645);
  nand g1688 (n_662, n_1991, n_1992, n_1993);
  xor g1689 (n_1994, n_646, n_647);
  xor g1690 (n_204, n_1994, n_648);
  nand g1691 (n_1995, n_646, n_647);
  nand g1692 (n_1996, n_648, n_647);
  nand g1693 (n_1997, n_646, n_648);
  nand g1694 (n_117, n_1995, n_1996, n_1997);
  xor g1695 (n_1998, A[36], A[34]);
  xor g1696 (n_653, n_1998, A[30]);
  nand g1697 (n_1999, A[36], A[34]);
  nand g1698 (n_2000, A[30], A[34]);
  nand g1699 (n_2001, A[36], A[30]);
  nand g1700 (n_663, n_1999, n_2000, n_2001);
  xor g1702 (n_654, n_1550, A[28]);
  nand g1704 (n_2004, A[28], A[20]);
  nand g1706 (n_664, n_1551, n_2004, n_1745);
  xor g1707 (n_2006, A[18], A[32]);
  xor g1708 (n_652, n_2006, A[26]);
  nand g1709 (n_2007, A[18], A[32]);
  nand g1712 (n_665, n_2007, n_1873, n_1940);
  xor g1713 (n_2010, A[24], n_649);
  xor g1714 (n_656, n_2010, n_650);
  nand g1715 (n_2011, A[24], n_649);
  nand g1716 (n_2012, n_650, n_649);
  nand g1717 (n_2013, A[24], n_650);
  nand g1718 (n_669, n_2011, n_2012, n_2013);
  xor g1719 (n_2014, n_651, n_652);
  xor g1720 (n_658, n_2014, n_653);
  nand g1721 (n_2015, n_651, n_652);
  nand g1722 (n_2016, n_653, n_652);
  nand g1723 (n_2017, n_651, n_653);
  nand g1724 (n_671, n_2015, n_2016, n_2017);
  xor g1725 (n_2018, n_654, n_655);
  xor g1726 (n_660, n_2018, n_656);
  nand g1727 (n_2019, n_654, n_655);
  nand g1728 (n_2020, n_656, n_655);
  nand g1729 (n_2021, n_654, n_656);
  nand g1730 (n_673, n_2019, n_2020, n_2021);
  xor g1731 (n_2022, n_657, n_658);
  xor g1732 (n_661, n_2022, n_659);
  nand g1733 (n_2023, n_657, n_658);
  nand g1734 (n_2024, n_659, n_658);
  nand g1735 (n_2025, n_657, n_659);
  nand g1736 (n_676, n_2023, n_2024, n_2025);
  xor g1737 (n_2026, n_660, n_661);
  xor g1738 (n_203, n_2026, n_662);
  nand g1739 (n_2027, n_660, n_661);
  nand g1740 (n_2028, n_662, n_661);
  nand g1741 (n_2029, n_660, n_662);
  nand g1742 (n_116, n_2027, n_2028, n_2029);
  xor g1743 (n_2030, A[37], A[35]);
  xor g1744 (n_667, n_2030, A[31]);
  nand g1745 (n_2031, A[37], A[35]);
  nand g1746 (n_2032, A[31], A[35]);
  nand g1747 (n_2033, A[37], A[31]);
  nand g1748 (n_677, n_2031, n_2032, n_2033);
  xor g1750 (n_668, n_1582, A[29]);
  nand g1752 (n_2036, A[29], A[21]);
  nand g1754 (n_678, n_1583, n_2036, n_1777);
  xor g1755 (n_2038, A[19], A[33]);
  xor g1756 (n_666, n_2038, A[27]);
  nand g1757 (n_2039, A[19], A[33]);
  nand g1760 (n_679, n_2039, n_1905, n_1972);
  xor g1761 (n_2042, A[25], n_663);
  xor g1762 (n_670, n_2042, n_664);
  nand g1763 (n_2043, A[25], n_663);
  nand g1764 (n_2044, n_664, n_663);
  nand g1765 (n_2045, A[25], n_664);
  nand g1766 (n_683, n_2043, n_2044, n_2045);
  xor g1767 (n_2046, n_665, n_666);
  xor g1768 (n_672, n_2046, n_667);
  nand g1769 (n_2047, n_665, n_666);
  nand g1770 (n_2048, n_667, n_666);
  nand g1771 (n_2049, n_665, n_667);
  nand g1772 (n_685, n_2047, n_2048, n_2049);
  xor g1773 (n_2050, n_668, n_669);
  xor g1774 (n_674, n_2050, n_670);
  nand g1775 (n_2051, n_668, n_669);
  nand g1776 (n_2052, n_670, n_669);
  nand g1777 (n_2053, n_668, n_670);
  nand g1778 (n_687, n_2051, n_2052, n_2053);
  xor g1779 (n_2054, n_671, n_672);
  xor g1780 (n_675, n_2054, n_673);
  nand g1781 (n_2055, n_671, n_672);
  nand g1782 (n_2056, n_673, n_672);
  nand g1783 (n_2057, n_671, n_673);
  nand g1784 (n_690, n_2055, n_2056, n_2057);
  xor g1785 (n_2058, n_674, n_675);
  xor g1786 (n_202, n_2058, n_676);
  nand g1787 (n_2059, n_674, n_675);
  nand g1788 (n_2060, n_676, n_675);
  nand g1789 (n_2061, n_674, n_676);
  nand g1790 (n_115, n_2059, n_2060, n_2061);
  xor g1791 (n_2062, A[38], A[36]);
  xor g1792 (n_681, n_2062, A[32]);
  nand g1793 (n_2063, A[38], A[36]);
  nand g1794 (n_2064, A[32], A[36]);
  nand g1795 (n_2065, A[38], A[32]);
  nand g1796 (n_691, n_2063, n_2064, n_2065);
  xor g1798 (n_682, n_1614, A[30]);
  nand g1800 (n_2068, A[30], A[22]);
  nand g1802 (n_692, n_1615, n_2068, n_1809);
  xor g1803 (n_2070, A[20], A[34]);
  xor g1804 (n_680, n_2070, A[28]);
  nand g1805 (n_2071, A[20], A[34]);
  nand g1808 (n_693, n_2071, n_1937, n_2004);
  xor g1809 (n_2074, A[26], n_677);
  xor g1810 (n_684, n_2074, n_678);
  nand g1811 (n_2075, A[26], n_677);
  nand g1812 (n_2076, n_678, n_677);
  nand g1813 (n_2077, A[26], n_678);
  nand g1814 (n_697, n_2075, n_2076, n_2077);
  xor g1815 (n_2078, n_679, n_680);
  xor g1816 (n_686, n_2078, n_681);
  nand g1817 (n_2079, n_679, n_680);
  nand g1818 (n_2080, n_681, n_680);
  nand g1819 (n_2081, n_679, n_681);
  nand g1820 (n_699, n_2079, n_2080, n_2081);
  xor g1821 (n_2082, n_682, n_683);
  xor g1822 (n_688, n_2082, n_684);
  nand g1823 (n_2083, n_682, n_683);
  nand g1824 (n_2084, n_684, n_683);
  nand g1825 (n_2085, n_682, n_684);
  nand g1826 (n_701, n_2083, n_2084, n_2085);
  xor g1827 (n_2086, n_685, n_686);
  xor g1828 (n_689, n_2086, n_687);
  nand g1829 (n_2087, n_685, n_686);
  nand g1830 (n_2088, n_687, n_686);
  nand g1831 (n_2089, n_685, n_687);
  nand g1832 (n_704, n_2087, n_2088, n_2089);
  xor g1833 (n_2090, n_688, n_689);
  xor g1834 (n_201, n_2090, n_690);
  nand g1835 (n_2091, n_688, n_689);
  nand g1836 (n_2092, n_690, n_689);
  nand g1837 (n_2093, n_688, n_690);
  nand g1838 (n_114, n_2091, n_2092, n_2093);
  xor g1839 (n_2094, A[39], A[37]);
  xor g1840 (n_695, n_2094, A[33]);
  nand g1841 (n_2095, A[39], A[37]);
  nand g1842 (n_2096, A[33], A[37]);
  nand g1843 (n_2097, A[39], A[33]);
  nand g1844 (n_705, n_2095, n_2096, n_2097);
  xor g1846 (n_696, n_1646, A[31]);
  nand g1848 (n_2100, A[31], A[23]);
  nand g1850 (n_706, n_1647, n_2100, n_1841);
  xor g1851 (n_2102, A[21], A[35]);
  xor g1852 (n_694, n_2102, A[29]);
  nand g1853 (n_2103, A[21], A[35]);
  nand g1856 (n_707, n_2103, n_1969, n_2036);
  xor g1857 (n_2106, A[27], n_691);
  xor g1858 (n_698, n_2106, n_692);
  nand g1859 (n_2107, A[27], n_691);
  nand g1860 (n_2108, n_692, n_691);
  nand g1861 (n_2109, A[27], n_692);
  nand g1862 (n_711, n_2107, n_2108, n_2109);
  xor g1863 (n_2110, n_693, n_694);
  xor g1864 (n_700, n_2110, n_695);
  nand g1865 (n_2111, n_693, n_694);
  nand g1866 (n_2112, n_695, n_694);
  nand g1867 (n_2113, n_693, n_695);
  nand g1868 (n_713, n_2111, n_2112, n_2113);
  xor g1869 (n_2114, n_696, n_697);
  xor g1870 (n_702, n_2114, n_698);
  nand g1871 (n_2115, n_696, n_697);
  nand g1872 (n_2116, n_698, n_697);
  nand g1873 (n_2117, n_696, n_698);
  nand g1874 (n_715, n_2115, n_2116, n_2117);
  xor g1875 (n_2118, n_699, n_700);
  xor g1876 (n_703, n_2118, n_701);
  nand g1877 (n_2119, n_699, n_700);
  nand g1878 (n_2120, n_701, n_700);
  nand g1879 (n_2121, n_699, n_701);
  nand g1880 (n_718, n_2119, n_2120, n_2121);
  xor g1881 (n_2122, n_702, n_703);
  xor g1882 (n_200, n_2122, n_704);
  nand g1883 (n_2123, n_702, n_703);
  nand g1884 (n_2124, n_704, n_703);
  nand g1885 (n_2125, n_702, n_704);
  nand g1886 (n_113, n_2123, n_2124, n_2125);
  xor g1887 (n_2126, A[40], A[38]);
  xor g1888 (n_709, n_2126, A[34]);
  nand g1889 (n_2127, A[40], A[38]);
  nand g1890 (n_2128, A[34], A[38]);
  nand g1891 (n_2129, A[40], A[34]);
  nand g1892 (n_719, n_2127, n_2128, n_2129);
  xor g1894 (n_710, n_1678, A[32]);
  nand g1896 (n_2132, A[32], A[24]);
  nand g1898 (n_720, n_1679, n_2132, n_1873);
  xor g1899 (n_2134, A[22], A[36]);
  xor g1900 (n_708, n_2134, A[30]);
  nand g1901 (n_2135, A[22], A[36]);
  nand g1904 (n_721, n_2135, n_2001, n_2068);
  xor g1905 (n_2138, A[28], n_705);
  xor g1906 (n_712, n_2138, n_706);
  nand g1907 (n_2139, A[28], n_705);
  nand g1908 (n_2140, n_706, n_705);
  nand g1909 (n_2141, A[28], n_706);
  nand g1910 (n_725, n_2139, n_2140, n_2141);
  xor g1911 (n_2142, n_707, n_708);
  xor g1912 (n_714, n_2142, n_709);
  nand g1913 (n_2143, n_707, n_708);
  nand g1914 (n_2144, n_709, n_708);
  nand g1915 (n_2145, n_707, n_709);
  nand g1916 (n_727, n_2143, n_2144, n_2145);
  xor g1917 (n_2146, n_710, n_711);
  xor g1918 (n_716, n_2146, n_712);
  nand g1919 (n_2147, n_710, n_711);
  nand g1920 (n_2148, n_712, n_711);
  nand g1921 (n_2149, n_710, n_712);
  nand g1922 (n_729, n_2147, n_2148, n_2149);
  xor g1923 (n_2150, n_713, n_714);
  xor g1924 (n_717, n_2150, n_715);
  nand g1925 (n_2151, n_713, n_714);
  nand g1926 (n_2152, n_715, n_714);
  nand g1927 (n_2153, n_713, n_715);
  nand g1928 (n_732, n_2151, n_2152, n_2153);
  xor g1929 (n_2154, n_716, n_717);
  xor g1930 (n_199, n_2154, n_718);
  nand g1931 (n_2155, n_716, n_717);
  nand g1932 (n_2156, n_718, n_717);
  nand g1933 (n_2157, n_716, n_718);
  nand g1934 (n_112, n_2155, n_2156, n_2157);
  xor g1935 (n_2158, A[41], A[39]);
  xor g1936 (n_723, n_2158, A[35]);
  nand g1937 (n_2159, A[41], A[39]);
  nand g1938 (n_2160, A[35], A[39]);
  nand g1939 (n_2161, A[41], A[35]);
  nand g1940 (n_733, n_2159, n_2160, n_2161);
  xor g1942 (n_724, n_1710, A[33]);
  nand g1944 (n_2164, A[33], A[25]);
  nand g1946 (n_734, n_1711, n_2164, n_1905);
  xor g1947 (n_2166, A[23], A[37]);
  xor g1948 (n_722, n_2166, A[31]);
  nand g1949 (n_2167, A[23], A[37]);
  nand g1952 (n_735, n_2167, n_2033, n_2100);
  xor g1953 (n_2170, A[29], n_719);
  xor g1954 (n_726, n_2170, n_720);
  nand g1955 (n_2171, A[29], n_719);
  nand g1956 (n_2172, n_720, n_719);
  nand g1957 (n_2173, A[29], n_720);
  nand g1958 (n_739, n_2171, n_2172, n_2173);
  xor g1959 (n_2174, n_721, n_722);
  xor g1960 (n_728, n_2174, n_723);
  nand g1961 (n_2175, n_721, n_722);
  nand g1962 (n_2176, n_723, n_722);
  nand g1963 (n_2177, n_721, n_723);
  nand g1964 (n_741, n_2175, n_2176, n_2177);
  xor g1965 (n_2178, n_724, n_725);
  xor g1966 (n_730, n_2178, n_726);
  nand g1967 (n_2179, n_724, n_725);
  nand g1968 (n_2180, n_726, n_725);
  nand g1969 (n_2181, n_724, n_726);
  nand g1970 (n_743, n_2179, n_2180, n_2181);
  xor g1971 (n_2182, n_727, n_728);
  xor g1972 (n_731, n_2182, n_729);
  nand g1973 (n_2183, n_727, n_728);
  nand g1974 (n_2184, n_729, n_728);
  nand g1975 (n_2185, n_727, n_729);
  nand g1976 (n_746, n_2183, n_2184, n_2185);
  xor g1977 (n_2186, n_730, n_731);
  xor g1978 (n_198, n_2186, n_732);
  nand g1979 (n_2187, n_730, n_731);
  nand g1980 (n_2188, n_732, n_731);
  nand g1981 (n_2189, n_730, n_732);
  nand g1982 (n_111, n_2187, n_2188, n_2189);
  xor g1983 (n_2190, A[42], A[40]);
  xor g1984 (n_737, n_2190, A[36]);
  nand g1985 (n_2191, A[42], A[40]);
  nand g1986 (n_2192, A[36], A[40]);
  nand g1987 (n_2193, A[42], A[36]);
  nand g1988 (n_747, n_2191, n_2192, n_2193);
  xor g1990 (n_738, n_1742, A[34]);
  nand g1992 (n_2196, A[34], A[26]);
  nand g1994 (n_748, n_1743, n_2196, n_1937);
  xor g1995 (n_2198, A[24], A[38]);
  xor g1996 (n_736, n_2198, A[32]);
  nand g1997 (n_2199, A[24], A[38]);
  nand g2000 (n_749, n_2199, n_2065, n_2132);
  xor g2001 (n_2202, A[30], n_733);
  xor g2002 (n_740, n_2202, n_734);
  nand g2003 (n_2203, A[30], n_733);
  nand g2004 (n_2204, n_734, n_733);
  nand g2005 (n_2205, A[30], n_734);
  nand g2006 (n_753, n_2203, n_2204, n_2205);
  xor g2007 (n_2206, n_735, n_736);
  xor g2008 (n_742, n_2206, n_737);
  nand g2009 (n_2207, n_735, n_736);
  nand g2010 (n_2208, n_737, n_736);
  nand g2011 (n_2209, n_735, n_737);
  nand g2012 (n_755, n_2207, n_2208, n_2209);
  xor g2013 (n_2210, n_738, n_739);
  xor g2014 (n_744, n_2210, n_740);
  nand g2015 (n_2211, n_738, n_739);
  nand g2016 (n_2212, n_740, n_739);
  nand g2017 (n_2213, n_738, n_740);
  nand g2018 (n_757, n_2211, n_2212, n_2213);
  xor g2019 (n_2214, n_741, n_742);
  xor g2020 (n_745, n_2214, n_743);
  nand g2021 (n_2215, n_741, n_742);
  nand g2022 (n_2216, n_743, n_742);
  nand g2023 (n_2217, n_741, n_743);
  nand g2024 (n_760, n_2215, n_2216, n_2217);
  xor g2025 (n_2218, n_744, n_745);
  xor g2026 (n_197, n_2218, n_746);
  nand g2027 (n_2219, n_744, n_745);
  nand g2028 (n_2220, n_746, n_745);
  nand g2029 (n_2221, n_744, n_746);
  nand g2030 (n_110, n_2219, n_2220, n_2221);
  xor g2031 (n_2222, A[43], A[41]);
  xor g2032 (n_751, n_2222, A[37]);
  nand g2033 (n_2223, A[43], A[41]);
  nand g2034 (n_2224, A[37], A[41]);
  nand g2035 (n_2225, A[43], A[37]);
  nand g2036 (n_761, n_2223, n_2224, n_2225);
  xor g2038 (n_752, n_1774, A[35]);
  nand g2040 (n_2228, A[35], A[27]);
  nand g2042 (n_762, n_1775, n_2228, n_1969);
  xor g2043 (n_2230, A[25], A[39]);
  xor g2044 (n_750, n_2230, A[33]);
  nand g2045 (n_2231, A[25], A[39]);
  nand g2048 (n_763, n_2231, n_2097, n_2164);
  xor g2049 (n_2234, A[31], n_747);
  xor g2050 (n_754, n_2234, n_748);
  nand g2051 (n_2235, A[31], n_747);
  nand g2052 (n_2236, n_748, n_747);
  nand g2053 (n_2237, A[31], n_748);
  nand g2054 (n_767, n_2235, n_2236, n_2237);
  xor g2055 (n_2238, n_749, n_750);
  xor g2056 (n_756, n_2238, n_751);
  nand g2057 (n_2239, n_749, n_750);
  nand g2058 (n_2240, n_751, n_750);
  nand g2059 (n_2241, n_749, n_751);
  nand g2060 (n_769, n_2239, n_2240, n_2241);
  xor g2061 (n_2242, n_752, n_753);
  xor g2062 (n_758, n_2242, n_754);
  nand g2063 (n_2243, n_752, n_753);
  nand g2064 (n_2244, n_754, n_753);
  nand g2065 (n_2245, n_752, n_754);
  nand g2066 (n_771, n_2243, n_2244, n_2245);
  xor g2067 (n_2246, n_755, n_756);
  xor g2068 (n_759, n_2246, n_757);
  nand g2069 (n_2247, n_755, n_756);
  nand g2070 (n_2248, n_757, n_756);
  nand g2071 (n_2249, n_755, n_757);
  nand g2072 (n_774, n_2247, n_2248, n_2249);
  xor g2073 (n_2250, n_758, n_759);
  xor g2074 (n_196, n_2250, n_760);
  nand g2075 (n_2251, n_758, n_759);
  nand g2076 (n_2252, n_760, n_759);
  nand g2077 (n_2253, n_758, n_760);
  nand g2078 (n_109, n_2251, n_2252, n_2253);
  xor g2079 (n_2254, A[44], A[42]);
  xor g2080 (n_765, n_2254, A[38]);
  nand g2081 (n_2255, A[44], A[42]);
  nand g2082 (n_2256, A[38], A[42]);
  nand g2083 (n_2257, A[44], A[38]);
  nand g2084 (n_775, n_2255, n_2256, n_2257);
  xor g2086 (n_766, n_1806, A[36]);
  nand g2088 (n_2260, A[36], A[28]);
  nand g2090 (n_776, n_1807, n_2260, n_2001);
  xor g2091 (n_2262, A[26], A[40]);
  xor g2092 (n_764, n_2262, A[34]);
  nand g2093 (n_2263, A[26], A[40]);
  nand g2096 (n_777, n_2263, n_2129, n_2196);
  xor g2097 (n_2266, A[32], n_761);
  xor g2098 (n_768, n_2266, n_762);
  nand g2099 (n_2267, A[32], n_761);
  nand g2100 (n_2268, n_762, n_761);
  nand g2101 (n_2269, A[32], n_762);
  nand g2102 (n_781, n_2267, n_2268, n_2269);
  xor g2103 (n_2270, n_763, n_764);
  xor g2104 (n_770, n_2270, n_765);
  nand g2105 (n_2271, n_763, n_764);
  nand g2106 (n_2272, n_765, n_764);
  nand g2107 (n_2273, n_763, n_765);
  nand g2108 (n_783, n_2271, n_2272, n_2273);
  xor g2109 (n_2274, n_766, n_767);
  xor g2110 (n_772, n_2274, n_768);
  nand g2111 (n_2275, n_766, n_767);
  nand g2112 (n_2276, n_768, n_767);
  nand g2113 (n_2277, n_766, n_768);
  nand g2114 (n_785, n_2275, n_2276, n_2277);
  xor g2115 (n_2278, n_769, n_770);
  xor g2116 (n_773, n_2278, n_771);
  nand g2117 (n_2279, n_769, n_770);
  nand g2118 (n_2280, n_771, n_770);
  nand g2119 (n_2281, n_769, n_771);
  nand g2120 (n_788, n_2279, n_2280, n_2281);
  xor g2121 (n_2282, n_772, n_773);
  xor g2122 (n_195, n_2282, n_774);
  nand g2123 (n_2283, n_772, n_773);
  nand g2124 (n_2284, n_774, n_773);
  nand g2125 (n_2285, n_772, n_774);
  nand g2126 (n_108, n_2283, n_2284, n_2285);
  xor g2127 (n_2286, A[45], A[43]);
  xor g2128 (n_779, n_2286, A[39]);
  nand g2129 (n_2287, A[45], A[43]);
  nand g2130 (n_2288, A[39], A[43]);
  nand g2131 (n_2289, A[45], A[39]);
  nand g2132 (n_789, n_2287, n_2288, n_2289);
  xor g2134 (n_780, n_1838, A[37]);
  nand g2136 (n_2292, A[37], A[29]);
  nand g2138 (n_790, n_1839, n_2292, n_2033);
  xor g2139 (n_2294, A[27], A[41]);
  xor g2140 (n_778, n_2294, A[35]);
  nand g2141 (n_2295, A[27], A[41]);
  nand g2144 (n_791, n_2295, n_2161, n_2228);
  xor g2145 (n_2298, A[33], n_775);
  xor g2146 (n_782, n_2298, n_776);
  nand g2147 (n_2299, A[33], n_775);
  nand g2148 (n_2300, n_776, n_775);
  nand g2149 (n_2301, A[33], n_776);
  nand g2150 (n_795, n_2299, n_2300, n_2301);
  xor g2151 (n_2302, n_777, n_778);
  xor g2152 (n_784, n_2302, n_779);
  nand g2153 (n_2303, n_777, n_778);
  nand g2154 (n_2304, n_779, n_778);
  nand g2155 (n_2305, n_777, n_779);
  nand g2156 (n_797, n_2303, n_2304, n_2305);
  xor g2157 (n_2306, n_780, n_781);
  xor g2158 (n_786, n_2306, n_782);
  nand g2159 (n_2307, n_780, n_781);
  nand g2160 (n_2308, n_782, n_781);
  nand g2161 (n_2309, n_780, n_782);
  nand g2162 (n_799, n_2307, n_2308, n_2309);
  xor g2163 (n_2310, n_783, n_784);
  xor g2164 (n_787, n_2310, n_785);
  nand g2165 (n_2311, n_783, n_784);
  nand g2166 (n_2312, n_785, n_784);
  nand g2167 (n_2313, n_783, n_785);
  nand g2168 (n_802, n_2311, n_2312, n_2313);
  xor g2169 (n_2314, n_786, n_787);
  xor g2170 (n_194, n_2314, n_788);
  nand g2171 (n_2315, n_786, n_787);
  nand g2172 (n_2316, n_788, n_787);
  nand g2173 (n_2317, n_786, n_788);
  nand g2174 (n_107, n_2315, n_2316, n_2317);
  xor g2175 (n_2318, A[46], A[44]);
  xor g2176 (n_793, n_2318, A[40]);
  nand g2177 (n_2319, A[46], A[44]);
  nand g2178 (n_2320, A[40], A[44]);
  nand g2179 (n_2321, A[46], A[40]);
  nand g2180 (n_803, n_2319, n_2320, n_2321);
  xor g2182 (n_794, n_1870, A[38]);
  nand g2184 (n_2324, A[38], A[30]);
  nand g2186 (n_804, n_1871, n_2324, n_2065);
  xor g2187 (n_2326, A[28], A[42]);
  xor g2188 (n_792, n_2326, A[36]);
  nand g2189 (n_2327, A[28], A[42]);
  nand g2192 (n_805, n_2327, n_2193, n_2260);
  xor g2193 (n_2330, A[34], n_789);
  xor g2194 (n_796, n_2330, n_790);
  nand g2195 (n_2331, A[34], n_789);
  nand g2196 (n_2332, n_790, n_789);
  nand g2197 (n_2333, A[34], n_790);
  nand g2198 (n_809, n_2331, n_2332, n_2333);
  xor g2199 (n_2334, n_791, n_792);
  xor g2200 (n_798, n_2334, n_793);
  nand g2201 (n_2335, n_791, n_792);
  nand g2202 (n_2336, n_793, n_792);
  nand g2203 (n_2337, n_791, n_793);
  nand g2204 (n_811, n_2335, n_2336, n_2337);
  xor g2205 (n_2338, n_794, n_795);
  xor g2206 (n_800, n_2338, n_796);
  nand g2207 (n_2339, n_794, n_795);
  nand g2208 (n_2340, n_796, n_795);
  nand g2209 (n_2341, n_794, n_796);
  nand g2210 (n_813, n_2339, n_2340, n_2341);
  xor g2211 (n_2342, n_797, n_798);
  xor g2212 (n_801, n_2342, n_799);
  nand g2213 (n_2343, n_797, n_798);
  nand g2214 (n_2344, n_799, n_798);
  nand g2215 (n_2345, n_797, n_799);
  nand g2216 (n_816, n_2343, n_2344, n_2345);
  xor g2217 (n_2346, n_800, n_801);
  xor g2218 (n_193, n_2346, n_802);
  nand g2219 (n_2347, n_800, n_801);
  nand g2220 (n_2348, n_802, n_801);
  nand g2221 (n_2349, n_800, n_802);
  nand g2222 (n_106, n_2347, n_2348, n_2349);
  xor g2223 (n_2350, A[47], A[45]);
  xor g2224 (n_807, n_2350, A[41]);
  nand g2225 (n_2351, A[47], A[45]);
  nand g2226 (n_2352, A[41], A[45]);
  nand g2227 (n_2353, A[47], A[41]);
  nand g2228 (n_817, n_2351, n_2352, n_2353);
  xor g2230 (n_808, n_1902, A[39]);
  nand g2232 (n_2356, A[39], A[31]);
  nand g2234 (n_818, n_1903, n_2356, n_2097);
  xor g2235 (n_2358, A[29], A[43]);
  xor g2236 (n_806, n_2358, A[37]);
  nand g2237 (n_2359, A[29], A[43]);
  nand g2240 (n_819, n_2359, n_2225, n_2292);
  xor g2241 (n_2362, A[35], n_803);
  xor g2242 (n_810, n_2362, n_804);
  nand g2243 (n_2363, A[35], n_803);
  nand g2244 (n_2364, n_804, n_803);
  nand g2245 (n_2365, A[35], n_804);
  nand g2246 (n_823, n_2363, n_2364, n_2365);
  xor g2247 (n_2366, n_805, n_806);
  xor g2248 (n_812, n_2366, n_807);
  nand g2249 (n_2367, n_805, n_806);
  nand g2250 (n_2368, n_807, n_806);
  nand g2251 (n_2369, n_805, n_807);
  nand g2252 (n_825, n_2367, n_2368, n_2369);
  xor g2253 (n_2370, n_808, n_809);
  xor g2254 (n_814, n_2370, n_810);
  nand g2255 (n_2371, n_808, n_809);
  nand g2256 (n_2372, n_810, n_809);
  nand g2257 (n_2373, n_808, n_810);
  nand g2258 (n_827, n_2371, n_2372, n_2373);
  xor g2259 (n_2374, n_811, n_812);
  xor g2260 (n_815, n_2374, n_813);
  nand g2261 (n_2375, n_811, n_812);
  nand g2262 (n_2376, n_813, n_812);
  nand g2263 (n_2377, n_811, n_813);
  nand g2264 (n_830, n_2375, n_2376, n_2377);
  xor g2265 (n_2378, n_814, n_815);
  xor g2266 (n_192, n_2378, n_816);
  nand g2267 (n_2379, n_814, n_815);
  nand g2268 (n_2380, n_816, n_815);
  nand g2269 (n_2381, n_814, n_816);
  nand g2270 (n_105, n_2379, n_2380, n_2381);
  xor g2271 (n_2382, A[48], A[46]);
  xor g2272 (n_821, n_2382, A[42]);
  nand g2273 (n_2383, A[48], A[46]);
  nand g2274 (n_2384, A[42], A[46]);
  nand g2275 (n_2385, A[48], A[42]);
  nand g2276 (n_831, n_2383, n_2384, n_2385);
  xor g2278 (n_822, n_1934, A[40]);
  nand g2280 (n_2388, A[40], A[32]);
  nand g2282 (n_832, n_1935, n_2388, n_2129);
  xor g2283 (n_2390, A[30], A[44]);
  xor g2284 (n_820, n_2390, A[38]);
  nand g2285 (n_2391, A[30], A[44]);
  nand g2288 (n_833, n_2391, n_2257, n_2324);
  xor g2289 (n_2394, A[36], n_817);
  xor g2290 (n_824, n_2394, n_818);
  nand g2291 (n_2395, A[36], n_817);
  nand g2292 (n_2396, n_818, n_817);
  nand g2293 (n_2397, A[36], n_818);
  nand g2294 (n_837, n_2395, n_2396, n_2397);
  xor g2295 (n_2398, n_819, n_820);
  xor g2296 (n_826, n_2398, n_821);
  nand g2297 (n_2399, n_819, n_820);
  nand g2298 (n_2400, n_821, n_820);
  nand g2299 (n_2401, n_819, n_821);
  nand g2300 (n_839, n_2399, n_2400, n_2401);
  xor g2301 (n_2402, n_822, n_823);
  xor g2302 (n_828, n_2402, n_824);
  nand g2303 (n_2403, n_822, n_823);
  nand g2304 (n_2404, n_824, n_823);
  nand g2305 (n_2405, n_822, n_824);
  nand g2306 (n_841, n_2403, n_2404, n_2405);
  xor g2307 (n_2406, n_825, n_826);
  xor g2308 (n_829, n_2406, n_827);
  nand g2309 (n_2407, n_825, n_826);
  nand g2310 (n_2408, n_827, n_826);
  nand g2311 (n_2409, n_825, n_827);
  nand g2312 (n_844, n_2407, n_2408, n_2409);
  xor g2313 (n_2410, n_828, n_829);
  xor g2314 (n_191, n_2410, n_830);
  nand g2315 (n_2411, n_828, n_829);
  nand g2316 (n_2412, n_830, n_829);
  nand g2317 (n_2413, n_828, n_830);
  nand g2318 (n_104, n_2411, n_2412, n_2413);
  xor g2319 (n_2414, A[49], A[47]);
  xor g2320 (n_835, n_2414, A[43]);
  nand g2321 (n_2415, A[49], A[47]);
  nand g2322 (n_2416, A[43], A[47]);
  nand g2323 (n_2417, A[49], A[43]);
  nand g2324 (n_845, n_2415, n_2416, n_2417);
  xor g2326 (n_836, n_1966, A[41]);
  nand g2328 (n_2420, A[41], A[33]);
  nand g2330 (n_846, n_1967, n_2420, n_2161);
  xor g2331 (n_2422, A[31], A[45]);
  xor g2332 (n_834, n_2422, A[39]);
  nand g2333 (n_2423, A[31], A[45]);
  nand g2336 (n_847, n_2423, n_2289, n_2356);
  xor g2337 (n_2426, A[37], n_831);
  xor g2338 (n_838, n_2426, n_832);
  nand g2339 (n_2427, A[37], n_831);
  nand g2340 (n_2428, n_832, n_831);
  nand g2341 (n_2429, A[37], n_832);
  nand g2342 (n_851, n_2427, n_2428, n_2429);
  xor g2343 (n_2430, n_833, n_834);
  xor g2344 (n_840, n_2430, n_835);
  nand g2345 (n_2431, n_833, n_834);
  nand g2346 (n_2432, n_835, n_834);
  nand g2347 (n_2433, n_833, n_835);
  nand g2348 (n_853, n_2431, n_2432, n_2433);
  xor g2349 (n_2434, n_836, n_837);
  xor g2350 (n_842, n_2434, n_838);
  nand g2351 (n_2435, n_836, n_837);
  nand g2352 (n_2436, n_838, n_837);
  nand g2353 (n_2437, n_836, n_838);
  nand g2354 (n_855, n_2435, n_2436, n_2437);
  xor g2355 (n_2438, n_839, n_840);
  xor g2356 (n_843, n_2438, n_841);
  nand g2357 (n_2439, n_839, n_840);
  nand g2358 (n_2440, n_841, n_840);
  nand g2359 (n_2441, n_839, n_841);
  nand g2360 (n_858, n_2439, n_2440, n_2441);
  xor g2361 (n_2442, n_842, n_843);
  xor g2362 (n_190, n_2442, n_844);
  nand g2363 (n_2443, n_842, n_843);
  nand g2364 (n_2444, n_844, n_843);
  nand g2365 (n_2445, n_842, n_844);
  nand g2366 (n_103, n_2443, n_2444, n_2445);
  xor g2367 (n_2446, A[50], A[48]);
  xor g2368 (n_849, n_2446, A[44]);
  nand g2369 (n_2447, A[50], A[48]);
  nand g2370 (n_2448, A[44], A[48]);
  nand g2371 (n_2449, A[50], A[44]);
  nand g2372 (n_859, n_2447, n_2448, n_2449);
  xor g2374 (n_850, n_1998, A[42]);
  nand g2376 (n_2452, A[42], A[34]);
  nand g2378 (n_860, n_1999, n_2452, n_2193);
  xor g2379 (n_2454, A[32], A[46]);
  xor g2380 (n_848, n_2454, A[40]);
  nand g2381 (n_2455, A[32], A[46]);
  nand g2384 (n_861, n_2455, n_2321, n_2388);
  xor g2385 (n_2458, A[38], n_845);
  xor g2386 (n_852, n_2458, n_846);
  nand g2387 (n_2459, A[38], n_845);
  nand g2388 (n_2460, n_846, n_845);
  nand g2389 (n_2461, A[38], n_846);
  nand g2390 (n_865, n_2459, n_2460, n_2461);
  xor g2391 (n_2462, n_847, n_848);
  xor g2392 (n_854, n_2462, n_849);
  nand g2393 (n_2463, n_847, n_848);
  nand g2394 (n_2464, n_849, n_848);
  nand g2395 (n_2465, n_847, n_849);
  nand g2396 (n_867, n_2463, n_2464, n_2465);
  xor g2397 (n_2466, n_850, n_851);
  xor g2398 (n_856, n_2466, n_852);
  nand g2399 (n_2467, n_850, n_851);
  nand g2400 (n_2468, n_852, n_851);
  nand g2401 (n_2469, n_850, n_852);
  nand g2402 (n_869, n_2467, n_2468, n_2469);
  xor g2403 (n_2470, n_853, n_854);
  xor g2404 (n_857, n_2470, n_855);
  nand g2405 (n_2471, n_853, n_854);
  nand g2406 (n_2472, n_855, n_854);
  nand g2407 (n_2473, n_853, n_855);
  nand g2408 (n_872, n_2471, n_2472, n_2473);
  xor g2409 (n_2474, n_856, n_857);
  xor g2410 (n_189, n_2474, n_858);
  nand g2411 (n_2475, n_856, n_857);
  nand g2412 (n_2476, n_858, n_857);
  nand g2413 (n_2477, n_856, n_858);
  nand g2414 (n_102, n_2475, n_2476, n_2477);
  xor g2415 (n_2478, A[51], A[49]);
  xor g2416 (n_863, n_2478, A[45]);
  nand g2417 (n_2479, A[51], A[49]);
  nand g2418 (n_2480, A[45], A[49]);
  nand g2419 (n_2481, A[51], A[45]);
  nand g2420 (n_873, n_2479, n_2480, n_2481);
  xor g2422 (n_864, n_2030, A[43]);
  nand g2424 (n_2484, A[43], A[35]);
  nand g2426 (n_874, n_2031, n_2484, n_2225);
  xor g2427 (n_2486, A[33], A[47]);
  xor g2428 (n_862, n_2486, A[41]);
  nand g2429 (n_2487, A[33], A[47]);
  nand g2432 (n_875, n_2487, n_2353, n_2420);
  xor g2433 (n_2490, A[39], n_859);
  xor g2434 (n_866, n_2490, n_860);
  nand g2435 (n_2491, A[39], n_859);
  nand g2436 (n_2492, n_860, n_859);
  nand g2437 (n_2493, A[39], n_860);
  nand g2438 (n_879, n_2491, n_2492, n_2493);
  xor g2439 (n_2494, n_861, n_862);
  xor g2440 (n_868, n_2494, n_863);
  nand g2441 (n_2495, n_861, n_862);
  nand g2442 (n_2496, n_863, n_862);
  nand g2443 (n_2497, n_861, n_863);
  nand g2444 (n_881, n_2495, n_2496, n_2497);
  xor g2445 (n_2498, n_864, n_865);
  xor g2446 (n_870, n_2498, n_866);
  nand g2447 (n_2499, n_864, n_865);
  nand g2448 (n_2500, n_866, n_865);
  nand g2449 (n_2501, n_864, n_866);
  nand g2450 (n_883, n_2499, n_2500, n_2501);
  xor g2451 (n_2502, n_867, n_868);
  xor g2452 (n_871, n_2502, n_869);
  nand g2453 (n_2503, n_867, n_868);
  nand g2454 (n_2504, n_869, n_868);
  nand g2455 (n_2505, n_867, n_869);
  nand g2456 (n_886, n_2503, n_2504, n_2505);
  xor g2457 (n_2506, n_870, n_871);
  xor g2458 (n_188, n_2506, n_872);
  nand g2459 (n_2507, n_870, n_871);
  nand g2460 (n_2508, n_872, n_871);
  nand g2461 (n_2509, n_870, n_872);
  nand g2462 (n_101, n_2507, n_2508, n_2509);
  xor g2463 (n_2510, A[52], A[50]);
  xor g2464 (n_877, n_2510, A[46]);
  nand g2465 (n_2511, A[52], A[50]);
  nand g2466 (n_2512, A[46], A[50]);
  nand g2467 (n_2513, A[52], A[46]);
  nand g2468 (n_887, n_2511, n_2512, n_2513);
  xor g2470 (n_878, n_2062, A[44]);
  nand g2472 (n_2516, A[44], A[36]);
  nand g2474 (n_888, n_2063, n_2516, n_2257);
  xor g2475 (n_2518, A[34], A[48]);
  xor g2476 (n_876, n_2518, A[42]);
  nand g2477 (n_2519, A[34], A[48]);
  nand g2480 (n_889, n_2519, n_2385, n_2452);
  xor g2481 (n_2522, A[40], n_873);
  xor g2482 (n_880, n_2522, n_874);
  nand g2483 (n_2523, A[40], n_873);
  nand g2484 (n_2524, n_874, n_873);
  nand g2485 (n_2525, A[40], n_874);
  nand g2486 (n_893, n_2523, n_2524, n_2525);
  xor g2487 (n_2526, n_875, n_876);
  xor g2488 (n_882, n_2526, n_877);
  nand g2489 (n_2527, n_875, n_876);
  nand g2490 (n_2528, n_877, n_876);
  nand g2491 (n_2529, n_875, n_877);
  nand g2492 (n_895, n_2527, n_2528, n_2529);
  xor g2493 (n_2530, n_878, n_879);
  xor g2494 (n_884, n_2530, n_880);
  nand g2495 (n_2531, n_878, n_879);
  nand g2496 (n_2532, n_880, n_879);
  nand g2497 (n_2533, n_878, n_880);
  nand g2498 (n_897, n_2531, n_2532, n_2533);
  xor g2499 (n_2534, n_881, n_882);
  xor g2500 (n_885, n_2534, n_883);
  nand g2501 (n_2535, n_881, n_882);
  nand g2502 (n_2536, n_883, n_882);
  nand g2503 (n_2537, n_881, n_883);
  nand g2504 (n_900, n_2535, n_2536, n_2537);
  xor g2505 (n_2538, n_884, n_885);
  xor g2506 (n_187, n_2538, n_886);
  nand g2507 (n_2539, n_884, n_885);
  nand g2508 (n_2540, n_886, n_885);
  nand g2509 (n_2541, n_884, n_886);
  nand g2510 (n_100, n_2539, n_2540, n_2541);
  xor g2511 (n_2542, A[53], A[51]);
  xor g2512 (n_891, n_2542, A[47]);
  nand g2513 (n_2543, A[53], A[51]);
  nand g2514 (n_2544, A[47], A[51]);
  nand g2515 (n_2545, A[53], A[47]);
  nand g2516 (n_901, n_2543, n_2544, n_2545);
  xor g2518 (n_892, n_2094, A[45]);
  nand g2520 (n_2548, A[45], A[37]);
  nand g2522 (n_902, n_2095, n_2548, n_2289);
  xor g2523 (n_2550, A[35], A[49]);
  xor g2524 (n_890, n_2550, A[43]);
  nand g2525 (n_2551, A[35], A[49]);
  nand g2528 (n_903, n_2551, n_2417, n_2484);
  xor g2529 (n_2554, A[41], n_887);
  xor g2530 (n_894, n_2554, n_888);
  nand g2531 (n_2555, A[41], n_887);
  nand g2532 (n_2556, n_888, n_887);
  nand g2533 (n_2557, A[41], n_888);
  nand g2534 (n_907, n_2555, n_2556, n_2557);
  xor g2535 (n_2558, n_889, n_890);
  xor g2536 (n_896, n_2558, n_891);
  nand g2537 (n_2559, n_889, n_890);
  nand g2538 (n_2560, n_891, n_890);
  nand g2539 (n_2561, n_889, n_891);
  nand g2540 (n_909, n_2559, n_2560, n_2561);
  xor g2541 (n_2562, n_892, n_893);
  xor g2542 (n_898, n_2562, n_894);
  nand g2543 (n_2563, n_892, n_893);
  nand g2544 (n_2564, n_894, n_893);
  nand g2545 (n_2565, n_892, n_894);
  nand g2546 (n_911, n_2563, n_2564, n_2565);
  xor g2547 (n_2566, n_895, n_896);
  xor g2548 (n_899, n_2566, n_897);
  nand g2549 (n_2567, n_895, n_896);
  nand g2550 (n_2568, n_897, n_896);
  nand g2551 (n_2569, n_895, n_897);
  nand g2552 (n_914, n_2567, n_2568, n_2569);
  xor g2553 (n_2570, n_898, n_899);
  xor g2554 (n_186, n_2570, n_900);
  nand g2555 (n_2571, n_898, n_899);
  nand g2556 (n_2572, n_900, n_899);
  nand g2557 (n_2573, n_898, n_900);
  nand g2558 (n_99, n_2571, n_2572, n_2573);
  xor g2559 (n_2574, A[54], A[52]);
  xor g2560 (n_905, n_2574, A[48]);
  nand g2561 (n_2575, A[54], A[52]);
  nand g2562 (n_2576, A[48], A[52]);
  nand g2563 (n_2577, A[54], A[48]);
  nand g2564 (n_915, n_2575, n_2576, n_2577);
  xor g2566 (n_906, n_2126, A[46]);
  nand g2568 (n_2580, A[46], A[38]);
  nand g2570 (n_916, n_2127, n_2580, n_2321);
  xor g2571 (n_2582, A[36], A[50]);
  xor g2572 (n_904, n_2582, A[44]);
  nand g2573 (n_2583, A[36], A[50]);
  nand g2576 (n_917, n_2583, n_2449, n_2516);
  xor g2577 (n_2586, A[42], n_901);
  xor g2578 (n_908, n_2586, n_902);
  nand g2579 (n_2587, A[42], n_901);
  nand g2580 (n_2588, n_902, n_901);
  nand g2581 (n_2589, A[42], n_902);
  nand g2582 (n_921, n_2587, n_2588, n_2589);
  xor g2583 (n_2590, n_903, n_904);
  xor g2584 (n_910, n_2590, n_905);
  nand g2585 (n_2591, n_903, n_904);
  nand g2586 (n_2592, n_905, n_904);
  nand g2587 (n_2593, n_903, n_905);
  nand g2588 (n_923, n_2591, n_2592, n_2593);
  xor g2589 (n_2594, n_906, n_907);
  xor g2590 (n_912, n_2594, n_908);
  nand g2591 (n_2595, n_906, n_907);
  nand g2592 (n_2596, n_908, n_907);
  nand g2593 (n_2597, n_906, n_908);
  nand g2594 (n_925, n_2595, n_2596, n_2597);
  xor g2595 (n_2598, n_909, n_910);
  xor g2596 (n_913, n_2598, n_911);
  nand g2597 (n_2599, n_909, n_910);
  nand g2598 (n_2600, n_911, n_910);
  nand g2599 (n_2601, n_909, n_911);
  nand g2600 (n_928, n_2599, n_2600, n_2601);
  xor g2601 (n_2602, n_912, n_913);
  xor g2602 (n_185, n_2602, n_914);
  nand g2603 (n_2603, n_912, n_913);
  nand g2604 (n_2604, n_914, n_913);
  nand g2605 (n_2605, n_912, n_914);
  nand g2606 (n_98, n_2603, n_2604, n_2605);
  xor g2607 (n_2606, A[55], A[53]);
  xor g2608 (n_919, n_2606, A[49]);
  nand g2609 (n_2607, A[55], A[53]);
  nand g2610 (n_2608, A[49], A[53]);
  nand g2611 (n_2609, A[55], A[49]);
  nand g2612 (n_929, n_2607, n_2608, n_2609);
  xor g2614 (n_920, n_2158, A[47]);
  nand g2616 (n_2612, A[47], A[39]);
  nand g2618 (n_930, n_2159, n_2612, n_2353);
  xor g2619 (n_2614, A[37], A[51]);
  xor g2620 (n_918, n_2614, A[45]);
  nand g2621 (n_2615, A[37], A[51]);
  nand g2624 (n_931, n_2615, n_2481, n_2548);
  xor g2625 (n_2618, A[43], n_915);
  xor g2626 (n_922, n_2618, n_916);
  nand g2627 (n_2619, A[43], n_915);
  nand g2628 (n_2620, n_916, n_915);
  nand g2629 (n_2621, A[43], n_916);
  nand g2630 (n_935, n_2619, n_2620, n_2621);
  xor g2631 (n_2622, n_917, n_918);
  xor g2632 (n_924, n_2622, n_919);
  nand g2633 (n_2623, n_917, n_918);
  nand g2634 (n_2624, n_919, n_918);
  nand g2635 (n_2625, n_917, n_919);
  nand g2636 (n_937, n_2623, n_2624, n_2625);
  xor g2637 (n_2626, n_920, n_921);
  xor g2638 (n_926, n_2626, n_922);
  nand g2639 (n_2627, n_920, n_921);
  nand g2640 (n_2628, n_922, n_921);
  nand g2641 (n_2629, n_920, n_922);
  nand g2642 (n_939, n_2627, n_2628, n_2629);
  xor g2643 (n_2630, n_923, n_924);
  xor g2644 (n_927, n_2630, n_925);
  nand g2645 (n_2631, n_923, n_924);
  nand g2646 (n_2632, n_925, n_924);
  nand g2647 (n_2633, n_923, n_925);
  nand g2648 (n_942, n_2631, n_2632, n_2633);
  xor g2649 (n_2634, n_926, n_927);
  xor g2650 (n_184, n_2634, n_928);
  nand g2651 (n_2635, n_926, n_927);
  nand g2652 (n_2636, n_928, n_927);
  nand g2653 (n_2637, n_926, n_928);
  nand g2654 (n_97, n_2635, n_2636, n_2637);
  xor g2655 (n_2638, A[56], A[54]);
  xor g2656 (n_933, n_2638, A[50]);
  nand g2657 (n_2639, A[56], A[54]);
  nand g2658 (n_2640, A[50], A[54]);
  nand g2659 (n_2641, A[56], A[50]);
  nand g2660 (n_943, n_2639, n_2640, n_2641);
  xor g2662 (n_934, n_2190, A[48]);
  nand g2664 (n_2644, A[48], A[40]);
  nand g2666 (n_944, n_2191, n_2644, n_2385);
  xor g2667 (n_2646, A[38], A[52]);
  xor g2668 (n_932, n_2646, A[46]);
  nand g2669 (n_2647, A[38], A[52]);
  nand g2672 (n_945, n_2647, n_2513, n_2580);
  xor g2673 (n_2650, A[44], n_929);
  xor g2674 (n_936, n_2650, n_930);
  nand g2675 (n_2651, A[44], n_929);
  nand g2676 (n_2652, n_930, n_929);
  nand g2677 (n_2653, A[44], n_930);
  nand g2678 (n_949, n_2651, n_2652, n_2653);
  xor g2679 (n_2654, n_931, n_932);
  xor g2680 (n_938, n_2654, n_933);
  nand g2681 (n_2655, n_931, n_932);
  nand g2682 (n_2656, n_933, n_932);
  nand g2683 (n_2657, n_931, n_933);
  nand g2684 (n_951, n_2655, n_2656, n_2657);
  xor g2685 (n_2658, n_934, n_935);
  xor g2686 (n_940, n_2658, n_936);
  nand g2687 (n_2659, n_934, n_935);
  nand g2688 (n_2660, n_936, n_935);
  nand g2689 (n_2661, n_934, n_936);
  nand g2690 (n_953, n_2659, n_2660, n_2661);
  xor g2691 (n_2662, n_937, n_938);
  xor g2692 (n_941, n_2662, n_939);
  nand g2693 (n_2663, n_937, n_938);
  nand g2694 (n_2664, n_939, n_938);
  nand g2695 (n_2665, n_937, n_939);
  nand g2696 (n_956, n_2663, n_2664, n_2665);
  xor g2697 (n_2666, n_940, n_941);
  xor g2698 (n_183, n_2666, n_942);
  nand g2699 (n_2667, n_940, n_941);
  nand g2700 (n_2668, n_942, n_941);
  nand g2701 (n_2669, n_940, n_942);
  nand g2702 (n_96, n_2667, n_2668, n_2669);
  xor g2703 (n_2670, A[57], A[55]);
  xor g2704 (n_947, n_2670, A[51]);
  nand g2705 (n_2671, A[57], A[55]);
  nand g2706 (n_2672, A[51], A[55]);
  nand g2707 (n_2673, A[57], A[51]);
  nand g2708 (n_957, n_2671, n_2672, n_2673);
  xor g2710 (n_948, n_2222, A[49]);
  nand g2712 (n_2676, A[49], A[41]);
  nand g2714 (n_958, n_2223, n_2676, n_2417);
  xor g2715 (n_2678, A[39], A[53]);
  xor g2716 (n_946, n_2678, A[47]);
  nand g2717 (n_2679, A[39], A[53]);
  nand g2720 (n_959, n_2679, n_2545, n_2612);
  xor g2721 (n_2682, A[45], n_943);
  xor g2722 (n_950, n_2682, n_944);
  nand g2723 (n_2683, A[45], n_943);
  nand g2724 (n_2684, n_944, n_943);
  nand g2725 (n_2685, A[45], n_944);
  nand g2726 (n_963, n_2683, n_2684, n_2685);
  xor g2727 (n_2686, n_945, n_946);
  xor g2728 (n_952, n_2686, n_947);
  nand g2729 (n_2687, n_945, n_946);
  nand g2730 (n_2688, n_947, n_946);
  nand g2731 (n_2689, n_945, n_947);
  nand g2732 (n_965, n_2687, n_2688, n_2689);
  xor g2733 (n_2690, n_948, n_949);
  xor g2734 (n_954, n_2690, n_950);
  nand g2735 (n_2691, n_948, n_949);
  nand g2736 (n_2692, n_950, n_949);
  nand g2737 (n_2693, n_948, n_950);
  nand g2738 (n_967, n_2691, n_2692, n_2693);
  xor g2739 (n_2694, n_951, n_952);
  xor g2740 (n_955, n_2694, n_953);
  nand g2741 (n_2695, n_951, n_952);
  nand g2742 (n_2696, n_953, n_952);
  nand g2743 (n_2697, n_951, n_953);
  nand g2744 (n_970, n_2695, n_2696, n_2697);
  xor g2745 (n_2698, n_954, n_955);
  xor g2746 (n_182, n_2698, n_956);
  nand g2747 (n_2699, n_954, n_955);
  nand g2748 (n_2700, n_956, n_955);
  nand g2749 (n_2701, n_954, n_956);
  nand g2750 (n_95, n_2699, n_2700, n_2701);
  xor g2751 (n_2702, A[58], A[56]);
  xor g2752 (n_961, n_2702, A[52]);
  nand g2753 (n_2703, A[58], A[56]);
  nand g2754 (n_2704, A[52], A[56]);
  nand g2755 (n_2705, A[58], A[52]);
  nand g2756 (n_971, n_2703, n_2704, n_2705);
  xor g2758 (n_962, n_2254, A[50]);
  nand g2760 (n_2708, A[50], A[42]);
  nand g2762 (n_972, n_2255, n_2708, n_2449);
  xor g2763 (n_2710, A[40], A[54]);
  xor g2764 (n_960, n_2710, A[48]);
  nand g2765 (n_2711, A[40], A[54]);
  nand g2768 (n_973, n_2711, n_2577, n_2644);
  xor g2769 (n_2714, A[46], n_957);
  xor g2770 (n_964, n_2714, n_958);
  nand g2771 (n_2715, A[46], n_957);
  nand g2772 (n_2716, n_958, n_957);
  nand g2773 (n_2717, A[46], n_958);
  nand g2774 (n_977, n_2715, n_2716, n_2717);
  xor g2775 (n_2718, n_959, n_960);
  xor g2776 (n_966, n_2718, n_961);
  nand g2777 (n_2719, n_959, n_960);
  nand g2778 (n_2720, n_961, n_960);
  nand g2779 (n_2721, n_959, n_961);
  nand g2780 (n_979, n_2719, n_2720, n_2721);
  xor g2781 (n_2722, n_962, n_963);
  xor g2782 (n_968, n_2722, n_964);
  nand g2783 (n_2723, n_962, n_963);
  nand g2784 (n_2724, n_964, n_963);
  nand g2785 (n_2725, n_962, n_964);
  nand g2786 (n_981, n_2723, n_2724, n_2725);
  xor g2787 (n_2726, n_965, n_966);
  xor g2788 (n_969, n_2726, n_967);
  nand g2789 (n_2727, n_965, n_966);
  nand g2790 (n_2728, n_967, n_966);
  nand g2791 (n_2729, n_965, n_967);
  nand g2792 (n_984, n_2727, n_2728, n_2729);
  xor g2793 (n_2730, n_968, n_969);
  xor g2794 (n_181, n_2730, n_970);
  nand g2795 (n_2731, n_968, n_969);
  nand g2796 (n_2732, n_970, n_969);
  nand g2797 (n_2733, n_968, n_970);
  nand g2798 (n_94, n_2731, n_2732, n_2733);
  xor g2799 (n_2734, A[59], A[57]);
  xor g2800 (n_975, n_2734, A[53]);
  nand g2801 (n_2735, A[59], A[57]);
  nand g2802 (n_2736, A[53], A[57]);
  nand g2803 (n_2737, A[59], A[53]);
  nand g2804 (n_985, n_2735, n_2736, n_2737);
  xor g2806 (n_976, n_2286, A[51]);
  nand g2808 (n_2740, A[51], A[43]);
  nand g2810 (n_987, n_2287, n_2740, n_2481);
  xor g2811 (n_2742, A[41], A[55]);
  xor g2812 (n_974, n_2742, A[49]);
  nand g2813 (n_2743, A[41], A[55]);
  nand g2816 (n_986, n_2743, n_2609, n_2676);
  xor g2817 (n_2746, A[47], n_971);
  xor g2818 (n_978, n_2746, n_972);
  nand g2819 (n_2747, A[47], n_971);
  nand g2820 (n_2748, n_972, n_971);
  nand g2821 (n_2749, A[47], n_972);
  nand g2822 (n_991, n_2747, n_2748, n_2749);
  xor g2823 (n_2750, n_973, n_974);
  xor g2824 (n_980, n_2750, n_975);
  nand g2825 (n_2751, n_973, n_974);
  nand g2826 (n_2752, n_975, n_974);
  nand g2827 (n_2753, n_973, n_975);
  nand g2828 (n_993, n_2751, n_2752, n_2753);
  xor g2829 (n_2754, n_976, n_977);
  xor g2830 (n_982, n_2754, n_978);
  nand g2831 (n_2755, n_976, n_977);
  nand g2832 (n_2756, n_978, n_977);
  nand g2833 (n_2757, n_976, n_978);
  nand g2834 (n_996, n_2755, n_2756, n_2757);
  xor g2835 (n_2758, n_979, n_980);
  xor g2836 (n_983, n_2758, n_981);
  nand g2837 (n_2759, n_979, n_980);
  nand g2838 (n_2760, n_981, n_980);
  nand g2839 (n_2761, n_979, n_981);
  nand g2840 (n_998, n_2759, n_2760, n_2761);
  xor g2841 (n_2762, n_982, n_983);
  xor g2842 (n_180, n_2762, n_984);
  nand g2843 (n_2763, n_982, n_983);
  nand g2844 (n_2764, n_984, n_983);
  nand g2845 (n_2765, n_982, n_984);
  nand g2846 (n_93, n_2763, n_2764, n_2765);
  xor g2847 (n_2766, A[58], A[54]);
  xor g2848 (n_989, n_2766, A[46]);
  nand g2849 (n_2767, A[58], A[54]);
  nand g2850 (n_2768, A[46], A[54]);
  nand g2851 (n_2769, A[58], A[46]);
  nand g2852 (n_999, n_2767, n_2768, n_2769);
  xor g2853 (n_2770, A[44], A[52]);
  xor g2854 (n_990, n_2770, A[42]);
  nand g2855 (n_2771, A[44], A[52]);
  nand g2856 (n_2772, A[42], A[52]);
  nand g2858 (n_1001, n_2771, n_2772, n_2255);
  xor g2859 (n_2774, A[56], A[50]);
  xor g2860 (n_988, n_2774, A[48]);
  nand g2863 (n_2777, A[56], A[48]);
  nand g2864 (n_1000, n_2641, n_2447, n_2777);
  xor g2865 (n_2778, A[60], n_985);
  xor g2866 (n_992, n_2778, n_986);
  nand g2867 (n_2779, A[60], n_985);
  nand g2868 (n_2780, n_986, n_985);
  nand g2869 (n_2781, A[60], n_986);
  nand g2870 (n_1005, n_2779, n_2780, n_2781);
  xor g2871 (n_2782, n_987, n_988);
  xor g2872 (n_994, n_2782, n_989);
  nand g2873 (n_2783, n_987, n_988);
  nand g2874 (n_2784, n_989, n_988);
  nand g2875 (n_2785, n_987, n_989);
  nand g2876 (n_1007, n_2783, n_2784, n_2785);
  xor g2877 (n_2786, n_990, n_991);
  xor g2878 (n_995, n_2786, n_992);
  nand g2879 (n_2787, n_990, n_991);
  nand g2880 (n_2788, n_992, n_991);
  nand g2881 (n_2789, n_990, n_992);
  nand g2882 (n_1010, n_2787, n_2788, n_2789);
  xor g2883 (n_2790, n_993, n_994);
  xor g2884 (n_997, n_2790, n_995);
  nand g2885 (n_2791, n_993, n_994);
  nand g2886 (n_2792, n_995, n_994);
  nand g2887 (n_2793, n_993, n_995);
  nand g2888 (n_1012, n_2791, n_2792, n_2793);
  xor g2889 (n_2794, n_996, n_997);
  xor g2890 (n_179, n_2794, n_998);
  nand g2891 (n_2795, n_996, n_997);
  nand g2892 (n_2796, n_998, n_997);
  nand g2893 (n_2797, n_996, n_998);
  nand g2894 (n_92, n_2795, n_2796, n_2797);
  xor g2895 (n_2798, A[59], A[55]);
  xor g2896 (n_1003, n_2798, A[47]);
  nand g2897 (n_2799, A[59], A[55]);
  nand g2898 (n_2800, A[47], A[55]);
  nand g2899 (n_2801, A[59], A[47]);
  nand g2900 (n_1014, n_2799, n_2800, n_2801);
  xor g2901 (n_2802, A[45], A[53]);
  xor g2902 (n_1004, n_2802, A[43]);
  nand g2903 (n_2803, A[45], A[53]);
  nand g2904 (n_2804, A[43], A[53]);
  nand g2906 (n_1015, n_2803, n_2804, n_2287);
  xor g2907 (n_2806, A[57], A[51]);
  xor g2908 (n_1002, n_2806, A[49]);
  nand g2911 (n_2809, A[57], A[49]);
  nand g2912 (n_1013, n_2673, n_2479, n_2809);
  xor g2913 (n_2810, A[61], n_999);
  xor g2914 (n_1006, n_2810, n_1000);
  nand g2915 (n_2811, A[61], n_999);
  nand g2916 (n_2812, n_1000, n_999);
  nand g2917 (n_2813, A[61], n_1000);
  nand g2918 (n_1019, n_2811, n_2812, n_2813);
  xor g2919 (n_2814, n_1001, n_1002);
  xor g2920 (n_1008, n_2814, n_1003);
  nand g2921 (n_2815, n_1001, n_1002);
  nand g2922 (n_2816, n_1003, n_1002);
  nand g2923 (n_2817, n_1001, n_1003);
  nand g2924 (n_1020, n_2815, n_2816, n_2817);
  xor g2925 (n_2818, n_1004, n_1005);
  xor g2926 (n_1009, n_2818, n_1006);
  nand g2927 (n_2819, n_1004, n_1005);
  nand g2928 (n_2820, n_1006, n_1005);
  nand g2929 (n_2821, n_1004, n_1006);
  nand g2930 (n_1024, n_2819, n_2820, n_2821);
  xor g2931 (n_2822, n_1007, n_1008);
  xor g2932 (n_1011, n_2822, n_1009);
  nand g2933 (n_2823, n_1007, n_1008);
  nand g2934 (n_2824, n_1009, n_1008);
  nand g2935 (n_2825, n_1007, n_1009);
  nand g2936 (n_1026, n_2823, n_2824, n_2825);
  xor g2937 (n_2826, n_1010, n_1011);
  xor g2938 (n_178, n_2826, n_1012);
  nand g2939 (n_2827, n_1010, n_1011);
  nand g2940 (n_2828, n_1012, n_1011);
  nand g2941 (n_2829, n_1010, n_1012);
  nand g2942 (n_91, n_2827, n_2828, n_2829);
  xor g2944 (n_1016, n_2702, A[48]);
  nand g2947 (n_2833, A[58], A[48]);
  nand g2948 (n_1027, n_2703, n_2777, n_2833);
  xor g2949 (n_2834, A[46], A[54]);
  xor g2950 (n_1018, n_2834, A[44]);
  nand g2952 (n_2836, A[44], A[54]);
  nand g2954 (n_1028, n_2768, n_2836, n_2319);
  xor g2956 (n_1017, n_2510, A[60]);
  nand g2958 (n_2840, A[60], A[50]);
  nand g2959 (n_2841, A[52], A[60]);
  nand g2960 (n_1030, n_2511, n_2840, n_2841);
  xor g2961 (n_2842, A[62], n_1013);
  xor g2962 (n_1021, n_2842, n_1014);
  nand g2963 (n_2843, A[62], n_1013);
  nand g2964 (n_2844, n_1014, n_1013);
  nand g2965 (n_2845, A[62], n_1014);
  nand g2966 (n_1033, n_2843, n_2844, n_2845);
  xor g2967 (n_2846, n_1015, n_1016);
  xor g2968 (n_1022, n_2846, n_1017);
  nand g2969 (n_2847, n_1015, n_1016);
  nand g2970 (n_2848, n_1017, n_1016);
  nand g2971 (n_2849, n_1015, n_1017);
  nand g2972 (n_1034, n_2847, n_2848, n_2849);
  xor g2973 (n_2850, n_1018, n_1019);
  xor g2974 (n_1023, n_2850, n_1020);
  nand g2975 (n_2851, n_1018, n_1019);
  nand g2976 (n_2852, n_1020, n_1019);
  nand g2977 (n_2853, n_1018, n_1020);
  nand g2978 (n_1038, n_2851, n_2852, n_2853);
  xor g2979 (n_2854, n_1021, n_1022);
  xor g2980 (n_1025, n_2854, n_1023);
  nand g2981 (n_2855, n_1021, n_1022);
  nand g2982 (n_2856, n_1023, n_1022);
  nand g2983 (n_2857, n_1021, n_1023);
  nand g2984 (n_1040, n_2855, n_2856, n_2857);
  xor g2985 (n_2858, n_1024, n_1025);
  xor g2986 (n_177, n_2858, n_1026);
  nand g2987 (n_2859, n_1024, n_1025);
  nand g2988 (n_2860, n_1026, n_1025);
  nand g2989 (n_2861, n_1024, n_1026);
  nand g2990 (n_90, n_2859, n_2860, n_2861);
  xor g2992 (n_1029, n_2734, A[49]);
  nand g2995 (n_2865, A[59], A[49]);
  nand g2996 (n_1041, n_2735, n_2809, n_2865);
  xor g2997 (n_2866, A[47], A[55]);
  xor g2998 (n_1032, n_2866, A[45]);
  nand g3000 (n_2868, A[45], A[55]);
  nand g3002 (n_1042, n_2800, n_2868, n_2351);
  xor g3004 (n_1031, n_2542, A[61]);
  nand g3006 (n_2872, A[61], A[51]);
  nand g3007 (n_2873, A[53], A[61]);
  nand g3008 (n_1044, n_2543, n_2872, n_2873);
  xor g3009 (n_2874, A[63], n_1027);
  xor g3010 (n_1035, n_2874, n_1028);
  nand g3011 (n_2875, A[63], n_1027);
  nand g3012 (n_2876, n_1028, n_1027);
  nand g3013 (n_2877, A[63], n_1028);
  nand g3014 (n_1047, n_2875, n_2876, n_2877);
  xor g3015 (n_2878, n_1029, n_1030);
  xor g3016 (n_1036, n_2878, n_1031);
  nand g3017 (n_2879, n_1029, n_1030);
  nand g3018 (n_2880, n_1031, n_1030);
  nand g3019 (n_2881, n_1029, n_1031);
  nand g3020 (n_1048, n_2879, n_2880, n_2881);
  xor g3021 (n_2882, n_1032, n_1033);
  xor g3022 (n_1037, n_2882, n_1034);
  nand g3023 (n_2883, n_1032, n_1033);
  nand g3024 (n_2884, n_1034, n_1033);
  nand g3025 (n_2885, n_1032, n_1034);
  nand g3026 (n_1052, n_2883, n_2884, n_2885);
  xor g3027 (n_2886, n_1035, n_1036);
  xor g3028 (n_1039, n_2886, n_1037);
  nand g3029 (n_2887, n_1035, n_1036);
  nand g3030 (n_2888, n_1037, n_1036);
  nand g3031 (n_2889, n_1035, n_1037);
  nand g3032 (n_1054, n_2887, n_2888, n_2889);
  xor g3033 (n_2890, n_1038, n_1039);
  xor g3034 (n_176, n_2890, n_1040);
  nand g3035 (n_2891, n_1038, n_1039);
  nand g3036 (n_2892, n_1040, n_1039);
  nand g3037 (n_2893, n_1038, n_1040);
  nand g3038 (n_89, n_2891, n_2892, n_2893);
  xor g3040 (n_1043, n_2702, A[50]);
  nand g3043 (n_2897, A[58], A[50]);
  nand g3044 (n_1055, n_2703, n_2641, n_2897);
  xor g3046 (n_1045, n_2382, A[54]);
  nand g3050 (n_1056, n_2383, n_2768, n_2577);
  xor g3051 (n_2902, A[52], A[62]);
  xor g3052 (n_1046, n_2902, A[64]);
  nand g3053 (n_2903, A[52], A[62]);
  nand g3054 (n_2904, A[64], A[62]);
  nand g3055 (n_2905, A[52], A[64]);
  nand g3056 (n_1058, n_2903, n_2904, n_2905);
  xor g3057 (n_2906, A[60], n_1041);
  xor g3058 (n_1049, n_2906, n_1042);
  nand g3059 (n_2907, A[60], n_1041);
  nand g3060 (n_2908, n_1042, n_1041);
  nand g3061 (n_2909, A[60], n_1042);
  nand g3062 (n_1061, n_2907, n_2908, n_2909);
  xor g3063 (n_2910, n_1043, n_1044);
  xor g3064 (n_1050, n_2910, n_1045);
  nand g3065 (n_2911, n_1043, n_1044);
  nand g3066 (n_2912, n_1045, n_1044);
  nand g3067 (n_2913, n_1043, n_1045);
  nand g3068 (n_1062, n_2911, n_2912, n_2913);
  xor g3069 (n_2914, n_1046, n_1047);
  xor g3070 (n_1051, n_2914, n_1048);
  nand g3071 (n_2915, n_1046, n_1047);
  nand g3072 (n_2916, n_1048, n_1047);
  nand g3073 (n_2917, n_1046, n_1048);
  nand g3074 (n_1066, n_2915, n_2916, n_2917);
  xor g3075 (n_2918, n_1049, n_1050);
  xor g3076 (n_1053, n_2918, n_1051);
  nand g3077 (n_2919, n_1049, n_1050);
  nand g3078 (n_2920, n_1051, n_1050);
  nand g3079 (n_2921, n_1049, n_1051);
  nand g3080 (n_1068, n_2919, n_2920, n_2921);
  xor g3081 (n_2922, n_1052, n_1053);
  xor g3082 (n_175, n_2922, n_1054);
  nand g3083 (n_2923, n_1052, n_1053);
  nand g3084 (n_2924, n_1054, n_1053);
  nand g3085 (n_2925, n_1052, n_1054);
  nand g3086 (n_88, n_2923, n_2924, n_2925);
  xor g3088 (n_1057, n_2734, A[51]);
  nand g3091 (n_2929, A[59], A[51]);
  nand g3092 (n_1072, n_2735, n_2673, n_2929);
  xor g3094 (n_1059, n_2414, A[55]);
  nand g3098 (n_1071, n_2415, n_2800, n_2609);
  xor g3099 (n_2934, A[53], A[63]);
  xor g3100 (n_1060, n_2934, A[65]);
  nand g3101 (n_2935, A[53], A[63]);
  nand g3102 (n_2936, A[65], A[63]);
  nand g3103 (n_2937, A[53], A[65]);
  nand g3104 (n_1075, n_2935, n_2936, n_2937);
  xor g3105 (n_2938, A[61], n_1055);
  xor g3106 (n_1063, n_2938, n_1056);
  nand g3107 (n_2939, A[61], n_1055);
  nand g3108 (n_2940, n_1056, n_1055);
  nand g3109 (n_2941, A[61], n_1056);
  nand g3110 (n_1077, n_2939, n_2940, n_2941);
  xor g3111 (n_2942, n_1057, n_1058);
  xor g3112 (n_1064, n_2942, n_1059);
  nand g3113 (n_2943, n_1057, n_1058);
  nand g3114 (n_2944, n_1059, n_1058);
  nand g3115 (n_2945, n_1057, n_1059);
  nand g3116 (n_1078, n_2943, n_2944, n_2945);
  xor g3117 (n_2946, n_1060, n_1061);
  xor g3118 (n_1065, n_2946, n_1062);
  nand g3119 (n_2947, n_1060, n_1061);
  nand g3120 (n_2948, n_1062, n_1061);
  nand g3121 (n_2949, n_1060, n_1062);
  nand g3122 (n_1082, n_2947, n_2948, n_2949);
  xor g3123 (n_2950, n_1063, n_1064);
  xor g3124 (n_1067, n_2950, n_1065);
  nand g3125 (n_2951, n_1063, n_1064);
  nand g3126 (n_2952, n_1065, n_1064);
  nand g3127 (n_2953, n_1063, n_1065);
  nand g3128 (n_1084, n_2951, n_2952, n_2953);
  xor g3129 (n_2954, n_1066, n_1067);
  xor g3130 (n_174, n_2954, n_1068);
  nand g3131 (n_2955, n_1066, n_1067);
  nand g3132 (n_2956, n_1068, n_1067);
  nand g3133 (n_2957, n_1066, n_1068);
  nand g3134 (n_87, n_2955, n_2956, n_2957);
  xor g3137 (n_2958, A[66], A[52]);
  xor g3138 (n_1073, n_2958, A[50]);
  nand g3139 (n_2959, A[66], A[52]);
  nand g3141 (n_2961, A[66], A[50]);
  nand g3142 (n_1089, n_2959, n_2511, n_2961);
  xor g3143 (n_2962, A[58], A[48]);
  xor g3144 (n_1074, n_2962, A[56]);
  xor g3149 (n_2966, A[54], A[60]);
  xor g3150 (n_1076, n_2966, A[64]);
  nand g3151 (n_2967, A[54], A[60]);
  nand g3152 (n_2968, A[64], A[60]);
  nand g3153 (n_2969, A[54], A[64]);
  nand g3154 (n_1092, n_2967, n_2968, n_2969);
  xor g3155 (n_2970, A[62], n_1071);
  xor g3156 (n_1079, n_2970, n_1072);
  nand g3157 (n_2971, A[62], n_1071);
  nand g3158 (n_2972, n_1072, n_1071);
  nand g3159 (n_2973, A[62], n_1072);
  nand g3160 (n_1094, n_2971, n_2972, n_2973);
  xor g3161 (n_2974, n_1073, n_1074);
  xor g3162 (n_1080, n_2974, n_1075);
  nand g3163 (n_2975, n_1073, n_1074);
  nand g3164 (n_2976, n_1075, n_1074);
  nand g3165 (n_2977, n_1073, n_1075);
  nand g3166 (n_1095, n_2975, n_2976, n_2977);
  xor g3167 (n_2978, n_1076, n_1077);
  xor g3168 (n_1081, n_2978, n_1078);
  nand g3169 (n_2979, n_1076, n_1077);
  nand g3170 (n_2980, n_1078, n_1077);
  nand g3171 (n_2981, n_1076, n_1078);
  nand g3172 (n_1099, n_2979, n_2980, n_2981);
  xor g3173 (n_2982, n_1079, n_1080);
  xor g3174 (n_1083, n_2982, n_1081);
  nand g3175 (n_2983, n_1079, n_1080);
  nand g3176 (n_2984, n_1081, n_1080);
  nand g3177 (n_2985, n_1079, n_1081);
  nand g3178 (n_1101, n_2983, n_2984, n_2985);
  xor g3179 (n_2986, n_1082, n_1083);
  xor g3180 (n_173, n_2986, n_1084);
  nand g3181 (n_2987, n_1082, n_1083);
  nand g3182 (n_2988, n_1084, n_1083);
  nand g3183 (n_2989, n_1082, n_1084);
  nand g3184 (n_86, n_2987, n_2988, n_2989);
  xor g3188 (n_1090, n_2478, A[66]);
  nand g3190 (n_2992, A[66], A[49]);
  nand g3191 (n_2993, A[51], A[66]);
  nand g3192 (n_1103, n_2479, n_2992, n_2993);
  xor g3194 (n_1091, n_2734, A[55]);
  nand g3198 (n_1104, n_2735, n_2671, n_2799);
  xor g3205 (n_3002, A[61], n_1027);
  xor g3206 (n_1096, n_3002, n_1089);
  nand g3207 (n_3003, A[61], n_1027);
  nand g3208 (n_3004, n_1089, n_1027);
  nand g3209 (n_3005, A[61], n_1089);
  nand g3210 (n_1109, n_3003, n_3004, n_3005);
  xor g3211 (n_3006, n_1090, n_1091);
  xor g3212 (n_1097, n_3006, n_1092);
  nand g3213 (n_3007, n_1090, n_1091);
  nand g3214 (n_3008, n_1092, n_1091);
  nand g3215 (n_3009, n_1090, n_1092);
  nand g3216 (n_1110, n_3007, n_3008, n_3009);
  xor g3217 (n_3010, n_1060, n_1094);
  xor g3218 (n_1098, n_3010, n_1095);
  nand g3219 (n_3011, n_1060, n_1094);
  nand g3220 (n_3012, n_1095, n_1094);
  nand g3221 (n_3013, n_1060, n_1095);
  nand g3222 (n_1114, n_3011, n_3012, n_3013);
  xor g3223 (n_3014, n_1096, n_1097);
  xor g3224 (n_1100, n_3014, n_1098);
  nand g3225 (n_3015, n_1096, n_1097);
  nand g3226 (n_3016, n_1098, n_1097);
  nand g3227 (n_3017, n_1096, n_1098);
  nand g3228 (n_1116, n_3015, n_3016, n_3017);
  xor g3229 (n_3018, n_1099, n_1100);
  xor g3230 (n_172, n_3018, n_1101);
  nand g3231 (n_3019, n_1099, n_1100);
  nand g3232 (n_3020, n_1101, n_1100);
  nand g3233 (n_3021, n_1099, n_1101);
  nand g3234 (n_85, n_3019, n_3020, n_3021);
  xor g3236 (n_1105, n_3022, A[52]);
  nand g3240 (n_1119, n_3023, n_2705, n_3025);
  xor g3242 (n_1107, n_3026, A[56]);
  nand g3246 (n_1120, n_3027, n_3028, n_2641);
  xor g3253 (n_3034, A[62], n_1103);
  xor g3254 (n_1111, n_3034, n_1104);
  nand g3255 (n_3035, A[62], n_1103);
  nand g3256 (n_3036, n_1104, n_1103);
  nand g3257 (n_3037, A[62], n_1104);
  nand g3258 (n_1124, n_3035, n_3036, n_3037);
  xor g3259 (n_3038, n_1105, n_1075);
  xor g3260 (n_1112, n_3038, n_1107);
  nand g3261 (n_3039, n_1105, n_1075);
  nand g3262 (n_3040, n_1107, n_1075);
  nand g3263 (n_3041, n_1105, n_1107);
  nand g3264 (n_1126, n_3039, n_3040, n_3041);
  xor g3265 (n_3042, n_1076, n_1109);
  xor g3266 (n_1113, n_3042, n_1110);
  nand g3267 (n_3043, n_1076, n_1109);
  nand g3268 (n_3044, n_1110, n_1109);
  nand g3269 (n_3045, n_1076, n_1110);
  nand g3270 (n_1128, n_3043, n_3044, n_3045);
  xor g3271 (n_3046, n_1111, n_1112);
  xor g3272 (n_1115, n_3046, n_1113);
  nand g3273 (n_3047, n_1111, n_1112);
  nand g3274 (n_3048, n_1113, n_1112);
  nand g3275 (n_3049, n_1111, n_1113);
  nand g3276 (n_1131, n_3047, n_3048, n_3049);
  xor g3277 (n_3050, n_1114, n_1115);
  xor g3278 (n_171, n_3050, n_1116);
  nand g3279 (n_3051, n_1114, n_1115);
  nand g3280 (n_3052, n_1116, n_1115);
  nand g3281 (n_3053, n_1114, n_1116);
  nand g3282 (n_84, n_3051, n_3052, n_3053);
  xor g3286 (n_1122, n_2806, A[55]);
  xor g3298 (n_1125, n_3062, n_1119);
  nand g3301 (n_3065, A[61], n_1119);
  nand g3302 (n_1138, n_3063, n_3064, n_3065);
  xor g3303 (n_3066, n_1120, n_1092);
  xor g3304 (n_1127, n_3066, n_1122);
  nand g3305 (n_3067, n_1120, n_1092);
  nand g3306 (n_3068, n_1122, n_1092);
  nand g3307 (n_3069, n_1120, n_1122);
  nand g3308 (n_1139, n_3067, n_3068, n_3069);
  xor g3309 (n_3070, n_1060, n_1124);
  xor g3310 (n_1129, n_3070, n_1125);
  nand g3311 (n_3071, n_1060, n_1124);
  nand g3312 (n_3072, n_1125, n_1124);
  nand g3313 (n_3073, n_1060, n_1125);
  nand g3314 (n_1141, n_3071, n_3072, n_3073);
  xor g3315 (n_3074, n_1126, n_1127);
  xor g3316 (n_1130, n_3074, n_1128);
  nand g3317 (n_3075, n_1126, n_1127);
  nand g3318 (n_3076, n_1128, n_1127);
  nand g3319 (n_3077, n_1126, n_1128);
  nand g3320 (n_1144, n_3075, n_3076, n_3077);
  xor g3321 (n_3078, n_1129, n_1130);
  xor g3322 (n_170, n_3078, n_1131);
  nand g3323 (n_3079, n_1129, n_1130);
  nand g3324 (n_3080, n_1131, n_1130);
  nand g3325 (n_3081, n_1129, n_1131);
  nand g3326 (n_83, n_3079, n_3080, n_3081);
  xor g3334 (n_1135, n_2638, A[60]);
  nand g3337 (n_3089, A[56], A[60]);
  nand g3338 (n_1148, n_2639, n_2967, n_3089);
  xor g3339 (n_3090, A[64], A[62]);
  xor g3340 (n_1137, n_3090, A[59]);
  nand g3342 (n_3092, A[59], A[62]);
  nand g3343 (n_3093, A[64], A[59]);
  nand g3344 (n_1151, n_2904, n_3092, n_3093);
  xor g3345 (n_3094, n_957, n_1075);
  xor g3346 (n_1140, n_3094, n_1135);
  nand g3347 (n_3095, n_957, n_1075);
  nand g3348 (n_3096, n_1135, n_1075);
  nand g3349 (n_3097, n_957, n_1135);
  nand g3350 (n_1153, n_3095, n_3096, n_3097);
  xor g3351 (n_3098, n_1105, n_1137);
  xor g3352 (n_1142, n_3098, n_1138);
  nand g3353 (n_3099, n_1105, n_1137);
  nand g3354 (n_3100, n_1138, n_1137);
  nand g3355 (n_3101, n_1105, n_1138);
  nand g3356 (n_1155, n_3099, n_3100, n_3101);
  xor g3357 (n_3102, n_1139, n_1140);
  xor g3358 (n_1143, n_3102, n_1141);
  nand g3359 (n_3103, n_1139, n_1140);
  nand g3360 (n_3104, n_1141, n_1140);
  nand g3361 (n_3105, n_1139, n_1141);
  nand g3362 (n_1157, n_3103, n_3104, n_3105);
  xor g3363 (n_3106, n_1142, n_1143);
  xor g3364 (n_169, n_3106, n_1144);
  nand g3365 (n_3107, n_1142, n_1143);
  nand g3366 (n_3108, n_1144, n_1143);
  nand g3367 (n_3109, n_1142, n_1144);
  nand g3368 (n_82, n_3107, n_3108, n_3109);
  xor g3372 (n_1149, n_2670, A[53]);
  nand g3376 (n_1159, n_2671, n_2607, n_2736);
  xor g3377 (n_3114, A[63], A[65]);
  xor g3378 (n_1150, n_3114, A[61]);
  nand g3380 (n_3116, A[61], A[65]);
  nand g3381 (n_3117, A[63], A[61]);
  nand g3382 (n_1160, n_2936, n_3116, n_3117);
  xor g3384 (n_1152, n_3118, n_1148);
  nand g3386 (n_3120, n_1148, n_1119);
  nand g3388 (n_1164, n_3064, n_3120, n_3121);
  xor g3389 (n_3122, n_1149, n_1150);
  xor g3390 (n_1154, n_3122, n_1151);
  nand g3391 (n_3123, n_1149, n_1150);
  nand g3392 (n_3124, n_1151, n_1150);
  nand g3393 (n_3125, n_1149, n_1151);
  nand g3394 (n_1166, n_3123, n_3124, n_3125);
  xor g3395 (n_3126, n_1152, n_1153);
  xor g3396 (n_1156, n_3126, n_1154);
  nand g3397 (n_3127, n_1152, n_1153);
  nand g3398 (n_3128, n_1154, n_1153);
  nand g3399 (n_3129, n_1152, n_1154);
  nand g3400 (n_1168, n_3127, n_3128, n_3129);
  xor g3401 (n_3130, n_1155, n_1156);
  xor g3402 (n_168, n_3130, n_1157);
  nand g3403 (n_3131, n_1155, n_1156);
  nand g3404 (n_3132, n_1157, n_1156);
  nand g3405 (n_3133, n_1155, n_1157);
  nand g3406 (n_81, n_3131, n_3132, n_3133);
  xor g3408 (n_1161, n_3022, A[56]);
  nand g3412 (n_1171, n_3023, n_2703, n_3028);
  xor g3419 (n_3142, A[62], A[59]);
  xor g3420 (n_1163, n_3142, n_1159);
  nand g3422 (n_3144, n_1159, A[59]);
  nand g3423 (n_3145, A[62], n_1159);
  nand g3424 (n_1175, n_3092, n_3144, n_3145);
  xor g3425 (n_3146, n_1160, n_1161);
  xor g3426 (n_1165, n_3146, n_1076);
  nand g3427 (n_3147, n_1160, n_1161);
  nand g3428 (n_3148, n_1076, n_1161);
  nand g3429 (n_3149, n_1160, n_1076);
  nand g3430 (n_1176, n_3147, n_3148, n_3149);
  xor g3431 (n_3150, n_1163, n_1164);
  xor g3432 (n_1167, n_3150, n_1165);
  nand g3433 (n_3151, n_1163, n_1164);
  nand g3434 (n_3152, n_1165, n_1164);
  nand g3435 (n_3153, n_1163, n_1165);
  nand g3436 (n_1179, n_3151, n_3152, n_3153);
  xor g3437 (n_3154, n_1166, n_1167);
  xor g3438 (n_167, n_3154, n_1168);
  nand g3439 (n_3155, n_1166, n_1167);
  nand g3440 (n_3156, n_1168, n_1167);
  nand g3441 (n_3157, n_1166, n_1168);
  nand g3442 (n_80, n_3155, n_3156, n_3157);
  xor g3446 (n_1173, n_2798, A[63]);
  nand g3448 (n_3160, A[63], A[55]);
  nand g3449 (n_3161, A[59], A[63]);
  nand g3450 (n_1181, n_2799, n_3160, n_3161);
  xor g3451 (n_3162, A[65], A[61]);
  nand g3456 (n_1183, n_3116, n_3164, n_3165);
  xor g3457 (n_3166, n_1171, n_1092);
  xor g3458 (n_1177, n_3166, n_1173);
  nand g3459 (n_3167, n_1171, n_1092);
  nand g3460 (n_3168, n_1173, n_1092);
  nand g3461 (n_3169, n_1171, n_1173);
  nand g3462 (n_1185, n_3167, n_3168, n_3169);
  xor g3463 (n_3170, n_1174, n_1175);
  xor g3464 (n_1178, n_3170, n_1176);
  nand g3465 (n_3171, n_1174, n_1175);
  nand g3466 (n_3172, n_1176, n_1175);
  nand g3467 (n_3173, n_1174, n_1176);
  nand g3468 (n_1188, n_3171, n_3172, n_3173);
  xor g3469 (n_3174, n_1177, n_1178);
  xor g3470 (n_166, n_3174, n_1179);
  nand g3471 (n_3175, n_1177, n_1178);
  nand g3472 (n_3176, n_1179, n_1178);
  nand g3473 (n_3177, n_1177, n_1179);
  nand g3474 (n_79, n_3175, n_3176, n_3177);
  xor g3481 (n_3182, A[60], A[64]);
  xor g3482 (n_1184, n_3182, A[62]);
  nand g3485 (n_3185, A[60], A[62]);
  nand g3486 (n_1192, n_2968, n_2904, n_3185);
  xor g3487 (n_3186, A[57], n_1181);
  xor g3488 (n_1186, n_3186, n_1161);
  nand g3489 (n_3187, A[57], n_1181);
  nand g3490 (n_3188, n_1161, n_1181);
  nand g3491 (n_3189, A[57], n_1161);
  nand g3492 (n_1195, n_3187, n_3188, n_3189);
  xor g3493 (n_3190, n_1183, n_1184);
  xor g3494 (n_1187, n_3190, n_1185);
  nand g3495 (n_3191, n_1183, n_1184);
  nand g3496 (n_3192, n_1185, n_1184);
  nand g3497 (n_3193, n_1183, n_1185);
  nand g3498 (n_1197, n_3191, n_3192, n_3193);
  xor g3499 (n_3194, n_1186, n_1187);
  xor g3500 (n_165, n_3194, n_1188);
  nand g3501 (n_3195, n_1186, n_1187);
  nand g3502 (n_3196, n_1188, n_1187);
  nand g3503 (n_3197, n_1186, n_1188);
  nand g3504 (n_164, n_3195, n_3196, n_3197);
  xor g3507 (n_3198, A[59], A[63]);
  xor g3508 (n_1193, n_3198, A[65]);
  nand g3511 (n_3201, A[59], A[65]);
  nand g3512 (n_1200, n_3161, n_2936, n_3201);
  xor g3514 (n_1194, n_3202, n_1171);
  nand g3517 (n_3205, A[61], n_1171);
  nand g3518 (n_1202, n_3164, n_3204, n_3205);
  xor g3519 (n_3206, n_1192, n_1193);
  xor g3520 (n_1196, n_3206, n_1194);
  nand g3521 (n_3207, n_1192, n_1193);
  nand g3522 (n_3208, n_1194, n_1193);
  nand g3523 (n_3209, n_1192, n_1194);
  nand g3524 (n_1204, n_3207, n_3208, n_3209);
  xor g3525 (n_3210, n_1195, n_1196);
  xor g3526 (n_78, n_3210, n_1197);
  nand g3527 (n_3211, n_1195, n_1196);
  nand g3528 (n_3212, n_1197, n_1196);
  nand g3529 (n_3213, n_1195, n_1197);
  nand g3530 (n_163, n_3211, n_3212, n_3213);
  xor g3532 (n_1199, n_3022, A[60]);
  nand g3534 (n_3216, A[60], A[58]);
  nand g3536 (n_1207, n_3023, n_3216, n_3217);
  xor g3538 (n_1201, n_3090, A[57]);
  nand g3540 (n_3220, A[57], A[62]);
  nand g3541 (n_3221, A[64], A[57]);
  nand g3542 (n_1208, n_2904, n_3220, n_3221);
  xor g3543 (n_3222, n_1199, n_1200);
  xor g3544 (n_1203, n_3222, n_1201);
  nand g3545 (n_3223, n_1199, n_1200);
  nand g3546 (n_3224, n_1201, n_1200);
  nand g3547 (n_3225, n_1199, n_1201);
  nand g3548 (n_1211, n_3223, n_3224, n_3225);
  xor g3549 (n_3226, n_1202, n_1203);
  xor g3550 (n_77, n_3226, n_1204);
  nand g3551 (n_3227, n_1202, n_1203);
  nand g3552 (n_3228, n_1204, n_1203);
  nand g3553 (n_3229, n_1202, n_1204);
  nand g3554 (n_76, n_3227, n_3228, n_3229);
  xor g3564 (n_1210, n_3234, n_1208);
  nand g3566 (n_3236, n_1208, n_1207);
  nand g3568 (n_1216, n_3235, n_3236, n_3237);
  xor g3569 (n_3238, n_1150, n_1210);
  xor g3570 (n_162, n_3238, n_1211);
  nand g3571 (n_3239, n_1150, n_1210);
  nand g3572 (n_3240, n_1211, n_1210);
  nand g3573 (n_3241, n_1150, n_1211);
  nand g3574 (n_75, n_3239, n_3240, n_3241);
  xor g3576 (n_1214, n_3242, A[60]);
  nand g3580 (n_1219, n_3243, n_2968, n_3217);
  xor g3582 (n_1215, n_3142, n_1160);
  nand g3584 (n_3248, n_1160, A[59]);
  nand g3585 (n_3249, A[62], n_1160);
  nand g3586 (n_1221, n_3092, n_3248, n_3249);
  xor g3587 (n_3250, n_1214, n_1215);
  xor g3588 (n_161, n_3250, n_1216);
  nand g3589 (n_3251, n_1214, n_1215);
  nand g3590 (n_3252, n_1216, n_1215);
  nand g3591 (n_3253, n_1214, n_1216);
  nand g3592 (n_160, n_3251, n_3252, n_3253);
  xor g3595 (n_3254, A[63], A[61]);
  nand g3600 (n_1224, n_3117, n_3256, n_3257);
  xor g3601 (n_3258, n_1219, n_1220);
  xor g3602 (n_74, n_3258, n_1221);
  nand g3603 (n_3259, n_1219, n_1220);
  nand g3604 (n_3260, n_1221, n_1220);
  nand g3605 (n_3261, n_1219, n_1221);
  nand g3606 (n_159, n_3259, n_3260, n_3261);
  xor g3608 (n_1223, n_3242, A[62]);
  nand g3612 (n_1227, n_3243, n_2904, n_3265);
  xor g3613 (n_3266, A[65], n_1223);
  xor g3614 (n_73, n_3266, n_1224);
  nand g3615 (n_3267, A[65], n_1223);
  nand g3616 (n_3268, n_1224, n_1223);
  nand g3617 (n_3269, A[65], n_1224);
  nand g3618 (n_158, n_3267, n_3268, n_3269);
  nand g3625 (n_3273, A[65], n_1227);
  nand g3626 (n_157, n_3271, n_3272, n_3273);
  xor g3628 (n_71, n_3242, A[63]);
  nand g3630 (n_3276, A[63], A[64]);
  nand g3632 (n_156, n_3243, n_3276, n_3277);
  nand g25 (n_3299, n_1232, n_3296, n_3297);
  nand g28 (n_3300, A[2], n_235);
  nand g29 (n_3301, A[2], n_3299);
  nand g30 (n_3302, n_235, n_3299);
  nand g31 (n_3304, n_3300, n_3301, n_3302);
  xor g33 (Z[4], n_3299, n_367);
  nand g34 (n_3305, n_148, n_234);
  nand g35 (n_3306, n_148, n_3304);
  nand g36 (n_3307, n_234, n_3304);
  nand g37 (n_3309, n_3305, n_3306, n_3307);
  xor g38 (n_3308, n_148, n_234);
  xor g39 (Z[5], n_3304, n_3308);
  nand g40 (n_3310, n_147, n_233);
  nand g41 (n_3311, n_147, n_3309);
  nand g42 (n_3312, n_233, n_3309);
  nand g43 (n_3314, n_3310, n_3311, n_3312);
  xor g44 (n_3313, n_147, n_233);
  xor g45 (Z[6], n_3309, n_3313);
  nand g46 (n_3315, n_146, n_232);
  nand g47 (n_3316, n_146, n_3314);
  nand g48 (n_3317, n_232, n_3314);
  nand g49 (n_3319, n_3315, n_3316, n_3317);
  xor g50 (n_3318, n_146, n_232);
  xor g51 (Z[7], n_3314, n_3318);
  nand g52 (n_3320, n_145, n_231);
  nand g53 (n_3321, n_145, n_3319);
  nand g54 (n_3322, n_231, n_3319);
  nand g55 (n_3324, n_3320, n_3321, n_3322);
  xor g56 (n_3323, n_145, n_231);
  xor g57 (Z[8], n_3319, n_3323);
  nand g58 (n_3325, n_144, n_230);
  nand g59 (n_3326, n_144, n_3324);
  nand g60 (n_3327, n_230, n_3324);
  nand g61 (n_3329, n_3325, n_3326, n_3327);
  xor g62 (n_3328, n_144, n_230);
  xor g63 (Z[9], n_3324, n_3328);
  nand g64 (n_3330, n_143, n_229);
  nand g65 (n_3331, n_143, n_3329);
  nand g66 (n_3332, n_229, n_3329);
  nand g67 (n_3334, n_3330, n_3331, n_3332);
  xor g68 (n_3333, n_143, n_229);
  xor g69 (Z[10], n_3329, n_3333);
  nand g70 (n_3335, n_142, n_228);
  nand g71 (n_3336, n_142, n_3334);
  nand g72 (n_3337, n_228, n_3334);
  nand g73 (n_3339, n_3335, n_3336, n_3337);
  xor g74 (n_3338, n_142, n_228);
  xor g75 (Z[11], n_3334, n_3338);
  nand g76 (n_3340, n_141, n_227);
  nand g77 (n_3341, n_141, n_3339);
  nand g78 (n_3342, n_227, n_3339);
  nand g79 (n_3344, n_3340, n_3341, n_3342);
  xor g80 (n_3343, n_141, n_227);
  xor g81 (Z[12], n_3339, n_3343);
  nand g82 (n_3345, n_140, n_226);
  nand g83 (n_3346, n_140, n_3344);
  nand g84 (n_3347, n_226, n_3344);
  nand g85 (n_3349, n_3345, n_3346, n_3347);
  xor g86 (n_3348, n_140, n_226);
  xor g87 (Z[13], n_3344, n_3348);
  nand g88 (n_3350, n_139, n_225);
  nand g89 (n_3351, n_139, n_3349);
  nand g90 (n_3352, n_225, n_3349);
  nand g91 (n_3354, n_3350, n_3351, n_3352);
  xor g92 (n_3353, n_139, n_225);
  xor g93 (Z[14], n_3349, n_3353);
  nand g94 (n_3355, n_138, n_224);
  nand g95 (n_3356, n_138, n_3354);
  nand g96 (n_3357, n_224, n_3354);
  nand g97 (n_3359, n_3355, n_3356, n_3357);
  xor g98 (n_3358, n_138, n_224);
  xor g99 (Z[15], n_3354, n_3358);
  nand g100 (n_3360, n_137, n_223);
  nand g101 (n_3361, n_137, n_3359);
  nand g102 (n_3362, n_223, n_3359);
  nand g103 (n_3364, n_3360, n_3361, n_3362);
  xor g104 (n_3363, n_137, n_223);
  xor g105 (Z[16], n_3359, n_3363);
  nand g106 (n_3365, n_136, n_222);
  nand g107 (n_3366, n_136, n_3364);
  nand g108 (n_3367, n_222, n_3364);
  nand g109 (n_3369, n_3365, n_3366, n_3367);
  xor g110 (n_3368, n_136, n_222);
  xor g111 (Z[17], n_3364, n_3368);
  nand g112 (n_3370, n_135, n_221);
  nand g113 (n_3371, n_135, n_3369);
  nand g114 (n_3372, n_221, n_3369);
  nand g115 (n_3374, n_3370, n_3371, n_3372);
  xor g116 (n_3373, n_135, n_221);
  xor g117 (Z[18], n_3369, n_3373);
  nand g118 (n_3375, n_134, n_220);
  nand g119 (n_3376, n_134, n_3374);
  nand g120 (n_3377, n_220, n_3374);
  nand g121 (n_3379, n_3375, n_3376, n_3377);
  xor g122 (n_3378, n_134, n_220);
  xor g123 (Z[19], n_3374, n_3378);
  nand g124 (n_3380, n_133, n_219);
  nand g125 (n_3381, n_133, n_3379);
  nand g126 (n_3382, n_219, n_3379);
  nand g127 (n_3384, n_3380, n_3381, n_3382);
  xor g128 (n_3383, n_133, n_219);
  xor g129 (Z[20], n_3379, n_3383);
  nand g130 (n_3385, n_132, n_218);
  nand g131 (n_3386, n_132, n_3384);
  nand g132 (n_3387, n_218, n_3384);
  nand g133 (n_3389, n_3385, n_3386, n_3387);
  xor g134 (n_3388, n_132, n_218);
  xor g135 (Z[21], n_3384, n_3388);
  nand g136 (n_3390, n_131, n_217);
  nand g137 (n_3391, n_131, n_3389);
  nand g138 (n_3392, n_217, n_3389);
  nand g139 (n_3394, n_3390, n_3391, n_3392);
  xor g140 (n_3393, n_131, n_217);
  xor g141 (Z[22], n_3389, n_3393);
  nand g142 (n_3395, n_130, n_216);
  nand g143 (n_3396, n_130, n_3394);
  nand g144 (n_3397, n_216, n_3394);
  nand g145 (n_3399, n_3395, n_3396, n_3397);
  xor g146 (n_3398, n_130, n_216);
  xor g147 (Z[23], n_3394, n_3398);
  nand g148 (n_3400, n_129, n_215);
  nand g149 (n_3401, n_129, n_3399);
  nand g150 (n_3402, n_215, n_3399);
  nand g151 (n_3404, n_3400, n_3401, n_3402);
  xor g152 (n_3403, n_129, n_215);
  xor g153 (Z[24], n_3399, n_3403);
  nand g154 (n_3405, n_128, n_214);
  nand g155 (n_3406, n_128, n_3404);
  nand g156 (n_3407, n_214, n_3404);
  nand g157 (n_3409, n_3405, n_3406, n_3407);
  xor g158 (n_3408, n_128, n_214);
  xor g159 (Z[25], n_3404, n_3408);
  nand g160 (n_3410, n_127, n_213);
  nand g161 (n_3411, n_127, n_3409);
  nand g162 (n_3412, n_213, n_3409);
  nand g163 (n_3414, n_3410, n_3411, n_3412);
  xor g164 (n_3413, n_127, n_213);
  xor g165 (Z[26], n_3409, n_3413);
  nand g166 (n_3415, n_126, n_212);
  nand g167 (n_3416, n_126, n_3414);
  nand g168 (n_3417, n_212, n_3414);
  nand g169 (n_3419, n_3415, n_3416, n_3417);
  xor g170 (n_3418, n_126, n_212);
  xor g171 (Z[27], n_3414, n_3418);
  nand g172 (n_3420, n_125, n_211);
  nand g173 (n_3421, n_125, n_3419);
  nand g174 (n_3422, n_211, n_3419);
  nand g175 (n_3424, n_3420, n_3421, n_3422);
  xor g176 (n_3423, n_125, n_211);
  xor g177 (Z[28], n_3419, n_3423);
  nand g178 (n_3425, n_124, n_210);
  nand g179 (n_3426, n_124, n_3424);
  nand g180 (n_3427, n_210, n_3424);
  nand g181 (n_3429, n_3425, n_3426, n_3427);
  xor g182 (n_3428, n_124, n_210);
  xor g183 (Z[29], n_3424, n_3428);
  nand g184 (n_3430, n_123, n_209);
  nand g185 (n_3431, n_123, n_3429);
  nand g186 (n_3432, n_209, n_3429);
  nand g187 (n_3434, n_3430, n_3431, n_3432);
  xor g188 (n_3433, n_123, n_209);
  xor g189 (Z[30], n_3429, n_3433);
  nand g190 (n_3435, n_122, n_208);
  nand g191 (n_3436, n_122, n_3434);
  nand g192 (n_3437, n_208, n_3434);
  nand g193 (n_3439, n_3435, n_3436, n_3437);
  xor g194 (n_3438, n_122, n_208);
  xor g195 (Z[31], n_3434, n_3438);
  nand g196 (n_3440, n_121, n_207);
  nand g197 (n_3441, n_121, n_3439);
  nand g198 (n_3442, n_207, n_3439);
  nand g199 (n_3444, n_3440, n_3441, n_3442);
  xor g200 (n_3443, n_121, n_207);
  xor g201 (Z[32], n_3439, n_3443);
  nand g202 (n_3445, n_120, n_206);
  nand g203 (n_3446, n_120, n_3444);
  nand g204 (n_3447, n_206, n_3444);
  nand g205 (n_3449, n_3445, n_3446, n_3447);
  xor g206 (n_3448, n_120, n_206);
  xor g207 (Z[33], n_3444, n_3448);
  nand g208 (n_3450, n_119, n_205);
  nand g209 (n_3451, n_119, n_3449);
  nand g210 (n_3452, n_205, n_3449);
  nand g211 (n_3454, n_3450, n_3451, n_3452);
  xor g212 (n_3453, n_119, n_205);
  xor g213 (Z[34], n_3449, n_3453);
  nand g214 (n_3455, n_118, n_204);
  nand g215 (n_3456, n_118, n_3454);
  nand g216 (n_3457, n_204, n_3454);
  nand g217 (n_3459, n_3455, n_3456, n_3457);
  xor g218 (n_3458, n_118, n_204);
  xor g219 (Z[35], n_3454, n_3458);
  nand g220 (n_3460, n_117, n_203);
  nand g221 (n_3461, n_117, n_3459);
  nand g222 (n_3462, n_203, n_3459);
  nand g223 (n_3464, n_3460, n_3461, n_3462);
  xor g224 (n_3463, n_117, n_203);
  xor g225 (Z[36], n_3459, n_3463);
  nand g226 (n_3465, n_116, n_202);
  nand g227 (n_3466, n_116, n_3464);
  nand g228 (n_3467, n_202, n_3464);
  nand g229 (n_3469, n_3465, n_3466, n_3467);
  xor g230 (n_3468, n_116, n_202);
  xor g231 (Z[37], n_3464, n_3468);
  nand g232 (n_3470, n_115, n_201);
  nand g233 (n_3471, n_115, n_3469);
  nand g234 (n_3472, n_201, n_3469);
  nand g235 (n_3474, n_3470, n_3471, n_3472);
  xor g236 (n_3473, n_115, n_201);
  xor g237 (Z[38], n_3469, n_3473);
  nand g238 (n_3475, n_114, n_200);
  nand g239 (n_3476, n_114, n_3474);
  nand g240 (n_3477, n_200, n_3474);
  nand g241 (n_3479, n_3475, n_3476, n_3477);
  xor g242 (n_3478, n_114, n_200);
  xor g243 (Z[39], n_3474, n_3478);
  nand g244 (n_3480, n_113, n_199);
  nand g245 (n_3481, n_113, n_3479);
  nand g246 (n_3482, n_199, n_3479);
  nand g247 (n_3484, n_3480, n_3481, n_3482);
  xor g248 (n_3483, n_113, n_199);
  xor g249 (Z[40], n_3479, n_3483);
  nand g250 (n_3485, n_112, n_198);
  nand g251 (n_3486, n_112, n_3484);
  nand g252 (n_3487, n_198, n_3484);
  nand g253 (n_3489, n_3485, n_3486, n_3487);
  xor g254 (n_3488, n_112, n_198);
  xor g255 (Z[41], n_3484, n_3488);
  nand g256 (n_3490, n_111, n_197);
  nand g257 (n_3491, n_111, n_3489);
  nand g258 (n_3492, n_197, n_3489);
  nand g259 (n_3494, n_3490, n_3491, n_3492);
  xor g260 (n_3493, n_111, n_197);
  xor g261 (Z[42], n_3489, n_3493);
  nand g262 (n_3495, n_110, n_196);
  nand g263 (n_3496, n_110, n_3494);
  nand g264 (n_3497, n_196, n_3494);
  nand g265 (n_3499, n_3495, n_3496, n_3497);
  xor g266 (n_3498, n_110, n_196);
  xor g267 (Z[43], n_3494, n_3498);
  nand g268 (n_3500, n_109, n_195);
  nand g269 (n_3501, n_109, n_3499);
  nand g270 (n_3502, n_195, n_3499);
  nand g271 (n_3504, n_3500, n_3501, n_3502);
  xor g272 (n_3503, n_109, n_195);
  xor g273 (Z[44], n_3499, n_3503);
  nand g274 (n_3505, n_108, n_194);
  nand g275 (n_3506, n_108, n_3504);
  nand g276 (n_3507, n_194, n_3504);
  nand g277 (n_3509, n_3505, n_3506, n_3507);
  xor g278 (n_3508, n_108, n_194);
  xor g279 (Z[45], n_3504, n_3508);
  nand g280 (n_3510, n_107, n_193);
  nand g281 (n_3511, n_107, n_3509);
  nand g282 (n_3512, n_193, n_3509);
  nand g283 (n_3514, n_3510, n_3511, n_3512);
  xor g284 (n_3513, n_107, n_193);
  xor g285 (Z[46], n_3509, n_3513);
  nand g286 (n_3515, n_106, n_192);
  nand g287 (n_3516, n_106, n_3514);
  nand g288 (n_3517, n_192, n_3514);
  nand g289 (n_3519, n_3515, n_3516, n_3517);
  xor g290 (n_3518, n_106, n_192);
  xor g291 (Z[47], n_3514, n_3518);
  nand g292 (n_3520, n_105, n_191);
  nand g293 (n_3521, n_105, n_3519);
  nand g294 (n_3522, n_191, n_3519);
  nand g295 (n_3524, n_3520, n_3521, n_3522);
  xor g296 (n_3523, n_105, n_191);
  xor g297 (Z[48], n_3519, n_3523);
  nand g298 (n_3525, n_104, n_190);
  nand g299 (n_3526, n_104, n_3524);
  nand g300 (n_3527, n_190, n_3524);
  nand g301 (n_3529, n_3525, n_3526, n_3527);
  xor g302 (n_3528, n_104, n_190);
  xor g303 (Z[49], n_3524, n_3528);
  nand g304 (n_3530, n_103, n_189);
  nand g305 (n_3531, n_103, n_3529);
  nand g306 (n_3532, n_189, n_3529);
  nand g307 (n_3534, n_3530, n_3531, n_3532);
  xor g308 (n_3533, n_103, n_189);
  xor g309 (Z[50], n_3529, n_3533);
  nand g310 (n_3535, n_102, n_188);
  nand g311 (n_3536, n_102, n_3534);
  nand g312 (n_3537, n_188, n_3534);
  nand g313 (n_3539, n_3535, n_3536, n_3537);
  xor g314 (n_3538, n_102, n_188);
  xor g315 (Z[51], n_3534, n_3538);
  nand g316 (n_3540, n_101, n_187);
  nand g317 (n_3541, n_101, n_3539);
  nand g318 (n_3542, n_187, n_3539);
  nand g319 (n_3544, n_3540, n_3541, n_3542);
  xor g320 (n_3543, n_101, n_187);
  xor g321 (Z[52], n_3539, n_3543);
  nand g322 (n_3545, n_100, n_186);
  nand g323 (n_3546, n_100, n_3544);
  nand g324 (n_3547, n_186, n_3544);
  nand g325 (n_3549, n_3545, n_3546, n_3547);
  xor g326 (n_3548, n_100, n_186);
  xor g327 (Z[53], n_3544, n_3548);
  nand g328 (n_3550, n_99, n_185);
  nand g329 (n_3551, n_99, n_3549);
  nand g330 (n_3552, n_185, n_3549);
  nand g331 (n_3554, n_3550, n_3551, n_3552);
  xor g332 (n_3553, n_99, n_185);
  xor g333 (Z[54], n_3549, n_3553);
  nand g334 (n_3555, n_98, n_184);
  nand g335 (n_3556, n_98, n_3554);
  nand g336 (n_3557, n_184, n_3554);
  nand g337 (n_3559, n_3555, n_3556, n_3557);
  xor g338 (n_3558, n_98, n_184);
  xor g339 (Z[55], n_3554, n_3558);
  nand g340 (n_3560, n_97, n_183);
  nand g341 (n_3561, n_97, n_3559);
  nand g342 (n_3562, n_183, n_3559);
  nand g343 (n_3564, n_3560, n_3561, n_3562);
  xor g344 (n_3563, n_97, n_183);
  xor g345 (Z[56], n_3559, n_3563);
  nand g346 (n_3565, n_96, n_182);
  nand g347 (n_3566, n_96, n_3564);
  nand g348 (n_3567, n_182, n_3564);
  nand g349 (n_3569, n_3565, n_3566, n_3567);
  xor g350 (n_3568, n_96, n_182);
  xor g351 (Z[57], n_3564, n_3568);
  nand g352 (n_3570, n_95, n_181);
  nand g353 (n_3571, n_95, n_3569);
  nand g354 (n_3572, n_181, n_3569);
  nand g355 (n_3574, n_3570, n_3571, n_3572);
  xor g356 (n_3573, n_95, n_181);
  xor g357 (Z[58], n_3569, n_3573);
  nand g358 (n_3575, n_94, n_180);
  nand g359 (n_3576, n_94, n_3574);
  nand g360 (n_3577, n_180, n_3574);
  nand g361 (n_3579, n_3575, n_3576, n_3577);
  xor g362 (n_3578, n_94, n_180);
  xor g363 (Z[59], n_3574, n_3578);
  nand g364 (n_3580, n_93, n_179);
  nand g365 (n_3581, n_93, n_3579);
  nand g366 (n_3582, n_179, n_3579);
  nand g367 (n_3584, n_3580, n_3581, n_3582);
  xor g368 (n_3583, n_93, n_179);
  xor g369 (Z[60], n_3579, n_3583);
  nand g370 (n_3585, n_92, n_178);
  nand g371 (n_3586, n_92, n_3584);
  nand g372 (n_3587, n_178, n_3584);
  nand g373 (n_3589, n_3585, n_3586, n_3587);
  xor g374 (n_3588, n_92, n_178);
  xor g375 (Z[61], n_3584, n_3588);
  nand g376 (n_3590, n_91, n_177);
  nand g377 (n_3591, n_91, n_3589);
  nand g378 (n_3592, n_177, n_3589);
  nand g379 (n_3594, n_3590, n_3591, n_3592);
  xor g380 (n_3593, n_91, n_177);
  xor g381 (Z[62], n_3589, n_3593);
  nand g382 (n_3595, n_90, n_176);
  nand g383 (n_3596, n_90, n_3594);
  nand g384 (n_3597, n_176, n_3594);
  nand g385 (n_3599, n_3595, n_3596, n_3597);
  xor g386 (n_3598, n_90, n_176);
  xor g387 (Z[63], n_3594, n_3598);
  nand g388 (n_3600, n_89, n_175);
  nand g389 (n_3601, n_89, n_3599);
  nand g390 (n_3602, n_175, n_3599);
  nand g391 (n_3604, n_3600, n_3601, n_3602);
  xor g392 (n_3603, n_89, n_175);
  xor g393 (Z[64], n_3599, n_3603);
  nand g394 (n_3605, n_88, n_174);
  nand g395 (n_3606, n_88, n_3604);
  nand g396 (n_3607, n_174, n_3604);
  nand g397 (n_3609, n_3605, n_3606, n_3607);
  xor g398 (n_3608, n_88, n_174);
  xor g399 (Z[65], n_3604, n_3608);
  nand g400 (n_3610, n_87, n_173);
  nand g401 (n_3611, n_87, n_3609);
  nand g402 (n_3612, n_173, n_3609);
  nand g403 (n_3614, n_3610, n_3611, n_3612);
  xor g404 (n_3613, n_87, n_173);
  xor g405 (Z[66], n_3609, n_3613);
  nand g406 (n_3615, n_86, n_172);
  nand g407 (n_3616, n_86, n_3614);
  nand g408 (n_3617, n_172, n_3614);
  nand g409 (n_3619, n_3615, n_3616, n_3617);
  xor g410 (n_3618, n_86, n_172);
  xor g411 (Z[67], n_3614, n_3618);
  nand g412 (n_3620, n_85, n_171);
  nand g413 (n_3621, n_85, n_3619);
  nand g414 (n_3622, n_171, n_3619);
  nand g415 (n_3624, n_3620, n_3621, n_3622);
  xor g416 (n_3623, n_85, n_171);
  xor g417 (Z[68], n_3619, n_3623);
  nand g418 (n_3625, n_84, n_170);
  nand g419 (n_3626, n_84, n_3624);
  nand g420 (n_3627, n_170, n_3624);
  nand g421 (n_3629, n_3625, n_3626, n_3627);
  xor g422 (n_3628, n_84, n_170);
  xor g423 (Z[69], n_3624, n_3628);
  nand g424 (n_3630, n_83, n_169);
  nand g425 (n_3631, n_83, n_3629);
  nand g426 (n_3632, n_169, n_3629);
  nand g427 (n_3634, n_3630, n_3631, n_3632);
  xor g428 (n_3633, n_83, n_169);
  xor g429 (Z[70], n_3629, n_3633);
  nand g430 (n_3635, n_82, n_168);
  nand g431 (n_3636, n_82, n_3634);
  nand g432 (n_3637, n_168, n_3634);
  nand g433 (n_3639, n_3635, n_3636, n_3637);
  xor g434 (n_3638, n_82, n_168);
  xor g435 (Z[71], n_3634, n_3638);
  nand g436 (n_3640, n_81, n_167);
  nand g437 (n_3641, n_81, n_3639);
  nand g438 (n_3642, n_167, n_3639);
  nand g439 (n_3644, n_3640, n_3641, n_3642);
  xor g440 (n_3643, n_81, n_167);
  xor g441 (Z[72], n_3639, n_3643);
  nand g442 (n_3645, n_80, n_166);
  nand g443 (n_3646, n_80, n_3644);
  nand g444 (n_3647, n_166, n_3644);
  nand g445 (n_3649, n_3645, n_3646, n_3647);
  xor g446 (n_3648, n_80, n_166);
  xor g447 (Z[73], n_3644, n_3648);
  nand g448 (n_3650, n_79, n_165);
  nand g449 (n_3651, n_79, n_3649);
  nand g450 (n_3652, n_165, n_3649);
  nand g451 (n_3654, n_3650, n_3651, n_3652);
  xor g452 (n_3653, n_79, n_165);
  xor g453 (Z[74], n_3649, n_3653);
  nand g454 (n_3655, n_78, n_164);
  nand g455 (n_3656, n_78, n_3654);
  nand g456 (n_3657, n_164, n_3654);
  nand g457 (n_3659, n_3655, n_3656, n_3657);
  xor g458 (n_3658, n_78, n_164);
  xor g459 (Z[75], n_3654, n_3658);
  nand g460 (n_3660, n_77, n_163);
  nand g461 (n_3661, n_77, n_3659);
  nand g462 (n_3662, n_163, n_3659);
  nand g463 (n_3664, n_3660, n_3661, n_3662);
  xor g464 (n_3663, n_77, n_163);
  xor g465 (Z[76], n_3659, n_3663);
  nand g466 (n_3665, n_76, n_162);
  nand g467 (n_3666, n_76, n_3664);
  nand g468 (n_3667, n_162, n_3664);
  nand g469 (n_3669, n_3665, n_3666, n_3667);
  xor g470 (n_3668, n_76, n_162);
  xor g471 (Z[77], n_3664, n_3668);
  nand g472 (n_3670, n_75, n_161);
  nand g473 (n_3671, n_75, n_3669);
  nand g474 (n_3672, n_161, n_3669);
  nand g475 (n_3674, n_3670, n_3671, n_3672);
  xor g476 (n_3673, n_75, n_161);
  xor g477 (Z[78], n_3669, n_3673);
  nand g478 (n_3675, n_74, n_160);
  nand g479 (n_3676, n_74, n_3674);
  nand g480 (n_3677, n_160, n_3674);
  nand g481 (n_3679, n_3675, n_3676, n_3677);
  xor g482 (n_3678, n_74, n_160);
  xor g483 (Z[79], n_3674, n_3678);
  nand g484 (n_3680, n_73, n_159);
  nand g485 (n_3681, n_73, n_3679);
  nand g486 (n_3682, n_159, n_3679);
  nand g487 (n_3684, n_3680, n_3681, n_3682);
  xor g488 (n_3683, n_73, n_159);
  xor g489 (Z[80], n_3679, n_3683);
  nand g490 (n_3685, n_72, n_158);
  nand g491 (n_3686, n_72, n_3684);
  nand g492 (n_3687, n_158, n_3684);
  nand g493 (n_3689, n_3685, n_3686, n_3687);
  xor g494 (n_3688, n_72, n_158);
  xor g495 (Z[81], n_3684, n_3688);
  nand g496 (n_3690, n_71, n_157);
  nand g497 (n_3691, n_71, n_3689);
  nand g498 (n_3692, n_157, n_3689);
  nand g499 (n_3694, n_3690, n_3691, n_3692);
  xor g500 (n_3693, n_71, n_157);
  xor g501 (Z[82], n_3689, n_3693);
  nand g504 (n_3697, n_156, n_3694);
  nand g505 (n_3699, n_3695, n_3696, n_3697);
  xor g507 (Z[83], n_3694, n_3698);
  nand g510 (n_3702, A[65], n_3699);
  nand g511 (n_3704, n_3700, n_3701, n_3702);
  xor g513 (Z[84], n_3699, n_3703);
  or g3652 (n_335, wc, wc0, n_148);
  not gc0 (wc0, n_1235);
  not gc (wc, n_1247);
  or g3653 (n_344, wc1, wc2, n_328);
  not gc2 (wc2, n_1247);
  not gc1 (wc1, n_1268);
  or g3654 (n_356, wc3, n_333, n_328);
  not gc3 (wc3, n_1296);
  or g3655 (n_373, wc4, n_342, n_333);
  not gc4 (wc4, n_1332);
  or g3656 (n_394, wc5, n_355, n_342);
  not gc5 (wc5, n_1376);
  or g3657 (n_419, wc6, wc7, n_355);
  not gc7 (wc7, n_1427);
  not gc6 (wc6, n_1428);
  or g3658 (n_420, wc8, wc9, n_333);
  not gc9 (wc9, n_1431);
  not gc8 (wc8, n_1433);
  or g3659 (n_448, wc10, wc11, n_328);
  not gc11 (wc11, n_1427);
  not gc10 (wc10, n_1493);
  or g3660 (n_447, wc12, wc13, n_342);
  not gc13 (wc13, n_1495);
  not gc12 (wc12, n_1497);
  or g3661 (n_526, wc14, wc15, n_355);
  not gc15 (wc15, n_1560);
  not gc14 (wc14, n_1684);
  or g3662 (n_552, wc16, wc17, n_372);
  not gc17 (wc17, n_1489);
  not gc16 (wc16, n_1748);
  or g3663 (n_580, wc18, wc19, n_393);
  not gc19 (wc19, n_1553);
  not gc18 (wc18, n_1812);
  or g3664 (n_608, wc20, wc21, n_418);
  not gc21 (wc21, n_1617);
  not gc20 (wc20, n_1876);
  xnor g3665 (n_3022, A[66], A[58]);
  or g3666 (n_3023, wc22, A[66]);
  not gc22 (wc22, A[58]);
  or g3667 (n_3025, wc23, A[66]);
  not gc23 (wc23, A[52]);
  xnor g3668 (n_3062, A[61], A[59]);
  or g3669 (n_3063, A[59], wc24);
  not gc24 (wc24, A[61]);
  or g3670 (n_3028, wc25, A[66]);
  not gc25 (wc25, A[56]);
  xnor g3671 (n_1174, n_3162, A[57]);
  or g3672 (n_3164, A[57], wc26);
  not gc26 (wc26, A[61]);
  or g3673 (n_3165, A[57], wc27);
  not gc27 (wc27, A[65]);
  xnor g3674 (n_3202, A[61], A[57]);
  or g3675 (n_3217, wc28, A[66]);
  not gc28 (wc28, A[60]);
  xnor g3676 (n_3242, A[66], A[64]);
  or g3677 (n_3243, wc29, A[66]);
  not gc29 (wc29, A[64]);
  xnor g3678 (n_1220, n_3254, A[65]);
  or g3679 (n_3256, wc30, A[65]);
  not gc30 (wc30, A[61]);
  or g3680 (n_3257, wc31, A[65]);
  not gc31 (wc31, A[63]);
  or g3681 (n_3265, wc32, A[66]);
  not gc32 (wc32, A[62]);
  or g3683 (n_3271, A[63], wc33);
  not gc33 (wc33, A[65]);
  or g3684 (n_3277, wc34, A[66]);
  not gc34 (wc34, A[63]);
  or g3685 (n_3700, wc35, A[66]);
  not gc35 (wc35, A[65]);
  xnor g3686 (n_3703, A[66], A[65]);
  or g3687 (n_3121, A[59], wc36);
  not gc36 (wc36, n_1148);
  xnor g3688 (n_3026, A[66], A[50]);
  or g3689 (n_3027, wc37, A[66]);
  not gc37 (wc37, A[50]);
  or g3690 (n_3064, A[59], wc38);
  not gc38 (wc38, n_1119);
  xnor g3691 (n_3118, n_1119, A[59]);
  or g3692 (n_3204, A[57], wc39);
  not gc39 (wc39, n_1171);
  xnor g3693 (n_3234, n_1207, A[59]);
  or g3694 (n_3235, A[59], wc40);
  not gc40 (wc40, n_1207);
  or g3695 (n_3237, A[59], wc41);
  not gc41 (wc41, n_1208);
  xnor g3696 (n_72, n_3114, n_1227);
  or g3697 (n_3272, A[63], wc42);
  not gc42 (wc42, n_1227);
  or g3698 (n_3695, A[65], wc43);
  not gc43 (wc43, n_156);
  xnor g3699 (n_3698, n_156, A[65]);
  or g3701 (n_3296, wc44, n_1235);
  not gc44 (wc44, A[3]);
  or g3702 (n_3297, wc45, n_1235);
  not gc45 (wc45, A[1]);
  xnor g3703 (Z[3], n_1235, n_1258);
  or g3704 (n_3696, A[65], wc46);
  not gc46 (wc46, n_3694);
  or g3705 (n_3701, A[66], wc47);
  not gc47 (wc47, n_3699);
  not g3706 (Z[85], n_3704);
endmodule

module mult_signed_const_16824_GENERIC(A, Z);
  input [66:0] A;
  output [85:0] Z;
  wire [66:0] A;
  wire [85:0] Z;
  mult_signed_const_16824_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_9979_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 349525;"
  input [44:0] A;
  output [63:0] Z;
  wire [44:0] A;
  wire [63:0] Z;
  wire n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72;
  wire n_73, n_74, n_75, n_76, n_77, n_78, n_79, n_80;
  wire n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88;
  wire n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96;
  wire n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104;
  wire n_105, n_106, n_107, n_108, n_109, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_239, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253;
  wire n_254, n_255, n_256, n_257, n_258, n_259, n_260, n_261;
  wire n_262, n_263, n_264, n_265, n_266, n_267, n_268, n_269;
  wire n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285;
  wire n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398;
  wire n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406;
  wire n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414;
  wire n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422;
  wire n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430;
  wire n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502;
  wire n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510;
  wire n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518;
  wire n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526;
  wire n_527, n_528, n_529, n_530, n_531, n_532, n_533, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550;
  wire n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558;
  wire n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566;
  wire n_567, n_568, n_569, n_570, n_571, n_572, n_573, n_574;
  wire n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582;
  wire n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590;
  wire n_591, n_592, n_593, n_594, n_595, n_596, n_597, n_598;
  wire n_599, n_600, n_601, n_602, n_603, n_604, n_605, n_606;
  wire n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614;
  wire n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_622;
  wire n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630;
  wire n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638;
  wire n_639, n_640, n_641, n_642, n_643, n_644, n_645, n_646;
  wire n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654;
  wire n_655, n_656, n_657, n_658, n_659, n_660, n_661, n_662;
  wire n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670;
  wire n_671, n_672, n_675, n_676, n_677, n_678, n_679, n_680;
  wire n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688;
  wire n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699;
  wire n_700, n_701, n_702, n_703, n_704, n_705, n_707, n_708;
  wire n_709, n_710, n_711, n_712, n_713, n_714, n_715, n_716;
  wire n_717, n_718, n_719, n_720, n_723, n_724, n_725, n_726;
  wire n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734;
  wire n_735, n_737, n_738, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_752, n_754, n_755, n_756;
  wire n_757, n_758, n_759, n_760, n_761, n_763, n_767, n_768;
  wire n_769, n_770, n_771, n_772, n_777, n_778, n_779, n_780;
  wire n_781, n_782, n_783, n_785, n_788, n_789, n_790, n_791;
  wire n_792, n_798, n_799, n_800, n_801, n_805, n_806, n_807;
  wire n_808, n_812, n_813, n_814, n_815, n_817, n_819, n_820;
  wire n_824, n_825, n_827, n_828, n_831, n_834, n_835, n_836;
  wire n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844;
  wire n_846, n_847, n_848, n_849, n_853, n_854, n_855, n_856;
  wire n_857, n_858, n_859, n_860, n_862, n_864, n_865, n_866;
  wire n_867, n_868, n_869, n_870, n_872, n_874, n_875, n_876;
  wire n_877, n_878, n_879, n_880, n_881, n_884, n_886, n_887;
  wire n_888, n_889, n_890, n_891, n_892, n_893, n_894, n_895;
  wire n_896, n_897, n_900, n_904, n_905, n_906, n_907, n_908;
  wire n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_918;
  wire n_919, n_920, n_922, n_923, n_924, n_925, n_926, n_927;
  wire n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935;
  wire n_936, n_938, n_939, n_941, n_942, n_943, n_944, n_945;
  wire n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953;
  wire n_954, n_955, n_956, n_957, n_958, n_959, n_961, n_962;
  wire n_964, n_965, n_966, n_967, n_968, n_969, n_970, n_971;
  wire n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_981;
  wire n_982, n_983, n_984, n_986, n_987, n_988, n_989, n_990;
  wire n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998;
  wire n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1010, n_1011;
  wire n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021;
  wire n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029;
  wire n_1030, n_1031, n_1033, n_1034, n_1036, n_1037, n_1040, n_1041;
  wire n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049;
  wire n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057;
  wire n_1058, n_1059, n_1060, n_1064, n_1065, n_1066, n_1067, n_1068;
  wire n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077;
  wire n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085;
  wire n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093;
  wire n_1098, n_1099, n_1100, n_1102, n_1103, n_1104, n_1105, n_1106;
  wire n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114;
  wire n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122;
  wire n_1123, n_1124, n_1125, n_1130, n_1132, n_1134, n_1135, n_1136;
  wire n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144;
  wire n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152;
  wire n_1153, n_1154, n_1155, n_1156, n_1157, n_1160, n_1161, n_1162;
  wire n_1163, n_1164, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171;
  wire n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179;
  wire n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187;
  wire n_1188, n_1189, n_1192, n_1194, n_1195, n_1198, n_1199, n_1200;
  wire n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208;
  wire n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216;
  wire n_1217, n_1218, n_1219, n_1220, n_1221, n_1224, n_1226, n_1227;
  wire n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237;
  wire n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
  wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253;
  wire n_1254, n_1256, n_1258, n_1259, n_1262, n_1263, n_1264, n_1265;
  wire n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273;
  wire n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281;
  wire n_1282, n_1283, n_1284, n_1285, n_1288, n_1290, n_1291, n_1294;
  wire n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302;
  wire n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310;
  wire n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318;
  wire n_1319, n_1320, n_1322, n_1323, n_1326, n_1327, n_1328, n_1329;
  wire n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337;
  wire n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345;
  wire n_1346, n_1347, n_1348, n_1349, n_1352, n_1354, n_1355, n_1358;
  wire n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366;
  wire n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374;
  wire n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382;
  wire n_1384, n_1386, n_1387, n_1390, n_1391, n_1392, n_1393, n_1394;
  wire n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402;
  wire n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410;
  wire n_1411, n_1412, n_1413, n_1416, n_1418, n_1419, n_1422, n_1423;
  wire n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431;
  wire n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439;
  wire n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1448;
  wire n_1450, n_1451, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467;
  wire n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475;
  wire n_1476, n_1477, n_1480, n_1482, n_1483, n_1486, n_1487, n_1488;
  wire n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496;
  wire n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504;
  wire n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512;
  wire n_1514, n_1515, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523;
  wire n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531;
  wire n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539;
  wire n_1540, n_1541, n_1544, n_1546, n_1547, n_1550, n_1551, n_1552;
  wire n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560;
  wire n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568;
  wire n_1569, n_1570, n_1571, n_1572, n_1573, n_1576, n_1578, n_1579;
  wire n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589;
  wire n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597;
  wire n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605;
  wire n_1608, n_1610, n_1611, n_1614, n_1615, n_1616, n_1617, n_1618;
  wire n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626;
  wire n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634;
  wire n_1635, n_1636, n_1637, n_1640, n_1642, n_1643, n_1646, n_1647;
  wire n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655;
  wire n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663;
  wire n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1672, n_1674;
  wire n_1675, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684;
  wire n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692;
  wire n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700;
  wire n_1701, n_1704, n_1706, n_1707, n_1710, n_1711, n_1712, n_1713;
  wire n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721;
  wire n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729;
  wire n_1730, n_1731, n_1732, n_1733, n_1736, n_1738, n_1739, n_1742;
  wire n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750;
  wire n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758;
  wire n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1768;
  wire n_1770, n_1771, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779;
  wire n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787;
  wire n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795;
  wire n_1796, n_1797, n_1800, n_1802, n_1803, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1832, n_1834, n_1835;
  wire n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845;
  wire n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853;
  wire n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861;
  wire n_1862, n_1863, n_1864, n_1866, n_1870, n_1871, n_1872, n_1873;
  wire n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881;
  wire n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889;
  wire n_1890, n_1891, n_1893, n_1894, n_1895, n_1898, n_1901, n_1902;
  wire n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910;
  wire n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918;
  wire n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1928;
  wire n_1930, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939;
  wire n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947;
  wire n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955;
  wire n_1958, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968;
  wire n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976;
  wire n_1977, n_1978, n_1979, n_1980, n_1981, n_1986, n_1989, n_1992;
  wire n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000;
  wire n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008;
  wire n_2009, n_2010, n_2018, n_2020, n_2021, n_2022, n_2023, n_2024;
  wire n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032;
  wire n_2033, n_2042, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049;
  wire n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057;
  wire n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071;
  wire n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2086, n_2087;
  wire n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095;
  wire n_2096, n_2097, n_2104, n_2105, n_2106, n_2108, n_2109, n_2110;
  wire n_2111, n_2112, n_2113, n_2120, n_2121, n_2122, n_2123, n_2124;
  wire n_2125, n_2126, n_2127, n_2128, n_2129, n_2136, n_2137, n_2138;
  wire n_2139, n_2140, n_2141, n_2146, n_2147, n_2148, n_2149, n_2150;
  wire n_2151, n_2152, n_2153, n_2156, n_2157, n_2158, n_2159, n_2160;
  wire n_2161, n_2165, n_2166, n_2167, n_2168, n_2169, n_2171, n_2172;
  wire n_2173, n_2176, n_2177, n_2189, n_2191, n_2193, n_2194, n_2195;
  wire n_2196, n_2197, n_2199, n_2200, n_2201, n_2202, n_2203, n_2205;
  wire n_2206, n_2207, n_2208, n_2209, n_2211, n_2212, n_2213, n_2214;
  wire n_2215, n_2217, n_2218, n_2219, n_2220, n_2221, n_2223, n_2224;
  wire n_2225, n_2226, n_2227, n_2229, n_2230, n_2231, n_2232, n_2233;
  wire n_2235, n_2236, n_2237, n_2238, n_2239, n_2241, n_2242, n_2243;
  wire n_2244, n_2245, n_2247, n_2248, n_2249, n_2250, n_2251, n_2253;
  wire n_2254, n_2255, n_2256, n_2257, n_2259, n_2260, n_2261, n_2262;
  wire n_2263, n_2265, n_2266, n_2267, n_2268, n_2269, n_2271, n_2272;
  wire n_2273, n_2274, n_2275, n_2277, n_2278, n_2279, n_2280, n_2281;
  wire n_2283, n_2284, n_2285, n_2286, n_2287, n_2289, n_2290, n_2291;
  wire n_2292, n_2293, n_2295, n_2296, n_2297, n_2298, n_2299, n_2301;
  wire n_2302, n_2303, n_2304, n_2305, n_2307, n_2308, n_2309, n_2310;
  wire n_2311, n_2313, n_2314, n_2315, n_2316, n_2317, n_2319, n_2320;
  wire n_2321, n_2322, n_2323, n_2325, n_2326, n_2327, n_2328, n_2329;
  wire n_2331, n_2332, n_2333, n_2334, n_2335, n_2337, n_2338, n_2339;
  wire n_2340, n_2341, n_2343, n_2344, n_2345, n_2346, n_2347, n_2349;
  wire n_2350, n_2351, n_2352, n_2353, n_2355, n_2356, n_2357, n_2358;
  wire n_2359, n_2361, n_2362, n_2363, n_2364, n_2365, n_2367, n_2368;
  wire n_2371, n_2376, n_2378, n_2379, n_2381, n_2383, n_2385, n_2386;
  wire n_2388, n_2389, n_2391, n_2393, n_2395, n_2396, n_2398, n_2399;
  wire n_2401, n_2403, n_2405, n_2406, n_2408, n_2409, n_2411, n_2413;
  wire n_2415, n_2416, n_2418, n_2419, n_2421, n_2423, n_2425, n_2426;
  wire n_2428, n_2429, n_2431, n_2433, n_2435, n_2436, n_2438, n_2439;
  wire n_2441, n_2443, n_2445, n_2446, n_2448, n_2449, n_2451, n_2453;
  wire n_2455, n_2456, n_2458, n_2459, n_2461, n_2463, n_2465, n_2466;
  wire n_2468, n_2469, n_2471, n_2473, n_2475, n_2476, n_2478, n_2479;
  wire n_2481, n_2483, n_2485, n_2486, n_2488, n_2489, n_2491, n_2493;
  wire n_2495, n_2496, n_2498, n_2499, n_2501, n_2503, n_2505, n_2506;
  wire n_2508, n_2509, n_2511, n_2513, n_2515, n_2516, n_2518, n_2519;
  wire n_2521, n_2525, n_2526, n_2527, n_2529, n_2530, n_2531, n_2533;
  wire n_2534, n_2535, n_2536, n_2538, n_2540, n_2542, n_2543, n_2544;
  wire n_2546, n_2547, n_2548, n_2550, n_2551, n_2553, n_2555, n_2557;
  wire n_2558, n_2559, n_2561, n_2562, n_2563, n_2565, n_2566, n_2568;
  wire n_2570, n_2572, n_2573, n_2574, n_2576, n_2577, n_2578, n_2580;
  wire n_2581, n_2583, n_2585, n_2587, n_2588, n_2589, n_2591, n_2592;
  wire n_2593, n_2595, n_2596, n_2598, n_2600, n_2602, n_2603, n_2604;
  wire n_2606, n_2607, n_2608, n_2610, n_2611, n_2613, n_2615, n_2617;
  wire n_2618, n_2619, n_2621, n_2622, n_2623, n_2625, n_2626, n_2628;
  wire n_2630, n_2632, n_2633, n_2634, n_2636, n_2638, n_2639, n_2640;
  wire n_2642, n_2643, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650;
  wire n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658;
  wire n_2659, n_2661, n_2664, n_2666, n_2667, n_2668, n_2671, n_2674;
  wire n_2676, n_2677, n_2679, n_2681, n_2682, n_2684, n_2686, n_2687;
  wire n_2689, n_2691, n_2692, n_2694, n_2695, n_2697, n_2700, n_2702;
  wire n_2703, n_2704, n_2707, n_2710, n_2712, n_2713, n_2715, n_2717;
  wire n_2718, n_2720, n_2722, n_2723, n_2725, n_2727, n_2728, n_2730;
  wire n_2731, n_2733, n_2736, n_2738, n_2739, n_2740, n_2743, n_2746;
  wire n_2748, n_2749, n_2751, n_2753, n_2754, n_2756, n_2758, n_2759;
  wire n_2761, n_2763, n_2764, n_2765, n_2767, n_2768, n_2770, n_2771;
  wire n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779;
  wire n_2780, n_2781, n_2783, n_2784, n_2785, n_2787, n_2788, n_2789;
  wire n_2791, n_2792, n_2793, n_2795, n_2796, n_2797, n_2799, n_2800;
  wire n_2801, n_2803, n_2804, n_2805, n_2807, n_2808, n_2809, n_2811;
  wire n_2812, n_2813, n_2814, n_2816, n_2818, n_2820, n_2821, n_2822;
  wire n_2824, n_2826, n_2828, n_2829, n_2831, n_2833, n_2834, n_2836;
  wire n_2838, n_2839, n_2842, n_2844, n_2845, n_2846, n_2848, n_2849;
  wire n_2850, n_2852, n_2853, n_2854, n_2856, n_2857, n_2858, n_2860;
  wire n_2861, n_2862, n_2864, n_2865, n_2866, n_2868, n_2869, n_2870;
  wire n_2872, n_2874, n_2875, n_2876, n_2878, n_2879, n_2881, n_2882;
  wire n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890;
  wire n_2891, n_2892, n_2894, n_2895, n_2896, n_2898, n_2899, n_2900;
  wire n_2902, n_2903, n_2904, n_2906, n_2907, n_2908, n_2910, n_2911;
  wire n_2912, n_2914, n_2915, n_2916, n_2918, n_2919, n_2921, n_2922;
  wire n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, n_2930;
  wire n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938;
  wire n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946;
  wire n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954;
  wire n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962;
  wire n_2963, n_2964, n_2965, n_2966, n_2968, n_2971, n_2972, n_2974;
  wire n_2975, n_2976, n_2977, n_2979, n_2980, n_2981, n_2983, n_2984;
  wire n_2985, n_2986, n_2988, n_2989, n_2991, n_2992, n_2994, n_2995;
  wire n_2996, n_2997, n_2999, n_3000, n_3001, n_3003, n_3004, n_3005;
  wire n_3006, n_3008, n_3009, n_3011, n_3012, n_3014, n_3015, n_3016;
  wire n_3017, n_3019, n_3020, n_3021, n_3022, n_3024, n_3025, n_3026;
  wire n_3027, n_3029, n_3030, n_3032, n_3033, n_3035, n_3036, n_3037;
  wire n_3038, n_3040, n_3041, n_3042, n_3044, n_3045, n_3046, n_3047;
  wire n_3049, n_3050, n_3052, n_3053, n_3055, n_3056, n_3057, n_3058;
  wire n_3060, n_3061, n_3062, n_3063, n_3065, n_3066, n_3067, n_3068;
  wire n_3070, n_3071, n_3073, n_3074, n_3076, n_3077, n_3078, n_3079;
  wire n_3081, n_3082, n_3084, n_3085, n_3087, n_3088, n_3089, n_3090;
  wire n_3092, n_3093, n_3095, n_3096, n_3098, n_3099, n_3100, n_3101;
  wire n_3103, n_3104, n_3105, n_3106, n_3108, n_3109, n_3110, n_3111;
  wire n_3113, n_3114, n_3116, n_3117, n_3119, n_3120, n_3121, n_3122;
  wire n_3124;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g356 (n_169, A[4], A[0]);
  and g2 (n_104, A[4], A[0]);
  xor g357 (n_834, A[1], A[3]);
  xor g358 (n_168, n_834, A[5]);
  nand g3 (n_835, A[1], A[3]);
  nand g359 (n_836, A[5], A[3]);
  nand g360 (n_837, A[1], A[5]);
  nand g361 (n_103, n_835, n_836, n_837);
  xor g362 (n_239, A[6], A[4]);
  and g363 (n_240, A[6], A[4]);
  xor g364 (n_838, A[0], A[2]);
  xor g365 (n_167, n_838, n_239);
  nand g366 (n_839, A[0], A[2]);
  nand g4 (n_840, n_239, A[2]);
  nand g5 (n_841, A[0], n_239);
  nand g367 (n_102, n_839, n_840, n_841);
  xor g368 (n_842, A[1], A[7]);
  xor g369 (n_241, n_842, A[5]);
  nand g370 (n_843, A[1], A[7]);
  nand g371 (n_844, A[5], A[7]);
  nand g6 (n_243, n_843, n_844, n_837);
  xor g373 (n_846, A[3], n_240);
  xor g374 (n_166, n_846, n_241);
  nand g375 (n_847, A[3], n_240);
  nand g376 (n_848, n_241, n_240);
  nand g377 (n_849, A[3], n_241);
  nand g378 (n_101, n_847, n_848, n_849);
  xor g379 (n_242, A[8], A[6]);
  and g380 (n_245, A[8], A[6]);
  xor g382 (n_244, n_838, A[4]);
  nand g385 (n_853, A[2], A[4]);
  xor g387 (n_854, n_242, n_243);
  xor g388 (n_165, n_854, n_244);
  nand g389 (n_855, n_242, n_243);
  nand g390 (n_856, n_244, n_243);
  nand g391 (n_857, n_242, n_244);
  nand g392 (n_100, n_855, n_856, n_857);
  xor g393 (n_858, A[1], A[9]);
  xor g394 (n_247, n_858, A[3]);
  nand g395 (n_859, A[1], A[9]);
  nand g396 (n_860, A[3], A[9]);
  nand g398 (n_250, n_859, n_860, n_835);
  xor g399 (n_862, A[7], A[5]);
  xor g400 (n_248, n_862, n_245);
  nand g402 (n_864, n_245, A[5]);
  nand g403 (n_865, A[7], n_245);
  nand g404 (n_252, n_844, n_864, n_865);
  xor g405 (n_866, n_246, n_247);
  xor g406 (n_164, n_866, n_248);
  nand g407 (n_867, n_246, n_247);
  nand g408 (n_868, n_248, n_247);
  nand g409 (n_869, n_246, n_248);
  nand g410 (n_99, n_867, n_868, n_869);
  xor g411 (n_249, A[10], A[8]);
  and g412 (n_254, A[10], A[8]);
  xor g413 (n_870, A[4], A[2]);
  xor g414 (n_251, n_870, A[6]);
  nand g416 (n_872, A[6], A[2]);
  xor g419 (n_874, A[0], n_249);
  xor g420 (n_253, n_874, n_250);
  nand g421 (n_875, A[0], n_249);
  nand g422 (n_876, n_250, n_249);
  nand g423 (n_877, A[0], n_250);
  nand g424 (n_258, n_875, n_876, n_877);
  xor g425 (n_878, n_251, n_252);
  xor g426 (n_163, n_878, n_253);
  nand g427 (n_879, n_251, n_252);
  nand g428 (n_880, n_253, n_252);
  nand g429 (n_881, n_251, n_253);
  nand g430 (n_98, n_879, n_880, n_881);
  xor g432 (n_256, n_858, A[5]);
  nand g434 (n_884, A[5], A[9]);
  nand g436 (n_261, n_859, n_884, n_837);
  xor g437 (n_886, A[3], A[11]);
  xor g438 (n_257, n_886, A[7]);
  nand g439 (n_887, A[3], A[11]);
  nand g440 (n_888, A[7], A[11]);
  nand g441 (n_889, A[3], A[7]);
  nand g442 (n_262, n_887, n_888, n_889);
  xor g443 (n_890, n_254, n_255);
  xor g444 (n_259, n_890, n_256);
  nand g445 (n_891, n_254, n_255);
  nand g446 (n_892, n_256, n_255);
  nand g447 (n_893, n_254, n_256);
  nand g448 (n_266, n_891, n_892, n_893);
  xor g449 (n_894, n_257, n_258);
  xor g450 (n_162, n_894, n_259);
  nand g451 (n_895, n_257, n_258);
  nand g452 (n_896, n_259, n_258);
  nand g453 (n_897, n_257, n_259);
  nand g454 (n_97, n_895, n_896, n_897);
  xor g455 (n_260, A[12], A[10]);
  and g456 (n_267, A[12], A[10]);
  xor g458 (n_263, n_239, A[8]);
  nand g460 (n_900, A[8], A[4]);
  xor g464 (n_264, n_838, n_260);
  nand g466 (n_904, n_260, A[0]);
  nand g467 (n_905, A[2], n_260);
  nand g468 (n_271, n_839, n_904, n_905);
  xor g469 (n_906, n_261, n_262);
  xor g470 (n_265, n_906, n_263);
  nand g471 (n_907, n_261, n_262);
  nand g472 (n_908, n_263, n_262);
  nand g473 (n_909, n_261, n_263);
  nand g474 (n_273, n_907, n_908, n_909);
  xor g475 (n_910, n_264, n_265);
  xor g476 (n_161, n_910, n_266);
  nand g477 (n_911, n_264, n_265);
  nand g478 (n_912, n_266, n_265);
  nand g479 (n_913, n_264, n_266);
  nand g480 (n_96, n_911, n_912, n_913);
  xor g481 (n_914, A[1], A[11]);
  xor g482 (n_270, n_914, A[7]);
  nand g483 (n_915, A[1], A[11]);
  nand g486 (n_276, n_915, n_888, n_843);
  xor g487 (n_918, A[5], A[13]);
  xor g488 (n_269, n_918, A[3]);
  nand g489 (n_919, A[5], A[13]);
  nand g490 (n_920, A[3], A[13]);
  nand g492 (n_277, n_919, n_920, n_836);
  xor g493 (n_922, A[9], n_267);
  xor g494 (n_272, n_922, n_268);
  nand g495 (n_923, A[9], n_267);
  nand g496 (n_924, n_268, n_267);
  nand g497 (n_925, A[9], n_268);
  nand g498 (n_280, n_923, n_924, n_925);
  xor g499 (n_926, n_269, n_270);
  xor g500 (n_274, n_926, n_271);
  nand g501 (n_927, n_269, n_270);
  nand g502 (n_928, n_271, n_270);
  nand g503 (n_929, n_269, n_271);
  nand g504 (n_282, n_927, n_928, n_929);
  xor g505 (n_930, n_272, n_273);
  xor g506 (n_160, n_930, n_274);
  nand g507 (n_931, n_272, n_273);
  nand g508 (n_932, n_274, n_273);
  nand g509 (n_933, n_272, n_274);
  nand g510 (n_95, n_931, n_932, n_933);
  xor g511 (n_275, A[14], A[12]);
  and g512 (n_284, A[14], A[12]);
  xor g513 (n_934, A[8], A[0]);
  xor g514 (n_279, n_934, A[6]);
  nand g515 (n_935, A[8], A[0]);
  nand g516 (n_936, A[6], A[0]);
  xor g519 (n_938, A[10], A[4]);
  xor g520 (n_278, n_938, A[2]);
  nand g521 (n_939, A[10], A[4]);
  nand g523 (n_941, A[10], A[2]);
  nand g524 (n_286, n_939, n_853, n_941);
  xor g525 (n_942, n_275, n_276);
  xor g526 (n_281, n_942, n_277);
  nand g527 (n_943, n_275, n_276);
  nand g528 (n_944, n_277, n_276);
  nand g529 (n_945, n_275, n_277);
  nand g530 (n_290, n_943, n_944, n_945);
  xor g531 (n_946, n_278, n_279);
  xor g532 (n_283, n_946, n_280);
  nand g533 (n_947, n_278, n_279);
  nand g534 (n_948, n_280, n_279);
  nand g535 (n_949, n_278, n_280);
  nand g536 (n_293, n_947, n_948, n_949);
  xor g537 (n_950, n_281, n_282);
  xor g538 (n_159, n_950, n_283);
  nand g539 (n_951, n_281, n_282);
  nand g540 (n_952, n_283, n_282);
  nand g541 (n_953, n_281, n_283);
  nand g542 (n_94, n_951, n_952, n_953);
  xor g543 (n_954, A[1], A[15]);
  xor g544 (n_287, n_954, A[13]);
  nand g545 (n_955, A[1], A[15]);
  nand g546 (n_956, A[13], A[15]);
  nand g547 (n_957, A[1], A[13]);
  nand g548 (n_295, n_955, n_956, n_957);
  xor g549 (n_958, A[9], A[7]);
  xor g550 (n_288, n_958, A[11]);
  nand g551 (n_959, A[9], A[7]);
  nand g553 (n_961, A[9], A[11]);
  nand g554 (n_296, n_959, n_888, n_961);
  xor g555 (n_962, A[5], A[3]);
  xor g556 (n_289, n_962, n_284);
  nand g558 (n_964, n_284, A[3]);
  nand g559 (n_965, A[5], n_284);
  nand g560 (n_299, n_836, n_964, n_965);
  xor g561 (n_966, n_285, n_286);
  xor g562 (n_291, n_966, n_287);
  nand g563 (n_967, n_285, n_286);
  nand g564 (n_968, n_287, n_286);
  nand g565 (n_969, n_285, n_287);
  nand g566 (n_301, n_967, n_968, n_969);
  xor g567 (n_970, n_288, n_289);
  xor g568 (n_292, n_970, n_290);
  nand g569 (n_971, n_288, n_289);
  nand g570 (n_972, n_290, n_289);
  nand g571 (n_973, n_288, n_290);
  nand g572 (n_303, n_971, n_972, n_973);
  xor g573 (n_974, n_291, n_292);
  xor g574 (n_158, n_974, n_293);
  nand g575 (n_975, n_291, n_292);
  nand g576 (n_976, n_293, n_292);
  nand g577 (n_977, n_291, n_293);
  nand g578 (n_93, n_975, n_976, n_977);
  xor g579 (n_294, A[16], A[14]);
  and g580 (n_305, A[16], A[14]);
  xor g581 (n_978, A[10], A[2]);
  xor g582 (n_298, n_978, A[0]);
  nand g585 (n_981, A[10], A[0]);
  nand g586 (n_306, n_941, n_839, n_981);
  xor g587 (n_982, A[8], A[12]);
  xor g588 (n_297, n_982, A[6]);
  nand g589 (n_983, A[8], A[12]);
  nand g590 (n_984, A[6], A[12]);
  xor g593 (n_986, A[4], n_294);
  xor g594 (n_300, n_986, n_295);
  nand g595 (n_987, A[4], n_294);
  nand g596 (n_988, n_295, n_294);
  nand g597 (n_989, A[4], n_295);
  nand g598 (n_311, n_987, n_988, n_989);
  xor g599 (n_990, n_296, n_297);
  xor g600 (n_302, n_990, n_298);
  nand g601 (n_991, n_296, n_297);
  nand g602 (n_992, n_298, n_297);
  nand g603 (n_993, n_296, n_298);
  nand g604 (n_313, n_991, n_992, n_993);
  xor g605 (n_994, n_299, n_300);
  xor g606 (n_304, n_994, n_301);
  nand g607 (n_995, n_299, n_300);
  nand g608 (n_996, n_301, n_300);
  nand g609 (n_997, n_299, n_301);
  nand g610 (n_315, n_995, n_996, n_997);
  xor g611 (n_998, n_302, n_303);
  xor g612 (n_157, n_998, n_304);
  nand g613 (n_999, n_302, n_303);
  nand g614 (n_1000, n_304, n_303);
  nand g615 (n_1001, n_302, n_304);
  nand g616 (n_92, n_999, n_1000, n_1001);
  xor g617 (n_1002, A[1], A[17]);
  xor g618 (n_309, n_1002, A[15]);
  nand g619 (n_1003, A[1], A[17]);
  nand g620 (n_1004, A[15], A[17]);
  nand g622 (n_318, n_1003, n_1004, n_955);
  xor g624 (n_310, n_886, A[9]);
  nand g628 (n_320, n_887, n_961, n_860);
  xor g629 (n_1010, A[13], A[7]);
  xor g630 (n_308, n_1010, A[5]);
  nand g631 (n_1011, A[13], A[7]);
  nand g634 (n_319, n_1011, n_844, n_919);
  xor g635 (n_1014, n_305, n_306);
  xor g636 (n_312, n_1014, n_307);
  nand g637 (n_1015, n_305, n_306);
  nand g638 (n_1016, n_307, n_306);
  nand g639 (n_1017, n_305, n_307);
  nand g640 (n_106, n_1015, n_1016, n_1017);
  xor g641 (n_1018, n_308, n_309);
  xor g642 (n_314, n_1018, n_310);
  nand g643 (n_1019, n_308, n_309);
  nand g644 (n_1020, n_310, n_309);
  nand g645 (n_1021, n_308, n_310);
  nand g646 (n_108, n_1019, n_1020, n_1021);
  xor g647 (n_1022, n_311, n_312);
  xor g648 (n_316, n_1022, n_313);
  nand g649 (n_1023, n_311, n_312);
  nand g650 (n_1024, n_313, n_312);
  nand g651 (n_1025, n_311, n_313);
  nand g652 (n_323, n_1023, n_1024, n_1025);
  xor g653 (n_1026, n_314, n_315);
  xor g654 (n_156, n_1026, n_316);
  nand g655 (n_1027, n_314, n_315);
  nand g656 (n_1028, n_316, n_315);
  nand g657 (n_1029, n_314, n_316);
  nand g658 (n_91, n_1027, n_1028, n_1029);
  xor g659 (n_317, A[18], A[16]);
  and g660 (n_325, A[18], A[16]);
  xor g661 (n_1030, A[12], A[4]);
  xor g662 (n_321, n_1030, A[2]);
  nand g663 (n_1031, A[12], A[4]);
  nand g665 (n_1033, A[12], A[2]);
  nand g666 (n_326, n_1031, n_853, n_1033);
  xor g667 (n_1034, A[10], A[0]);
  xor g668 (n_322, n_1034, A[14]);
  nand g670 (n_1036, A[14], A[0]);
  nand g671 (n_1037, A[10], A[14]);
  nand g672 (n_327, n_981, n_1036, n_1037);
  xor g674 (n_105, n_242, n_317);
  nand g676 (n_1040, n_317, A[6]);
  nand g677 (n_1041, A[8], n_317);
  xor g679 (n_1042, n_318, n_319);
  xor g680 (n_107, n_1042, n_320);
  nand g681 (n_1043, n_318, n_319);
  nand g682 (n_1044, n_320, n_319);
  nand g683 (n_1045, n_318, n_320);
  nand g684 (n_333, n_1043, n_1044, n_1045);
  xor g685 (n_1046, n_321, n_322);
  xor g686 (n_109, n_1046, n_105);
  nand g687 (n_1047, n_321, n_322);
  nand g688 (n_1048, n_105, n_322);
  nand g689 (n_1049, n_321, n_105);
  nand g690 (n_334, n_1047, n_1048, n_1049);
  xor g691 (n_1050, n_106, n_107);
  xor g692 (n_324, n_1050, n_108);
  nand g693 (n_1051, n_106, n_107);
  nand g694 (n_1052, n_108, n_107);
  nand g695 (n_1053, n_106, n_108);
  nand g696 (n_337, n_1051, n_1052, n_1053);
  xor g697 (n_1054, n_109, n_323);
  xor g698 (n_155, n_1054, n_324);
  nand g699 (n_1055, n_109, n_323);
  nand g700 (n_1056, n_324, n_323);
  nand g701 (n_1057, n_109, n_324);
  nand g702 (n_90, n_1055, n_1056, n_1057);
  xor g703 (n_1058, A[1], A[19]);
  xor g704 (n_329, n_1058, A[13]);
  nand g705 (n_1059, A[1], A[19]);
  nand g706 (n_1060, A[13], A[19]);
  nand g708 (n_339, n_1059, n_1060, n_957);
  xor g710 (n_330, n_962, A[17]);
  nand g712 (n_1064, A[17], A[3]);
  nand g713 (n_1065, A[5], A[17]);
  nand g714 (n_340, n_836, n_1064, n_1065);
  xor g715 (n_1066, A[11], A[15]);
  xor g716 (n_328, n_1066, A[9]);
  nand g717 (n_1067, A[11], A[15]);
  nand g718 (n_1068, A[9], A[15]);
  nand g720 (n_341, n_1067, n_1068, n_961);
  xor g721 (n_1070, A[7], n_325);
  xor g722 (n_332, n_1070, n_326);
  nand g723 (n_1071, A[7], n_325);
  nand g724 (n_1072, n_326, n_325);
  nand g725 (n_1073, A[7], n_326);
  nand g726 (n_345, n_1071, n_1072, n_1073);
  xor g727 (n_1074, n_327, n_328);
  xor g728 (n_335, n_1074, n_329);
  nand g729 (n_1075, n_327, n_328);
  nand g730 (n_1076, n_329, n_328);
  nand g731 (n_1077, n_327, n_329);
  nand g732 (n_347, n_1075, n_1076, n_1077);
  xor g733 (n_1078, n_330, n_331);
  xor g734 (n_336, n_1078, n_332);
  nand g735 (n_1079, n_330, n_331);
  nand g736 (n_1080, n_332, n_331);
  nand g737 (n_1081, n_330, n_332);
  nand g738 (n_349, n_1079, n_1080, n_1081);
  xor g739 (n_1082, n_333, n_334);
  xor g740 (n_338, n_1082, n_335);
  nand g741 (n_1083, n_333, n_334);
  nand g742 (n_1084, n_335, n_334);
  nand g743 (n_1085, n_333, n_335);
  nand g744 (n_351, n_1083, n_1084, n_1085);
  xor g745 (n_1086, n_336, n_337);
  xor g746 (n_154, n_1086, n_338);
  nand g747 (n_1087, n_336, n_337);
  nand g748 (n_1088, n_338, n_337);
  nand g749 (n_1089, n_336, n_338);
  nand g750 (n_89, n_1087, n_1088, n_1089);
  xor g751 (n_1090, A[20], A[18]);
  xor g752 (n_343, n_1090, A[14]);
  nand g753 (n_1091, A[20], A[18]);
  nand g754 (n_1092, A[14], A[18]);
  nand g755 (n_1093, A[20], A[14]);
  nand g756 (n_353, n_1091, n_1092, n_1093);
  xor g758 (n_344, n_239, A[12]);
  xor g763 (n_1098, A[2], A[16]);
  xor g764 (n_342, n_1098, A[10]);
  nand g765 (n_1099, A[2], A[16]);
  nand g766 (n_1100, A[10], A[16]);
  nand g768 (n_355, n_1099, n_1100, n_941);
  xor g769 (n_1102, A[8], n_339);
  xor g770 (n_346, n_1102, n_340);
  nand g771 (n_1103, A[8], n_339);
  nand g772 (n_1104, n_340, n_339);
  nand g773 (n_1105, A[8], n_340);
  nand g774 (n_359, n_1103, n_1104, n_1105);
  xor g775 (n_1106, n_341, n_342);
  xor g776 (n_348, n_1106, n_343);
  nand g777 (n_1107, n_341, n_342);
  nand g778 (n_1108, n_343, n_342);
  nand g779 (n_1109, n_341, n_343);
  nand g780 (n_361, n_1107, n_1108, n_1109);
  xor g781 (n_1110, n_344, n_345);
  xor g782 (n_350, n_1110, n_346);
  nand g783 (n_1111, n_344, n_345);
  nand g784 (n_1112, n_346, n_345);
  nand g785 (n_1113, n_344, n_346);
  nand g786 (n_363, n_1111, n_1112, n_1113);
  xor g787 (n_1114, n_347, n_348);
  xor g788 (n_352, n_1114, n_349);
  nand g789 (n_1115, n_347, n_348);
  nand g790 (n_1116, n_349, n_348);
  nand g791 (n_1117, n_347, n_349);
  nand g792 (n_365, n_1115, n_1116, n_1117);
  xor g793 (n_1118, n_350, n_351);
  xor g794 (n_153, n_1118, n_352);
  nand g795 (n_1119, n_350, n_351);
  nand g796 (n_1120, n_352, n_351);
  nand g797 (n_1121, n_350, n_352);
  nand g798 (n_88, n_1119, n_1120, n_1121);
  xor g799 (n_1122, A[21], A[19]);
  xor g800 (n_357, n_1122, A[15]);
  nand g801 (n_1123, A[21], A[19]);
  nand g802 (n_1124, A[15], A[19]);
  nand g803 (n_1125, A[21], A[15]);
  nand g804 (n_367, n_1123, n_1124, n_1125);
  xor g806 (n_358, n_862, A[13]);
  xor g811 (n_1130, A[3], A[17]);
  xor g812 (n_356, n_1130, A[11]);
  nand g814 (n_1132, A[11], A[17]);
  nand g816 (n_369, n_1064, n_1132, n_887);
  xor g817 (n_1134, A[9], n_353);
  xor g818 (n_360, n_1134, n_354);
  nand g819 (n_1135, A[9], n_353);
  nand g820 (n_1136, n_354, n_353);
  nand g821 (n_1137, A[9], n_354);
  nand g822 (n_373, n_1135, n_1136, n_1137);
  xor g823 (n_1138, n_355, n_356);
  xor g824 (n_362, n_1138, n_357);
  nand g825 (n_1139, n_355, n_356);
  nand g826 (n_1140, n_357, n_356);
  nand g827 (n_1141, n_355, n_357);
  nand g828 (n_375, n_1139, n_1140, n_1141);
  xor g829 (n_1142, n_358, n_359);
  xor g830 (n_364, n_1142, n_360);
  nand g831 (n_1143, n_358, n_359);
  nand g832 (n_1144, n_360, n_359);
  nand g833 (n_1145, n_358, n_360);
  nand g834 (n_377, n_1143, n_1144, n_1145);
  xor g835 (n_1146, n_361, n_362);
  xor g836 (n_366, n_1146, n_363);
  nand g837 (n_1147, n_361, n_362);
  nand g838 (n_1148, n_363, n_362);
  nand g839 (n_1149, n_361, n_363);
  nand g840 (n_171, n_1147, n_1148, n_1149);
  xor g841 (n_1150, n_364, n_365);
  xor g842 (n_152, n_1150, n_366);
  nand g843 (n_1151, n_364, n_365);
  nand g844 (n_1152, n_366, n_365);
  nand g845 (n_1153, n_364, n_366);
  nand g846 (n_87, n_1151, n_1152, n_1153);
  xor g847 (n_1154, A[22], A[20]);
  xor g848 (n_371, n_1154, A[16]);
  nand g849 (n_1155, A[22], A[20]);
  nand g850 (n_1156, A[16], A[20]);
  nand g851 (n_1157, A[22], A[16]);
  nand g852 (n_379, n_1155, n_1156, n_1157);
  xor g854 (n_372, n_242, A[14]);
  nand g856 (n_1160, A[14], A[6]);
  nand g857 (n_1161, A[8], A[14]);
  xor g859 (n_1162, A[4], A[18]);
  xor g860 (n_370, n_1162, A[12]);
  nand g861 (n_1163, A[4], A[18]);
  nand g862 (n_1164, A[12], A[18]);
  nand g864 (n_381, n_1163, n_1164, n_1031);
  xor g865 (n_1166, A[10], n_367);
  xor g866 (n_374, n_1166, n_319);
  nand g867 (n_1167, A[10], n_367);
  nand g868 (n_1168, n_319, n_367);
  nand g869 (n_1169, A[10], n_319);
  nand g870 (n_385, n_1167, n_1168, n_1169);
  xor g871 (n_1170, n_369, n_370);
  xor g872 (n_376, n_1170, n_371);
  nand g873 (n_1171, n_369, n_370);
  nand g874 (n_1172, n_371, n_370);
  nand g875 (n_1173, n_369, n_371);
  nand g876 (n_387, n_1171, n_1172, n_1173);
  xor g877 (n_1174, n_372, n_373);
  xor g878 (n_378, n_1174, n_374);
  nand g879 (n_1175, n_372, n_373);
  nand g880 (n_1176, n_374, n_373);
  nand g881 (n_1177, n_372, n_374);
  nand g882 (n_389, n_1175, n_1176, n_1177);
  xor g883 (n_1178, n_375, n_376);
  xor g884 (n_170, n_1178, n_377);
  nand g885 (n_1179, n_375, n_376);
  nand g886 (n_1180, n_377, n_376);
  nand g887 (n_1181, n_375, n_377);
  nand g888 (n_392, n_1179, n_1180, n_1181);
  xor g889 (n_1182, n_378, n_170);
  xor g890 (n_151, n_1182, n_171);
  nand g891 (n_1183, n_378, n_170);
  nand g892 (n_1184, n_171, n_170);
  nand g893 (n_1185, n_378, n_171);
  nand g894 (n_86, n_1183, n_1184, n_1185);
  xor g895 (n_1186, A[23], A[21]);
  xor g896 (n_383, n_1186, A[17]);
  nand g897 (n_1187, A[23], A[21]);
  nand g898 (n_1188, A[17], A[21]);
  nand g899 (n_1189, A[23], A[17]);
  nand g900 (n_393, n_1187, n_1188, n_1189);
  xor g902 (n_384, n_958, A[15]);
  nand g904 (n_1192, A[15], A[7]);
  nand g906 (n_394, n_959, n_1192, n_1068);
  xor g907 (n_1194, A[5], A[19]);
  xor g908 (n_382, n_1194, A[13]);
  nand g909 (n_1195, A[5], A[19]);
  nand g912 (n_395, n_1195, n_1060, n_919);
  xor g913 (n_1198, A[11], n_379);
  xor g914 (n_386, n_1198, n_380);
  nand g915 (n_1199, A[11], n_379);
  nand g916 (n_1200, n_380, n_379);
  nand g917 (n_1201, A[11], n_380);
  nand g918 (n_399, n_1199, n_1200, n_1201);
  xor g919 (n_1202, n_381, n_382);
  xor g920 (n_388, n_1202, n_383);
  nand g921 (n_1203, n_381, n_382);
  nand g922 (n_1204, n_383, n_382);
  nand g923 (n_1205, n_381, n_383);
  nand g924 (n_401, n_1203, n_1204, n_1205);
  xor g925 (n_1206, n_384, n_385);
  xor g926 (n_390, n_1206, n_386);
  nand g927 (n_1207, n_384, n_385);
  nand g928 (n_1208, n_386, n_385);
  nand g929 (n_1209, n_384, n_386);
  nand g930 (n_403, n_1207, n_1208, n_1209);
  xor g931 (n_1210, n_387, n_388);
  xor g932 (n_391, n_1210, n_389);
  nand g933 (n_1211, n_387, n_388);
  nand g934 (n_1212, n_389, n_388);
  nand g935 (n_1213, n_387, n_389);
  nand g936 (n_406, n_1211, n_1212, n_1213);
  xor g937 (n_1214, n_390, n_391);
  xor g938 (n_150, n_1214, n_392);
  nand g939 (n_1215, n_390, n_391);
  nand g940 (n_1216, n_392, n_391);
  nand g941 (n_1217, n_390, n_392);
  nand g942 (n_85, n_1215, n_1216, n_1217);
  xor g943 (n_1218, A[24], A[22]);
  xor g944 (n_397, n_1218, A[18]);
  nand g945 (n_1219, A[24], A[22]);
  nand g946 (n_1220, A[18], A[22]);
  nand g947 (n_1221, A[24], A[18]);
  nand g948 (n_407, n_1219, n_1220, n_1221);
  xor g950 (n_398, n_249, A[16]);
  nand g952 (n_1224, A[16], A[8]);
  xor g955 (n_1226, A[6], A[20]);
  xor g956 (n_396, n_1226, A[14]);
  nand g957 (n_1227, A[6], A[20]);
  nand g960 (n_409, n_1227, n_1093, n_1160);
  xor g961 (n_1230, A[12], n_393);
  xor g962 (n_400, n_1230, n_394);
  nand g963 (n_1231, A[12], n_393);
  nand g964 (n_1232, n_394, n_393);
  nand g965 (n_1233, A[12], n_394);
  nand g966 (n_413, n_1231, n_1232, n_1233);
  xor g967 (n_1234, n_395, n_396);
  xor g968 (n_402, n_1234, n_397);
  nand g969 (n_1235, n_395, n_396);
  nand g970 (n_1236, n_397, n_396);
  nand g971 (n_1237, n_395, n_397);
  nand g972 (n_415, n_1235, n_1236, n_1237);
  xor g973 (n_1238, n_398, n_399);
  xor g974 (n_404, n_1238, n_400);
  nand g975 (n_1239, n_398, n_399);
  nand g976 (n_1240, n_400, n_399);
  nand g977 (n_1241, n_398, n_400);
  nand g978 (n_417, n_1239, n_1240, n_1241);
  xor g979 (n_1242, n_401, n_402);
  xor g980 (n_405, n_1242, n_403);
  nand g981 (n_1243, n_401, n_402);
  nand g982 (n_1244, n_403, n_402);
  nand g983 (n_1245, n_401, n_403);
  nand g984 (n_420, n_1243, n_1244, n_1245);
  xor g985 (n_1246, n_404, n_405);
  xor g986 (n_149, n_1246, n_406);
  nand g987 (n_1247, n_404, n_405);
  nand g988 (n_1248, n_406, n_405);
  nand g989 (n_1249, n_404, n_406);
  nand g990 (n_84, n_1247, n_1248, n_1249);
  xor g991 (n_1250, A[25], A[23]);
  xor g992 (n_411, n_1250, A[19]);
  nand g993 (n_1251, A[25], A[23]);
  nand g994 (n_1252, A[19], A[23]);
  nand g995 (n_1253, A[25], A[19]);
  nand g996 (n_421, n_1251, n_1252, n_1253);
  xor g997 (n_1254, A[11], A[9]);
  xor g998 (n_412, n_1254, A[17]);
  nand g1000 (n_1256, A[17], A[9]);
  nand g1002 (n_422, n_961, n_1256, n_1132);
  xor g1003 (n_1258, A[7], A[21]);
  xor g1004 (n_410, n_1258, A[15]);
  nand g1005 (n_1259, A[7], A[21]);
  nand g1008 (n_423, n_1259, n_1125, n_1192);
  xor g1009 (n_1262, A[13], n_407);
  xor g1010 (n_414, n_1262, n_408);
  nand g1011 (n_1263, A[13], n_407);
  nand g1012 (n_1264, n_408, n_407);
  nand g1013 (n_1265, A[13], n_408);
  nand g1014 (n_427, n_1263, n_1264, n_1265);
  xor g1015 (n_1266, n_409, n_410);
  xor g1016 (n_416, n_1266, n_411);
  nand g1017 (n_1267, n_409, n_410);
  nand g1018 (n_1268, n_411, n_410);
  nand g1019 (n_1269, n_409, n_411);
  nand g1020 (n_429, n_1267, n_1268, n_1269);
  xor g1021 (n_1270, n_412, n_413);
  xor g1022 (n_418, n_1270, n_414);
  nand g1023 (n_1271, n_412, n_413);
  nand g1024 (n_1272, n_414, n_413);
  nand g1025 (n_1273, n_412, n_414);
  nand g1026 (n_431, n_1271, n_1272, n_1273);
  xor g1027 (n_1274, n_415, n_416);
  xor g1028 (n_419, n_1274, n_417);
  nand g1029 (n_1275, n_415, n_416);
  nand g1030 (n_1276, n_417, n_416);
  nand g1031 (n_1277, n_415, n_417);
  nand g1032 (n_434, n_1275, n_1276, n_1277);
  xor g1033 (n_1278, n_418, n_419);
  xor g1034 (n_148, n_1278, n_420);
  nand g1035 (n_1279, n_418, n_419);
  nand g1036 (n_1280, n_420, n_419);
  nand g1037 (n_1281, n_418, n_420);
  nand g1038 (n_83, n_1279, n_1280, n_1281);
  xor g1039 (n_1282, A[26], A[24]);
  xor g1040 (n_425, n_1282, A[20]);
  nand g1041 (n_1283, A[26], A[24]);
  nand g1042 (n_1284, A[20], A[24]);
  nand g1043 (n_1285, A[26], A[20]);
  nand g1044 (n_435, n_1283, n_1284, n_1285);
  xor g1046 (n_426, n_260, A[18]);
  nand g1048 (n_1288, A[18], A[10]);
  xor g1051 (n_1290, A[8], A[22]);
  xor g1052 (n_424, n_1290, A[16]);
  nand g1053 (n_1291, A[8], A[22]);
  nand g1056 (n_437, n_1291, n_1157, n_1224);
  xor g1057 (n_1294, A[14], n_421);
  xor g1058 (n_428, n_1294, n_422);
  nand g1059 (n_1295, A[14], n_421);
  nand g1060 (n_1296, n_422, n_421);
  nand g1061 (n_1297, A[14], n_422);
  nand g1062 (n_441, n_1295, n_1296, n_1297);
  xor g1063 (n_1298, n_423, n_424);
  xor g1064 (n_430, n_1298, n_425);
  nand g1065 (n_1299, n_423, n_424);
  nand g1066 (n_1300, n_425, n_424);
  nand g1067 (n_1301, n_423, n_425);
  nand g1068 (n_443, n_1299, n_1300, n_1301);
  xor g1069 (n_1302, n_426, n_427);
  xor g1070 (n_432, n_1302, n_428);
  nand g1071 (n_1303, n_426, n_427);
  nand g1072 (n_1304, n_428, n_427);
  nand g1073 (n_1305, n_426, n_428);
  nand g1074 (n_445, n_1303, n_1304, n_1305);
  xor g1075 (n_1306, n_429, n_430);
  xor g1076 (n_433, n_1306, n_431);
  nand g1077 (n_1307, n_429, n_430);
  nand g1078 (n_1308, n_431, n_430);
  nand g1079 (n_1309, n_429, n_431);
  nand g1080 (n_448, n_1307, n_1308, n_1309);
  xor g1081 (n_1310, n_432, n_433);
  xor g1082 (n_147, n_1310, n_434);
  nand g1083 (n_1311, n_432, n_433);
  nand g1084 (n_1312, n_434, n_433);
  nand g1085 (n_1313, n_432, n_434);
  nand g1086 (n_82, n_1311, n_1312, n_1313);
  xor g1087 (n_1314, A[27], A[25]);
  xor g1088 (n_439, n_1314, A[21]);
  nand g1089 (n_1315, A[27], A[25]);
  nand g1090 (n_1316, A[21], A[25]);
  nand g1091 (n_1317, A[27], A[21]);
  nand g1092 (n_449, n_1315, n_1316, n_1317);
  xor g1093 (n_1318, A[13], A[11]);
  xor g1094 (n_440, n_1318, A[19]);
  nand g1095 (n_1319, A[13], A[11]);
  nand g1096 (n_1320, A[19], A[11]);
  nand g1098 (n_450, n_1319, n_1320, n_1060);
  xor g1099 (n_1322, A[9], A[23]);
  xor g1100 (n_438, n_1322, A[17]);
  nand g1101 (n_1323, A[9], A[23]);
  nand g1104 (n_451, n_1323, n_1189, n_1256);
  xor g1105 (n_1326, A[15], n_435);
  xor g1106 (n_442, n_1326, n_436);
  nand g1107 (n_1327, A[15], n_435);
  nand g1108 (n_1328, n_436, n_435);
  nand g1109 (n_1329, A[15], n_436);
  nand g1110 (n_455, n_1327, n_1328, n_1329);
  xor g1111 (n_1330, n_437, n_438);
  xor g1112 (n_444, n_1330, n_439);
  nand g1113 (n_1331, n_437, n_438);
  nand g1114 (n_1332, n_439, n_438);
  nand g1115 (n_1333, n_437, n_439);
  nand g1116 (n_457, n_1331, n_1332, n_1333);
  xor g1117 (n_1334, n_440, n_441);
  xor g1118 (n_446, n_1334, n_442);
  nand g1119 (n_1335, n_440, n_441);
  nand g1120 (n_1336, n_442, n_441);
  nand g1121 (n_1337, n_440, n_442);
  nand g1122 (n_459, n_1335, n_1336, n_1337);
  xor g1123 (n_1338, n_443, n_444);
  xor g1124 (n_447, n_1338, n_445);
  nand g1125 (n_1339, n_443, n_444);
  nand g1126 (n_1340, n_445, n_444);
  nand g1127 (n_1341, n_443, n_445);
  nand g1128 (n_462, n_1339, n_1340, n_1341);
  xor g1129 (n_1342, n_446, n_447);
  xor g1130 (n_146, n_1342, n_448);
  nand g1131 (n_1343, n_446, n_447);
  nand g1132 (n_1344, n_448, n_447);
  nand g1133 (n_1345, n_446, n_448);
  nand g1134 (n_81, n_1343, n_1344, n_1345);
  xor g1135 (n_1346, A[28], A[26]);
  xor g1136 (n_453, n_1346, A[22]);
  nand g1137 (n_1347, A[28], A[26]);
  nand g1138 (n_1348, A[22], A[26]);
  nand g1139 (n_1349, A[28], A[22]);
  nand g1140 (n_463, n_1347, n_1348, n_1349);
  xor g1142 (n_454, n_275, A[20]);
  nand g1144 (n_1352, A[20], A[12]);
  xor g1147 (n_1354, A[10], A[24]);
  xor g1148 (n_452, n_1354, A[18]);
  nand g1149 (n_1355, A[10], A[24]);
  nand g1152 (n_465, n_1355, n_1221, n_1288);
  xor g1153 (n_1358, A[16], n_449);
  xor g1154 (n_456, n_1358, n_450);
  nand g1155 (n_1359, A[16], n_449);
  nand g1156 (n_1360, n_450, n_449);
  nand g1157 (n_1361, A[16], n_450);
  nand g1158 (n_469, n_1359, n_1360, n_1361);
  xor g1159 (n_1362, n_451, n_452);
  xor g1160 (n_458, n_1362, n_453);
  nand g1161 (n_1363, n_451, n_452);
  nand g1162 (n_1364, n_453, n_452);
  nand g1163 (n_1365, n_451, n_453);
  nand g1164 (n_471, n_1363, n_1364, n_1365);
  xor g1165 (n_1366, n_454, n_455);
  xor g1166 (n_460, n_1366, n_456);
  nand g1167 (n_1367, n_454, n_455);
  nand g1168 (n_1368, n_456, n_455);
  nand g1169 (n_1369, n_454, n_456);
  nand g1170 (n_473, n_1367, n_1368, n_1369);
  xor g1171 (n_1370, n_457, n_458);
  xor g1172 (n_461, n_1370, n_459);
  nand g1173 (n_1371, n_457, n_458);
  nand g1174 (n_1372, n_459, n_458);
  nand g1175 (n_1373, n_457, n_459);
  nand g1176 (n_476, n_1371, n_1372, n_1373);
  xor g1177 (n_1374, n_460, n_461);
  xor g1178 (n_145, n_1374, n_462);
  nand g1179 (n_1375, n_460, n_461);
  nand g1180 (n_1376, n_462, n_461);
  nand g1181 (n_1377, n_460, n_462);
  nand g1182 (n_80, n_1375, n_1376, n_1377);
  xor g1183 (n_1378, A[29], A[27]);
  xor g1184 (n_467, n_1378, A[23]);
  nand g1185 (n_1379, A[29], A[27]);
  nand g1186 (n_1380, A[23], A[27]);
  nand g1187 (n_1381, A[29], A[23]);
  nand g1188 (n_477, n_1379, n_1380, n_1381);
  xor g1189 (n_1382, A[15], A[13]);
  xor g1190 (n_468, n_1382, A[21]);
  nand g1192 (n_1384, A[21], A[13]);
  nand g1194 (n_478, n_956, n_1384, n_1125);
  xor g1195 (n_1386, A[11], A[25]);
  xor g1196 (n_466, n_1386, A[19]);
  nand g1197 (n_1387, A[11], A[25]);
  nand g1200 (n_479, n_1387, n_1253, n_1320);
  xor g1201 (n_1390, A[17], n_463);
  xor g1202 (n_470, n_1390, n_464);
  nand g1203 (n_1391, A[17], n_463);
  nand g1204 (n_1392, n_464, n_463);
  nand g1205 (n_1393, A[17], n_464);
  nand g1206 (n_483, n_1391, n_1392, n_1393);
  xor g1207 (n_1394, n_465, n_466);
  xor g1208 (n_472, n_1394, n_467);
  nand g1209 (n_1395, n_465, n_466);
  nand g1210 (n_1396, n_467, n_466);
  nand g1211 (n_1397, n_465, n_467);
  nand g1212 (n_485, n_1395, n_1396, n_1397);
  xor g1213 (n_1398, n_468, n_469);
  xor g1214 (n_474, n_1398, n_470);
  nand g1215 (n_1399, n_468, n_469);
  nand g1216 (n_1400, n_470, n_469);
  nand g1217 (n_1401, n_468, n_470);
  nand g1218 (n_487, n_1399, n_1400, n_1401);
  xor g1219 (n_1402, n_471, n_472);
  xor g1220 (n_475, n_1402, n_473);
  nand g1221 (n_1403, n_471, n_472);
  nand g1222 (n_1404, n_473, n_472);
  nand g1223 (n_1405, n_471, n_473);
  nand g1224 (n_490, n_1403, n_1404, n_1405);
  xor g1225 (n_1406, n_474, n_475);
  xor g1226 (n_144, n_1406, n_476);
  nand g1227 (n_1407, n_474, n_475);
  nand g1228 (n_1408, n_476, n_475);
  nand g1229 (n_1409, n_474, n_476);
  nand g1230 (n_79, n_1407, n_1408, n_1409);
  xor g1231 (n_1410, A[30], A[28]);
  xor g1232 (n_481, n_1410, A[24]);
  nand g1233 (n_1411, A[30], A[28]);
  nand g1234 (n_1412, A[24], A[28]);
  nand g1235 (n_1413, A[30], A[24]);
  nand g1236 (n_491, n_1411, n_1412, n_1413);
  xor g1238 (n_482, n_294, A[22]);
  nand g1240 (n_1416, A[22], A[14]);
  xor g1243 (n_1418, A[12], A[26]);
  xor g1244 (n_480, n_1418, A[20]);
  nand g1245 (n_1419, A[12], A[26]);
  nand g1248 (n_493, n_1419, n_1285, n_1352);
  xor g1249 (n_1422, A[18], n_477);
  xor g1250 (n_484, n_1422, n_478);
  nand g1251 (n_1423, A[18], n_477);
  nand g1252 (n_1424, n_478, n_477);
  nand g1253 (n_1425, A[18], n_478);
  nand g1254 (n_497, n_1423, n_1424, n_1425);
  xor g1255 (n_1426, n_479, n_480);
  xor g1256 (n_486, n_1426, n_481);
  nand g1257 (n_1427, n_479, n_480);
  nand g1258 (n_1428, n_481, n_480);
  nand g1259 (n_1429, n_479, n_481);
  nand g1260 (n_499, n_1427, n_1428, n_1429);
  xor g1261 (n_1430, n_482, n_483);
  xor g1262 (n_488, n_1430, n_484);
  nand g1263 (n_1431, n_482, n_483);
  nand g1264 (n_1432, n_484, n_483);
  nand g1265 (n_1433, n_482, n_484);
  nand g1266 (n_501, n_1431, n_1432, n_1433);
  xor g1267 (n_1434, n_485, n_486);
  xor g1268 (n_489, n_1434, n_487);
  nand g1269 (n_1435, n_485, n_486);
  nand g1270 (n_1436, n_487, n_486);
  nand g1271 (n_1437, n_485, n_487);
  nand g1272 (n_504, n_1435, n_1436, n_1437);
  xor g1273 (n_1438, n_488, n_489);
  xor g1274 (n_143, n_1438, n_490);
  nand g1275 (n_1439, n_488, n_489);
  nand g1276 (n_1440, n_490, n_489);
  nand g1277 (n_1441, n_488, n_490);
  nand g1278 (n_78, n_1439, n_1440, n_1441);
  xor g1279 (n_1442, A[31], A[29]);
  xor g1280 (n_495, n_1442, A[25]);
  nand g1281 (n_1443, A[31], A[29]);
  nand g1282 (n_1444, A[25], A[29]);
  nand g1283 (n_1445, A[31], A[25]);
  nand g1284 (n_505, n_1443, n_1444, n_1445);
  xor g1285 (n_1446, A[17], A[15]);
  xor g1286 (n_496, n_1446, A[23]);
  nand g1288 (n_1448, A[23], A[15]);
  nand g1290 (n_506, n_1004, n_1448, n_1189);
  xor g1291 (n_1450, A[13], A[27]);
  xor g1292 (n_494, n_1450, A[21]);
  nand g1293 (n_1451, A[13], A[27]);
  nand g1296 (n_507, n_1451, n_1317, n_1384);
  xor g1297 (n_1454, A[19], n_491);
  xor g1298 (n_498, n_1454, n_492);
  nand g1299 (n_1455, A[19], n_491);
  nand g1300 (n_1456, n_492, n_491);
  nand g1301 (n_1457, A[19], n_492);
  nand g1302 (n_511, n_1455, n_1456, n_1457);
  xor g1303 (n_1458, n_493, n_494);
  xor g1304 (n_500, n_1458, n_495);
  nand g1305 (n_1459, n_493, n_494);
  nand g1306 (n_1460, n_495, n_494);
  nand g1307 (n_1461, n_493, n_495);
  nand g1308 (n_513, n_1459, n_1460, n_1461);
  xor g1309 (n_1462, n_496, n_497);
  xor g1310 (n_502, n_1462, n_498);
  nand g1311 (n_1463, n_496, n_497);
  nand g1312 (n_1464, n_498, n_497);
  nand g1313 (n_1465, n_496, n_498);
  nand g1314 (n_515, n_1463, n_1464, n_1465);
  xor g1315 (n_1466, n_499, n_500);
  xor g1316 (n_503, n_1466, n_501);
  nand g1317 (n_1467, n_499, n_500);
  nand g1318 (n_1468, n_501, n_500);
  nand g1319 (n_1469, n_499, n_501);
  nand g1320 (n_518, n_1467, n_1468, n_1469);
  xor g1321 (n_1470, n_502, n_503);
  xor g1322 (n_142, n_1470, n_504);
  nand g1323 (n_1471, n_502, n_503);
  nand g1324 (n_1472, n_504, n_503);
  nand g1325 (n_1473, n_502, n_504);
  nand g1326 (n_77, n_1471, n_1472, n_1473);
  xor g1327 (n_1474, A[32], A[30]);
  xor g1328 (n_509, n_1474, A[26]);
  nand g1329 (n_1475, A[32], A[30]);
  nand g1330 (n_1476, A[26], A[30]);
  nand g1331 (n_1477, A[32], A[26]);
  nand g1332 (n_519, n_1475, n_1476, n_1477);
  xor g1334 (n_510, n_317, A[24]);
  nand g1336 (n_1480, A[24], A[16]);
  xor g1339 (n_1482, A[14], A[28]);
  xor g1340 (n_508, n_1482, A[22]);
  nand g1341 (n_1483, A[14], A[28]);
  nand g1344 (n_521, n_1483, n_1349, n_1416);
  xor g1345 (n_1486, A[20], n_505);
  xor g1346 (n_512, n_1486, n_506);
  nand g1347 (n_1487, A[20], n_505);
  nand g1348 (n_1488, n_506, n_505);
  nand g1349 (n_1489, A[20], n_506);
  nand g1350 (n_525, n_1487, n_1488, n_1489);
  xor g1351 (n_1490, n_507, n_508);
  xor g1352 (n_514, n_1490, n_509);
  nand g1353 (n_1491, n_507, n_508);
  nand g1354 (n_1492, n_509, n_508);
  nand g1355 (n_1493, n_507, n_509);
  nand g1356 (n_527, n_1491, n_1492, n_1493);
  xor g1357 (n_1494, n_510, n_511);
  xor g1358 (n_516, n_1494, n_512);
  nand g1359 (n_1495, n_510, n_511);
  nand g1360 (n_1496, n_512, n_511);
  nand g1361 (n_1497, n_510, n_512);
  nand g1362 (n_529, n_1495, n_1496, n_1497);
  xor g1363 (n_1498, n_513, n_514);
  xor g1364 (n_517, n_1498, n_515);
  nand g1365 (n_1499, n_513, n_514);
  nand g1366 (n_1500, n_515, n_514);
  nand g1367 (n_1501, n_513, n_515);
  nand g1368 (n_532, n_1499, n_1500, n_1501);
  xor g1369 (n_1502, n_516, n_517);
  xor g1370 (n_141, n_1502, n_518);
  nand g1371 (n_1503, n_516, n_517);
  nand g1372 (n_1504, n_518, n_517);
  nand g1373 (n_1505, n_516, n_518);
  nand g1374 (n_76, n_1503, n_1504, n_1505);
  xor g1375 (n_1506, A[33], A[31]);
  xor g1376 (n_523, n_1506, A[27]);
  nand g1377 (n_1507, A[33], A[31]);
  nand g1378 (n_1508, A[27], A[31]);
  nand g1379 (n_1509, A[33], A[27]);
  nand g1380 (n_533, n_1507, n_1508, n_1509);
  xor g1381 (n_1510, A[19], A[17]);
  xor g1382 (n_524, n_1510, A[25]);
  nand g1383 (n_1511, A[19], A[17]);
  nand g1384 (n_1512, A[25], A[17]);
  nand g1386 (n_534, n_1511, n_1512, n_1253);
  xor g1387 (n_1514, A[15], A[29]);
  xor g1388 (n_522, n_1514, A[23]);
  nand g1389 (n_1515, A[15], A[29]);
  nand g1392 (n_535, n_1515, n_1381, n_1448);
  xor g1393 (n_1518, A[21], n_519);
  xor g1394 (n_526, n_1518, n_520);
  nand g1395 (n_1519, A[21], n_519);
  nand g1396 (n_1520, n_520, n_519);
  nand g1397 (n_1521, A[21], n_520);
  nand g1398 (n_539, n_1519, n_1520, n_1521);
  xor g1399 (n_1522, n_521, n_522);
  xor g1400 (n_528, n_1522, n_523);
  nand g1401 (n_1523, n_521, n_522);
  nand g1402 (n_1524, n_523, n_522);
  nand g1403 (n_1525, n_521, n_523);
  nand g1404 (n_541, n_1523, n_1524, n_1525);
  xor g1405 (n_1526, n_524, n_525);
  xor g1406 (n_530, n_1526, n_526);
  nand g1407 (n_1527, n_524, n_525);
  nand g1408 (n_1528, n_526, n_525);
  nand g1409 (n_1529, n_524, n_526);
  nand g1410 (n_543, n_1527, n_1528, n_1529);
  xor g1411 (n_1530, n_527, n_528);
  xor g1412 (n_531, n_1530, n_529);
  nand g1413 (n_1531, n_527, n_528);
  nand g1414 (n_1532, n_529, n_528);
  nand g1415 (n_1533, n_527, n_529);
  nand g1416 (n_546, n_1531, n_1532, n_1533);
  xor g1417 (n_1534, n_530, n_531);
  xor g1418 (n_140, n_1534, n_532);
  nand g1419 (n_1535, n_530, n_531);
  nand g1420 (n_1536, n_532, n_531);
  nand g1421 (n_1537, n_530, n_532);
  nand g1422 (n_75, n_1535, n_1536, n_1537);
  xor g1423 (n_1538, A[34], A[32]);
  xor g1424 (n_537, n_1538, A[28]);
  nand g1425 (n_1539, A[34], A[32]);
  nand g1426 (n_1540, A[28], A[32]);
  nand g1427 (n_1541, A[34], A[28]);
  nand g1428 (n_547, n_1539, n_1540, n_1541);
  xor g1430 (n_538, n_1090, A[26]);
  nand g1432 (n_1544, A[26], A[18]);
  nand g1434 (n_548, n_1091, n_1544, n_1285);
  xor g1435 (n_1546, A[16], A[30]);
  xor g1436 (n_536, n_1546, A[24]);
  nand g1437 (n_1547, A[16], A[30]);
  nand g1440 (n_549, n_1547, n_1413, n_1480);
  xor g1441 (n_1550, A[22], n_533);
  xor g1442 (n_540, n_1550, n_534);
  nand g1443 (n_1551, A[22], n_533);
  nand g1444 (n_1552, n_534, n_533);
  nand g1445 (n_1553, A[22], n_534);
  nand g1446 (n_553, n_1551, n_1552, n_1553);
  xor g1447 (n_1554, n_535, n_536);
  xor g1448 (n_542, n_1554, n_537);
  nand g1449 (n_1555, n_535, n_536);
  nand g1450 (n_1556, n_537, n_536);
  nand g1451 (n_1557, n_535, n_537);
  nand g1452 (n_555, n_1555, n_1556, n_1557);
  xor g1453 (n_1558, n_538, n_539);
  xor g1454 (n_544, n_1558, n_540);
  nand g1455 (n_1559, n_538, n_539);
  nand g1456 (n_1560, n_540, n_539);
  nand g1457 (n_1561, n_538, n_540);
  nand g1458 (n_557, n_1559, n_1560, n_1561);
  xor g1459 (n_1562, n_541, n_542);
  xor g1460 (n_545, n_1562, n_543);
  nand g1461 (n_1563, n_541, n_542);
  nand g1462 (n_1564, n_543, n_542);
  nand g1463 (n_1565, n_541, n_543);
  nand g1464 (n_560, n_1563, n_1564, n_1565);
  xor g1465 (n_1566, n_544, n_545);
  xor g1466 (n_139, n_1566, n_546);
  nand g1467 (n_1567, n_544, n_545);
  nand g1468 (n_1568, n_546, n_545);
  nand g1469 (n_1569, n_544, n_546);
  nand g1470 (n_74, n_1567, n_1568, n_1569);
  xor g1471 (n_1570, A[35], A[33]);
  xor g1472 (n_551, n_1570, A[29]);
  nand g1473 (n_1571, A[35], A[33]);
  nand g1474 (n_1572, A[29], A[33]);
  nand g1475 (n_1573, A[35], A[29]);
  nand g1476 (n_561, n_1571, n_1572, n_1573);
  xor g1478 (n_552, n_1122, A[27]);
  nand g1480 (n_1576, A[27], A[19]);
  nand g1482 (n_562, n_1123, n_1576, n_1317);
  xor g1483 (n_1578, A[17], A[31]);
  xor g1484 (n_550, n_1578, A[25]);
  nand g1485 (n_1579, A[17], A[31]);
  nand g1488 (n_563, n_1579, n_1445, n_1512);
  xor g1489 (n_1582, A[23], n_547);
  xor g1490 (n_554, n_1582, n_548);
  nand g1491 (n_1583, A[23], n_547);
  nand g1492 (n_1584, n_548, n_547);
  nand g1493 (n_1585, A[23], n_548);
  nand g1494 (n_567, n_1583, n_1584, n_1585);
  xor g1495 (n_1586, n_549, n_550);
  xor g1496 (n_556, n_1586, n_551);
  nand g1497 (n_1587, n_549, n_550);
  nand g1498 (n_1588, n_551, n_550);
  nand g1499 (n_1589, n_549, n_551);
  nand g1500 (n_569, n_1587, n_1588, n_1589);
  xor g1501 (n_1590, n_552, n_553);
  xor g1502 (n_558, n_1590, n_554);
  nand g1503 (n_1591, n_552, n_553);
  nand g1504 (n_1592, n_554, n_553);
  nand g1505 (n_1593, n_552, n_554);
  nand g1506 (n_571, n_1591, n_1592, n_1593);
  xor g1507 (n_1594, n_555, n_556);
  xor g1508 (n_559, n_1594, n_557);
  nand g1509 (n_1595, n_555, n_556);
  nand g1510 (n_1596, n_557, n_556);
  nand g1511 (n_1597, n_555, n_557);
  nand g1512 (n_574, n_1595, n_1596, n_1597);
  xor g1513 (n_1598, n_558, n_559);
  xor g1514 (n_138, n_1598, n_560);
  nand g1515 (n_1599, n_558, n_559);
  nand g1516 (n_1600, n_560, n_559);
  nand g1517 (n_1601, n_558, n_560);
  nand g1518 (n_73, n_1599, n_1600, n_1601);
  xor g1519 (n_1602, A[36], A[34]);
  xor g1520 (n_565, n_1602, A[30]);
  nand g1521 (n_1603, A[36], A[34]);
  nand g1522 (n_1604, A[30], A[34]);
  nand g1523 (n_1605, A[36], A[30]);
  nand g1524 (n_575, n_1603, n_1604, n_1605);
  xor g1526 (n_566, n_1154, A[28]);
  nand g1528 (n_1608, A[28], A[20]);
  nand g1530 (n_576, n_1155, n_1608, n_1349);
  xor g1531 (n_1610, A[18], A[32]);
  xor g1532 (n_564, n_1610, A[26]);
  nand g1533 (n_1611, A[18], A[32]);
  nand g1536 (n_577, n_1611, n_1477, n_1544);
  xor g1537 (n_1614, A[24], n_561);
  xor g1538 (n_568, n_1614, n_562);
  nand g1539 (n_1615, A[24], n_561);
  nand g1540 (n_1616, n_562, n_561);
  nand g1541 (n_1617, A[24], n_562);
  nand g1542 (n_581, n_1615, n_1616, n_1617);
  xor g1543 (n_1618, n_563, n_564);
  xor g1544 (n_570, n_1618, n_565);
  nand g1545 (n_1619, n_563, n_564);
  nand g1546 (n_1620, n_565, n_564);
  nand g1547 (n_1621, n_563, n_565);
  nand g1548 (n_583, n_1619, n_1620, n_1621);
  xor g1549 (n_1622, n_566, n_567);
  xor g1550 (n_572, n_1622, n_568);
  nand g1551 (n_1623, n_566, n_567);
  nand g1552 (n_1624, n_568, n_567);
  nand g1553 (n_1625, n_566, n_568);
  nand g1554 (n_585, n_1623, n_1624, n_1625);
  xor g1555 (n_1626, n_569, n_570);
  xor g1556 (n_573, n_1626, n_571);
  nand g1557 (n_1627, n_569, n_570);
  nand g1558 (n_1628, n_571, n_570);
  nand g1559 (n_1629, n_569, n_571);
  nand g1560 (n_588, n_1627, n_1628, n_1629);
  xor g1561 (n_1630, n_572, n_573);
  xor g1562 (n_137, n_1630, n_574);
  nand g1563 (n_1631, n_572, n_573);
  nand g1564 (n_1632, n_574, n_573);
  nand g1565 (n_1633, n_572, n_574);
  nand g1566 (n_72, n_1631, n_1632, n_1633);
  xor g1567 (n_1634, A[37], A[35]);
  xor g1568 (n_579, n_1634, A[31]);
  nand g1569 (n_1635, A[37], A[35]);
  nand g1570 (n_1636, A[31], A[35]);
  nand g1571 (n_1637, A[37], A[31]);
  nand g1572 (n_589, n_1635, n_1636, n_1637);
  xor g1574 (n_580, n_1186, A[29]);
  nand g1576 (n_1640, A[29], A[21]);
  nand g1578 (n_590, n_1187, n_1640, n_1381);
  xor g1579 (n_1642, A[19], A[33]);
  xor g1580 (n_578, n_1642, A[27]);
  nand g1581 (n_1643, A[19], A[33]);
  nand g1584 (n_591, n_1643, n_1509, n_1576);
  xor g1585 (n_1646, A[25], n_575);
  xor g1586 (n_582, n_1646, n_576);
  nand g1587 (n_1647, A[25], n_575);
  nand g1588 (n_1648, n_576, n_575);
  nand g1589 (n_1649, A[25], n_576);
  nand g1590 (n_595, n_1647, n_1648, n_1649);
  xor g1591 (n_1650, n_577, n_578);
  xor g1592 (n_584, n_1650, n_579);
  nand g1593 (n_1651, n_577, n_578);
  nand g1594 (n_1652, n_579, n_578);
  nand g1595 (n_1653, n_577, n_579);
  nand g1596 (n_597, n_1651, n_1652, n_1653);
  xor g1597 (n_1654, n_580, n_581);
  xor g1598 (n_586, n_1654, n_582);
  nand g1599 (n_1655, n_580, n_581);
  nand g1600 (n_1656, n_582, n_581);
  nand g1601 (n_1657, n_580, n_582);
  nand g1602 (n_599, n_1655, n_1656, n_1657);
  xor g1603 (n_1658, n_583, n_584);
  xor g1604 (n_587, n_1658, n_585);
  nand g1605 (n_1659, n_583, n_584);
  nand g1606 (n_1660, n_585, n_584);
  nand g1607 (n_1661, n_583, n_585);
  nand g1608 (n_602, n_1659, n_1660, n_1661);
  xor g1609 (n_1662, n_586, n_587);
  xor g1610 (n_136, n_1662, n_588);
  nand g1611 (n_1663, n_586, n_587);
  nand g1612 (n_1664, n_588, n_587);
  nand g1613 (n_1665, n_586, n_588);
  nand g1614 (n_71, n_1663, n_1664, n_1665);
  xor g1615 (n_1666, A[38], A[36]);
  xor g1616 (n_593, n_1666, A[32]);
  nand g1617 (n_1667, A[38], A[36]);
  nand g1618 (n_1668, A[32], A[36]);
  nand g1619 (n_1669, A[38], A[32]);
  nand g1620 (n_603, n_1667, n_1668, n_1669);
  xor g1622 (n_594, n_1218, A[30]);
  nand g1624 (n_1672, A[30], A[22]);
  nand g1626 (n_604, n_1219, n_1672, n_1413);
  xor g1627 (n_1674, A[20], A[34]);
  xor g1628 (n_592, n_1674, A[28]);
  nand g1629 (n_1675, A[20], A[34]);
  nand g1632 (n_605, n_1675, n_1541, n_1608);
  xor g1633 (n_1678, A[26], n_589);
  xor g1634 (n_596, n_1678, n_590);
  nand g1635 (n_1679, A[26], n_589);
  nand g1636 (n_1680, n_590, n_589);
  nand g1637 (n_1681, A[26], n_590);
  nand g1638 (n_609, n_1679, n_1680, n_1681);
  xor g1639 (n_1682, n_591, n_592);
  xor g1640 (n_598, n_1682, n_593);
  nand g1641 (n_1683, n_591, n_592);
  nand g1642 (n_1684, n_593, n_592);
  nand g1643 (n_1685, n_591, n_593);
  nand g1644 (n_611, n_1683, n_1684, n_1685);
  xor g1645 (n_1686, n_594, n_595);
  xor g1646 (n_600, n_1686, n_596);
  nand g1647 (n_1687, n_594, n_595);
  nand g1648 (n_1688, n_596, n_595);
  nand g1649 (n_1689, n_594, n_596);
  nand g1650 (n_613, n_1687, n_1688, n_1689);
  xor g1651 (n_1690, n_597, n_598);
  xor g1652 (n_601, n_1690, n_599);
  nand g1653 (n_1691, n_597, n_598);
  nand g1654 (n_1692, n_599, n_598);
  nand g1655 (n_1693, n_597, n_599);
  nand g1656 (n_616, n_1691, n_1692, n_1693);
  xor g1657 (n_1694, n_600, n_601);
  xor g1658 (n_135, n_1694, n_602);
  nand g1659 (n_1695, n_600, n_601);
  nand g1660 (n_1696, n_602, n_601);
  nand g1661 (n_1697, n_600, n_602);
  nand g1662 (n_70, n_1695, n_1696, n_1697);
  xor g1663 (n_1698, A[39], A[37]);
  xor g1664 (n_607, n_1698, A[33]);
  nand g1665 (n_1699, A[39], A[37]);
  nand g1666 (n_1700, A[33], A[37]);
  nand g1667 (n_1701, A[39], A[33]);
  nand g1668 (n_617, n_1699, n_1700, n_1701);
  xor g1670 (n_608, n_1250, A[31]);
  nand g1672 (n_1704, A[31], A[23]);
  nand g1674 (n_618, n_1251, n_1704, n_1445);
  xor g1675 (n_1706, A[21], A[35]);
  xor g1676 (n_606, n_1706, A[29]);
  nand g1677 (n_1707, A[21], A[35]);
  nand g1680 (n_619, n_1707, n_1573, n_1640);
  xor g1681 (n_1710, A[27], n_603);
  xor g1682 (n_610, n_1710, n_604);
  nand g1683 (n_1711, A[27], n_603);
  nand g1684 (n_1712, n_604, n_603);
  nand g1685 (n_1713, A[27], n_604);
  nand g1686 (n_623, n_1711, n_1712, n_1713);
  xor g1687 (n_1714, n_605, n_606);
  xor g1688 (n_612, n_1714, n_607);
  nand g1689 (n_1715, n_605, n_606);
  nand g1690 (n_1716, n_607, n_606);
  nand g1691 (n_1717, n_605, n_607);
  nand g1692 (n_625, n_1715, n_1716, n_1717);
  xor g1693 (n_1718, n_608, n_609);
  xor g1694 (n_614, n_1718, n_610);
  nand g1695 (n_1719, n_608, n_609);
  nand g1696 (n_1720, n_610, n_609);
  nand g1697 (n_1721, n_608, n_610);
  nand g1698 (n_627, n_1719, n_1720, n_1721);
  xor g1699 (n_1722, n_611, n_612);
  xor g1700 (n_615, n_1722, n_613);
  nand g1701 (n_1723, n_611, n_612);
  nand g1702 (n_1724, n_613, n_612);
  nand g1703 (n_1725, n_611, n_613);
  nand g1704 (n_630, n_1723, n_1724, n_1725);
  xor g1705 (n_1726, n_614, n_615);
  xor g1706 (n_134, n_1726, n_616);
  nand g1707 (n_1727, n_614, n_615);
  nand g1708 (n_1728, n_616, n_615);
  nand g1709 (n_1729, n_614, n_616);
  nand g1710 (n_69, n_1727, n_1728, n_1729);
  xor g1711 (n_1730, A[40], A[38]);
  xor g1712 (n_621, n_1730, A[34]);
  nand g1713 (n_1731, A[40], A[38]);
  nand g1714 (n_1732, A[34], A[38]);
  nand g1715 (n_1733, A[40], A[34]);
  nand g1716 (n_631, n_1731, n_1732, n_1733);
  xor g1718 (n_622, n_1282, A[32]);
  nand g1720 (n_1736, A[32], A[24]);
  nand g1722 (n_632, n_1283, n_1736, n_1477);
  xor g1723 (n_1738, A[22], A[36]);
  xor g1724 (n_620, n_1738, A[30]);
  nand g1725 (n_1739, A[22], A[36]);
  nand g1728 (n_633, n_1739, n_1605, n_1672);
  xor g1729 (n_1742, A[28], n_617);
  xor g1730 (n_624, n_1742, n_618);
  nand g1731 (n_1743, A[28], n_617);
  nand g1732 (n_1744, n_618, n_617);
  nand g1733 (n_1745, A[28], n_618);
  nand g1734 (n_637, n_1743, n_1744, n_1745);
  xor g1735 (n_1746, n_619, n_620);
  xor g1736 (n_626, n_1746, n_621);
  nand g1737 (n_1747, n_619, n_620);
  nand g1738 (n_1748, n_621, n_620);
  nand g1739 (n_1749, n_619, n_621);
  nand g1740 (n_639, n_1747, n_1748, n_1749);
  xor g1741 (n_1750, n_622, n_623);
  xor g1742 (n_628, n_1750, n_624);
  nand g1743 (n_1751, n_622, n_623);
  nand g1744 (n_1752, n_624, n_623);
  nand g1745 (n_1753, n_622, n_624);
  nand g1746 (n_641, n_1751, n_1752, n_1753);
  xor g1747 (n_1754, n_625, n_626);
  xor g1748 (n_629, n_1754, n_627);
  nand g1749 (n_1755, n_625, n_626);
  nand g1750 (n_1756, n_627, n_626);
  nand g1751 (n_1757, n_625, n_627);
  nand g1752 (n_644, n_1755, n_1756, n_1757);
  xor g1753 (n_1758, n_628, n_629);
  xor g1754 (n_133, n_1758, n_630);
  nand g1755 (n_1759, n_628, n_629);
  nand g1756 (n_1760, n_630, n_629);
  nand g1757 (n_1761, n_628, n_630);
  nand g1758 (n_68, n_1759, n_1760, n_1761);
  xor g1759 (n_1762, A[41], A[39]);
  xor g1760 (n_635, n_1762, A[35]);
  nand g1761 (n_1763, A[41], A[39]);
  nand g1762 (n_1764, A[35], A[39]);
  nand g1763 (n_1765, A[41], A[35]);
  nand g1764 (n_645, n_1763, n_1764, n_1765);
  xor g1766 (n_636, n_1314, A[33]);
  nand g1768 (n_1768, A[33], A[25]);
  nand g1770 (n_646, n_1315, n_1768, n_1509);
  xor g1771 (n_1770, A[23], A[37]);
  xor g1772 (n_634, n_1770, A[31]);
  nand g1773 (n_1771, A[23], A[37]);
  nand g1776 (n_647, n_1771, n_1637, n_1704);
  xor g1777 (n_1774, A[29], n_631);
  xor g1778 (n_638, n_1774, n_632);
  nand g1779 (n_1775, A[29], n_631);
  nand g1780 (n_1776, n_632, n_631);
  nand g1781 (n_1777, A[29], n_632);
  nand g1782 (n_651, n_1775, n_1776, n_1777);
  xor g1783 (n_1778, n_633, n_634);
  xor g1784 (n_640, n_1778, n_635);
  nand g1785 (n_1779, n_633, n_634);
  nand g1786 (n_1780, n_635, n_634);
  nand g1787 (n_1781, n_633, n_635);
  nand g1788 (n_653, n_1779, n_1780, n_1781);
  xor g1789 (n_1782, n_636, n_637);
  xor g1790 (n_642, n_1782, n_638);
  nand g1791 (n_1783, n_636, n_637);
  nand g1792 (n_1784, n_638, n_637);
  nand g1793 (n_1785, n_636, n_638);
  nand g1794 (n_655, n_1783, n_1784, n_1785);
  xor g1795 (n_1786, n_639, n_640);
  xor g1796 (n_643, n_1786, n_641);
  nand g1797 (n_1787, n_639, n_640);
  nand g1798 (n_1788, n_641, n_640);
  nand g1799 (n_1789, n_639, n_641);
  nand g1800 (n_658, n_1787, n_1788, n_1789);
  xor g1801 (n_1790, n_642, n_643);
  xor g1802 (n_132, n_1790, n_644);
  nand g1803 (n_1791, n_642, n_643);
  nand g1804 (n_1792, n_644, n_643);
  nand g1805 (n_1793, n_642, n_644);
  nand g1806 (n_67, n_1791, n_1792, n_1793);
  xor g1807 (n_1794, A[42], A[40]);
  xor g1808 (n_649, n_1794, A[36]);
  nand g1809 (n_1795, A[42], A[40]);
  nand g1810 (n_1796, A[36], A[40]);
  nand g1811 (n_1797, A[42], A[36]);
  nand g1812 (n_659, n_1795, n_1796, n_1797);
  xor g1814 (n_650, n_1346, A[34]);
  nand g1816 (n_1800, A[34], A[26]);
  nand g1818 (n_660, n_1347, n_1800, n_1541);
  xor g1819 (n_1802, A[24], A[38]);
  xor g1820 (n_648, n_1802, A[32]);
  nand g1821 (n_1803, A[24], A[38]);
  nand g1824 (n_661, n_1803, n_1669, n_1736);
  xor g1825 (n_1806, A[30], n_645);
  xor g1826 (n_652, n_1806, n_646);
  nand g1827 (n_1807, A[30], n_645);
  nand g1828 (n_1808, n_646, n_645);
  nand g1829 (n_1809, A[30], n_646);
  nand g1830 (n_665, n_1807, n_1808, n_1809);
  xor g1831 (n_1810, n_647, n_648);
  xor g1832 (n_654, n_1810, n_649);
  nand g1833 (n_1811, n_647, n_648);
  nand g1834 (n_1812, n_649, n_648);
  nand g1835 (n_1813, n_647, n_649);
  nand g1836 (n_667, n_1811, n_1812, n_1813);
  xor g1837 (n_1814, n_650, n_651);
  xor g1838 (n_656, n_1814, n_652);
  nand g1839 (n_1815, n_650, n_651);
  nand g1840 (n_1816, n_652, n_651);
  nand g1841 (n_1817, n_650, n_652);
  nand g1842 (n_669, n_1815, n_1816, n_1817);
  xor g1843 (n_1818, n_653, n_654);
  xor g1844 (n_657, n_1818, n_655);
  nand g1845 (n_1819, n_653, n_654);
  nand g1846 (n_1820, n_655, n_654);
  nand g1847 (n_1821, n_653, n_655);
  nand g1848 (n_672, n_1819, n_1820, n_1821);
  xor g1849 (n_1822, n_656, n_657);
  xor g1850 (n_131, n_1822, n_658);
  nand g1851 (n_1823, n_656, n_657);
  nand g1852 (n_1824, n_658, n_657);
  nand g1853 (n_1825, n_656, n_658);
  nand g1854 (n_66, n_1823, n_1824, n_1825);
  xor g1855 (n_1826, A[43], A[41]);
  xor g1856 (n_663, n_1826, A[37]);
  nand g1857 (n_1827, A[43], A[41]);
  nand g1858 (n_1828, A[37], A[41]);
  nand g1859 (n_1829, A[43], A[37]);
  nand g1860 (n_676, n_1827, n_1828, n_1829);
  xor g1862 (n_664, n_1378, A[35]);
  nand g1864 (n_1832, A[35], A[27]);
  nand g1866 (n_677, n_1379, n_1832, n_1573);
  xor g1867 (n_1834, A[25], A[39]);
  xor g1868 (n_662, n_1834, A[33]);
  nand g1869 (n_1835, A[25], A[39]);
  nand g1872 (n_675, n_1835, n_1701, n_1768);
  xor g1873 (n_1838, A[31], n_659);
  xor g1874 (n_666, n_1838, n_660);
  nand g1875 (n_1839, A[31], n_659);
  nand g1876 (n_1840, n_660, n_659);
  nand g1877 (n_1841, A[31], n_660);
  nand g1878 (n_681, n_1839, n_1840, n_1841);
  xor g1879 (n_1842, n_661, n_662);
  xor g1880 (n_668, n_1842, n_663);
  nand g1881 (n_1843, n_661, n_662);
  nand g1882 (n_1844, n_663, n_662);
  nand g1883 (n_1845, n_661, n_663);
  nand g1884 (n_683, n_1843, n_1844, n_1845);
  xor g1885 (n_1846, n_664, n_665);
  xor g1886 (n_670, n_1846, n_666);
  nand g1887 (n_1847, n_664, n_665);
  nand g1888 (n_1848, n_666, n_665);
  nand g1889 (n_1849, n_664, n_666);
  nand g1890 (n_685, n_1847, n_1848, n_1849);
  xor g1891 (n_1850, n_667, n_668);
  xor g1892 (n_671, n_1850, n_669);
  nand g1893 (n_1851, n_667, n_668);
  nand g1894 (n_1852, n_669, n_668);
  nand g1895 (n_1853, n_667, n_669);
  nand g1896 (n_688, n_1851, n_1852, n_1853);
  xor g1897 (n_1854, n_670, n_671);
  xor g1898 (n_130, n_1854, n_672);
  nand g1899 (n_1855, n_670, n_671);
  nand g1900 (n_1856, n_672, n_671);
  nand g1901 (n_1857, n_670, n_672);
  nand g1902 (n_65, n_1855, n_1856, n_1857);
  xor g1905 (n_1858, A[44], A[38]);
  xor g1906 (n_679, n_1858, A[30]);
  nand g1907 (n_1859, A[44], A[38]);
  nand g1908 (n_1860, A[30], A[38]);
  nand g1909 (n_1861, A[44], A[30]);
  nand g1910 (n_692, n_1859, n_1860, n_1861);
  xor g1911 (n_1862, A[28], A[42]);
  xor g1912 (n_680, n_1862, A[26]);
  nand g1913 (n_1863, A[28], A[42]);
  nand g1914 (n_1864, A[26], A[42]);
  nand g1916 (n_693, n_1863, n_1864, n_1347);
  xor g1917 (n_1866, A[36], A[40]);
  xor g1918 (n_678, n_1866, A[34]);
  nand g1922 (n_694, n_1796, n_1733, n_1603);
  xor g1923 (n_1870, A[32], n_675);
  xor g1924 (n_682, n_1870, n_676);
  nand g1925 (n_1871, A[32], n_675);
  nand g1926 (n_1872, n_676, n_675);
  nand g1927 (n_1873, A[32], n_676);
  nand g1928 (n_698, n_1871, n_1872, n_1873);
  xor g1929 (n_1874, n_677, n_678);
  xor g1930 (n_684, n_1874, n_679);
  nand g1931 (n_1875, n_677, n_678);
  nand g1932 (n_1876, n_679, n_678);
  nand g1933 (n_1877, n_677, n_679);
  nand g1934 (n_700, n_1875, n_1876, n_1877);
  xor g1935 (n_1878, n_680, n_681);
  xor g1936 (n_686, n_1878, n_682);
  nand g1937 (n_1879, n_680, n_681);
  nand g1938 (n_1880, n_682, n_681);
  nand g1939 (n_1881, n_680, n_682);
  nand g1940 (n_703, n_1879, n_1880, n_1881);
  xor g1941 (n_1882, n_683, n_684);
  xor g1942 (n_687, n_1882, n_685);
  nand g1943 (n_1883, n_683, n_684);
  nand g1944 (n_1884, n_685, n_684);
  nand g1945 (n_1885, n_683, n_685);
  nand g1946 (n_705, n_1883, n_1884, n_1885);
  xor g1947 (n_1886, n_686, n_687);
  xor g1948 (n_129, n_1886, n_688);
  nand g1949 (n_1887, n_686, n_687);
  nand g1950 (n_1888, n_688, n_687);
  nand g1951 (n_1889, n_686, n_688);
  nand g1952 (n_64, n_1887, n_1888, n_1889);
  xor g1955 (n_1890, A[37], A[29]);
  xor g1956 (n_696, n_1890, A[27]);
  nand g1957 (n_1891, A[37], A[29]);
  nand g1959 (n_1893, A[37], A[27]);
  nand g1960 (n_707, n_1891, n_1379, n_1893);
  xor g1961 (n_1894, A[43], A[35]);
  xor g1962 (n_697, n_1894, A[41]);
  nand g1963 (n_1895, A[43], A[35]);
  nand g1966 (n_709, n_1895, n_1765, n_1827);
  xor g1967 (n_1898, A[39], A[33]);
  xor g1968 (n_695, n_1898, A[31]);
  nand g1971 (n_1901, A[39], A[31]);
  nand g1972 (n_708, n_1701, n_1507, n_1901);
  xor g1973 (n_1902, A[44], n_692);
  xor g1974 (n_699, n_1902, n_693);
  nand g1975 (n_1903, A[44], n_692);
  nand g1976 (n_1904, n_693, n_692);
  nand g1977 (n_1905, A[44], n_693);
  nand g1978 (n_713, n_1903, n_1904, n_1905);
  xor g1979 (n_1906, n_694, n_695);
  xor g1980 (n_701, n_1906, n_696);
  nand g1981 (n_1907, n_694, n_695);
  nand g1982 (n_1908, n_696, n_695);
  nand g1983 (n_1909, n_694, n_696);
  nand g1984 (n_715, n_1907, n_1908, n_1909);
  xor g1985 (n_1910, n_697, n_698);
  xor g1986 (n_702, n_1910, n_699);
  nand g1987 (n_1911, n_697, n_698);
  nand g1988 (n_1912, n_699, n_698);
  nand g1989 (n_1913, n_697, n_699);
  nand g1990 (n_718, n_1911, n_1912, n_1913);
  xor g1991 (n_1914, n_700, n_701);
  xor g1992 (n_704, n_1914, n_702);
  nand g1993 (n_1915, n_700, n_701);
  nand g1994 (n_1916, n_702, n_701);
  nand g1995 (n_1917, n_700, n_702);
  nand g1996 (n_720, n_1915, n_1916, n_1917);
  xor g1997 (n_1918, n_703, n_704);
  xor g1998 (n_128, n_1918, n_705);
  nand g1999 (n_1919, n_703, n_704);
  nand g2000 (n_1920, n_705, n_704);
  nand g2001 (n_1921, n_703, n_705);
  nand g2002 (n_63, n_1919, n_1920, n_1921);
  xor g2004 (n_711, n_1922, A[38]);
  nand g2006 (n_1924, A[38], A[42]);
  nand g2008 (n_723, n_1923, n_1924, n_1925);
  xor g2010 (n_712, n_1410, A[36]);
  nand g2012 (n_1928, A[36], A[28]);
  nand g2014 (n_724, n_1411, n_1928, n_1605);
  xor g2015 (n_1930, A[40], A[34]);
  xor g2016 (n_710, n_1930, A[32]);
  nand g2019 (n_1933, A[40], A[32]);
  nand g2020 (n_725, n_1733, n_1539, n_1933);
  xor g2022 (n_714, n_1934, n_708);
  nand g2024 (n_1936, n_708, n_707);
  nand g2026 (n_729, n_1935, n_1936, n_1937);
  xor g2027 (n_1938, n_709, n_710);
  xor g2028 (n_716, n_1938, n_711);
  nand g2029 (n_1939, n_709, n_710);
  nand g2030 (n_1940, n_711, n_710);
  nand g2031 (n_1941, n_709, n_711);
  nand g2032 (n_731, n_1939, n_1940, n_1941);
  xor g2033 (n_1942, n_712, n_713);
  xor g2034 (n_717, n_1942, n_714);
  nand g2035 (n_1943, n_712, n_713);
  nand g2036 (n_1944, n_714, n_713);
  nand g2037 (n_1945, n_712, n_714);
  nand g2038 (n_733, n_1943, n_1944, n_1945);
  xor g2039 (n_1946, n_715, n_716);
  xor g2040 (n_719, n_1946, n_717);
  nand g2041 (n_1947, n_715, n_716);
  nand g2042 (n_1948, n_717, n_716);
  nand g2043 (n_1949, n_715, n_717);
  nand g2044 (n_735, n_1947, n_1948, n_1949);
  xor g2045 (n_1950, n_718, n_719);
  xor g2046 (n_127, n_1950, n_720);
  nand g2047 (n_1951, n_718, n_719);
  nand g2048 (n_1952, n_720, n_719);
  nand g2049 (n_1953, n_718, n_720);
  nand g2050 (n_62, n_1951, n_1952, n_1953);
  xor g2053 (n_1954, A[41], A[29]);
  xor g2054 (n_727, n_1954, A[37]);
  nand g2055 (n_1955, A[41], A[29]);
  nand g2058 (n_738, n_1955, n_1891, n_1828);
  xor g2059 (n_1958, A[35], A[39]);
  xor g2060 (n_726, n_1958, A[33]);
  nand g2064 (n_737, n_1764, n_1701, n_1571);
  xor g2066 (n_728, n_1962, n_723);
  nand g2069 (n_1965, A[31], n_723);
  nand g2070 (n_742, n_1963, n_1964, n_1965);
  xor g2071 (n_1966, n_724, n_725);
  xor g2072 (n_730, n_1966, n_726);
  nand g2073 (n_1967, n_724, n_725);
  nand g2074 (n_1968, n_726, n_725);
  nand g2075 (n_1969, n_724, n_726);
  nand g2076 (n_744, n_1967, n_1968, n_1969);
  xor g2077 (n_1970, n_727, n_728);
  xor g2078 (n_732, n_1970, n_729);
  nand g2079 (n_1971, n_727, n_728);
  nand g2080 (n_1972, n_729, n_728);
  nand g2081 (n_1973, n_727, n_729);
  nand g2082 (n_745, n_1971, n_1972, n_1973);
  xor g2083 (n_1974, n_730, n_731);
  xor g2084 (n_734, n_1974, n_732);
  nand g2085 (n_1975, n_730, n_731);
  nand g2086 (n_1976, n_732, n_731);
  nand g2087 (n_1977, n_730, n_732);
  nand g2088 (n_748, n_1975, n_1976, n_1977);
  xor g2089 (n_1978, n_733, n_734);
  xor g2090 (n_126, n_1978, n_735);
  nand g2091 (n_1979, n_733, n_734);
  nand g2092 (n_1980, n_735, n_734);
  nand g2093 (n_1981, n_733, n_735);
  nand g2094 (n_61, n_1979, n_1980, n_1981);
  xor g2101 (n_1986, A[30], A[36]);
  xor g2102 (n_740, n_1986, A[40]);
  nand g2105 (n_1989, A[30], A[40]);
  nand g2106 (n_752, n_1605, n_1796, n_1989);
  xor g2108 (n_741, n_1538, A[43]);
  nand g2110 (n_1992, A[43], A[32]);
  nand g2111 (n_1993, A[34], A[43]);
  nand g2112 (n_755, n_1539, n_1992, n_1993);
  xor g2113 (n_1994, n_737, n_738);
  xor g2114 (n_743, n_1994, n_711);
  nand g2115 (n_1995, n_737, n_738);
  nand g2116 (n_1996, n_711, n_738);
  nand g2117 (n_1997, n_737, n_711);
  nand g2118 (n_757, n_1995, n_1996, n_1997);
  xor g2119 (n_1998, n_740, n_741);
  xor g2120 (n_746, n_1998, n_742);
  nand g2121 (n_1999, n_740, n_741);
  nand g2122 (n_2000, n_742, n_741);
  nand g2123 (n_2001, n_740, n_742);
  nand g2124 (n_759, n_1999, n_2000, n_2001);
  xor g2125 (n_2002, n_743, n_744);
  xor g2126 (n_747, n_2002, n_745);
  nand g2127 (n_2003, n_743, n_744);
  nand g2128 (n_2004, n_745, n_744);
  nand g2129 (n_2005, n_743, n_745);
  nand g2130 (n_761, n_2003, n_2004, n_2005);
  xor g2131 (n_2006, n_746, n_747);
  xor g2132 (n_125, n_2006, n_748);
  nand g2133 (n_2007, n_746, n_747);
  nand g2134 (n_2008, n_748, n_747);
  nand g2135 (n_2009, n_746, n_748);
  nand g2136 (n_124, n_2007, n_2008, n_2009);
  xor g2139 (n_2010, A[41], A[37]);
  xor g2140 (n_754, n_2010, A[35]);
  nand g2144 (n_763, n_1828, n_1635, n_1765);
  xor g2152 (n_756, n_2018, n_752);
  nand g2154 (n_2020, n_752, n_723);
  nand g2156 (n_768, n_1964, n_2020, n_2021);
  xor g2157 (n_2022, n_695, n_754);
  xor g2158 (n_758, n_2022, n_755);
  nand g2159 (n_2023, n_695, n_754);
  nand g2160 (n_2024, n_755, n_754);
  nand g2161 (n_2025, n_695, n_755);
  nand g2162 (n_769, n_2023, n_2024, n_2025);
  xor g2163 (n_2026, n_756, n_757);
  xor g2164 (n_760, n_2026, n_758);
  nand g2165 (n_2027, n_756, n_757);
  nand g2166 (n_2028, n_758, n_757);
  nand g2167 (n_2029, n_756, n_758);
  nand g2168 (n_772, n_2027, n_2028, n_2029);
  xor g2169 (n_2030, n_759, n_760);
  xor g2170 (n_60, n_2030, n_761);
  nand g2171 (n_2031, n_759, n_760);
  nand g2172 (n_2032, n_761, n_760);
  nand g2173 (n_2033, n_759, n_761);
  nand g2174 (n_59, n_2031, n_2032, n_2033);
  xor g2187 (n_2042, A[32], A[43]);
  xor g2188 (n_767, n_2042, n_763);
  nand g2190 (n_2044, n_763, A[43]);
  nand g2191 (n_2045, A[32], n_763);
  nand g2192 (n_779, n_1992, n_2044, n_2045);
  xor g2193 (n_2046, n_708, n_678);
  xor g2194 (n_770, n_2046, n_711);
  nand g2195 (n_2047, n_708, n_678);
  nand g2196 (n_2048, n_711, n_678);
  nand g2197 (n_2049, n_708, n_711);
  nand g2198 (n_780, n_2047, n_2048, n_2049);
  xor g2199 (n_2050, n_767, n_768);
  xor g2200 (n_771, n_2050, n_769);
  nand g2201 (n_2051, n_767, n_768);
  nand g2202 (n_2052, n_769, n_768);
  nand g2203 (n_2053, n_767, n_769);
  nand g2204 (n_783, n_2051, n_2052, n_2053);
  xor g2205 (n_2054, n_770, n_771);
  xor g2206 (n_123, n_2054, n_772);
  nand g2207 (n_2055, n_770, n_771);
  nand g2208 (n_2056, n_772, n_771);
  nand g2209 (n_2057, n_770, n_772);
  nand g2210 (n_58, n_2055, n_2056, n_2057);
  xor g2214 (n_777, n_1634, A[43]);
  nand g2218 (n_785, n_1635, n_1895, n_1829);
  nand g2224 (n_788, n_1701, n_2064, n_2065);
  xor g2225 (n_2066, n_694, n_723);
  xor g2226 (n_781, n_2066, n_777);
  nand g2227 (n_2067, n_694, n_723);
  nand g2228 (n_2068, n_777, n_723);
  nand g2229 (n_2069, n_694, n_777);
  nand g2230 (n_790, n_2067, n_2068, n_2069);
  xor g2231 (n_2070, n_778, n_779);
  xor g2232 (n_782, n_2070, n_780);
  nand g2233 (n_2071, n_778, n_779);
  nand g2234 (n_2072, n_780, n_779);
  nand g2235 (n_2073, n_778, n_780);
  nand g2236 (n_792, n_2071, n_2072, n_2073);
  xor g2237 (n_2074, n_781, n_782);
  xor g2238 (n_122, n_2074, n_783);
  nand g2239 (n_2075, n_781, n_782);
  nand g2240 (n_2076, n_783, n_782);
  nand g2241 (n_2077, n_781, n_783);
  nand g2242 (n_57, n_2075, n_2076, n_2077);
  xor g2255 (n_2086, A[41], n_785);
  xor g2256 (n_789, n_2086, n_678);
  nand g2257 (n_2087, A[41], n_785);
  nand g2258 (n_2088, n_678, n_785);
  nand g2259 (n_2089, A[41], n_678);
  nand g2260 (n_799, n_2087, n_2088, n_2089);
  xor g2261 (n_2090, n_711, n_788);
  xor g2262 (n_791, n_2090, n_789);
  nand g2263 (n_2091, n_711, n_788);
  nand g2264 (n_2092, n_789, n_788);
  nand g2265 (n_2093, n_711, n_789);
  nand g2266 (n_801, n_2091, n_2092, n_2093);
  xor g2267 (n_2094, n_790, n_791);
  xor g2268 (n_121, n_2094, n_792);
  nand g2269 (n_2095, n_790, n_791);
  nand g2270 (n_2096, n_792, n_791);
  nand g2271 (n_2097, n_790, n_792);
  nand g2272 (n_56, n_2095, n_2096, n_2097);
  nand g2285 (n_2105, A[39], n_694);
  nand g2286 (n_806, n_2064, n_2104, n_2105);
  xor g2287 (n_2106, n_723, n_777);
  xor g2288 (n_800, n_2106, n_798);
  nand g2290 (n_2108, n_798, n_777);
  nand g2291 (n_2109, n_723, n_798);
  nand g2292 (n_808, n_2068, n_2108, n_2109);
  xor g2293 (n_2110, n_799, n_800);
  xor g2294 (n_120, n_2110, n_801);
  nand g2295 (n_2111, n_799, n_800);
  nand g2296 (n_2112, n_801, n_800);
  nand g2297 (n_2113, n_799, n_801);
  nand g2298 (n_119, n_2111, n_2112, n_2113);
  xor g2306 (n_805, n_1866, A[41]);
  nand g2308 (n_2120, A[41], A[40]);
  nand g2309 (n_2121, A[36], A[41]);
  nand g2310 (n_813, n_1796, n_2120, n_2121);
  xor g2311 (n_2122, n_785, n_711);
  xor g2312 (n_807, n_2122, n_805);
  nand g2313 (n_2123, n_785, n_711);
  nand g2314 (n_2124, n_805, n_711);
  nand g2315 (n_2125, n_785, n_805);
  nand g2316 (n_815, n_2123, n_2124, n_2125);
  xor g2317 (n_2126, n_806, n_807);
  xor g2318 (n_55, n_2126, n_808);
  nand g2319 (n_2127, n_806, n_807);
  nand g2320 (n_2128, n_808, n_807);
  nand g2321 (n_2129, n_806, n_808);
  nand g2322 (n_118, n_2127, n_2128, n_2129);
  xor g2326 (n_812, n_2010, A[39]);
  nand g2330 (n_817, n_1828, n_1763, n_1699);
  xor g2332 (n_814, n_2018, n_812);
  nand g2334 (n_2136, n_812, n_723);
  nand g2336 (n_820, n_1964, n_2136, n_2137);
  xor g2337 (n_2138, n_813, n_814);
  xor g2338 (n_54, n_2138, n_815);
  nand g2339 (n_2139, n_813, n_814);
  nand g2340 (n_2140, n_815, n_814);
  nand g2341 (n_2141, n_813, n_815);
  nand g2342 (n_117, n_2139, n_2140, n_2141);
  xor g2349 (n_2146, A[40], A[43]);
  xor g2350 (n_819, n_2146, n_817);
  nand g2351 (n_2147, A[40], A[43]);
  nand g2352 (n_2148, n_817, A[43]);
  nand g2353 (n_2149, A[40], n_817);
  nand g2354 (n_825, n_2147, n_2148, n_2149);
  xor g2355 (n_2150, n_711, n_819);
  xor g2356 (n_53, n_2150, n_820);
  nand g2357 (n_2151, n_711, n_819);
  nand g2358 (n_2152, n_820, n_819);
  nand g2359 (n_2153, n_711, n_820);
  nand g2360 (n_116, n_2151, n_2152, n_2153);
  nand g2368 (n_828, n_1763, n_2156, n_2157);
  xor g2369 (n_2158, n_723, n_824);
  xor g2370 (n_52, n_2158, n_825);
  nand g2371 (n_2159, n_723, n_824);
  nand g2372 (n_2160, n_825, n_824);
  nand g2373 (n_2161, n_723, n_825);
  nand g2374 (n_115, n_2159, n_2160, n_2161);
  xor g2376 (n_827, n_1922, A[40]);
  nand g2380 (n_831, n_1923, n_1795, n_2165);
  xor g2381 (n_2166, A[43], n_827);
  xor g2382 (n_51, n_2166, n_828);
  nand g2383 (n_2167, A[43], n_827);
  nand g2384 (n_2168, n_828, n_827);
  nand g2385 (n_2169, A[43], n_828);
  nand g2386 (n_114, n_2167, n_2168, n_2169);
  nand g2393 (n_2173, A[43], n_831);
  nand g2394 (n_113, n_2171, n_2172, n_2173);
  xor g2396 (n_49, n_1922, A[41]);
  nand g2398 (n_2176, A[41], A[42]);
  nand g2400 (n_112, n_1923, n_2176, n_2177);
  nor g11 (n_2193, A[2], A[0]);
  nor g13 (n_2189, A[1], A[3]);
  nor g15 (n_2199, A[2], n_169);
  nand g16 (n_2194, A[2], n_169);
  nor g17 (n_2195, n_104, n_168);
  nand g18 (n_2196, n_104, n_168);
  nor g19 (n_2205, n_103, n_167);
  nand g20 (n_2200, n_103, n_167);
  nor g21 (n_2201, n_102, n_166);
  nand g22 (n_2202, n_102, n_166);
  nor g23 (n_2211, n_101, n_165);
  nand g24 (n_2206, n_101, n_165);
  nor g25 (n_2207, n_100, n_164);
  nand g26 (n_2208, n_100, n_164);
  nor g27 (n_2217, n_99, n_163);
  nand g28 (n_2212, n_99, n_163);
  nor g29 (n_2213, n_98, n_162);
  nand g30 (n_2214, n_98, n_162);
  nor g31 (n_2223, n_97, n_161);
  nand g32 (n_2218, n_97, n_161);
  nor g33 (n_2219, n_96, n_160);
  nand g34 (n_2220, n_96, n_160);
  nor g35 (n_2229, n_95, n_159);
  nand g36 (n_2224, n_95, n_159);
  nor g37 (n_2225, n_94, n_158);
  nand g38 (n_2226, n_94, n_158);
  nor g39 (n_2235, n_93, n_157);
  nand g40 (n_2230, n_93, n_157);
  nor g41 (n_2231, n_92, n_156);
  nand g42 (n_2232, n_92, n_156);
  nor g43 (n_2241, n_91, n_155);
  nand g44 (n_2236, n_91, n_155);
  nor g45 (n_2237, n_90, n_154);
  nand g46 (n_2238, n_90, n_154);
  nor g47 (n_2247, n_89, n_153);
  nand g48 (n_2242, n_89, n_153);
  nor g49 (n_2243, n_88, n_152);
  nand g50 (n_2244, n_88, n_152);
  nor g51 (n_2253, n_87, n_151);
  nand g52 (n_2248, n_87, n_151);
  nor g53 (n_2249, n_86, n_150);
  nand g54 (n_2250, n_86, n_150);
  nor g55 (n_2259, n_85, n_149);
  nand g56 (n_2254, n_85, n_149);
  nor g57 (n_2255, n_84, n_148);
  nand g58 (n_2256, n_84, n_148);
  nor g59 (n_2265, n_83, n_147);
  nand g60 (n_2260, n_83, n_147);
  nor g61 (n_2261, n_82, n_146);
  nand g62 (n_2262, n_82, n_146);
  nor g63 (n_2271, n_81, n_145);
  nand g64 (n_2266, n_81, n_145);
  nor g65 (n_2267, n_80, n_144);
  nand g66 (n_2268, n_80, n_144);
  nor g67 (n_2277, n_79, n_143);
  nand g68 (n_2272, n_79, n_143);
  nor g69 (n_2273, n_78, n_142);
  nand g70 (n_2274, n_78, n_142);
  nor g71 (n_2283, n_77, n_141);
  nand g72 (n_2278, n_77, n_141);
  nor g73 (n_2279, n_76, n_140);
  nand g74 (n_2280, n_76, n_140);
  nor g75 (n_2289, n_75, n_139);
  nand g76 (n_2284, n_75, n_139);
  nor g77 (n_2285, n_74, n_138);
  nand g78 (n_2286, n_74, n_138);
  nor g79 (n_2295, n_73, n_137);
  nand g80 (n_2290, n_73, n_137);
  nor g81 (n_2291, n_72, n_136);
  nand g82 (n_2292, n_72, n_136);
  nor g83 (n_2301, n_71, n_135);
  nand g84 (n_2296, n_71, n_135);
  nor g85 (n_2297, n_70, n_134);
  nand g86 (n_2298, n_70, n_134);
  nor g87 (n_2307, n_69, n_133);
  nand g88 (n_2302, n_69, n_133);
  nor g89 (n_2303, n_68, n_132);
  nand g90 (n_2304, n_68, n_132);
  nor g91 (n_2313, n_67, n_131);
  nand g92 (n_2308, n_67, n_131);
  nor g93 (n_2309, n_66, n_130);
  nand g94 (n_2310, n_66, n_130);
  nor g95 (n_2319, n_65, n_129);
  nand g96 (n_2314, n_65, n_129);
  nor g97 (n_2315, n_64, n_128);
  nand g98 (n_2316, n_64, n_128);
  nor g99 (n_2325, n_63, n_127);
  nand g100 (n_2320, n_63, n_127);
  nor g101 (n_2321, n_62, n_126);
  nand g102 (n_2322, n_62, n_126);
  nor g103 (n_2331, n_61, n_125);
  nand g104 (n_2326, n_61, n_125);
  nor g105 (n_2327, n_60, n_124);
  nand g106 (n_2328, n_60, n_124);
  nor g107 (n_2337, n_59, n_123);
  nand g108 (n_2332, n_59, n_123);
  nor g109 (n_2333, n_58, n_122);
  nand g110 (n_2334, n_58, n_122);
  nor g111 (n_2343, n_57, n_121);
  nand g112 (n_2338, n_57, n_121);
  nor g113 (n_2339, n_56, n_120);
  nand g114 (n_2340, n_56, n_120);
  nor g115 (n_2349, n_55, n_119);
  nand g116 (n_2344, n_55, n_119);
  nor g117 (n_2345, n_54, n_118);
  nand g118 (n_2346, n_54, n_118);
  nor g119 (n_2355, n_53, n_117);
  nand g120 (n_2350, n_53, n_117);
  nor g121 (n_2351, n_52, n_116);
  nand g122 (n_2352, n_52, n_116);
  nor g123 (n_2361, n_51, n_115);
  nand g124 (n_2356, n_51, n_115);
  nor g125 (n_2357, n_50, n_114);
  nand g126 (n_2358, n_50, n_114);
  nor g127 (n_2367, n_49, n_113);
  nand g128 (n_2362, n_49, n_113);
  nor g138 (n_2191, n_839, n_2189);
  nor g142 (n_2197, n_2194, n_2195);
  nor g145 (n_2381, n_2199, n_2195);
  nor g146 (n_2203, n_2200, n_2201);
  nor g149 (n_2383, n_2205, n_2201);
  nor g150 (n_2209, n_2206, n_2207);
  nor g153 (n_2391, n_2211, n_2207);
  nor g154 (n_2215, n_2212, n_2213);
  nor g157 (n_2393, n_2217, n_2213);
  nor g158 (n_2221, n_2218, n_2219);
  nor g161 (n_2401, n_2223, n_2219);
  nor g162 (n_2227, n_2224, n_2225);
  nor g165 (n_2403, n_2229, n_2225);
  nor g166 (n_2233, n_2230, n_2231);
  nor g169 (n_2411, n_2235, n_2231);
  nor g170 (n_2239, n_2236, n_2237);
  nor g173 (n_2413, n_2241, n_2237);
  nor g174 (n_2245, n_2242, n_2243);
  nor g177 (n_2421, n_2247, n_2243);
  nor g178 (n_2251, n_2248, n_2249);
  nor g181 (n_2423, n_2253, n_2249);
  nor g182 (n_2257, n_2254, n_2255);
  nor g185 (n_2431, n_2259, n_2255);
  nor g186 (n_2263, n_2260, n_2261);
  nor g189 (n_2433, n_2265, n_2261);
  nor g190 (n_2269, n_2266, n_2267);
  nor g193 (n_2441, n_2271, n_2267);
  nor g194 (n_2275, n_2272, n_2273);
  nor g197 (n_2443, n_2277, n_2273);
  nor g198 (n_2281, n_2278, n_2279);
  nor g201 (n_2451, n_2283, n_2279);
  nor g202 (n_2287, n_2284, n_2285);
  nor g205 (n_2453, n_2289, n_2285);
  nor g206 (n_2293, n_2290, n_2291);
  nor g209 (n_2461, n_2295, n_2291);
  nor g210 (n_2299, n_2296, n_2297);
  nor g213 (n_2463, n_2301, n_2297);
  nor g214 (n_2305, n_2302, n_2303);
  nor g217 (n_2471, n_2307, n_2303);
  nor g218 (n_2311, n_2308, n_2309);
  nor g221 (n_2473, n_2313, n_2309);
  nor g222 (n_2317, n_2314, n_2315);
  nor g225 (n_2481, n_2319, n_2315);
  nor g226 (n_2323, n_2320, n_2321);
  nor g229 (n_2483, n_2325, n_2321);
  nor g230 (n_2329, n_2326, n_2327);
  nor g233 (n_2491, n_2331, n_2327);
  nor g234 (n_2335, n_2332, n_2333);
  nor g237 (n_2493, n_2337, n_2333);
  nor g238 (n_2341, n_2338, n_2339);
  nor g241 (n_2501, n_2343, n_2339);
  nor g242 (n_2347, n_2344, n_2345);
  nor g245 (n_2503, n_2349, n_2345);
  nor g246 (n_2353, n_2350, n_2351);
  nor g249 (n_2511, n_2355, n_2351);
  nor g250 (n_2359, n_2356, n_2357);
  nor g253 (n_2513, n_2361, n_2357);
  nor g254 (n_2365, n_2362, n_2363);
  nor g257 (n_2521, n_2367, n_2363);
  nor g267 (n_2379, n_2205, n_2378);
  nand g276 (n_2531, n_2381, n_2383);
  nor g277 (n_2389, n_2217, n_2388);
  nand g286 (n_2538, n_2391, n_2393);
  nor g287 (n_2399, n_2229, n_2398);
  nand g296 (n_2546, n_2401, n_2403);
  nor g297 (n_2409, n_2241, n_2408);
  nand g306 (n_2553, n_2411, n_2413);
  nor g307 (n_2419, n_2253, n_2418);
  nand g316 (n_2561, n_2421, n_2423);
  nor g317 (n_2429, n_2265, n_2428);
  nand g326 (n_2568, n_2431, n_2433);
  nor g327 (n_2439, n_2277, n_2438);
  nand g336 (n_2576, n_2441, n_2443);
  nor g337 (n_2449, n_2289, n_2448);
  nand g346 (n_2583, n_2451, n_2453);
  nor g347 (n_2459, n_2301, n_2458);
  nand g2408 (n_2591, n_2461, n_2463);
  nor g2409 (n_2469, n_2313, n_2468);
  nand g2418 (n_2598, n_2471, n_2473);
  nor g2419 (n_2479, n_2325, n_2478);
  nand g2428 (n_2606, n_2481, n_2483);
  nor g2429 (n_2489, n_2337, n_2488);
  nand g2438 (n_2613, n_2491, n_2493);
  nor g2439 (n_2499, n_2349, n_2498);
  nand g2448 (n_2621, n_2501, n_2503);
  nor g2449 (n_2509, n_2361, n_2508);
  nand g2458 (n_2628, n_2511, n_2513);
  nor g2459 (n_2519, n_2371, n_2518);
  nand g2466 (n_2974, n_2194, n_2525);
  nand g2468 (n_2976, n_2378, n_2526);
  nand g2471 (n_2979, n_2529, n_2530);
  nand g2474 (n_2636, n_2533, n_2534);
  nor g2475 (n_2536, n_2223, n_2535);
  nor g2478 (n_2646, n_2223, n_2538);
  nor g2484 (n_2544, n_2542, n_2535);
  nor g2487 (n_2652, n_2538, n_2542);
  nor g2488 (n_2548, n_2546, n_2535);
  nor g2491 (n_2655, n_2538, n_2546);
  nor g2492 (n_2551, n_2247, n_2550);
  nor g2495 (n_2771, n_2247, n_2553);
  nor g2501 (n_2559, n_2557, n_2550);
  nor g2504 (n_2777, n_2553, n_2557);
  nor g2505 (n_2563, n_2561, n_2550);
  nor g2508 (n_2661, n_2553, n_2561);
  nor g2509 (n_2566, n_2271, n_2565);
  nor g2512 (n_2674, n_2271, n_2568);
  nor g2518 (n_2574, n_2572, n_2565);
  nor g2521 (n_2684, n_2568, n_2572);
  nor g2522 (n_2578, n_2576, n_2565);
  nor g2525 (n_2689, n_2568, n_2576);
  nor g2526 (n_2581, n_2295, n_2580);
  nor g2529 (n_2882, n_2295, n_2583);
  nor g2535 (n_2589, n_2587, n_2580);
  nor g2538 (n_2888, n_2583, n_2587);
  nor g2539 (n_2593, n_2591, n_2580);
  nor g2542 (n_2697, n_2583, n_2591);
  nor g2543 (n_2596, n_2319, n_2595);
  nor g2546 (n_2710, n_2319, n_2598);
  nor g2552 (n_2604, n_2602, n_2595);
  nor g2555 (n_2720, n_2598, n_2602);
  nor g2556 (n_2608, n_2606, n_2595);
  nor g2559 (n_2725, n_2598, n_2606);
  nor g2560 (n_2611, n_2343, n_2610);
  nor g2563 (n_2826, n_2343, n_2613);
  nor g2569 (n_2619, n_2617, n_2610);
  nor g2572 (n_2836, n_2613, n_2617);
  nor g2573 (n_2623, n_2621, n_2610);
  nor g2576 (n_2733, n_2613, n_2621);
  nor g2577 (n_2626, n_2367, n_2625);
  nor g2580 (n_2746, n_2367, n_2628);
  nor g2586 (n_2634, n_2632, n_2625);
  nor g2589 (n_2756, n_2628, n_2632);
  nand g2592 (n_2983, n_2206, n_2638);
  nand g2593 (n_2639, n_2391, n_2636);
  nand g2594 (n_2985, n_2388, n_2639);
  nand g2597 (n_2988, n_2642, n_2643);
  nand g2600 (n_2991, n_2535, n_2645);
  nand g2601 (n_2648, n_2646, n_2636);
  nand g2602 (n_2994, n_2647, n_2648);
  nand g2603 (n_2651, n_2649, n_2636);
  nand g2604 (n_2996, n_2650, n_2651);
  nand g2605 (n_2654, n_2652, n_2636);
  nand g2606 (n_2999, n_2653, n_2654);
  nand g2607 (n_2657, n_2655, n_2636);
  nand g2608 (n_2761, n_2656, n_2657);
  nor g2609 (n_2659, n_2259, n_2658);
  nand g2618 (n_2785, n_2431, n_2661);
  nor g2619 (n_2668, n_2666, n_2658);
  nor g2624 (n_2671, n_2568, n_2658);
  nand g2633 (n_2797, n_2661, n_2674);
  nand g2638 (n_2801, n_2661, n_2679);
  nand g2643 (n_2805, n_2661, n_2684);
  nand g2648 (n_2809, n_2661, n_2689);
  nor g2649 (n_2695, n_2307, n_2694);
  nand g2658 (n_2896, n_2471, n_2697);
  nor g2659 (n_2704, n_2702, n_2694);
  nor g2664 (n_2707, n_2598, n_2694);
  nand g2673 (n_2908, n_2697, n_2710);
  nand g2678 (n_2912, n_2697, n_2715);
  nand g2683 (n_2916, n_2697, n_2720);
  nand g2688 (n_2816, n_2697, n_2725);
  nor g2689 (n_2731, n_2355, n_2730);
  nand g2698 (n_2848, n_2511, n_2733);
  nor g2699 (n_2740, n_2738, n_2730);
  nor g2704 (n_2743, n_2628, n_2730);
  nand g2713 (n_2860, n_2733, n_2746);
  nand g2718 (n_2864, n_2733, n_2751);
  nand g2723 (n_2868, n_2733, n_2756);
  nand g2726 (n_3003, n_2230, n_2763);
  nand g2727 (n_2764, n_2411, n_2761);
  nand g2728 (n_3005, n_2408, n_2764);
  nand g2731 (n_3008, n_2767, n_2768);
  nand g2734 (n_3011, n_2550, n_2770);
  nand g2735 (n_2773, n_2771, n_2761);
  nand g2736 (n_3014, n_2772, n_2773);
  nand g2737 (n_2776, n_2774, n_2761);
  nand g2738 (n_3016, n_2775, n_2776);
  nand g2739 (n_2779, n_2777, n_2761);
  nand g2740 (n_3019, n_2778, n_2779);
  nand g2741 (n_2780, n_2661, n_2761);
  nand g2742 (n_3021, n_2658, n_2780);
  nand g2745 (n_3024, n_2783, n_2784);
  nand g2748 (n_3026, n_2787, n_2788);
  nand g2751 (n_3029, n_2791, n_2792);
  nand g2754 (n_3032, n_2795, n_2796);
  nand g2757 (n_3035, n_2799, n_2800);
  nand g2760 (n_3037, n_2803, n_2804);
  nand g2763 (n_3040, n_2807, n_2808);
  nand g2766 (n_2872, n_2811, n_2812);
  nor g2767 (n_2814, n_2331, n_2813);
  nor g2770 (n_2922, n_2331, n_2816);
  nor g2776 (n_2822, n_2820, n_2813);
  nor g2779 (n_2928, n_2820, n_2816);
  nor g2780 (n_2824, n_2613, n_2813);
  nor g2783 (n_2931, n_2613, n_2816);
  nor g2804 (n_2846, n_2844, n_2813);
  nor g2807 (n_2946, n_2816, n_2844);
  nor g2808 (n_2850, n_2848, n_2813);
  nor g2811 (n_2949, n_2816, n_2848);
  nor g2812 (n_2854, n_2852, n_2813);
  nor g2815 (n_2952, n_2816, n_2852);
  nor g2816 (n_2858, n_2856, n_2813);
  nor g2819 (n_2955, n_2816, n_2856);
  nor g2820 (n_2862, n_2860, n_2813);
  nor g2823 (n_2958, n_2816, n_2860);
  nor g2824 (n_2866, n_2864, n_2813);
  nor g2827 (n_2961, n_2816, n_2864);
  nor g2828 (n_2870, n_2868, n_2813);
  nor g2831 (n_2964, n_2816, n_2868);
  nand g2834 (n_3044, n_2278, n_2874);
  nand g2835 (n_2875, n_2451, n_2872);
  nand g2836 (n_3046, n_2448, n_2875);
  nand g2839 (n_3049, n_2878, n_2879);
  nand g2842 (n_3052, n_2580, n_2881);
  nand g2843 (n_2884, n_2882, n_2872);
  nand g2844 (n_3055, n_2883, n_2884);
  nand g2845 (n_2887, n_2885, n_2872);
  nand g2846 (n_3057, n_2886, n_2887);
  nand g2847 (n_2890, n_2888, n_2872);
  nand g2848 (n_3060, n_2889, n_2890);
  nand g2849 (n_2891, n_2697, n_2872);
  nand g2850 (n_3062, n_2694, n_2891);
  nand g2853 (n_3065, n_2894, n_2895);
  nand g2856 (n_3067, n_2898, n_2899);
  nand g2859 (n_3070, n_2902, n_2903);
  nand g2862 (n_3073, n_2906, n_2907);
  nand g2865 (n_3076, n_2910, n_2911);
  nand g2868 (n_3078, n_2914, n_2915);
  nand g2871 (n_3081, n_2918, n_2919);
  nand g2874 (n_3084, n_2813, n_2921);
  nand g2875 (n_2924, n_2922, n_2872);
  nand g2876 (n_3087, n_2923, n_2924);
  nand g2877 (n_2927, n_2925, n_2872);
  nand g2878 (n_3089, n_2926, n_2927);
  nand g2879 (n_2930, n_2928, n_2872);
  nand g2880 (n_3092, n_2929, n_2930);
  nand g2881 (n_2933, n_2931, n_2872);
  nand g2882 (n_3095, n_2932, n_2933);
  nand g2883 (n_2936, n_2934, n_2872);
  nand g2884 (n_3098, n_2935, n_2936);
  nand g2885 (n_2939, n_2937, n_2872);
  nand g2886 (n_3100, n_2938, n_2939);
  nand g2887 (n_2942, n_2940, n_2872);
  nand g2888 (n_3103, n_2941, n_2942);
  nand g2889 (n_2945, n_2943, n_2872);
  nand g2890 (n_3105, n_2944, n_2945);
  nand g2891 (n_2948, n_2946, n_2872);
  nand g2892 (n_3108, n_2947, n_2948);
  nand g2893 (n_2951, n_2949, n_2872);
  nand g2894 (n_3110, n_2950, n_2951);
  nand g2895 (n_2954, n_2952, n_2872);
  nand g2896 (n_3113, n_2953, n_2954);
  nand g2897 (n_2957, n_2955, n_2872);
  nand g2898 (n_3116, n_2956, n_2957);
  nand g2899 (n_2960, n_2958, n_2872);
  nand g2900 (n_3119, n_2959, n_2960);
  nand g2901 (n_2963, n_2961, n_2872);
  nand g2902 (n_3121, n_2962, n_2963);
  nand g2903 (n_2966, n_2964, n_2872);
  nand g2904 (n_3124, n_2965, n_2966);
  xnor g2916 (Z[5], n_2974, n_2975);
  xnor g2918 (Z[6], n_2976, n_2977);
  xnor g2921 (Z[7], n_2979, n_2980);
  xnor g2923 (Z[8], n_2636, n_2981);
  xnor g2926 (Z[9], n_2983, n_2984);
  xnor g2928 (Z[10], n_2985, n_2986);
  xnor g2931 (Z[11], n_2988, n_2989);
  xnor g2934 (Z[12], n_2991, n_2992);
  xnor g2937 (Z[13], n_2994, n_2995);
  xnor g2939 (Z[14], n_2996, n_2997);
  xnor g2942 (Z[15], n_2999, n_3000);
  xnor g2944 (Z[16], n_2761, n_3001);
  xnor g2947 (Z[17], n_3003, n_3004);
  xnor g2949 (Z[18], n_3005, n_3006);
  xnor g2952 (Z[19], n_3008, n_3009);
  xnor g2955 (Z[20], n_3011, n_3012);
  xnor g2958 (Z[21], n_3014, n_3015);
  xnor g2960 (Z[22], n_3016, n_3017);
  xnor g2963 (Z[23], n_3019, n_3020);
  xnor g2965 (Z[24], n_3021, n_3022);
  xnor g2968 (Z[25], n_3024, n_3025);
  xnor g2970 (Z[26], n_3026, n_3027);
  xnor g2973 (Z[27], n_3029, n_3030);
  xnor g2976 (Z[28], n_3032, n_3033);
  xnor g2979 (Z[29], n_3035, n_3036);
  xnor g2981 (Z[30], n_3037, n_3038);
  xnor g2984 (Z[31], n_3040, n_3041);
  xnor g2986 (Z[32], n_2872, n_3042);
  xnor g2989 (Z[33], n_3044, n_3045);
  xnor g2991 (Z[34], n_3046, n_3047);
  xnor g2994 (Z[35], n_3049, n_3050);
  xnor g2997 (Z[36], n_3052, n_3053);
  xnor g3000 (Z[37], n_3055, n_3056);
  xnor g3002 (Z[38], n_3057, n_3058);
  xnor g3005 (Z[39], n_3060, n_3061);
  xnor g3007 (Z[40], n_3062, n_3063);
  xnor g3010 (Z[41], n_3065, n_3066);
  xnor g3012 (Z[42], n_3067, n_3068);
  xnor g3015 (Z[43], n_3070, n_3071);
  xnor g3018 (Z[44], n_3073, n_3074);
  xnor g3021 (Z[45], n_3076, n_3077);
  xnor g3023 (Z[46], n_3078, n_3079);
  xnor g3026 (Z[47], n_3081, n_3082);
  xnor g3029 (Z[48], n_3084, n_3085);
  xnor g3032 (Z[49], n_3087, n_3088);
  xnor g3034 (Z[50], n_3089, n_3090);
  xnor g3037 (Z[51], n_3092, n_3093);
  xnor g3040 (Z[52], n_3095, n_3096);
  xnor g3043 (Z[53], n_3098, n_3099);
  xnor g3045 (Z[54], n_3100, n_3101);
  xnor g3048 (Z[55], n_3103, n_3104);
  xnor g3050 (Z[56], n_3105, n_3106);
  xnor g3053 (Z[57], n_3108, n_3109);
  xnor g3055 (Z[58], n_3110, n_3111);
  xnor g3058 (Z[59], n_3113, n_3114);
  xnor g3061 (Z[60], n_3116, n_3117);
  xnor g3064 (Z[61], n_3119, n_3120);
  xnor g3066 (Z[62], n_3121, n_3122);
  or g3082 (n_246, wc, wc0, n_104);
  not gc0 (wc0, n_839);
  not gc (wc, n_853);
  or g3083 (n_255, wc1, wc2, n_240);
  not gc2 (wc2, n_853);
  not gc1 (wc1, n_872);
  or g3084 (n_268, wc3, n_245, n_240);
  not gc3 (wc3, n_900);
  or g3085 (n_285, wc4, wc5, n_245);
  not gc5 (wc5, n_935);
  not gc4 (wc4, n_936);
  or g3086 (n_307, wc6, wc7, n_245);
  not gc7 (wc7, n_983);
  not gc6 (wc6, n_984);
  or g3087 (n_354, wc8, wc9, n_240);
  not gc9 (wc9, n_984);
  not gc8 (wc8, n_1031);
  or g3088 (n_380, wc10, wc11, n_245);
  not gc11 (wc11, n_1160);
  not gc10 (wc10, n_1161);
  or g3089 (n_408, wc12, wc13, n_254);
  not gc13 (wc13, n_1100);
  not gc12 (wc12, n_1224);
  or g3090 (n_436, wc14, wc15, n_267);
  not gc15 (wc15, n_1164);
  not gc14 (wc14, n_1288);
  or g3091 (n_464, wc16, wc17, n_284);
  not gc17 (wc17, n_1093);
  not gc16 (wc16, n_1352);
  or g3092 (n_492, wc18, wc19, n_305);
  not gc19 (wc19, n_1157);
  not gc18 (wc18, n_1416);
  or g3093 (n_520, wc20, wc21, n_325);
  not gc21 (wc21, n_1221);
  not gc20 (wc20, n_1480);
  xnor g3094 (n_1922, A[44], A[42]);
  or g3095 (n_1923, wc22, A[44]);
  not gc22 (wc22, A[42]);
  or g3096 (n_1925, wc23, A[44]);
  not gc23 (wc23, A[38]);
  xnor g3097 (n_1962, A[43], A[31]);
  or g3098 (n_1963, wc24, A[43]);
  not gc24 (wc24, A[31]);
  xnor g3099 (n_778, n_1898, A[41]);
  or g3100 (n_2064, wc25, A[41]);
  not gc25 (wc25, A[39]);
  or g3101 (n_2065, wc26, A[41]);
  not gc26 (wc26, A[33]);
  xnor g3103 (n_824, n_1762, A[43]);
  or g3104 (n_2156, wc27, A[43]);
  not gc27 (wc27, A[39]);
  or g3105 (n_2157, wc28, A[43]);
  not gc28 (wc28, A[41]);
  or g3106 (n_2165, wc29, A[44]);
  not gc29 (wc29, A[40]);
  or g3108 (n_2171, A[41], wc30);
  not gc30 (wc30, A[43]);
  or g3109 (n_2177, wc31, A[44]);
  not gc31 (wc31, A[41]);
  and g3110 (n_2371, wc32, A[44]);
  not gc32 (wc32, A[43]);
  or g3111 (n_2368, wc33, A[44]);
  not gc33 (wc33, A[43]);
  or g3112 (n_331, wc34, wc35, n_245);
  not gc35 (wc35, n_1040);
  not gc34 (wc34, n_1041);
  or g3113 (n_2021, A[43], wc36);
  not gc36 (wc36, n_752);
  xnor g3114 (n_798, n_1762, n_694);
  or g3115 (n_2104, A[41], wc37);
  not gc37 (wc37, n_694);
  or g3116 (n_2137, A[43], wc38);
  not gc38 (wc38, n_812);
  and g3117 (n_2376, wc39, n_835);
  not gc39 (wc39, n_2191);
  or g3119 (n_2968, n_2193, wc40);
  not gc40 (wc40, n_839);
  or g3120 (n_2971, n_2189, wc41);
  not gc41 (wc41, n_835);
  xnor g3121 (n_1934, n_707, A[44]);
  or g3122 (n_1935, A[44], wc42);
  not gc42 (wc42, n_707);
  or g3123 (n_1937, A[44], wc43);
  not gc43 (wc43, n_708);
  or g3124 (n_1964, A[43], wc44);
  not gc44 (wc44, n_723);
  xnor g3125 (n_2018, n_723, A[43]);
  xnor g3126 (n_50, n_1826, n_831);
  or g3127 (n_2172, A[41], wc45);
  not gc45 (wc45, n_831);
  and g3128 (n_2363, A[43], wc46);
  not gc46 (wc46, n_112);
  or g3129 (n_2364, A[43], wc47);
  not gc47 (wc47, n_112);
  or g3130 (n_2972, wc48, n_2199);
  not gc48 (wc48, n_2194);
  or g3131 (n_3122, wc49, n_2371);
  not gc49 (wc49, n_2368);
  and g3132 (n_2378, wc50, n_2196);
  not gc50 (wc50, n_2197);
  or g3133 (n_2527, wc51, n_2205);
  not gc51 (wc51, n_2381);
  not g3134 (Z[2], n_2968);
  or g3135 (n_2975, wc52, n_2195);
  not gc52 (wc52, n_2196);
  or g3136 (n_2977, wc53, n_2205);
  not gc53 (wc53, n_2200);
  and g3137 (n_2385, wc54, n_2202);
  not gc54 (wc54, n_2203);
  or g3140 (n_2980, wc55, n_2201);
  not gc55 (wc55, n_2202);
  or g3141 (n_3120, wc56, n_2363);
  not gc56 (wc56, n_2364);
  and g3142 (n_2388, wc57, n_2208);
  not gc57 (wc57, n_2209);
  and g3143 (n_2529, wc58, n_2200);
  not gc58 (wc58, n_2379);
  and g3144 (n_2386, wc59, n_2383);
  not gc59 (wc59, n_2378);
  or g3145 (n_2525, n_2199, n_2376);
  or g3146 (n_2526, n_2376, wc60);
  not gc60 (wc60, n_2381);
  or g3147 (n_2530, n_2376, n_2527);
  xor g3148 (Z[3], n_839, n_2971);
  xor g3149 (Z[4], n_2376, n_2972);
  or g3150 (n_2981, wc61, n_2211);
  not gc61 (wc61, n_2206);
  or g3151 (n_2984, wc62, n_2207);
  not gc62 (wc62, n_2208);
  and g3152 (n_2518, n_2364, wc63);
  not gc63 (wc63, n_2365);
  and g3153 (n_2533, wc64, n_2385);
  not gc64 (wc64, n_2386);
  or g3154 (n_2640, wc65, n_2217);
  not gc65 (wc65, n_2391);
  or g3155 (n_2632, n_2371, wc66);
  not gc66 (wc66, n_2521);
  or g3156 (n_2534, n_2531, n_2376);
  or g3157 (n_2986, wc67, n_2217);
  not gc67 (wc67, n_2212);
  or g3158 (n_3114, wc68, n_2357);
  not gc68 (wc68, n_2358);
  or g3159 (n_3117, wc69, n_2367);
  not gc69 (wc69, n_2362);
  and g3160 (n_2395, wc70, n_2214);
  not gc70 (wc70, n_2215);
  and g3161 (n_2398, wc71, n_2220);
  not gc71 (wc71, n_2221);
  and g3162 (n_2515, wc72, n_2358);
  not gc72 (wc72, n_2359);
  and g3163 (n_2642, wc73, n_2212);
  not gc73 (wc73, n_2389);
  or g3164 (n_2989, wc74, n_2213);
  not gc74 (wc74, n_2214);
  or g3165 (n_2992, wc75, n_2223);
  not gc75 (wc75, n_2218);
  or g3166 (n_2995, wc76, n_2219);
  not gc76 (wc76, n_2220);
  or g3167 (n_3111, wc77, n_2361);
  not gc77 (wc77, n_2356);
  and g3168 (n_2405, wc78, n_2226);
  not gc78 (wc78, n_2227);
  and g3169 (n_2508, wc79, n_2352);
  not gc79 (wc79, n_2353);
  and g3170 (n_2396, wc80, n_2393);
  not gc80 (wc80, n_2388);
  or g3171 (n_2542, wc81, n_2229);
  not gc81 (wc81, n_2401);
  or g3172 (n_2738, wc82, n_2361);
  not gc82 (wc82, n_2511);
  and g3173 (n_2633, n_2368, wc83);
  not gc83 (wc83, n_2519);
  and g3174 (n_2649, wc84, n_2401);
  not gc84 (wc84, n_2538);
  or g3175 (n_2638, wc85, n_2211);
  not gc85 (wc85, n_2636);
  or g3176 (n_2643, n_2640, wc86);
  not gc86 (wc86, n_2636);
  or g3177 (n_2997, wc87, n_2229);
  not gc87 (wc87, n_2224);
  or g3178 (n_3000, wc88, n_2225);
  not gc88 (wc88, n_2226);
  or g3179 (n_3104, wc89, n_2345);
  not gc89 (wc89, n_2346);
  or g3180 (n_3106, wc90, n_2355);
  not gc90 (wc90, n_2350);
  or g3181 (n_3109, wc91, n_2351);
  not gc91 (wc91, n_2352);
  and g3182 (n_2408, wc92, n_2232);
  not gc92 (wc92, n_2233);
  and g3183 (n_2415, wc93, n_2238);
  not gc93 (wc93, n_2239);
  and g3184 (n_2505, wc94, n_2346);
  not gc94 (wc94, n_2347);
  and g3185 (n_2535, wc95, n_2395);
  not gc95 (wc95, n_2396);
  and g3186 (n_2543, wc96, n_2224);
  not gc96 (wc96, n_2399);
  and g3187 (n_2406, wc97, n_2403);
  not gc97 (wc97, n_2398);
  or g3188 (n_2765, wc98, n_2241);
  not gc98 (wc98, n_2411);
  and g3189 (n_2516, wc99, n_2513);
  not gc99 (wc99, n_2508);
  and g3190 (n_2751, wc100, n_2521);
  not gc100 (wc100, n_2628);
  or g3191 (n_2645, wc101, n_2538);
  not gc101 (wc101, n_2636);
  or g3192 (n_3001, wc102, n_2235);
  not gc102 (wc102, n_2230);
  or g3193 (n_3004, wc103, n_2231);
  not gc103 (wc103, n_2232);
  or g3194 (n_3006, wc104, n_2241);
  not gc104 (wc104, n_2236);
  or g3195 (n_3009, wc105, n_2237);
  not gc105 (wc105, n_2238);
  or g3196 (n_3012, wc106, n_2247);
  not gc106 (wc106, n_2242);
  or g3197 (n_3101, wc107, n_2349);
  not gc107 (wc107, n_2344);
  and g3198 (n_2418, wc108, n_2244);
  not gc108 (wc108, n_2245);
  and g3199 (n_2498, wc109, n_2340);
  not gc109 (wc109, n_2341);
  and g3200 (n_2547, wc110, n_2405);
  not gc110 (wc110, n_2406);
  and g3201 (n_2416, wc111, n_2413);
  not gc111 (wc111, n_2408);
  or g3202 (n_2557, wc112, n_2253);
  not gc112 (wc112, n_2421);
  or g3203 (n_2617, wc113, n_2349);
  not gc113 (wc113, n_2501);
  and g3204 (n_2739, wc114, n_2356);
  not gc114 (wc114, n_2509);
  and g3205 (n_2625, wc115, n_2515);
  not gc115 (wc115, n_2516);
  and g3206 (n_2540, wc116, n_2401);
  not gc116 (wc116, n_2535);
  or g3207 (n_3015, wc117, n_2243);
  not gc117 (wc117, n_2244);
  or g3208 (n_3017, wc118, n_2253);
  not gc118 (wc118, n_2248);
  or g3209 (n_3093, wc119, n_2333);
  not gc119 (wc119, n_2334);
  or g3210 (n_3096, wc120, n_2343);
  not gc120 (wc120, n_2338);
  or g3211 (n_3099, wc121, n_2339);
  not gc121 (wc121, n_2340);
  and g3212 (n_2425, wc122, n_2250);
  not gc122 (wc122, n_2251);
  and g3213 (n_2428, wc123, n_2256);
  not gc123 (wc123, n_2257);
  and g3214 (n_2435, wc124, n_2262);
  not gc124 (wc124, n_2263);
  and g3215 (n_2438, wc125, n_2268);
  not gc125 (wc125, n_2269);
  and g3216 (n_2445, wc126, n_2274);
  not gc126 (wc126, n_2275);
  and g3217 (n_2448, wc127, n_2280);
  not gc127 (wc127, n_2281);
  and g3218 (n_2455, wc128, n_2286);
  not gc128 (wc128, n_2287);
  and g3219 (n_2458, wc129, n_2292);
  not gc129 (wc129, n_2293);
  and g3220 (n_2465, wc130, n_2298);
  not gc130 (wc130, n_2299);
  and g3221 (n_2468, wc131, n_2304);
  not gc131 (wc131, n_2305);
  and g3222 (n_2475, wc132, n_2310);
  not gc132 (wc132, n_2311);
  and g3223 (n_2478, wc133, n_2316);
  not gc133 (wc133, n_2317);
  and g3224 (n_2767, wc134, n_2236);
  not gc134 (wc134, n_2409);
  and g3225 (n_2550, wc135, n_2415);
  not gc135 (wc135, n_2416);
  or g3226 (n_2666, wc136, n_2265);
  not gc136 (wc136, n_2431);
  or g3227 (n_2572, wc137, n_2277);
  not gc137 (wc137, n_2441);
  or g3228 (n_2876, wc138, n_2289);
  not gc138 (wc138, n_2451);
  or g3229 (n_2587, wc139, n_2301);
  not gc139 (wc139, n_2461);
  or g3230 (n_2702, wc140, n_2313);
  not gc140 (wc140, n_2471);
  and g3231 (n_2506, wc141, n_2503);
  not gc141 (wc141, n_2498);
  and g3232 (n_2647, wc142, n_2218);
  not gc142 (wc142, n_2536);
  and g3233 (n_2650, wc143, n_2398);
  not gc143 (wc143, n_2540);
  and g3234 (n_2653, n_2543, wc144);
  not gc144 (wc144, n_2544);
  and g3235 (n_2774, wc145, n_2421);
  not gc145 (wc145, n_2553);
  and g3236 (n_2630, wc146, n_2521);
  not gc146 (wc146, n_2625);
  or g3237 (n_3020, wc147, n_2249);
  not gc147 (wc147, n_2250);
  or g3238 (n_3022, wc148, n_2259);
  not gc148 (wc148, n_2254);
  or g3239 (n_3025, wc149, n_2255);
  not gc149 (wc149, n_2256);
  or g3240 (n_3027, wc150, n_2265);
  not gc150 (wc150, n_2260);
  or g3241 (n_3030, wc151, n_2261);
  not gc151 (wc151, n_2262);
  or g3242 (n_3033, wc152, n_2271);
  not gc152 (wc152, n_2266);
  or g3243 (n_3036, wc153, n_2267);
  not gc153 (wc153, n_2268);
  or g3244 (n_3038, wc154, n_2277);
  not gc154 (wc154, n_2272);
  or g3245 (n_3041, wc155, n_2273);
  not gc155 (wc155, n_2274);
  or g3246 (n_3042, wc156, n_2283);
  not gc156 (wc156, n_2278);
  or g3247 (n_3045, wc157, n_2279);
  not gc157 (wc157, n_2280);
  or g3248 (n_3047, wc158, n_2289);
  not gc158 (wc158, n_2284);
  or g3249 (n_3050, wc159, n_2285);
  not gc159 (wc159, n_2286);
  or g3250 (n_3053, wc160, n_2295);
  not gc160 (wc160, n_2290);
  or g3251 (n_3056, wc161, n_2291);
  not gc161 (wc161, n_2292);
  or g3252 (n_3058, wc162, n_2301);
  not gc162 (wc162, n_2296);
  or g3253 (n_3061, wc163, n_2297);
  not gc163 (wc163, n_2298);
  or g3254 (n_3063, wc164, n_2307);
  not gc164 (wc164, n_2302);
  or g3255 (n_3066, wc165, n_2303);
  not gc165 (wc165, n_2304);
  or g3256 (n_3068, wc166, n_2313);
  not gc166 (wc166, n_2308);
  or g3257 (n_3071, wc167, n_2309);
  not gc167 (wc167, n_2310);
  or g3258 (n_3074, wc168, n_2319);
  not gc168 (wc168, n_2314);
  or g3259 (n_3077, wc169, n_2315);
  not gc169 (wc169, n_2316);
  or g3260 (n_3088, wc170, n_2327);
  not gc170 (wc170, n_2328);
  and g3261 (n_2485, wc171, n_2322);
  not gc171 (wc171, n_2323);
  and g3262 (n_2495, wc172, n_2334);
  not gc172 (wc172, n_2335);
  and g3263 (n_2558, wc173, n_2248);
  not gc173 (wc173, n_2419);
  and g3264 (n_2426, wc174, n_2423);
  not gc174 (wc174, n_2418);
  and g3265 (n_2436, wc175, n_2433);
  not gc175 (wc175, n_2428);
  and g3266 (n_2446, wc176, n_2443);
  not gc176 (wc176, n_2438);
  and g3267 (n_2456, wc177, n_2453);
  not gc177 (wc177, n_2448);
  and g3268 (n_2466, wc178, n_2463);
  not gc178 (wc178, n_2458);
  and g3269 (n_2476, wc179, n_2473);
  not gc179 (wc179, n_2468);
  or g3270 (n_2602, wc180, n_2325);
  not gc180 (wc180, n_2481);
  and g3271 (n_2618, wc181, n_2344);
  not gc181 (wc181, n_2499);
  and g3272 (n_2622, wc182, n_2505);
  not gc182 (wc182, n_2506);
  and g3273 (n_2656, n_2547, wc183);
  not gc183 (wc183, n_2548);
  and g3274 (n_2555, wc184, n_2421);
  not gc184 (wc184, n_2550);
  and g3275 (n_2679, wc185, n_2441);
  not gc185 (wc185, n_2568);
  and g3276 (n_2885, wc186, n_2461);
  not gc186 (wc186, n_2583);
  and g3277 (n_2715, wc187, n_2481);
  not gc187 (wc187, n_2598);
  and g3278 (n_2748, wc188, n_2362);
  not gc188 (wc188, n_2626);
  and g3279 (n_2753, wc189, n_2518);
  not gc189 (wc189, n_2630);
  and g3280 (n_2758, n_2633, wc190);
  not gc190 (wc190, n_2634);
  or g3281 (n_3079, wc191, n_2325);
  not gc191 (wc191, n_2320);
  or g3282 (n_3082, wc192, n_2321);
  not gc192 (wc192, n_2322);
  or g3283 (n_3090, wc193, n_2337);
  not gc193 (wc193, n_2332);
  and g3284 (n_2488, wc194, n_2328);
  not gc194 (wc194, n_2329);
  and g3285 (n_2562, wc195, n_2425);
  not gc195 (wc195, n_2426);
  and g3286 (n_2667, wc196, n_2260);
  not gc196 (wc196, n_2429);
  and g3287 (n_2565, wc197, n_2435);
  not gc197 (wc197, n_2436);
  and g3288 (n_2573, wc198, n_2272);
  not gc198 (wc198, n_2439);
  and g3289 (n_2577, wc199, n_2445);
  not gc199 (wc199, n_2446);
  and g3290 (n_2878, wc200, n_2284);
  not gc200 (wc200, n_2449);
  and g3291 (n_2580, wc201, n_2455);
  not gc201 (wc201, n_2456);
  and g3292 (n_2588, wc202, n_2296);
  not gc202 (wc202, n_2459);
  and g3293 (n_2592, wc203, n_2465);
  not gc203 (wc203, n_2466);
  and g3294 (n_2703, wc204, n_2308);
  not gc204 (wc204, n_2469);
  and g3295 (n_2595, wc205, n_2475);
  not gc205 (wc205, n_2476);
  and g3296 (n_2603, wc206, n_2320);
  not gc206 (wc206, n_2479);
  and g3297 (n_2486, wc207, n_2483);
  not gc207 (wc207, n_2478);
  or g3298 (n_2820, wc208, n_2337);
  not gc208 (wc208, n_2491);
  and g3299 (n_2772, wc209, n_2242);
  not gc209 (wc209, n_2551);
  and g3300 (n_2775, wc210, n_2418);
  not gc210 (wc210, n_2555);
  or g3301 (n_2781, wc211, n_2259);
  not gc211 (wc211, n_2661);
  or g3302 (n_2789, n_2666, wc212);
  not gc212 (wc212, n_2661);
  or g3303 (n_2793, wc213, n_2568);
  not gc213 (wc213, n_2661);
  or g3304 (n_2892, wc214, n_2307);
  not gc214 (wc214, n_2697);
  or g3305 (n_2900, n_2702, wc215);
  not gc215 (wc215, n_2697);
  or g3306 (n_2904, wc216, n_2598);
  not gc216 (wc216, n_2697);
  or g3307 (n_3085, wc217, n_2331);
  not gc217 (wc217, n_2326);
  and g3308 (n_2607, wc218, n_2485);
  not gc218 (wc218, n_2486);
  and g3309 (n_2496, wc219, n_2493);
  not gc219 (wc219, n_2488);
  and g3310 (n_2778, n_2558, wc220);
  not gc220 (wc220, n_2559);
  and g3311 (n_2570, wc221, n_2441);
  not gc221 (wc221, n_2565);
  and g3312 (n_2585, wc222, n_2461);
  not gc222 (wc222, n_2580);
  and g3313 (n_2600, wc223, n_2481);
  not gc223 (wc223, n_2595);
  and g3314 (n_2831, wc224, n_2501);
  not gc224 (wc224, n_2613);
  or g3315 (n_2763, wc225, n_2235);
  not gc225 (wc225, n_2761);
  or g3316 (n_2768, n_2765, wc226);
  not gc226 (wc226, n_2761);
  or g3317 (n_2770, wc227, n_2553);
  not gc227 (wc227, n_2761);
  and g3318 (n_2821, wc228, n_2332);
  not gc228 (wc228, n_2489);
  and g3319 (n_2610, wc229, n_2495);
  not gc229 (wc229, n_2496);
  and g3320 (n_2658, n_2562, wc230);
  not gc230 (wc230, n_2563);
  and g3321 (n_2676, wc231, n_2266);
  not gc231 (wc231, n_2566);
  and g3322 (n_2681, wc232, n_2438);
  not gc232 (wc232, n_2570);
  and g3323 (n_2686, n_2573, wc233);
  not gc233 (wc233, n_2574);
  and g3324 (n_2691, n_2577, wc234);
  not gc234 (wc234, n_2578);
  and g3325 (n_2883, wc235, n_2290);
  not gc235 (wc235, n_2581);
  and g3326 (n_2886, wc236, n_2458);
  not gc236 (wc236, n_2585);
  and g3327 (n_2889, n_2588, wc237);
  not gc237 (wc237, n_2589);
  and g3328 (n_2694, n_2592, wc238);
  not gc238 (wc238, n_2593);
  and g3329 (n_2712, wc239, n_2314);
  not gc239 (wc239, n_2596);
  and g3330 (n_2717, wc240, n_2478);
  not gc240 (wc240, n_2600);
  and g3331 (n_2722, n_2603, wc241);
  not gc241 (wc241, n_2604);
  or g3332 (n_2844, wc242, n_2355);
  not gc242 (wc242, n_2733);
  or g3333 (n_2852, n_2738, wc243);
  not gc243 (wc243, n_2733);
  or g3334 (n_2856, wc244, n_2628);
  not gc244 (wc244, n_2733);
  or g3335 (n_2784, n_2781, wc245);
  not gc245 (wc245, n_2761);
  or g3336 (n_2788, n_2785, wc246);
  not gc246 (wc246, n_2761);
  or g3337 (n_2792, n_2789, wc247);
  not gc247 (wc247, n_2761);
  or g3338 (n_2796, n_2793, wc248);
  not gc248 (wc248, n_2761);
  or g3339 (n_2800, n_2797, wc249);
  not gc249 (wc249, n_2761);
  or g3340 (n_2804, n_2801, wc250);
  not gc250 (wc250, n_2761);
  or g3341 (n_2808, n_2805, wc251);
  not gc251 (wc251, n_2761);
  or g3342 (n_2812, n_2809, wc252);
  not gc252 (wc252, n_2761);
  and g3343 (n_2925, wc253, n_2491);
  not gc253 (wc253, n_2816);
  and g3344 (n_2727, n_2607, wc254);
  not gc254 (wc254, n_2608);
  and g3345 (n_2615, wc255, n_2501);
  not gc255 (wc255, n_2610);
  and g3346 (n_2664, wc256, n_2431);
  not gc256 (wc256, n_2658);
  and g3347 (n_2677, wc257, n_2674);
  not gc257 (wc257, n_2658);
  and g3348 (n_2682, wc258, n_2679);
  not gc258 (wc258, n_2658);
  and g3349 (n_2687, wc259, n_2684);
  not gc259 (wc259, n_2658);
  and g3350 (n_2692, wc260, n_2689);
  not gc260 (wc260, n_2658);
  and g3351 (n_2700, wc261, n_2471);
  not gc261 (wc261, n_2694);
  and g3352 (n_2713, wc262, n_2710);
  not gc262 (wc262, n_2694);
  and g3353 (n_2718, wc263, n_2715);
  not gc263 (wc263, n_2694);
  and g3354 (n_2723, wc264, n_2720);
  not gc264 (wc264, n_2694);
  and g3355 (n_2728, wc265, n_2725);
  not gc265 (wc265, n_2694);
  and g3356 (n_2934, wc266, n_2826);
  not gc266 (wc266, n_2816);
  and g3357 (n_2937, n_2831, wc267);
  not gc267 (wc267, n_2816);
  and g3358 (n_2940, wc268, n_2836);
  not gc268 (wc268, n_2816);
  and g3359 (n_2943, wc269, n_2733);
  not gc269 (wc269, n_2816);
  and g3360 (n_2828, wc270, n_2338);
  not gc270 (wc270, n_2611);
  and g3361 (n_2833, wc271, n_2498);
  not gc271 (wc271, n_2615);
  and g3362 (n_2838, n_2618, wc272);
  not gc272 (wc272, n_2619);
  and g3363 (n_2730, n_2622, wc273);
  not gc273 (wc273, n_2623);
  and g3364 (n_2783, wc274, n_2254);
  not gc274 (wc274, n_2659);
  and g3365 (n_2787, wc275, n_2428);
  not gc275 (wc275, n_2664);
  and g3366 (n_2791, n_2667, wc276);
  not gc276 (wc276, n_2668);
  and g3367 (n_2795, n_2565, wc277);
  not gc277 (wc277, n_2671);
  and g3368 (n_2799, wc278, n_2676);
  not gc278 (wc278, n_2677);
  and g3369 (n_2803, wc279, n_2681);
  not gc279 (wc279, n_2682);
  and g3370 (n_2807, wc280, n_2686);
  not gc280 (wc280, n_2687);
  and g3371 (n_2811, wc281, n_2691);
  not gc281 (wc281, n_2692);
  and g3372 (n_2894, wc282, n_2302);
  not gc282 (wc282, n_2695);
  and g3373 (n_2898, wc283, n_2468);
  not gc283 (wc283, n_2700);
  and g3374 (n_2902, n_2703, wc284);
  not gc284 (wc284, n_2704);
  and g3375 (n_2906, n_2595, wc285);
  not gc285 (wc285, n_2707);
  and g3376 (n_2910, wc286, n_2712);
  not gc286 (wc286, n_2713);
  and g3377 (n_2914, wc287, n_2717);
  not gc287 (wc287, n_2718);
  and g3378 (n_2918, wc288, n_2722);
  not gc288 (wc288, n_2723);
  and g3379 (n_2813, wc289, n_2727);
  not gc289 (wc289, n_2728);
  and g3380 (n_2736, wc290, n_2511);
  not gc290 (wc290, n_2730);
  and g3381 (n_2749, wc291, n_2746);
  not gc291 (wc291, n_2730);
  and g3382 (n_2754, wc292, n_2751);
  not gc292 (wc292, n_2730);
  and g3383 (n_2759, wc293, n_2756);
  not gc293 (wc293, n_2730);
  and g3384 (n_2845, wc294, n_2350);
  not gc294 (wc294, n_2731);
  and g3385 (n_2849, wc295, n_2508);
  not gc295 (wc295, n_2736);
  and g3386 (n_2853, n_2739, wc296);
  not gc296 (wc296, n_2740);
  and g3387 (n_2857, n_2625, wc297);
  not gc297 (wc297, n_2743);
  and g3388 (n_2861, wc298, n_2748);
  not gc298 (wc298, n_2749);
  and g3389 (n_2865, wc299, n_2753);
  not gc299 (wc299, n_2754);
  and g3390 (n_2869, wc300, n_2758);
  not gc300 (wc300, n_2759);
  and g3391 (n_2818, wc301, n_2491);
  not gc301 (wc301, n_2813);
  and g3392 (n_2829, wc302, n_2826);
  not gc302 (wc302, n_2813);
  and g3393 (n_2834, wc303, n_2831);
  not gc303 (wc303, n_2813);
  and g3394 (n_2839, wc304, n_2836);
  not gc304 (wc304, n_2813);
  and g3395 (n_2842, wc305, n_2733);
  not gc305 (wc305, n_2813);
  or g3396 (n_2874, wc306, n_2283);
  not gc306 (wc306, n_2872);
  or g3397 (n_2879, n_2876, wc307);
  not gc307 (wc307, n_2872);
  or g3398 (n_2881, wc308, n_2583);
  not gc308 (wc308, n_2872);
  or g3399 (n_2895, n_2892, wc309);
  not gc309 (wc309, n_2872);
  or g3400 (n_2899, wc310, n_2896);
  not gc310 (wc310, n_2872);
  or g3401 (n_2903, n_2900, wc311);
  not gc311 (wc311, n_2872);
  or g3402 (n_2907, n_2904, wc312);
  not gc312 (wc312, n_2872);
  or g3403 (n_2911, wc313, n_2908);
  not gc313 (wc313, n_2872);
  or g3404 (n_2915, wc314, n_2912);
  not gc314 (wc314, n_2872);
  or g3405 (n_2919, wc315, n_2916);
  not gc315 (wc315, n_2872);
  or g3406 (n_2921, wc316, n_2816);
  not gc316 (wc316, n_2872);
  and g3407 (n_2923, wc317, n_2326);
  not gc317 (wc317, n_2814);
  and g3408 (n_2926, wc318, n_2488);
  not gc318 (wc318, n_2818);
  and g3409 (n_2929, n_2821, wc319);
  not gc319 (wc319, n_2822);
  and g3410 (n_2932, n_2610, wc320);
  not gc320 (wc320, n_2824);
  and g3411 (n_2935, wc321, n_2828);
  not gc321 (wc321, n_2829);
  and g3412 (n_2938, wc322, n_2833);
  not gc322 (wc322, n_2834);
  and g3413 (n_2941, wc323, n_2838);
  not gc323 (wc323, n_2839);
  and g3414 (n_2944, wc324, n_2730);
  not gc324 (wc324, n_2842);
  and g3415 (n_2947, n_2845, wc325);
  not gc325 (wc325, n_2846);
  and g3416 (n_2950, n_2849, wc326);
  not gc326 (wc326, n_2850);
  and g3417 (n_2953, n_2853, wc327);
  not gc327 (wc327, n_2854);
  and g3418 (n_2956, n_2857, wc328);
  not gc328 (wc328, n_2858);
  and g3419 (n_2959, n_2861, wc329);
  not gc329 (wc329, n_2862);
  and g3420 (n_2962, n_2865, wc330);
  not gc330 (wc330, n_2866);
  and g3421 (n_2965, n_2869, wc331);
  not gc331 (wc331, n_2870);
  not g3422 (Z[63], n_3124);
endmodule

module mult_signed_const_9979_GENERIC(A, Z);
  input [44:0] A;
  output [63:0] Z;
  wire [44:0] A;
  wire [63:0] Z;
  mult_signed_const_9979_GENERIC_REAL g1(.A ({A[44:2], A[0], A[0]}), .Z
       (Z));
endmodule

