module add_signed_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [23:0] A, B;
  output [21:0] Z;
  wire [23:0] A, B;
  wire [21:0] Z;
  wire n_73, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163;
  wire n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171;
  wire n_172, n_173, n_174, n_175, n_176, n_180;
  nand g4 (n_73, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_77, A[1], B[1]);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_117, A[9], B[9]);
  nand g59 (n_118, A[9], n_116);
  nand g60 (n_119, B[9], n_116);
  nand g61 (n_121, n_117, n_118, n_119);
  xor g62 (n_120, A[9], B[9]);
  xor g63 (Z[9], n_116, n_120);
  nand g64 (n_122, A[10], B[10]);
  nand g65 (n_123, A[10], n_121);
  nand g66 (n_124, B[10], n_121);
  nand g67 (n_126, n_122, n_123, n_124);
  xor g68 (n_125, A[10], B[10]);
  xor g69 (Z[10], n_121, n_125);
  nand g70 (n_127, A[11], B[11]);
  nand g71 (n_128, A[11], n_126);
  nand g72 (n_129, B[11], n_126);
  nand g73 (n_131, n_127, n_128, n_129);
  xor g74 (n_130, A[11], B[11]);
  xor g75 (Z[11], n_126, n_130);
  nand g76 (n_132, A[12], B[12]);
  nand g77 (n_133, A[12], n_131);
  nand g78 (n_134, B[12], n_131);
  nand g79 (n_136, n_132, n_133, n_134);
  xor g80 (n_135, A[12], B[12]);
  xor g81 (Z[12], n_131, n_135);
  nand g82 (n_137, A[13], B[13]);
  nand g83 (n_138, A[13], n_136);
  nand g84 (n_139, B[13], n_136);
  nand g85 (n_141, n_137, n_138, n_139);
  xor g86 (n_140, A[13], B[13]);
  xor g87 (Z[13], n_136, n_140);
  nand g88 (n_142, A[14], B[14]);
  nand g89 (n_143, A[14], n_141);
  nand g90 (n_144, B[14], n_141);
  nand g91 (n_146, n_142, n_143, n_144);
  xor g92 (n_145, A[14], B[14]);
  xor g93 (Z[14], n_141, n_145);
  nand g94 (n_147, A[15], B[15]);
  nand g95 (n_148, A[15], n_146);
  nand g96 (n_149, B[15], n_146);
  nand g97 (n_151, n_147, n_148, n_149);
  xor g98 (n_150, A[15], B[15]);
  xor g99 (Z[15], n_146, n_150);
  nand g100 (n_152, A[16], B[16]);
  nand g101 (n_153, A[16], n_151);
  nand g102 (n_154, B[16], n_151);
  nand g103 (n_156, n_152, n_153, n_154);
  xor g104 (n_155, A[16], B[16]);
  xor g105 (Z[16], n_151, n_155);
  nand g106 (n_157, A[17], B[17]);
  nand g107 (n_158, A[17], n_156);
  nand g108 (n_159, B[17], n_156);
  nand g109 (n_161, n_157, n_158, n_159);
  xor g110 (n_160, A[17], B[17]);
  xor g111 (Z[17], n_156, n_160);
  nand g112 (n_162, A[18], B[18]);
  nand g113 (n_163, A[18], n_161);
  nand g114 (n_164, B[18], n_161);
  nand g115 (n_166, n_162, n_163, n_164);
  xor g116 (n_165, A[18], B[18]);
  xor g117 (Z[18], n_161, n_165);
  nand g118 (n_167, A[19], B[19]);
  nand g119 (n_168, A[19], n_166);
  nand g120 (n_169, B[19], n_166);
  nand g121 (n_171, n_167, n_168, n_169);
  xor g122 (n_170, A[19], B[19]);
  xor g123 (Z[19], n_166, n_170);
  nand g124 (n_172, A[20], B[20]);
  nand g125 (n_173, A[20], n_171);
  nand g126 (n_174, B[20], n_171);
  nand g127 (n_176, n_172, n_173, n_174);
  xor g128 (n_175, A[20], B[20]);
  xor g129 (Z[20], n_171, n_175);
  xor g135 (Z[21], n_176, n_180);
  xor g137 (n_180, A[21], B[21]);
  or g138 (n_78, wc, n_73);
  not gc (wc, A[1]);
  or g139 (n_79, wc0, n_73);
  not gc0 (wc0, B[1]);
  xnor g140 (Z[1], n_73, n_80);
endmodule

module add_signed_GENERIC(A, B, Z);
  input [23:0] A, B;
  output [21:0] Z;
  wire [23:0] A, B;
  wire [21:0] Z;
  add_signed_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3150_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  wire n_76, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_188;
  nand g4 (n_76, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_120, A[9], B[9]);
  nand g59 (n_121, A[9], n_119);
  nand g60 (n_122, B[9], n_119);
  nand g61 (n_124, n_120, n_121, n_122);
  xor g62 (n_123, A[9], B[9]);
  xor g63 (Z[9], n_119, n_123);
  nand g64 (n_125, A[10], B[10]);
  nand g65 (n_126, A[10], n_124);
  nand g66 (n_127, B[10], n_124);
  nand g67 (n_129, n_125, n_126, n_127);
  xor g68 (n_128, A[10], B[10]);
  xor g69 (Z[10], n_124, n_128);
  nand g70 (n_130, A[11], B[11]);
  nand g71 (n_131, A[11], n_129);
  nand g72 (n_132, B[11], n_129);
  nand g73 (n_134, n_130, n_131, n_132);
  xor g74 (n_133, A[11], B[11]);
  xor g75 (Z[11], n_129, n_133);
  nand g76 (n_135, A[12], B[12]);
  nand g77 (n_136, A[12], n_134);
  nand g78 (n_137, B[12], n_134);
  nand g79 (n_139, n_135, n_136, n_137);
  xor g80 (n_138, A[12], B[12]);
  xor g81 (Z[12], n_134, n_138);
  nand g82 (n_140, A[13], B[13]);
  nand g83 (n_141, A[13], n_139);
  nand g84 (n_142, B[13], n_139);
  nand g85 (n_144, n_140, n_141, n_142);
  xor g86 (n_143, A[13], B[13]);
  xor g87 (Z[13], n_139, n_143);
  nand g88 (n_145, A[14], B[14]);
  nand g89 (n_146, A[14], n_144);
  nand g90 (n_147, B[14], n_144);
  nand g91 (n_149, n_145, n_146, n_147);
  xor g92 (n_148, A[14], B[14]);
  xor g93 (Z[14], n_144, n_148);
  nand g94 (n_150, A[15], B[15]);
  nand g95 (n_151, A[15], n_149);
  nand g96 (n_152, B[15], n_149);
  nand g97 (n_154, n_150, n_151, n_152);
  xor g98 (n_153, A[15], B[15]);
  xor g99 (Z[15], n_149, n_153);
  nand g100 (n_155, A[16], B[16]);
  nand g101 (n_156, A[16], n_154);
  nand g102 (n_157, B[16], n_154);
  nand g103 (n_159, n_155, n_156, n_157);
  xor g104 (n_158, A[16], B[16]);
  xor g105 (Z[16], n_154, n_158);
  nand g106 (n_160, A[17], B[17]);
  nand g107 (n_161, A[17], n_159);
  nand g108 (n_162, B[17], n_159);
  nand g109 (n_164, n_160, n_161, n_162);
  xor g110 (n_163, A[17], B[17]);
  xor g111 (Z[17], n_159, n_163);
  nand g112 (n_165, A[18], B[18]);
  nand g113 (n_166, A[18], n_164);
  nand g114 (n_167, B[18], n_164);
  nand g115 (n_169, n_165, n_166, n_167);
  xor g116 (n_168, A[18], B[18]);
  xor g117 (Z[18], n_164, n_168);
  nand g118 (n_170, A[19], B[19]);
  nand g119 (n_171, A[19], n_169);
  nand g120 (n_172, B[19], n_169);
  nand g121 (n_174, n_170, n_171, n_172);
  xor g122 (n_173, A[19], B[19]);
  xor g123 (Z[19], n_169, n_173);
  nand g124 (n_175, A[20], B[20]);
  nand g125 (n_176, A[20], n_174);
  nand g126 (n_177, B[20], n_174);
  nand g127 (n_179, n_175, n_176, n_177);
  xor g128 (n_178, A[20], B[20]);
  xor g129 (Z[20], n_174, n_178);
  nand g130 (n_180, A[21], B[21]);
  nand g131 (n_181, A[21], n_179);
  nand g132 (n_182, B[21], n_179);
  nand g133 (n_184, n_180, n_181, n_182);
  xor g134 (n_183, A[21], B[21]);
  xor g135 (Z[21], n_179, n_183);
  xor g141 (Z[22], n_184, n_188);
  xor g143 (n_188, A[22], B[22]);
  or g144 (n_81, wc, n_76);
  not gc (wc, A[1]);
  or g145 (n_82, wc0, n_76);
  not gc0 (wc0, B[1]);
  xnor g146 (Z[1], n_76, n_83);
endmodule

module add_signed_3150_GENERIC(A, B, Z);
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  add_signed_3150_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3150_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  wire n_76, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_188;
  nand g4 (n_76, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_120, A[9], B[9]);
  nand g59 (n_121, A[9], n_119);
  nand g60 (n_122, B[9], n_119);
  nand g61 (n_124, n_120, n_121, n_122);
  xor g62 (n_123, A[9], B[9]);
  xor g63 (Z[9], n_119, n_123);
  nand g64 (n_125, A[10], B[10]);
  nand g65 (n_126, A[10], n_124);
  nand g66 (n_127, B[10], n_124);
  nand g67 (n_129, n_125, n_126, n_127);
  xor g68 (n_128, A[10], B[10]);
  xor g69 (Z[10], n_124, n_128);
  nand g70 (n_130, A[11], B[11]);
  nand g71 (n_131, A[11], n_129);
  nand g72 (n_132, B[11], n_129);
  nand g73 (n_134, n_130, n_131, n_132);
  xor g74 (n_133, A[11], B[11]);
  xor g75 (Z[11], n_129, n_133);
  nand g76 (n_135, A[12], B[12]);
  nand g77 (n_136, A[12], n_134);
  nand g78 (n_137, B[12], n_134);
  nand g79 (n_139, n_135, n_136, n_137);
  xor g80 (n_138, A[12], B[12]);
  xor g81 (Z[12], n_134, n_138);
  nand g82 (n_140, A[13], B[13]);
  nand g83 (n_141, A[13], n_139);
  nand g84 (n_142, B[13], n_139);
  nand g85 (n_144, n_140, n_141, n_142);
  xor g86 (n_143, A[13], B[13]);
  xor g87 (Z[13], n_139, n_143);
  nand g88 (n_145, A[14], B[14]);
  nand g89 (n_146, A[14], n_144);
  nand g90 (n_147, B[14], n_144);
  nand g91 (n_149, n_145, n_146, n_147);
  xor g92 (n_148, A[14], B[14]);
  xor g93 (Z[14], n_144, n_148);
  nand g94 (n_150, A[15], B[15]);
  nand g95 (n_151, A[15], n_149);
  nand g96 (n_152, B[15], n_149);
  nand g97 (n_154, n_150, n_151, n_152);
  xor g98 (n_153, A[15], B[15]);
  xor g99 (Z[15], n_149, n_153);
  nand g100 (n_155, A[16], B[16]);
  nand g101 (n_156, A[16], n_154);
  nand g102 (n_157, B[16], n_154);
  nand g103 (n_159, n_155, n_156, n_157);
  xor g104 (n_158, A[16], B[16]);
  xor g105 (Z[16], n_154, n_158);
  nand g106 (n_160, A[17], B[17]);
  nand g107 (n_161, A[17], n_159);
  nand g108 (n_162, B[17], n_159);
  nand g109 (n_164, n_160, n_161, n_162);
  xor g110 (n_163, A[17], B[17]);
  xor g111 (Z[17], n_159, n_163);
  nand g112 (n_165, A[18], B[18]);
  nand g113 (n_166, A[18], n_164);
  nand g114 (n_167, B[18], n_164);
  nand g115 (n_169, n_165, n_166, n_167);
  xor g116 (n_168, A[18], B[18]);
  xor g117 (Z[18], n_164, n_168);
  nand g118 (n_170, A[19], B[19]);
  nand g119 (n_171, A[19], n_169);
  nand g120 (n_172, B[19], n_169);
  nand g121 (n_174, n_170, n_171, n_172);
  xor g122 (n_173, A[19], B[19]);
  xor g123 (Z[19], n_169, n_173);
  nand g124 (n_175, A[20], B[20]);
  nand g125 (n_176, A[20], n_174);
  nand g126 (n_177, B[20], n_174);
  nand g127 (n_179, n_175, n_176, n_177);
  xor g128 (n_178, A[20], B[20]);
  xor g129 (Z[20], n_174, n_178);
  nand g130 (n_180, A[21], B[21]);
  nand g131 (n_181, A[21], n_179);
  nand g132 (n_182, B[21], n_179);
  nand g133 (n_184, n_180, n_181, n_182);
  xor g134 (n_183, A[21], B[21]);
  xor g135 (Z[21], n_179, n_183);
  xor g141 (Z[22], n_184, n_188);
  xor g143 (n_188, A[22], B[22]);
  or g144 (n_81, wc, n_76);
  not gc (wc, A[1]);
  or g145 (n_82, wc0, n_76);
  not gc0 (wc0, B[1]);
  xnor g146 (Z[1], n_76, n_83);
endmodule

module add_signed_3150_1_GENERIC(A, B, Z);
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  add_signed_3150_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3150_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  wire n_76, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_188;
  nand g4 (n_76, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_120, A[9], B[9]);
  nand g59 (n_121, A[9], n_119);
  nand g60 (n_122, B[9], n_119);
  nand g61 (n_124, n_120, n_121, n_122);
  xor g62 (n_123, A[9], B[9]);
  xor g63 (Z[9], n_119, n_123);
  nand g64 (n_125, A[10], B[10]);
  nand g65 (n_126, A[10], n_124);
  nand g66 (n_127, B[10], n_124);
  nand g67 (n_129, n_125, n_126, n_127);
  xor g68 (n_128, A[10], B[10]);
  xor g69 (Z[10], n_124, n_128);
  nand g70 (n_130, A[11], B[11]);
  nand g71 (n_131, A[11], n_129);
  nand g72 (n_132, B[11], n_129);
  nand g73 (n_134, n_130, n_131, n_132);
  xor g74 (n_133, A[11], B[11]);
  xor g75 (Z[11], n_129, n_133);
  nand g76 (n_135, A[12], B[12]);
  nand g77 (n_136, A[12], n_134);
  nand g78 (n_137, B[12], n_134);
  nand g79 (n_139, n_135, n_136, n_137);
  xor g80 (n_138, A[12], B[12]);
  xor g81 (Z[12], n_134, n_138);
  nand g82 (n_140, A[13], B[13]);
  nand g83 (n_141, A[13], n_139);
  nand g84 (n_142, B[13], n_139);
  nand g85 (n_144, n_140, n_141, n_142);
  xor g86 (n_143, A[13], B[13]);
  xor g87 (Z[13], n_139, n_143);
  nand g88 (n_145, A[14], B[14]);
  nand g89 (n_146, A[14], n_144);
  nand g90 (n_147, B[14], n_144);
  nand g91 (n_149, n_145, n_146, n_147);
  xor g92 (n_148, A[14], B[14]);
  xor g93 (Z[14], n_144, n_148);
  nand g94 (n_150, A[15], B[15]);
  nand g95 (n_151, A[15], n_149);
  nand g96 (n_152, B[15], n_149);
  nand g97 (n_154, n_150, n_151, n_152);
  xor g98 (n_153, A[15], B[15]);
  xor g99 (Z[15], n_149, n_153);
  nand g100 (n_155, A[16], B[16]);
  nand g101 (n_156, A[16], n_154);
  nand g102 (n_157, B[16], n_154);
  nand g103 (n_159, n_155, n_156, n_157);
  xor g104 (n_158, A[16], B[16]);
  xor g105 (Z[16], n_154, n_158);
  nand g106 (n_160, A[17], B[17]);
  nand g107 (n_161, A[17], n_159);
  nand g108 (n_162, B[17], n_159);
  nand g109 (n_164, n_160, n_161, n_162);
  xor g110 (n_163, A[17], B[17]);
  xor g111 (Z[17], n_159, n_163);
  nand g112 (n_165, A[18], B[18]);
  nand g113 (n_166, A[18], n_164);
  nand g114 (n_167, B[18], n_164);
  nand g115 (n_169, n_165, n_166, n_167);
  xor g116 (n_168, A[18], B[18]);
  xor g117 (Z[18], n_164, n_168);
  nand g118 (n_170, A[19], B[19]);
  nand g119 (n_171, A[19], n_169);
  nand g120 (n_172, B[19], n_169);
  nand g121 (n_174, n_170, n_171, n_172);
  xor g122 (n_173, A[19], B[19]);
  xor g123 (Z[19], n_169, n_173);
  nand g124 (n_175, A[20], B[20]);
  nand g125 (n_176, A[20], n_174);
  nand g126 (n_177, B[20], n_174);
  nand g127 (n_179, n_175, n_176, n_177);
  xor g128 (n_178, A[20], B[20]);
  xor g129 (Z[20], n_174, n_178);
  nand g130 (n_180, A[21], B[21]);
  nand g131 (n_181, A[21], n_179);
  nand g132 (n_182, B[21], n_179);
  nand g133 (n_184, n_180, n_181, n_182);
  xor g134 (n_183, A[21], B[21]);
  xor g135 (Z[21], n_179, n_183);
  xor g141 (Z[22], n_184, n_188);
  xor g143 (n_188, A[22], B[22]);
  or g144 (n_81, wc, n_76);
  not gc (wc, A[1]);
  or g145 (n_82, wc0, n_76);
  not gc0 (wc0, B[1]);
  xnor g146 (Z[1], n_76, n_83);
endmodule

module add_signed_3150_2_GENERIC(A, B, Z);
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  add_signed_3150_2_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3179_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  wire n_79, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_196;
  nand g4 (n_79, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_83, A[1], B[1]);
  nand g13 (n_87, n_83, n_84, n_85);
  xor g14 (n_86, A[1], B[1]);
  nand g16 (n_88, A[2], B[2]);
  nand g17 (n_89, A[2], n_87);
  nand g18 (n_90, B[2], n_87);
  nand g19 (n_92, n_88, n_89, n_90);
  xor g20 (n_91, A[2], B[2]);
  xor g21 (Z[2], n_87, n_91);
  nand g22 (n_93, A[3], B[3]);
  nand g23 (n_94, A[3], n_92);
  nand g24 (n_95, B[3], n_92);
  nand g25 (n_97, n_93, n_94, n_95);
  xor g26 (n_96, A[3], B[3]);
  xor g27 (Z[3], n_92, n_96);
  nand g28 (n_98, A[4], B[4]);
  nand g29 (n_99, A[4], n_97);
  nand g30 (n_100, B[4], n_97);
  nand g31 (n_102, n_98, n_99, n_100);
  xor g32 (n_101, A[4], B[4]);
  xor g33 (Z[4], n_97, n_101);
  nand g34 (n_103, A[5], B[5]);
  nand g35 (n_104, A[5], n_102);
  nand g36 (n_105, B[5], n_102);
  nand g37 (n_107, n_103, n_104, n_105);
  xor g38 (n_106, A[5], B[5]);
  xor g39 (Z[5], n_102, n_106);
  nand g40 (n_108, A[6], B[6]);
  nand g41 (n_109, A[6], n_107);
  nand g42 (n_110, B[6], n_107);
  nand g43 (n_112, n_108, n_109, n_110);
  xor g44 (n_111, A[6], B[6]);
  xor g45 (Z[6], n_107, n_111);
  nand g46 (n_113, A[7], B[7]);
  nand g47 (n_114, A[7], n_112);
  nand g48 (n_115, B[7], n_112);
  nand g49 (n_117, n_113, n_114, n_115);
  xor g50 (n_116, A[7], B[7]);
  xor g51 (Z[7], n_112, n_116);
  nand g52 (n_118, A[8], B[8]);
  nand g53 (n_119, A[8], n_117);
  nand g54 (n_120, B[8], n_117);
  nand g55 (n_122, n_118, n_119, n_120);
  xor g56 (n_121, A[8], B[8]);
  xor g57 (Z[8], n_117, n_121);
  nand g58 (n_123, A[9], B[9]);
  nand g59 (n_124, A[9], n_122);
  nand g60 (n_125, B[9], n_122);
  nand g61 (n_127, n_123, n_124, n_125);
  xor g62 (n_126, A[9], B[9]);
  xor g63 (Z[9], n_122, n_126);
  nand g64 (n_128, A[10], B[10]);
  nand g65 (n_129, A[10], n_127);
  nand g66 (n_130, B[10], n_127);
  nand g67 (n_132, n_128, n_129, n_130);
  xor g68 (n_131, A[10], B[10]);
  xor g69 (Z[10], n_127, n_131);
  nand g70 (n_133, A[11], B[11]);
  nand g71 (n_134, A[11], n_132);
  nand g72 (n_135, B[11], n_132);
  nand g73 (n_137, n_133, n_134, n_135);
  xor g74 (n_136, A[11], B[11]);
  xor g75 (Z[11], n_132, n_136);
  nand g76 (n_138, A[12], B[12]);
  nand g77 (n_139, A[12], n_137);
  nand g78 (n_140, B[12], n_137);
  nand g79 (n_142, n_138, n_139, n_140);
  xor g80 (n_141, A[12], B[12]);
  xor g81 (Z[12], n_137, n_141);
  nand g82 (n_143, A[13], B[13]);
  nand g83 (n_144, A[13], n_142);
  nand g84 (n_145, B[13], n_142);
  nand g85 (n_147, n_143, n_144, n_145);
  xor g86 (n_146, A[13], B[13]);
  xor g87 (Z[13], n_142, n_146);
  nand g88 (n_148, A[14], B[14]);
  nand g89 (n_149, A[14], n_147);
  nand g90 (n_150, B[14], n_147);
  nand g91 (n_152, n_148, n_149, n_150);
  xor g92 (n_151, A[14], B[14]);
  xor g93 (Z[14], n_147, n_151);
  nand g94 (n_153, A[15], B[15]);
  nand g95 (n_154, A[15], n_152);
  nand g96 (n_155, B[15], n_152);
  nand g97 (n_157, n_153, n_154, n_155);
  xor g98 (n_156, A[15], B[15]);
  xor g99 (Z[15], n_152, n_156);
  nand g100 (n_158, A[16], B[16]);
  nand g101 (n_159, A[16], n_157);
  nand g102 (n_160, B[16], n_157);
  nand g103 (n_162, n_158, n_159, n_160);
  xor g104 (n_161, A[16], B[16]);
  xor g105 (Z[16], n_157, n_161);
  nand g106 (n_163, A[17], B[17]);
  nand g107 (n_164, A[17], n_162);
  nand g108 (n_165, B[17], n_162);
  nand g109 (n_167, n_163, n_164, n_165);
  xor g110 (n_166, A[17], B[17]);
  xor g111 (Z[17], n_162, n_166);
  nand g112 (n_168, A[18], B[18]);
  nand g113 (n_169, A[18], n_167);
  nand g114 (n_170, B[18], n_167);
  nand g115 (n_172, n_168, n_169, n_170);
  xor g116 (n_171, A[18], B[18]);
  xor g117 (Z[18], n_167, n_171);
  nand g118 (n_173, A[19], B[19]);
  nand g119 (n_174, A[19], n_172);
  nand g120 (n_175, B[19], n_172);
  nand g121 (n_177, n_173, n_174, n_175);
  xor g122 (n_176, A[19], B[19]);
  xor g123 (Z[19], n_172, n_176);
  nand g124 (n_178, A[20], B[20]);
  nand g125 (n_179, A[20], n_177);
  nand g126 (n_180, B[20], n_177);
  nand g127 (n_182, n_178, n_179, n_180);
  xor g128 (n_181, A[20], B[20]);
  xor g129 (Z[20], n_177, n_181);
  nand g130 (n_183, A[21], B[21]);
  nand g131 (n_184, A[21], n_182);
  nand g132 (n_185, B[21], n_182);
  nand g133 (n_187, n_183, n_184, n_185);
  xor g134 (n_186, A[21], B[21]);
  xor g135 (Z[21], n_182, n_186);
  nand g136 (n_188, A[22], B[22]);
  nand g137 (n_189, A[22], n_187);
  nand g138 (n_190, B[22], n_187);
  nand g139 (n_192, n_188, n_189, n_190);
  xor g140 (n_191, A[22], B[22]);
  xor g141 (Z[22], n_187, n_191);
  xor g147 (Z[23], n_192, n_196);
  xor g149 (n_196, A[23], B[23]);
  or g150 (n_84, wc, n_79);
  not gc (wc, A[1]);
  or g151 (n_85, wc0, n_79);
  not gc0 (wc0, B[1]);
  xnor g152 (Z[1], n_79, n_86);
endmodule

module add_signed_3179_GENERIC(A, B, Z);
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  add_signed_3179_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3179_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  wire n_79, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_196;
  nand g4 (n_79, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_83, A[1], B[1]);
  nand g13 (n_87, n_83, n_84, n_85);
  xor g14 (n_86, A[1], B[1]);
  nand g16 (n_88, A[2], B[2]);
  nand g17 (n_89, A[2], n_87);
  nand g18 (n_90, B[2], n_87);
  nand g19 (n_92, n_88, n_89, n_90);
  xor g20 (n_91, A[2], B[2]);
  xor g21 (Z[2], n_87, n_91);
  nand g22 (n_93, A[3], B[3]);
  nand g23 (n_94, A[3], n_92);
  nand g24 (n_95, B[3], n_92);
  nand g25 (n_97, n_93, n_94, n_95);
  xor g26 (n_96, A[3], B[3]);
  xor g27 (Z[3], n_92, n_96);
  nand g28 (n_98, A[4], B[4]);
  nand g29 (n_99, A[4], n_97);
  nand g30 (n_100, B[4], n_97);
  nand g31 (n_102, n_98, n_99, n_100);
  xor g32 (n_101, A[4], B[4]);
  xor g33 (Z[4], n_97, n_101);
  nand g34 (n_103, A[5], B[5]);
  nand g35 (n_104, A[5], n_102);
  nand g36 (n_105, B[5], n_102);
  nand g37 (n_107, n_103, n_104, n_105);
  xor g38 (n_106, A[5], B[5]);
  xor g39 (Z[5], n_102, n_106);
  nand g40 (n_108, A[6], B[6]);
  nand g41 (n_109, A[6], n_107);
  nand g42 (n_110, B[6], n_107);
  nand g43 (n_112, n_108, n_109, n_110);
  xor g44 (n_111, A[6], B[6]);
  xor g45 (Z[6], n_107, n_111);
  nand g46 (n_113, A[7], B[7]);
  nand g47 (n_114, A[7], n_112);
  nand g48 (n_115, B[7], n_112);
  nand g49 (n_117, n_113, n_114, n_115);
  xor g50 (n_116, A[7], B[7]);
  xor g51 (Z[7], n_112, n_116);
  nand g52 (n_118, A[8], B[8]);
  nand g53 (n_119, A[8], n_117);
  nand g54 (n_120, B[8], n_117);
  nand g55 (n_122, n_118, n_119, n_120);
  xor g56 (n_121, A[8], B[8]);
  xor g57 (Z[8], n_117, n_121);
  nand g58 (n_123, A[9], B[9]);
  nand g59 (n_124, A[9], n_122);
  nand g60 (n_125, B[9], n_122);
  nand g61 (n_127, n_123, n_124, n_125);
  xor g62 (n_126, A[9], B[9]);
  xor g63 (Z[9], n_122, n_126);
  nand g64 (n_128, A[10], B[10]);
  nand g65 (n_129, A[10], n_127);
  nand g66 (n_130, B[10], n_127);
  nand g67 (n_132, n_128, n_129, n_130);
  xor g68 (n_131, A[10], B[10]);
  xor g69 (Z[10], n_127, n_131);
  nand g70 (n_133, A[11], B[11]);
  nand g71 (n_134, A[11], n_132);
  nand g72 (n_135, B[11], n_132);
  nand g73 (n_137, n_133, n_134, n_135);
  xor g74 (n_136, A[11], B[11]);
  xor g75 (Z[11], n_132, n_136);
  nand g76 (n_138, A[12], B[12]);
  nand g77 (n_139, A[12], n_137);
  nand g78 (n_140, B[12], n_137);
  nand g79 (n_142, n_138, n_139, n_140);
  xor g80 (n_141, A[12], B[12]);
  xor g81 (Z[12], n_137, n_141);
  nand g82 (n_143, A[13], B[13]);
  nand g83 (n_144, A[13], n_142);
  nand g84 (n_145, B[13], n_142);
  nand g85 (n_147, n_143, n_144, n_145);
  xor g86 (n_146, A[13], B[13]);
  xor g87 (Z[13], n_142, n_146);
  nand g88 (n_148, A[14], B[14]);
  nand g89 (n_149, A[14], n_147);
  nand g90 (n_150, B[14], n_147);
  nand g91 (n_152, n_148, n_149, n_150);
  xor g92 (n_151, A[14], B[14]);
  xor g93 (Z[14], n_147, n_151);
  nand g94 (n_153, A[15], B[15]);
  nand g95 (n_154, A[15], n_152);
  nand g96 (n_155, B[15], n_152);
  nand g97 (n_157, n_153, n_154, n_155);
  xor g98 (n_156, A[15], B[15]);
  xor g99 (Z[15], n_152, n_156);
  nand g100 (n_158, A[16], B[16]);
  nand g101 (n_159, A[16], n_157);
  nand g102 (n_160, B[16], n_157);
  nand g103 (n_162, n_158, n_159, n_160);
  xor g104 (n_161, A[16], B[16]);
  xor g105 (Z[16], n_157, n_161);
  nand g106 (n_163, A[17], B[17]);
  nand g107 (n_164, A[17], n_162);
  nand g108 (n_165, B[17], n_162);
  nand g109 (n_167, n_163, n_164, n_165);
  xor g110 (n_166, A[17], B[17]);
  xor g111 (Z[17], n_162, n_166);
  nand g112 (n_168, A[18], B[18]);
  nand g113 (n_169, A[18], n_167);
  nand g114 (n_170, B[18], n_167);
  nand g115 (n_172, n_168, n_169, n_170);
  xor g116 (n_171, A[18], B[18]);
  xor g117 (Z[18], n_167, n_171);
  nand g118 (n_173, A[19], B[19]);
  nand g119 (n_174, A[19], n_172);
  nand g120 (n_175, B[19], n_172);
  nand g121 (n_177, n_173, n_174, n_175);
  xor g122 (n_176, A[19], B[19]);
  xor g123 (Z[19], n_172, n_176);
  nand g124 (n_178, A[20], B[20]);
  nand g125 (n_179, A[20], n_177);
  nand g126 (n_180, B[20], n_177);
  nand g127 (n_182, n_178, n_179, n_180);
  xor g128 (n_181, A[20], B[20]);
  xor g129 (Z[20], n_177, n_181);
  nand g130 (n_183, A[21], B[21]);
  nand g131 (n_184, A[21], n_182);
  nand g132 (n_185, B[21], n_182);
  nand g133 (n_187, n_183, n_184, n_185);
  xor g134 (n_186, A[21], B[21]);
  xor g135 (Z[21], n_182, n_186);
  nand g136 (n_188, A[22], B[22]);
  nand g137 (n_189, A[22], n_187);
  nand g138 (n_190, B[22], n_187);
  nand g139 (n_192, n_188, n_189, n_190);
  xor g140 (n_191, A[22], B[22]);
  xor g141 (Z[22], n_187, n_191);
  xor g147 (Z[23], n_192, n_196);
  xor g149 (n_196, A[23], B[23]);
  or g150 (n_84, wc, n_79);
  not gc (wc, A[1]);
  or g151 (n_85, wc0, n_79);
  not gc0 (wc0, B[1]);
  xnor g152 (Z[1], n_79, n_86);
endmodule

module add_signed_3179_1_GENERIC(A, B, Z);
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  add_signed_3179_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3179_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  wire n_79, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_196;
  nand g4 (n_79, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_83, A[1], B[1]);
  nand g13 (n_87, n_83, n_84, n_85);
  xor g14 (n_86, A[1], B[1]);
  nand g16 (n_88, A[2], B[2]);
  nand g17 (n_89, A[2], n_87);
  nand g18 (n_90, B[2], n_87);
  nand g19 (n_92, n_88, n_89, n_90);
  xor g20 (n_91, A[2], B[2]);
  xor g21 (Z[2], n_87, n_91);
  nand g22 (n_93, A[3], B[3]);
  nand g23 (n_94, A[3], n_92);
  nand g24 (n_95, B[3], n_92);
  nand g25 (n_97, n_93, n_94, n_95);
  xor g26 (n_96, A[3], B[3]);
  xor g27 (Z[3], n_92, n_96);
  nand g28 (n_98, A[4], B[4]);
  nand g29 (n_99, A[4], n_97);
  nand g30 (n_100, B[4], n_97);
  nand g31 (n_102, n_98, n_99, n_100);
  xor g32 (n_101, A[4], B[4]);
  xor g33 (Z[4], n_97, n_101);
  nand g34 (n_103, A[5], B[5]);
  nand g35 (n_104, A[5], n_102);
  nand g36 (n_105, B[5], n_102);
  nand g37 (n_107, n_103, n_104, n_105);
  xor g38 (n_106, A[5], B[5]);
  xor g39 (Z[5], n_102, n_106);
  nand g40 (n_108, A[6], B[6]);
  nand g41 (n_109, A[6], n_107);
  nand g42 (n_110, B[6], n_107);
  nand g43 (n_112, n_108, n_109, n_110);
  xor g44 (n_111, A[6], B[6]);
  xor g45 (Z[6], n_107, n_111);
  nand g46 (n_113, A[7], B[7]);
  nand g47 (n_114, A[7], n_112);
  nand g48 (n_115, B[7], n_112);
  nand g49 (n_117, n_113, n_114, n_115);
  xor g50 (n_116, A[7], B[7]);
  xor g51 (Z[7], n_112, n_116);
  nand g52 (n_118, A[8], B[8]);
  nand g53 (n_119, A[8], n_117);
  nand g54 (n_120, B[8], n_117);
  nand g55 (n_122, n_118, n_119, n_120);
  xor g56 (n_121, A[8], B[8]);
  xor g57 (Z[8], n_117, n_121);
  nand g58 (n_123, A[9], B[9]);
  nand g59 (n_124, A[9], n_122);
  nand g60 (n_125, B[9], n_122);
  nand g61 (n_127, n_123, n_124, n_125);
  xor g62 (n_126, A[9], B[9]);
  xor g63 (Z[9], n_122, n_126);
  nand g64 (n_128, A[10], B[10]);
  nand g65 (n_129, A[10], n_127);
  nand g66 (n_130, B[10], n_127);
  nand g67 (n_132, n_128, n_129, n_130);
  xor g68 (n_131, A[10], B[10]);
  xor g69 (Z[10], n_127, n_131);
  nand g70 (n_133, A[11], B[11]);
  nand g71 (n_134, A[11], n_132);
  nand g72 (n_135, B[11], n_132);
  nand g73 (n_137, n_133, n_134, n_135);
  xor g74 (n_136, A[11], B[11]);
  xor g75 (Z[11], n_132, n_136);
  nand g76 (n_138, A[12], B[12]);
  nand g77 (n_139, A[12], n_137);
  nand g78 (n_140, B[12], n_137);
  nand g79 (n_142, n_138, n_139, n_140);
  xor g80 (n_141, A[12], B[12]);
  xor g81 (Z[12], n_137, n_141);
  nand g82 (n_143, A[13], B[13]);
  nand g83 (n_144, A[13], n_142);
  nand g84 (n_145, B[13], n_142);
  nand g85 (n_147, n_143, n_144, n_145);
  xor g86 (n_146, A[13], B[13]);
  xor g87 (Z[13], n_142, n_146);
  nand g88 (n_148, A[14], B[14]);
  nand g89 (n_149, A[14], n_147);
  nand g90 (n_150, B[14], n_147);
  nand g91 (n_152, n_148, n_149, n_150);
  xor g92 (n_151, A[14], B[14]);
  xor g93 (Z[14], n_147, n_151);
  nand g94 (n_153, A[15], B[15]);
  nand g95 (n_154, A[15], n_152);
  nand g96 (n_155, B[15], n_152);
  nand g97 (n_157, n_153, n_154, n_155);
  xor g98 (n_156, A[15], B[15]);
  xor g99 (Z[15], n_152, n_156);
  nand g100 (n_158, A[16], B[16]);
  nand g101 (n_159, A[16], n_157);
  nand g102 (n_160, B[16], n_157);
  nand g103 (n_162, n_158, n_159, n_160);
  xor g104 (n_161, A[16], B[16]);
  xor g105 (Z[16], n_157, n_161);
  nand g106 (n_163, A[17], B[17]);
  nand g107 (n_164, A[17], n_162);
  nand g108 (n_165, B[17], n_162);
  nand g109 (n_167, n_163, n_164, n_165);
  xor g110 (n_166, A[17], B[17]);
  xor g111 (Z[17], n_162, n_166);
  nand g112 (n_168, A[18], B[18]);
  nand g113 (n_169, A[18], n_167);
  nand g114 (n_170, B[18], n_167);
  nand g115 (n_172, n_168, n_169, n_170);
  xor g116 (n_171, A[18], B[18]);
  xor g117 (Z[18], n_167, n_171);
  nand g118 (n_173, A[19], B[19]);
  nand g119 (n_174, A[19], n_172);
  nand g120 (n_175, B[19], n_172);
  nand g121 (n_177, n_173, n_174, n_175);
  xor g122 (n_176, A[19], B[19]);
  xor g123 (Z[19], n_172, n_176);
  nand g124 (n_178, A[20], B[20]);
  nand g125 (n_179, A[20], n_177);
  nand g126 (n_180, B[20], n_177);
  nand g127 (n_182, n_178, n_179, n_180);
  xor g128 (n_181, A[20], B[20]);
  xor g129 (Z[20], n_177, n_181);
  nand g130 (n_183, A[21], B[21]);
  nand g131 (n_184, A[21], n_182);
  nand g132 (n_185, B[21], n_182);
  nand g133 (n_187, n_183, n_184, n_185);
  xor g134 (n_186, A[21], B[21]);
  xor g135 (Z[21], n_182, n_186);
  nand g136 (n_188, A[22], B[22]);
  nand g137 (n_189, A[22], n_187);
  nand g138 (n_190, B[22], n_187);
  nand g139 (n_192, n_188, n_189, n_190);
  xor g140 (n_191, A[22], B[22]);
  xor g141 (Z[22], n_187, n_191);
  xor g147 (Z[23], n_192, n_196);
  xor g149 (n_196, A[23], B[23]);
  or g150 (n_84, wc, n_79);
  not gc (wc, A[1]);
  or g151 (n_85, wc0, n_79);
  not gc0 (wc0, B[1]);
  xnor g152 (Z[1], n_79, n_86);
endmodule

module add_signed_3179_2_GENERIC(A, B, Z);
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  add_signed_3179_2_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3179_3_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  wire n_79, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_196;
  nand g4 (n_79, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_83, A[1], B[1]);
  nand g13 (n_87, n_83, n_84, n_85);
  xor g14 (n_86, A[1], B[1]);
  nand g16 (n_88, A[2], B[2]);
  nand g17 (n_89, A[2], n_87);
  nand g18 (n_90, B[2], n_87);
  nand g19 (n_92, n_88, n_89, n_90);
  xor g20 (n_91, A[2], B[2]);
  xor g21 (Z[2], n_87, n_91);
  nand g22 (n_93, A[3], B[3]);
  nand g23 (n_94, A[3], n_92);
  nand g24 (n_95, B[3], n_92);
  nand g25 (n_97, n_93, n_94, n_95);
  xor g26 (n_96, A[3], B[3]);
  xor g27 (Z[3], n_92, n_96);
  nand g28 (n_98, A[4], B[4]);
  nand g29 (n_99, A[4], n_97);
  nand g30 (n_100, B[4], n_97);
  nand g31 (n_102, n_98, n_99, n_100);
  xor g32 (n_101, A[4], B[4]);
  xor g33 (Z[4], n_97, n_101);
  nand g34 (n_103, A[5], B[5]);
  nand g35 (n_104, A[5], n_102);
  nand g36 (n_105, B[5], n_102);
  nand g37 (n_107, n_103, n_104, n_105);
  xor g38 (n_106, A[5], B[5]);
  xor g39 (Z[5], n_102, n_106);
  nand g40 (n_108, A[6], B[6]);
  nand g41 (n_109, A[6], n_107);
  nand g42 (n_110, B[6], n_107);
  nand g43 (n_112, n_108, n_109, n_110);
  xor g44 (n_111, A[6], B[6]);
  xor g45 (Z[6], n_107, n_111);
  nand g46 (n_113, A[7], B[7]);
  nand g47 (n_114, A[7], n_112);
  nand g48 (n_115, B[7], n_112);
  nand g49 (n_117, n_113, n_114, n_115);
  xor g50 (n_116, A[7], B[7]);
  xor g51 (Z[7], n_112, n_116);
  nand g52 (n_118, A[8], B[8]);
  nand g53 (n_119, A[8], n_117);
  nand g54 (n_120, B[8], n_117);
  nand g55 (n_122, n_118, n_119, n_120);
  xor g56 (n_121, A[8], B[8]);
  xor g57 (Z[8], n_117, n_121);
  nand g58 (n_123, A[9], B[9]);
  nand g59 (n_124, A[9], n_122);
  nand g60 (n_125, B[9], n_122);
  nand g61 (n_127, n_123, n_124, n_125);
  xor g62 (n_126, A[9], B[9]);
  xor g63 (Z[9], n_122, n_126);
  nand g64 (n_128, A[10], B[10]);
  nand g65 (n_129, A[10], n_127);
  nand g66 (n_130, B[10], n_127);
  nand g67 (n_132, n_128, n_129, n_130);
  xor g68 (n_131, A[10], B[10]);
  xor g69 (Z[10], n_127, n_131);
  nand g70 (n_133, A[11], B[11]);
  nand g71 (n_134, A[11], n_132);
  nand g72 (n_135, B[11], n_132);
  nand g73 (n_137, n_133, n_134, n_135);
  xor g74 (n_136, A[11], B[11]);
  xor g75 (Z[11], n_132, n_136);
  nand g76 (n_138, A[12], B[12]);
  nand g77 (n_139, A[12], n_137);
  nand g78 (n_140, B[12], n_137);
  nand g79 (n_142, n_138, n_139, n_140);
  xor g80 (n_141, A[12], B[12]);
  xor g81 (Z[12], n_137, n_141);
  nand g82 (n_143, A[13], B[13]);
  nand g83 (n_144, A[13], n_142);
  nand g84 (n_145, B[13], n_142);
  nand g85 (n_147, n_143, n_144, n_145);
  xor g86 (n_146, A[13], B[13]);
  xor g87 (Z[13], n_142, n_146);
  nand g88 (n_148, A[14], B[14]);
  nand g89 (n_149, A[14], n_147);
  nand g90 (n_150, B[14], n_147);
  nand g91 (n_152, n_148, n_149, n_150);
  xor g92 (n_151, A[14], B[14]);
  xor g93 (Z[14], n_147, n_151);
  nand g94 (n_153, A[15], B[15]);
  nand g95 (n_154, A[15], n_152);
  nand g96 (n_155, B[15], n_152);
  nand g97 (n_157, n_153, n_154, n_155);
  xor g98 (n_156, A[15], B[15]);
  xor g99 (Z[15], n_152, n_156);
  nand g100 (n_158, A[16], B[16]);
  nand g101 (n_159, A[16], n_157);
  nand g102 (n_160, B[16], n_157);
  nand g103 (n_162, n_158, n_159, n_160);
  xor g104 (n_161, A[16], B[16]);
  xor g105 (Z[16], n_157, n_161);
  nand g106 (n_163, A[17], B[17]);
  nand g107 (n_164, A[17], n_162);
  nand g108 (n_165, B[17], n_162);
  nand g109 (n_167, n_163, n_164, n_165);
  xor g110 (n_166, A[17], B[17]);
  xor g111 (Z[17], n_162, n_166);
  nand g112 (n_168, A[18], B[18]);
  nand g113 (n_169, A[18], n_167);
  nand g114 (n_170, B[18], n_167);
  nand g115 (n_172, n_168, n_169, n_170);
  xor g116 (n_171, A[18], B[18]);
  xor g117 (Z[18], n_167, n_171);
  nand g118 (n_173, A[19], B[19]);
  nand g119 (n_174, A[19], n_172);
  nand g120 (n_175, B[19], n_172);
  nand g121 (n_177, n_173, n_174, n_175);
  xor g122 (n_176, A[19], B[19]);
  xor g123 (Z[19], n_172, n_176);
  nand g124 (n_178, A[20], B[20]);
  nand g125 (n_179, A[20], n_177);
  nand g126 (n_180, B[20], n_177);
  nand g127 (n_182, n_178, n_179, n_180);
  xor g128 (n_181, A[20], B[20]);
  xor g129 (Z[20], n_177, n_181);
  nand g130 (n_183, A[21], B[21]);
  nand g131 (n_184, A[21], n_182);
  nand g132 (n_185, B[21], n_182);
  nand g133 (n_187, n_183, n_184, n_185);
  xor g134 (n_186, A[21], B[21]);
  xor g135 (Z[21], n_182, n_186);
  nand g136 (n_188, A[22], B[22]);
  nand g137 (n_189, A[22], n_187);
  nand g138 (n_190, B[22], n_187);
  nand g139 (n_192, n_188, n_189, n_190);
  xor g140 (n_191, A[22], B[22]);
  xor g141 (Z[22], n_187, n_191);
  xor g147 (Z[23], n_192, n_196);
  xor g149 (n_196, A[23], B[23]);
  or g150 (n_84, wc, n_79);
  not gc (wc, A[1]);
  or g151 (n_85, wc0, n_79);
  not gc0 (wc0, B[1]);
  xnor g152 (Z[1], n_79, n_86);
endmodule

module add_signed_3179_3_GENERIC(A, B, Z);
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  add_signed_3179_3_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_33_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [21:0] A, B;
  output [22:0] Z;
  wire [21:0] A, B;
  wire [22:0] Z;
  wire n_71, n_72, n_75, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_85, n_86, n_87, n_88, n_89, n_91, n_92;
  wire n_93, n_94, n_95, n_97, n_98, n_99, n_100, n_101;
  wire n_103, n_104, n_105, n_106, n_107, n_109, n_110, n_111;
  wire n_112, n_113, n_115, n_116, n_117, n_118, n_119, n_121;
  wire n_122, n_123, n_124, n_125, n_127, n_128, n_129, n_130;
  wire n_131, n_133, n_134, n_135, n_136, n_137, n_139, n_140;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_149, n_151;
  wire n_153, n_154, n_156, n_157, n_159, n_161, n_163, n_164;
  wire n_166, n_167, n_169, n_171, n_173, n_174, n_176, n_177;
  wire n_179, n_181, n_183, n_184, n_186, n_188, n_189, n_190;
  wire n_192, n_193, n_194, n_196, n_197, n_198, n_199, n_201;
  wire n_203, n_205, n_206, n_207, n_209, n_210, n_211, n_213;
  wire n_214, n_216, n_217, n_219, n_220, n_222, n_224, n_225;
  wire n_226, n_228, n_229, n_231, n_232, n_233, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_246, n_247, n_248, n_250, n_251, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_263;
  wire n_264, n_265, n_267, n_268, n_269, n_270, n_272, n_273;
  wire n_274, n_276, n_277, n_278, n_279, n_281, n_282, n_284;
  wire n_285, n_287, n_288, n_289, n_290, n_292, n_293, n_294;
  wire n_296, n_297, n_298, n_299, n_301, n_302, n_304, n_305;
  wire n_307, n_308;
  not g3 (Z[22], n_71);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_72, A[0], B[0]);
  nor g9 (n_75, A[1], B[1]);
  nand g10 (n_78, A[1], B[1]);
  nor g11 (n_85, A[2], B[2]);
  nand g12 (n_80, A[2], B[2]);
  nor g13 (n_81, A[3], B[3]);
  nand g14 (n_82, A[3], B[3]);
  nor g15 (n_91, A[4], B[4]);
  nand g16 (n_86, A[4], B[4]);
  nor g17 (n_87, A[5], B[5]);
  nand g18 (n_88, A[5], B[5]);
  nor g19 (n_97, A[6], B[6]);
  nand g20 (n_92, A[6], B[6]);
  nor g21 (n_93, A[7], B[7]);
  nand g22 (n_94, A[7], B[7]);
  nor g23 (n_103, A[8], B[8]);
  nand g24 (n_98, A[8], B[8]);
  nor g25 (n_99, A[9], B[9]);
  nand g26 (n_100, A[9], B[9]);
  nor g27 (n_109, A[10], B[10]);
  nand g28 (n_104, A[10], B[10]);
  nor g29 (n_105, A[11], B[11]);
  nand g30 (n_106, A[11], B[11]);
  nor g31 (n_115, A[12], B[12]);
  nand g32 (n_110, A[12], B[12]);
  nor g33 (n_111, A[13], B[13]);
  nand g34 (n_112, A[13], B[13]);
  nor g35 (n_121, A[14], B[14]);
  nand g36 (n_116, A[14], B[14]);
  nor g37 (n_117, A[15], B[15]);
  nand g38 (n_118, A[15], B[15]);
  nor g39 (n_127, A[16], B[16]);
  nand g40 (n_122, A[16], B[16]);
  nor g41 (n_123, A[17], B[17]);
  nand g42 (n_124, A[17], B[17]);
  nor g43 (n_133, A[18], B[18]);
  nand g44 (n_128, A[18], B[18]);
  nor g45 (n_129, A[19], B[19]);
  nand g46 (n_130, A[19], B[19]);
  nor g47 (n_139, A[20], B[20]);
  nand g48 (n_134, A[20], B[20]);
  nand g53 (n_140, n_78, n_79);
  nor g54 (n_83, n_80, n_81);
  nor g57 (n_143, n_85, n_81);
  nor g58 (n_89, n_86, n_87);
  nor g61 (n_149, n_91, n_87);
  nor g62 (n_95, n_92, n_93);
  nor g65 (n_151, n_97, n_93);
  nor g66 (n_101, n_98, n_99);
  nor g69 (n_159, n_103, n_99);
  nor g70 (n_107, n_104, n_105);
  nor g73 (n_161, n_109, n_105);
  nor g74 (n_113, n_110, n_111);
  nor g77 (n_169, n_115, n_111);
  nor g78 (n_119, n_116, n_117);
  nor g81 (n_171, n_121, n_117);
  nor g82 (n_125, n_122, n_123);
  nor g85 (n_179, n_127, n_123);
  nor g86 (n_131, n_128, n_129);
  nor g89 (n_181, n_133, n_129);
  nor g90 (n_137, n_134, n_135);
  nor g93 (n_217, n_139, n_135);
  nand g96 (n_263, n_80, n_142);
  nand g97 (n_145, n_143, n_140);
  nand g98 (n_186, n_144, n_145);
  nor g99 (n_147, n_97, n_146);
  nand g108 (n_194, n_149, n_151);
  nor g109 (n_157, n_109, n_156);
  nand g118 (n_201, n_159, n_161);
  nor g119 (n_167, n_121, n_166);
  nand g128 (n_209, n_169, n_171);
  nor g129 (n_177, n_133, n_176);
  nand g138 (n_216, n_179, n_181);
  nand g141 (n_267, n_86, n_188);
  nand g142 (n_189, n_149, n_186);
  nand g143 (n_269, n_146, n_189);
  nand g146 (n_272, n_192, n_193);
  nand g149 (n_222, n_196, n_197);
  nor g150 (n_199, n_115, n_198);
  nor g153 (n_232, n_115, n_201);
  nor g159 (n_207, n_205, n_198);
  nor g162 (n_238, n_201, n_205);
  nor g163 (n_211, n_209, n_198);
  nor g166 (n_241, n_201, n_209);
  nor g167 (n_214, n_139, n_213);
  nor g170 (n_254, n_139, n_216);
  nand g178 (n_276, n_98, n_224);
  nand g179 (n_225, n_159, n_222);
  nand g180 (n_278, n_156, n_225);
  nand g183 (n_281, n_228, n_229);
  nand g186 (n_284, n_198, n_231);
  nand g187 (n_234, n_232, n_222);
  nand g188 (n_287, n_233, n_234);
  nand g189 (n_237, n_235, n_222);
  nand g190 (n_289, n_236, n_237);
  nand g191 (n_240, n_238, n_222);
  nand g192 (n_292, n_239, n_240);
  nand g193 (n_243, n_241, n_222);
  nand g194 (n_244, n_242, n_243);
  nand g197 (n_296, n_122, n_246);
  nand g198 (n_247, n_179, n_244);
  nand g199 (n_298, n_176, n_247);
  nand g202 (n_301, n_250, n_251);
  nand g205 (n_304, n_213, n_253);
  nand g206 (n_256, n_254, n_244);
  nand g207 (n_307, n_255, n_256);
  nand g208 (n_259, n_257, n_244);
  nand g209 (n_71, n_258, n_259);
  xnor g213 (Z[2], n_140, n_261);
  xnor g216 (Z[3], n_263, n_264);
  xnor g218 (Z[4], n_186, n_265);
  xnor g221 (Z[5], n_267, n_268);
  xnor g223 (Z[6], n_269, n_270);
  xnor g226 (Z[7], n_272, n_273);
  xnor g228 (Z[8], n_222, n_274);
  xnor g231 (Z[9], n_276, n_277);
  xnor g233 (Z[10], n_278, n_279);
  xnor g236 (Z[11], n_281, n_282);
  xnor g239 (Z[12], n_284, n_285);
  xnor g242 (Z[13], n_287, n_288);
  xnor g244 (Z[14], n_289, n_290);
  xnor g247 (Z[15], n_292, n_293);
  xnor g249 (Z[16], n_244, n_294);
  xnor g252 (Z[17], n_296, n_297);
  xnor g254 (Z[18], n_298, n_299);
  xnor g257 (Z[19], n_301, n_302);
  xnor g260 (Z[20], n_304, n_305);
  xnor g263 (Z[21], n_307, n_308);
  and g266 (n_135, A[21], B[21]);
  or g267 (n_136, A[21], B[21]);
  and g268 (n_176, wc, n_124);
  not gc (wc, n_125);
  and g269 (n_183, wc0, n_130);
  not gc0 (wc0, n_131);
  and g270 (n_156, wc1, n_100);
  not gc1 (wc1, n_101);
  and g271 (n_163, wc2, n_106);
  not gc2 (wc2, n_107);
  and g272 (n_166, wc3, n_112);
  not gc3 (wc3, n_113);
  and g273 (n_173, wc4, n_118);
  not gc4 (wc4, n_119);
  and g274 (n_146, wc5, n_88);
  not gc5 (wc5, n_89);
  and g275 (n_153, wc6, n_94);
  not gc6 (wc6, n_95);
  and g276 (n_144, wc7, n_82);
  not gc7 (wc7, n_83);
  or g277 (n_79, n_72, n_75);
  or g278 (n_190, wc8, n_97);
  not gc8 (wc8, n_149);
  or g279 (n_226, wc9, n_109);
  not gc9 (wc9, n_159);
  or g280 (n_205, wc10, n_121);
  not gc10 (wc10, n_169);
  or g281 (n_248, wc11, n_133);
  not gc11 (wc11, n_179);
  or g282 (n_260, wc12, n_75);
  not gc12 (wc12, n_78);
  or g283 (n_261, wc13, n_85);
  not gc13 (wc13, n_80);
  or g284 (n_264, wc14, n_81);
  not gc14 (wc14, n_82);
  or g285 (n_265, wc15, n_91);
  not gc15 (wc15, n_86);
  or g286 (n_268, wc16, n_87);
  not gc16 (wc16, n_88);
  or g287 (n_270, wc17, n_97);
  not gc17 (wc17, n_92);
  or g288 (n_273, wc18, n_93);
  not gc18 (wc18, n_94);
  or g289 (n_274, wc19, n_103);
  not gc19 (wc19, n_98);
  or g290 (n_277, wc20, n_99);
  not gc20 (wc20, n_100);
  or g291 (n_279, wc21, n_109);
  not gc21 (wc21, n_104);
  or g292 (n_282, wc22, n_105);
  not gc22 (wc22, n_106);
  or g293 (n_285, wc23, n_115);
  not gc23 (wc23, n_110);
  or g294 (n_288, wc24, n_111);
  not gc24 (wc24, n_112);
  or g295 (n_290, wc25, n_121);
  not gc25 (wc25, n_116);
  or g296 (n_293, wc26, n_117);
  not gc26 (wc26, n_118);
  or g297 (n_294, wc27, n_127);
  not gc27 (wc27, n_122);
  or g298 (n_297, wc28, n_123);
  not gc28 (wc28, n_124);
  or g299 (n_299, wc29, n_133);
  not gc29 (wc29, n_128);
  or g300 (n_302, wc30, n_129);
  not gc30 (wc30, n_130);
  or g301 (n_305, wc31, n_139);
  not gc31 (wc31, n_134);
  and g302 (n_184, wc32, n_181);
  not gc32 (wc32, n_176);
  and g303 (n_219, n_136, wc33);
  not gc33 (wc33, n_137);
  and g304 (n_164, wc34, n_161);
  not gc34 (wc34, n_156);
  and g305 (n_174, wc35, n_171);
  not gc35 (wc35, n_166);
  and g306 (n_154, wc36, n_151);
  not gc36 (wc36, n_146);
  and g307 (n_235, wc37, n_169);
  not gc37 (wc37, n_201);
  xor g308 (Z[1], n_72, n_260);
  or g309 (n_308, wc38, n_135);
  not gc38 (wc38, n_136);
  and g310 (n_213, wc39, n_183);
  not gc39 (wc39, n_184);
  and g311 (n_257, wc40, n_217);
  not gc40 (wc40, n_216);
  and g312 (n_198, wc41, n_163);
  not gc41 (wc41, n_164);
  and g313 (n_210, wc42, n_173);
  not gc42 (wc42, n_174);
  and g314 (n_196, wc43, n_153);
  not gc43 (wc43, n_154);
  or g315 (n_142, wc44, n_85);
  not gc44 (wc44, n_140);
  and g316 (n_192, wc45, n_92);
  not gc45 (wc45, n_147);
  and g317 (n_228, wc46, n_104);
  not gc46 (wc46, n_157);
  and g318 (n_206, wc47, n_116);
  not gc47 (wc47, n_167);
  and g319 (n_250, wc48, n_128);
  not gc48 (wc48, n_177);
  and g320 (n_220, wc49, n_217);
  not gc49 (wc49, n_213);
  and g321 (n_203, wc50, n_169);
  not gc50 (wc50, n_198);
  and g322 (n_258, wc51, n_219);
  not gc51 (wc51, n_220);
  and g323 (n_242, n_210, wc52);
  not gc52 (wc52, n_211);
  or g324 (n_197, n_194, wc53);
  not gc53 (wc53, n_186);
  or g325 (n_188, wc54, n_91);
  not gc54 (wc54, n_186);
  or g326 (n_193, n_190, wc55);
  not gc55 (wc55, n_186);
  and g327 (n_233, wc56, n_110);
  not gc56 (wc56, n_199);
  and g328 (n_236, wc57, n_166);
  not gc57 (wc57, n_203);
  and g329 (n_239, n_206, wc58);
  not gc58 (wc58, n_207);
  and g330 (n_255, wc59, n_134);
  not gc59 (wc59, n_214);
  or g331 (n_224, wc60, n_103);
  not gc60 (wc60, n_222);
  or g332 (n_229, n_226, wc61);
  not gc61 (wc61, n_222);
  or g333 (n_231, wc62, n_201);
  not gc62 (wc62, n_222);
  or g334 (n_246, wc63, n_127);
  not gc63 (wc63, n_244);
  or g335 (n_251, n_248, wc64);
  not gc64 (wc64, n_244);
  or g336 (n_253, wc65, n_216);
  not gc65 (wc65, n_244);
endmodule

module add_signed_33_GENERIC(A, B, Z);
  input [21:0] A, B;
  output [22:0] Z;
  wire [21:0] A, B;
  wire [22:0] Z;
  add_signed_33_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_62_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [20:0] A, B;
  output [21:0] Z;
  wire [20:0] A, B;
  wire [21:0] Z;
  wire n_68, n_69, n_72, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_82, n_83, n_84, n_85, n_86, n_88, n_89;
  wire n_90, n_91, n_92, n_94, n_95, n_96, n_97, n_98;
  wire n_100, n_101, n_102, n_103, n_104, n_106, n_107, n_108;
  wire n_109, n_110, n_112, n_113, n_114, n_115, n_116, n_118;
  wire n_119, n_120, n_121, n_122, n_124, n_125, n_126, n_127;
  wire n_128, n_130, n_131, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_140, n_142, n_144, n_145, n_147, n_148, n_150;
  wire n_152, n_154, n_155, n_157, n_158, n_160, n_162, n_164;
  wire n_165, n_167, n_168, n_170, n_172, n_174, n_175, n_177;
  wire n_179, n_180, n_181, n_183, n_184, n_185, n_187, n_188;
  wire n_189, n_190, n_192, n_194, n_196, n_197, n_198, n_200;
  wire n_201, n_202, n_204, n_205, n_206, n_207, n_209, n_210;
  wire n_212, n_213, n_214, n_216, n_217, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_234, n_235, n_236, n_238, n_239;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_248, n_249;
  wire n_250, n_252, n_253, n_254, n_255, n_257, n_258, n_259;
  wire n_261, n_262, n_263, n_264, n_266, n_267, n_269, n_270;
  wire n_272, n_273, n_274, n_275, n_277, n_278, n_279, n_281;
  wire n_282, n_283, n_284, n_286, n_287, n_289, n_290;
  not g3 (Z[21], n_68);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_69, A[0], B[0]);
  nor g9 (n_72, A[1], B[1]);
  nand g10 (n_75, A[1], B[1]);
  nor g11 (n_82, A[2], B[2]);
  nand g12 (n_77, A[2], B[2]);
  nor g13 (n_78, A[3], B[3]);
  nand g14 (n_79, A[3], B[3]);
  nor g15 (n_88, A[4], B[4]);
  nand g16 (n_83, A[4], B[4]);
  nor g17 (n_84, A[5], B[5]);
  nand g18 (n_85, A[5], B[5]);
  nor g19 (n_94, A[6], B[6]);
  nand g20 (n_89, A[6], B[6]);
  nor g21 (n_90, A[7], B[7]);
  nand g22 (n_91, A[7], B[7]);
  nor g23 (n_100, A[8], B[8]);
  nand g24 (n_95, A[8], B[8]);
  nor g25 (n_96, A[9], B[9]);
  nand g26 (n_97, A[9], B[9]);
  nor g27 (n_106, A[10], B[10]);
  nand g28 (n_101, A[10], B[10]);
  nor g29 (n_102, A[11], B[11]);
  nand g30 (n_103, A[11], B[11]);
  nor g31 (n_112, A[12], B[12]);
  nand g32 (n_107, A[12], B[12]);
  nor g33 (n_108, A[13], B[13]);
  nand g34 (n_109, A[13], B[13]);
  nor g35 (n_118, A[14], B[14]);
  nand g36 (n_113, A[14], B[14]);
  nor g37 (n_114, A[15], B[15]);
  nand g38 (n_115, A[15], B[15]);
  nor g39 (n_124, A[16], B[16]);
  nand g40 (n_119, A[16], B[16]);
  nor g41 (n_120, A[17], B[17]);
  nand g42 (n_121, A[17], B[17]);
  nor g43 (n_130, A[18], B[18]);
  nand g44 (n_125, A[18], B[18]);
  nor g45 (n_126, A[19], B[19]);
  nand g46 (n_127, A[19], B[19]);
  nand g51 (n_131, n_75, n_76);
  nor g52 (n_80, n_77, n_78);
  nor g55 (n_134, n_82, n_78);
  nor g56 (n_86, n_83, n_84);
  nor g59 (n_140, n_88, n_84);
  nor g60 (n_92, n_89, n_90);
  nor g63 (n_142, n_94, n_90);
  nor g64 (n_98, n_95, n_96);
  nor g67 (n_150, n_100, n_96);
  nor g68 (n_104, n_101, n_102);
  nor g71 (n_152, n_106, n_102);
  nor g72 (n_110, n_107, n_108);
  nor g75 (n_160, n_112, n_108);
  nor g76 (n_116, n_113, n_114);
  nor g79 (n_162, n_118, n_114);
  nor g80 (n_122, n_119, n_120);
  nor g83 (n_170, n_124, n_120);
  nor g84 (n_128, n_125, n_126);
  nor g87 (n_172, n_130, n_126);
  nand g90 (n_248, n_77, n_133);
  nand g91 (n_136, n_134, n_131);
  nand g92 (n_177, n_135, n_136);
  nor g93 (n_138, n_94, n_137);
  nand g102 (n_185, n_140, n_142);
  nor g103 (n_148, n_106, n_147);
  nand g112 (n_192, n_150, n_152);
  nor g113 (n_158, n_118, n_157);
  nand g122 (n_200, n_160, n_162);
  nor g123 (n_168, n_130, n_167);
  nand g132 (n_209, n_170, n_172);
  nand g135 (n_252, n_83, n_179);
  nand g136 (n_180, n_140, n_177);
  nand g137 (n_254, n_137, n_180);
  nand g140 (n_257, n_183, n_184);
  nand g143 (n_210, n_187, n_188);
  nor g144 (n_190, n_112, n_189);
  nor g147 (n_220, n_112, n_192);
  nor g153 (n_198, n_196, n_189);
  nor g156 (n_226, n_192, n_196);
  nor g157 (n_202, n_200, n_189);
  nor g160 (n_229, n_192, n_200);
  nor g161 (n_207, n_204, n_205);
  nor g164 (n_242, n_204, n_209);
  nand g167 (n_261, n_95, n_212);
  nand g168 (n_213, n_150, n_210);
  nand g169 (n_263, n_147, n_213);
  nand g172 (n_266, n_216, n_217);
  nand g175 (n_269, n_189, n_219);
  nand g176 (n_222, n_220, n_210);
  nand g177 (n_272, n_221, n_222);
  nand g178 (n_225, n_223, n_210);
  nand g179 (n_274, n_224, n_225);
  nand g180 (n_228, n_226, n_210);
  nand g181 (n_277, n_227, n_228);
  nand g182 (n_231, n_229, n_210);
  nand g183 (n_232, n_230, n_231);
  nand g186 (n_281, n_119, n_234);
  nand g187 (n_235, n_170, n_232);
  nand g188 (n_283, n_167, n_235);
  nand g191 (n_286, n_238, n_239);
  nand g194 (n_289, n_205, n_241);
  nand g195 (n_244, n_242, n_232);
  nand g196 (n_68, n_243, n_244);
  xnor g200 (Z[2], n_131, n_246);
  xnor g203 (Z[3], n_248, n_249);
  xnor g205 (Z[4], n_177, n_250);
  xnor g208 (Z[5], n_252, n_253);
  xnor g210 (Z[6], n_254, n_255);
  xnor g213 (Z[7], n_257, n_258);
  xnor g215 (Z[8], n_210, n_259);
  xnor g218 (Z[9], n_261, n_262);
  xnor g220 (Z[10], n_263, n_264);
  xnor g223 (Z[11], n_266, n_267);
  xnor g226 (Z[12], n_269, n_270);
  xnor g229 (Z[13], n_272, n_273);
  xnor g231 (Z[14], n_274, n_275);
  xnor g234 (Z[15], n_277, n_278);
  xnor g236 (Z[16], n_232, n_279);
  xnor g239 (Z[17], n_281, n_282);
  xnor g241 (Z[18], n_283, n_284);
  xnor g244 (Z[19], n_286, n_287);
  xnor g247 (Z[20], n_289, n_290);
  and g250 (n_204, A[20], B[20]);
  or g251 (n_206, A[20], B[20]);
  and g252 (n_167, wc, n_121);
  not gc (wc, n_122);
  and g253 (n_174, wc0, n_127);
  not gc0 (wc0, n_128);
  and g254 (n_147, wc1, n_97);
  not gc1 (wc1, n_98);
  and g255 (n_154, wc2, n_103);
  not gc2 (wc2, n_104);
  and g256 (n_157, wc3, n_109);
  not gc3 (wc3, n_110);
  and g257 (n_164, wc4, n_115);
  not gc4 (wc4, n_116);
  and g258 (n_137, wc5, n_85);
  not gc5 (wc5, n_86);
  and g259 (n_144, wc6, n_91);
  not gc6 (wc6, n_92);
  and g260 (n_135, wc7, n_79);
  not gc7 (wc7, n_80);
  or g261 (n_76, n_69, n_72);
  or g262 (n_181, wc8, n_94);
  not gc8 (wc8, n_140);
  or g263 (n_214, wc9, n_106);
  not gc9 (wc9, n_150);
  or g264 (n_196, wc10, n_118);
  not gc10 (wc10, n_160);
  or g265 (n_236, wc11, n_130);
  not gc11 (wc11, n_170);
  or g266 (n_245, wc12, n_72);
  not gc12 (wc12, n_75);
  or g267 (n_246, wc13, n_82);
  not gc13 (wc13, n_77);
  or g268 (n_249, wc14, n_78);
  not gc14 (wc14, n_79);
  or g269 (n_250, wc15, n_88);
  not gc15 (wc15, n_83);
  or g270 (n_253, wc16, n_84);
  not gc16 (wc16, n_85);
  or g271 (n_255, wc17, n_94);
  not gc17 (wc17, n_89);
  or g272 (n_258, wc18, n_90);
  not gc18 (wc18, n_91);
  or g273 (n_259, wc19, n_100);
  not gc19 (wc19, n_95);
  or g274 (n_262, wc20, n_96);
  not gc20 (wc20, n_97);
  or g275 (n_264, wc21, n_106);
  not gc21 (wc21, n_101);
  or g276 (n_267, wc22, n_102);
  not gc22 (wc22, n_103);
  or g277 (n_270, wc23, n_112);
  not gc23 (wc23, n_107);
  or g278 (n_273, wc24, n_108);
  not gc24 (wc24, n_109);
  or g279 (n_275, wc25, n_118);
  not gc25 (wc25, n_113);
  or g280 (n_278, wc26, n_114);
  not gc26 (wc26, n_115);
  or g281 (n_279, wc27, n_124);
  not gc27 (wc27, n_119);
  or g282 (n_282, wc28, n_120);
  not gc28 (wc28, n_121);
  or g283 (n_284, wc29, n_130);
  not gc29 (wc29, n_125);
  or g284 (n_287, wc30, n_126);
  not gc30 (wc30, n_127);
  and g285 (n_175, wc31, n_172);
  not gc31 (wc31, n_167);
  and g286 (n_155, wc32, n_152);
  not gc32 (wc32, n_147);
  and g287 (n_165, wc33, n_162);
  not gc33 (wc33, n_157);
  and g288 (n_145, wc34, n_142);
  not gc34 (wc34, n_137);
  and g289 (n_223, wc35, n_160);
  not gc35 (wc35, n_192);
  xor g290 (Z[1], n_69, n_245);
  or g291 (n_290, wc36, n_204);
  not gc36 (wc36, n_206);
  and g292 (n_205, wc37, n_174);
  not gc37 (wc37, n_175);
  and g293 (n_189, wc38, n_154);
  not gc38 (wc38, n_155);
  and g294 (n_201, wc39, n_164);
  not gc39 (wc39, n_165);
  and g295 (n_187, wc40, n_144);
  not gc40 (wc40, n_145);
  or g296 (n_133, wc41, n_82);
  not gc41 (wc41, n_131);
  and g297 (n_183, wc42, n_89);
  not gc42 (wc42, n_138);
  and g298 (n_216, wc43, n_101);
  not gc43 (wc43, n_148);
  and g299 (n_197, wc44, n_113);
  not gc44 (wc44, n_158);
  and g300 (n_238, wc45, n_125);
  not gc45 (wc45, n_168);
  and g301 (n_194, wc46, n_160);
  not gc46 (wc46, n_189);
  and g302 (n_243, n_206, wc47);
  not gc47 (wc47, n_207);
  and g303 (n_230, n_201, wc48);
  not gc48 (wc48, n_202);
  or g304 (n_188, n_185, wc49);
  not gc49 (wc49, n_177);
  or g305 (n_179, wc50, n_88);
  not gc50 (wc50, n_177);
  or g306 (n_184, n_181, wc51);
  not gc51 (wc51, n_177);
  and g307 (n_221, wc52, n_107);
  not gc52 (wc52, n_190);
  and g308 (n_224, wc53, n_157);
  not gc53 (wc53, n_194);
  and g309 (n_227, n_197, wc54);
  not gc54 (wc54, n_198);
  or g310 (n_212, wc55, n_100);
  not gc55 (wc55, n_210);
  or g311 (n_217, n_214, wc56);
  not gc56 (wc56, n_210);
  or g312 (n_219, wc57, n_192);
  not gc57 (wc57, n_210);
  or g313 (n_234, wc58, n_124);
  not gc58 (wc58, n_232);
  or g314 (n_239, n_236, wc59);
  not gc59 (wc59, n_232);
  or g315 (n_241, wc60, n_209);
  not gc60 (wc60, n_232);
endmodule

module add_signed_62_GENERIC(A, B, Z);
  input [20:0] A, B;
  output [21:0] Z;
  wire [20:0] A, B;
  wire [21:0] Z;
  add_signed_62_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_65_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [21:0] A, B;
  output [22:0] Z;
  wire [21:0] A, B;
  wire [22:0] Z;
  wire n_71, n_72, n_75, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_85, n_86, n_87, n_88, n_89, n_91, n_92;
  wire n_93, n_94, n_95, n_97, n_98, n_99, n_100, n_101;
  wire n_103, n_104, n_105, n_106, n_107, n_109, n_110, n_111;
  wire n_112, n_113, n_115, n_116, n_117, n_118, n_119, n_121;
  wire n_122, n_123, n_124, n_125, n_127, n_128, n_129, n_130;
  wire n_131, n_133, n_134, n_135, n_136, n_137, n_139, n_140;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_149, n_151;
  wire n_153, n_154, n_156, n_157, n_159, n_161, n_163, n_164;
  wire n_166, n_167, n_169, n_171, n_173, n_174, n_176, n_177;
  wire n_179, n_181, n_183, n_184, n_186, n_188, n_189, n_190;
  wire n_192, n_193, n_194, n_196, n_197, n_198, n_199, n_201;
  wire n_203, n_205, n_206, n_207, n_209, n_210, n_211, n_213;
  wire n_214, n_216, n_217, n_219, n_220, n_222, n_224, n_225;
  wire n_226, n_228, n_229, n_231, n_232, n_233, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_246, n_247, n_248, n_250, n_251, n_253, n_254;
  wire n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_263;
  wire n_264, n_265, n_267, n_268, n_269, n_270, n_272, n_273;
  wire n_274, n_276, n_277, n_278, n_279, n_281, n_282, n_284;
  wire n_285, n_287, n_288, n_289, n_290, n_292, n_293, n_294;
  wire n_296, n_297, n_298, n_299, n_301, n_302, n_304, n_305;
  wire n_307, n_308;
  not g3 (Z[22], n_71);
  xor g4 (Z[0], A[0], B[0]);
  nand g5 (n_72, A[0], B[0]);
  nor g9 (n_75, A[1], B[1]);
  nand g10 (n_78, A[1], B[1]);
  nor g11 (n_85, A[2], B[2]);
  nand g12 (n_80, A[2], B[2]);
  nor g13 (n_81, A[3], B[3]);
  nand g14 (n_82, A[3], B[3]);
  nor g15 (n_91, A[4], B[4]);
  nand g16 (n_86, A[4], B[4]);
  nor g17 (n_87, A[5], B[5]);
  nand g18 (n_88, A[5], B[5]);
  nor g19 (n_97, A[6], B[6]);
  nand g20 (n_92, A[6], B[6]);
  nor g21 (n_93, A[7], B[7]);
  nand g22 (n_94, A[7], B[7]);
  nor g23 (n_103, A[8], B[8]);
  nand g24 (n_98, A[8], B[8]);
  nor g25 (n_99, A[9], B[9]);
  nand g26 (n_100, A[9], B[9]);
  nor g27 (n_109, A[10], B[10]);
  nand g28 (n_104, A[10], B[10]);
  nor g29 (n_105, A[11], B[11]);
  nand g30 (n_106, A[11], B[11]);
  nor g31 (n_115, A[12], B[12]);
  nand g32 (n_110, A[12], B[12]);
  nor g33 (n_111, A[13], B[13]);
  nand g34 (n_112, A[13], B[13]);
  nor g35 (n_121, A[14], B[14]);
  nand g36 (n_116, A[14], B[14]);
  nor g37 (n_117, A[15], B[15]);
  nand g38 (n_118, A[15], B[15]);
  nor g39 (n_127, A[16], B[16]);
  nand g40 (n_122, A[16], B[16]);
  nor g41 (n_123, A[17], B[17]);
  nand g42 (n_124, A[17], B[17]);
  nor g43 (n_133, A[18], B[18]);
  nand g44 (n_128, A[18], B[18]);
  nor g45 (n_129, A[19], B[19]);
  nand g46 (n_130, A[19], B[19]);
  nor g47 (n_139, A[20], B[20]);
  nand g48 (n_134, A[20], B[20]);
  nand g53 (n_140, n_78, n_79);
  nor g54 (n_83, n_80, n_81);
  nor g57 (n_143, n_85, n_81);
  nor g58 (n_89, n_86, n_87);
  nor g61 (n_149, n_91, n_87);
  nor g62 (n_95, n_92, n_93);
  nor g65 (n_151, n_97, n_93);
  nor g66 (n_101, n_98, n_99);
  nor g69 (n_159, n_103, n_99);
  nor g70 (n_107, n_104, n_105);
  nor g73 (n_161, n_109, n_105);
  nor g74 (n_113, n_110, n_111);
  nor g77 (n_169, n_115, n_111);
  nor g78 (n_119, n_116, n_117);
  nor g81 (n_171, n_121, n_117);
  nor g82 (n_125, n_122, n_123);
  nor g85 (n_179, n_127, n_123);
  nor g86 (n_131, n_128, n_129);
  nor g89 (n_181, n_133, n_129);
  nor g90 (n_137, n_134, n_135);
  nor g93 (n_217, n_139, n_135);
  nand g96 (n_263, n_80, n_142);
  nand g97 (n_145, n_143, n_140);
  nand g98 (n_186, n_144, n_145);
  nor g99 (n_147, n_97, n_146);
  nand g108 (n_194, n_149, n_151);
  nor g109 (n_157, n_109, n_156);
  nand g118 (n_201, n_159, n_161);
  nor g119 (n_167, n_121, n_166);
  nand g128 (n_209, n_169, n_171);
  nor g129 (n_177, n_133, n_176);
  nand g138 (n_216, n_179, n_181);
  nand g141 (n_267, n_86, n_188);
  nand g142 (n_189, n_149, n_186);
  nand g143 (n_269, n_146, n_189);
  nand g146 (n_272, n_192, n_193);
  nand g149 (n_222, n_196, n_197);
  nor g150 (n_199, n_115, n_198);
  nor g153 (n_232, n_115, n_201);
  nor g159 (n_207, n_205, n_198);
  nor g162 (n_238, n_201, n_205);
  nor g163 (n_211, n_209, n_198);
  nor g166 (n_241, n_201, n_209);
  nor g167 (n_214, n_139, n_213);
  nor g170 (n_254, n_139, n_216);
  nand g178 (n_276, n_98, n_224);
  nand g179 (n_225, n_159, n_222);
  nand g180 (n_278, n_156, n_225);
  nand g183 (n_281, n_228, n_229);
  nand g186 (n_284, n_198, n_231);
  nand g187 (n_234, n_232, n_222);
  nand g188 (n_287, n_233, n_234);
  nand g189 (n_237, n_235, n_222);
  nand g190 (n_289, n_236, n_237);
  nand g191 (n_240, n_238, n_222);
  nand g192 (n_292, n_239, n_240);
  nand g193 (n_243, n_241, n_222);
  nand g194 (n_244, n_242, n_243);
  nand g197 (n_296, n_122, n_246);
  nand g198 (n_247, n_179, n_244);
  nand g199 (n_298, n_176, n_247);
  nand g202 (n_301, n_250, n_251);
  nand g205 (n_304, n_213, n_253);
  nand g206 (n_256, n_254, n_244);
  nand g207 (n_307, n_255, n_256);
  nand g208 (n_259, n_257, n_244);
  nand g209 (n_71, n_258, n_259);
  xnor g213 (Z[2], n_140, n_261);
  xnor g216 (Z[3], n_263, n_264);
  xnor g218 (Z[4], n_186, n_265);
  xnor g221 (Z[5], n_267, n_268);
  xnor g223 (Z[6], n_269, n_270);
  xnor g226 (Z[7], n_272, n_273);
  xnor g228 (Z[8], n_222, n_274);
  xnor g231 (Z[9], n_276, n_277);
  xnor g233 (Z[10], n_278, n_279);
  xnor g236 (Z[11], n_281, n_282);
  xnor g239 (Z[12], n_284, n_285);
  xnor g242 (Z[13], n_287, n_288);
  xnor g244 (Z[14], n_289, n_290);
  xnor g247 (Z[15], n_292, n_293);
  xnor g249 (Z[16], n_244, n_294);
  xnor g252 (Z[17], n_296, n_297);
  xnor g254 (Z[18], n_298, n_299);
  xnor g257 (Z[19], n_301, n_302);
  xnor g260 (Z[20], n_304, n_305);
  xnor g263 (Z[21], n_307, n_308);
  and g266 (n_135, A[21], B[21]);
  or g267 (n_136, A[21], B[21]);
  and g268 (n_176, wc, n_124);
  not gc (wc, n_125);
  and g269 (n_183, wc0, n_130);
  not gc0 (wc0, n_131);
  and g270 (n_156, wc1, n_100);
  not gc1 (wc1, n_101);
  and g271 (n_163, wc2, n_106);
  not gc2 (wc2, n_107);
  and g272 (n_166, wc3, n_112);
  not gc3 (wc3, n_113);
  and g273 (n_173, wc4, n_118);
  not gc4 (wc4, n_119);
  and g274 (n_146, wc5, n_88);
  not gc5 (wc5, n_89);
  and g275 (n_153, wc6, n_94);
  not gc6 (wc6, n_95);
  and g276 (n_144, wc7, n_82);
  not gc7 (wc7, n_83);
  or g277 (n_79, n_72, n_75);
  or g278 (n_190, wc8, n_97);
  not gc8 (wc8, n_149);
  or g279 (n_226, wc9, n_109);
  not gc9 (wc9, n_159);
  or g280 (n_205, wc10, n_121);
  not gc10 (wc10, n_169);
  or g281 (n_248, wc11, n_133);
  not gc11 (wc11, n_179);
  or g282 (n_260, wc12, n_75);
  not gc12 (wc12, n_78);
  or g283 (n_261, wc13, n_85);
  not gc13 (wc13, n_80);
  or g284 (n_264, wc14, n_81);
  not gc14 (wc14, n_82);
  or g285 (n_265, wc15, n_91);
  not gc15 (wc15, n_86);
  or g286 (n_268, wc16, n_87);
  not gc16 (wc16, n_88);
  or g287 (n_270, wc17, n_97);
  not gc17 (wc17, n_92);
  or g288 (n_273, wc18, n_93);
  not gc18 (wc18, n_94);
  or g289 (n_274, wc19, n_103);
  not gc19 (wc19, n_98);
  or g290 (n_277, wc20, n_99);
  not gc20 (wc20, n_100);
  or g291 (n_279, wc21, n_109);
  not gc21 (wc21, n_104);
  or g292 (n_282, wc22, n_105);
  not gc22 (wc22, n_106);
  or g293 (n_285, wc23, n_115);
  not gc23 (wc23, n_110);
  or g294 (n_288, wc24, n_111);
  not gc24 (wc24, n_112);
  or g295 (n_290, wc25, n_121);
  not gc25 (wc25, n_116);
  or g296 (n_293, wc26, n_117);
  not gc26 (wc26, n_118);
  or g297 (n_294, wc27, n_127);
  not gc27 (wc27, n_122);
  or g298 (n_297, wc28, n_123);
  not gc28 (wc28, n_124);
  or g299 (n_299, wc29, n_133);
  not gc29 (wc29, n_128);
  or g300 (n_302, wc30, n_129);
  not gc30 (wc30, n_130);
  or g301 (n_305, wc31, n_139);
  not gc31 (wc31, n_134);
  and g302 (n_184, wc32, n_181);
  not gc32 (wc32, n_176);
  and g303 (n_219, n_136, wc33);
  not gc33 (wc33, n_137);
  and g304 (n_164, wc34, n_161);
  not gc34 (wc34, n_156);
  and g305 (n_174, wc35, n_171);
  not gc35 (wc35, n_166);
  and g306 (n_154, wc36, n_151);
  not gc36 (wc36, n_146);
  and g307 (n_235, wc37, n_169);
  not gc37 (wc37, n_201);
  xor g308 (Z[1], n_72, n_260);
  or g309 (n_308, wc38, n_135);
  not gc38 (wc38, n_136);
  and g310 (n_213, wc39, n_183);
  not gc39 (wc39, n_184);
  and g311 (n_257, wc40, n_217);
  not gc40 (wc40, n_216);
  and g312 (n_198, wc41, n_163);
  not gc41 (wc41, n_164);
  and g313 (n_210, wc42, n_173);
  not gc42 (wc42, n_174);
  and g314 (n_196, wc43, n_153);
  not gc43 (wc43, n_154);
  or g315 (n_142, wc44, n_85);
  not gc44 (wc44, n_140);
  and g316 (n_192, wc45, n_92);
  not gc45 (wc45, n_147);
  and g317 (n_228, wc46, n_104);
  not gc46 (wc46, n_157);
  and g318 (n_206, wc47, n_116);
  not gc47 (wc47, n_167);
  and g319 (n_250, wc48, n_128);
  not gc48 (wc48, n_177);
  and g320 (n_220, wc49, n_217);
  not gc49 (wc49, n_213);
  and g321 (n_203, wc50, n_169);
  not gc50 (wc50, n_198);
  and g322 (n_258, wc51, n_219);
  not gc51 (wc51, n_220);
  and g323 (n_242, n_210, wc52);
  not gc52 (wc52, n_211);
  or g324 (n_197, n_194, wc53);
  not gc53 (wc53, n_186);
  or g325 (n_188, wc54, n_91);
  not gc54 (wc54, n_186);
  or g326 (n_193, n_190, wc55);
  not gc55 (wc55, n_186);
  and g327 (n_233, wc56, n_110);
  not gc56 (wc56, n_199);
  and g328 (n_236, wc57, n_166);
  not gc57 (wc57, n_203);
  and g329 (n_239, n_206, wc58);
  not gc58 (wc58, n_207);
  and g330 (n_255, wc59, n_134);
  not gc59 (wc59, n_214);
  or g331 (n_224, wc60, n_103);
  not gc60 (wc60, n_222);
  or g332 (n_229, n_226, wc61);
  not gc61 (wc61, n_222);
  or g333 (n_231, wc62, n_201);
  not gc62 (wc62, n_222);
  or g334 (n_246, wc63, n_127);
  not gc63 (wc63, n_244);
  or g335 (n_251, n_248, wc64);
  not gc64 (wc64, n_244);
  or g336 (n_253, wc65, n_216);
  not gc65 (wc65, n_244);
endmodule

module add_signed_65_GENERIC(A, B, Z);
  input [21:0] A, B;
  output [22:0] Z;
  wire [21:0] A, B;
  wire [22:0] Z;
  add_signed_65_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_6773_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [26:0] A, B;
  output [24:0] Z;
  wire [26:0] A, B;
  wire [24:0] Z;
  wire n_82, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_204;
  nand g4 (n_82, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_86, A[1], B[1]);
  nand g13 (n_90, n_86, n_87, n_88);
  xor g14 (n_89, A[1], B[1]);
  nand g16 (n_91, A[2], B[2]);
  nand g17 (n_92, A[2], n_90);
  nand g18 (n_93, B[2], n_90);
  nand g19 (n_95, n_91, n_92, n_93);
  xor g20 (n_94, A[2], B[2]);
  xor g21 (Z[2], n_90, n_94);
  nand g22 (n_96, A[3], B[3]);
  nand g23 (n_97, A[3], n_95);
  nand g24 (n_98, B[3], n_95);
  nand g25 (n_100, n_96, n_97, n_98);
  xor g26 (n_99, A[3], B[3]);
  xor g27 (Z[3], n_95, n_99);
  nand g28 (n_101, A[4], B[4]);
  nand g29 (n_102, A[4], n_100);
  nand g30 (n_103, B[4], n_100);
  nand g31 (n_105, n_101, n_102, n_103);
  xor g32 (n_104, A[4], B[4]);
  xor g33 (Z[4], n_100, n_104);
  nand g34 (n_106, A[5], B[5]);
  nand g35 (n_107, A[5], n_105);
  nand g36 (n_108, B[5], n_105);
  nand g37 (n_110, n_106, n_107, n_108);
  xor g38 (n_109, A[5], B[5]);
  xor g39 (Z[5], n_105, n_109);
  nand g40 (n_111, A[6], B[6]);
  nand g41 (n_112, A[6], n_110);
  nand g42 (n_113, B[6], n_110);
  nand g43 (n_115, n_111, n_112, n_113);
  xor g44 (n_114, A[6], B[6]);
  xor g45 (Z[6], n_110, n_114);
  nand g46 (n_116, A[7], B[7]);
  nand g47 (n_117, A[7], n_115);
  nand g48 (n_118, B[7], n_115);
  nand g49 (n_120, n_116, n_117, n_118);
  xor g50 (n_119, A[7], B[7]);
  xor g51 (Z[7], n_115, n_119);
  nand g52 (n_121, A[8], B[8]);
  nand g53 (n_122, A[8], n_120);
  nand g54 (n_123, B[8], n_120);
  nand g55 (n_125, n_121, n_122, n_123);
  xor g56 (n_124, A[8], B[8]);
  xor g57 (Z[8], n_120, n_124);
  nand g58 (n_126, A[9], B[9]);
  nand g59 (n_127, A[9], n_125);
  nand g60 (n_128, B[9], n_125);
  nand g61 (n_130, n_126, n_127, n_128);
  xor g62 (n_129, A[9], B[9]);
  xor g63 (Z[9], n_125, n_129);
  nand g64 (n_131, A[10], B[10]);
  nand g65 (n_132, A[10], n_130);
  nand g66 (n_133, B[10], n_130);
  nand g67 (n_135, n_131, n_132, n_133);
  xor g68 (n_134, A[10], B[10]);
  xor g69 (Z[10], n_130, n_134);
  nand g70 (n_136, A[11], B[11]);
  nand g71 (n_137, A[11], n_135);
  nand g72 (n_138, B[11], n_135);
  nand g73 (n_140, n_136, n_137, n_138);
  xor g74 (n_139, A[11], B[11]);
  xor g75 (Z[11], n_135, n_139);
  nand g76 (n_141, A[12], B[12]);
  nand g77 (n_142, A[12], n_140);
  nand g78 (n_143, B[12], n_140);
  nand g79 (n_145, n_141, n_142, n_143);
  xor g80 (n_144, A[12], B[12]);
  xor g81 (Z[12], n_140, n_144);
  nand g82 (n_146, A[13], B[13]);
  nand g83 (n_147, A[13], n_145);
  nand g84 (n_148, B[13], n_145);
  nand g85 (n_150, n_146, n_147, n_148);
  xor g86 (n_149, A[13], B[13]);
  xor g87 (Z[13], n_145, n_149);
  nand g88 (n_151, A[14], B[14]);
  nand g89 (n_152, A[14], n_150);
  nand g90 (n_153, B[14], n_150);
  nand g91 (n_155, n_151, n_152, n_153);
  xor g92 (n_154, A[14], B[14]);
  xor g93 (Z[14], n_150, n_154);
  nand g94 (n_156, A[15], B[15]);
  nand g95 (n_157, A[15], n_155);
  nand g96 (n_158, B[15], n_155);
  nand g97 (n_160, n_156, n_157, n_158);
  xor g98 (n_159, A[15], B[15]);
  xor g99 (Z[15], n_155, n_159);
  nand g100 (n_161, A[16], B[16]);
  nand g101 (n_162, A[16], n_160);
  nand g102 (n_163, B[16], n_160);
  nand g103 (n_165, n_161, n_162, n_163);
  xor g104 (n_164, A[16], B[16]);
  xor g105 (Z[16], n_160, n_164);
  nand g106 (n_166, A[17], B[17]);
  nand g107 (n_167, A[17], n_165);
  nand g108 (n_168, B[17], n_165);
  nand g109 (n_170, n_166, n_167, n_168);
  xor g110 (n_169, A[17], B[17]);
  xor g111 (Z[17], n_165, n_169);
  nand g112 (n_171, A[18], B[18]);
  nand g113 (n_172, A[18], n_170);
  nand g114 (n_173, B[18], n_170);
  nand g115 (n_175, n_171, n_172, n_173);
  xor g116 (n_174, A[18], B[18]);
  xor g117 (Z[18], n_170, n_174);
  nand g118 (n_176, A[19], B[19]);
  nand g119 (n_177, A[19], n_175);
  nand g120 (n_178, B[19], n_175);
  nand g121 (n_180, n_176, n_177, n_178);
  xor g122 (n_179, A[19], B[19]);
  xor g123 (Z[19], n_175, n_179);
  nand g124 (n_181, A[20], B[20]);
  nand g125 (n_182, A[20], n_180);
  nand g126 (n_183, B[20], n_180);
  nand g127 (n_185, n_181, n_182, n_183);
  xor g128 (n_184, A[20], B[20]);
  xor g129 (Z[20], n_180, n_184);
  nand g130 (n_186, A[21], B[21]);
  nand g131 (n_187, A[21], n_185);
  nand g132 (n_188, B[21], n_185);
  nand g133 (n_190, n_186, n_187, n_188);
  xor g134 (n_189, A[21], B[21]);
  xor g135 (Z[21], n_185, n_189);
  nand g136 (n_191, A[22], B[22]);
  nand g137 (n_192, A[22], n_190);
  nand g138 (n_193, B[22], n_190);
  nand g139 (n_195, n_191, n_192, n_193);
  xor g140 (n_194, A[22], B[22]);
  xor g141 (Z[22], n_190, n_194);
  nand g142 (n_196, A[23], B[23]);
  nand g143 (n_197, A[23], n_195);
  nand g144 (n_198, B[23], n_195);
  nand g145 (n_200, n_196, n_197, n_198);
  xor g146 (n_199, A[23], B[23]);
  xor g147 (Z[23], n_195, n_199);
  xor g153 (Z[24], n_200, n_204);
  xor g155 (n_204, A[24], B[24]);
  or g156 (n_87, wc, n_82);
  not gc (wc, A[1]);
  or g157 (n_88, wc0, n_82);
  not gc0 (wc0, B[1]);
  xnor g158 (Z[1], n_82, n_89);
endmodule

module add_signed_6773_GENERIC(A, B, Z);
  input [26:0] A, B;
  output [24:0] Z;
  wire [26:0] A, B;
  wire [24:0] Z;
  add_signed_6773_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_carry_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_signed_carry
  input [20:0] A, B;
  input CI;
  output [20:0] Z;
  wire [20:0] A, B;
  wire CI;
  wire [20:0] Z;
  wire n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_172;
  nand g4 (n_69, A[0], B[0]);
  nand g5 (n_70, A[0], CI);
  nand g6 (n_71, B[0], CI);
  nand g7 (n_73, n_69, n_70, n_71);
  xor g8 (n_72, A[0], B[0]);
  xor g9 (Z[0], CI, n_72);
  nand g10 (n_74, A[1], B[1]);
  nand g11 (n_75, A[1], n_73);
  nand g12 (n_76, B[1], n_73);
  nand g13 (n_78, n_74, n_75, n_76);
  xor g14 (n_77, A[1], B[1]);
  xor g15 (Z[1], n_73, n_77);
  nand g16 (n_79, A[2], B[2]);
  nand g17 (n_80, A[2], n_78);
  nand g18 (n_81, B[2], n_78);
  nand g19 (n_83, n_79, n_80, n_81);
  xor g20 (n_82, A[2], B[2]);
  xor g21 (Z[2], n_78, n_82);
  nand g22 (n_84, A[3], B[3]);
  nand g23 (n_85, A[3], n_83);
  nand g24 (n_86, B[3], n_83);
  nand g25 (n_88, n_84, n_85, n_86);
  xor g26 (n_87, A[3], B[3]);
  xor g27 (Z[3], n_83, n_87);
  nand g28 (n_89, A[4], B[4]);
  nand g29 (n_90, A[4], n_88);
  nand g30 (n_91, B[4], n_88);
  nand g31 (n_93, n_89, n_90, n_91);
  xor g32 (n_92, A[4], B[4]);
  xor g33 (Z[4], n_88, n_92);
  nand g34 (n_94, A[5], B[5]);
  nand g35 (n_95, A[5], n_93);
  nand g36 (n_96, B[5], n_93);
  nand g37 (n_98, n_94, n_95, n_96);
  xor g38 (n_97, A[5], B[5]);
  xor g39 (Z[5], n_93, n_97);
  nand g40 (n_99, A[6], B[6]);
  nand g41 (n_100, A[6], n_98);
  nand g42 (n_101, B[6], n_98);
  nand g43 (n_103, n_99, n_100, n_101);
  xor g44 (n_102, A[6], B[6]);
  xor g45 (Z[6], n_98, n_102);
  nand g46 (n_104, A[7], B[7]);
  nand g47 (n_105, A[7], n_103);
  nand g48 (n_106, B[7], n_103);
  nand g49 (n_108, n_104, n_105, n_106);
  xor g50 (n_107, A[7], B[7]);
  xor g51 (Z[7], n_103, n_107);
  nand g52 (n_109, A[8], B[8]);
  nand g53 (n_110, A[8], n_108);
  nand g54 (n_111, B[8], n_108);
  nand g55 (n_113, n_109, n_110, n_111);
  xor g56 (n_112, A[8], B[8]);
  xor g57 (Z[8], n_108, n_112);
  nand g58 (n_114, A[9], B[9]);
  nand g59 (n_115, A[9], n_113);
  nand g60 (n_116, B[9], n_113);
  nand g61 (n_118, n_114, n_115, n_116);
  xor g62 (n_117, A[9], B[9]);
  xor g63 (Z[9], n_113, n_117);
  nand g64 (n_119, A[10], B[10]);
  nand g65 (n_120, A[10], n_118);
  nand g66 (n_121, B[10], n_118);
  nand g67 (n_123, n_119, n_120, n_121);
  xor g68 (n_122, A[10], B[10]);
  xor g69 (Z[10], n_118, n_122);
  nand g70 (n_124, A[11], B[11]);
  nand g71 (n_125, A[11], n_123);
  nand g72 (n_126, B[11], n_123);
  nand g73 (n_128, n_124, n_125, n_126);
  xor g74 (n_127, A[11], B[11]);
  xor g75 (Z[11], n_123, n_127);
  nand g76 (n_129, A[12], B[12]);
  nand g77 (n_130, A[12], n_128);
  nand g78 (n_131, B[12], n_128);
  nand g79 (n_133, n_129, n_130, n_131);
  xor g80 (n_132, A[12], B[12]);
  xor g81 (Z[12], n_128, n_132);
  nand g82 (n_134, A[13], B[13]);
  nand g83 (n_135, A[13], n_133);
  nand g84 (n_136, B[13], n_133);
  nand g85 (n_138, n_134, n_135, n_136);
  xor g86 (n_137, A[13], B[13]);
  xor g87 (Z[13], n_133, n_137);
  nand g88 (n_139, A[14], B[14]);
  nand g89 (n_140, A[14], n_138);
  nand g90 (n_141, B[14], n_138);
  nand g91 (n_143, n_139, n_140, n_141);
  xor g92 (n_142, A[14], B[14]);
  xor g93 (Z[14], n_138, n_142);
  nand g94 (n_144, A[15], B[15]);
  nand g95 (n_145, A[15], n_143);
  nand g96 (n_146, B[15], n_143);
  nand g97 (n_148, n_144, n_145, n_146);
  xor g98 (n_147, A[15], B[15]);
  xor g99 (Z[15], n_143, n_147);
  nand g100 (n_149, A[16], B[16]);
  nand g101 (n_150, A[16], n_148);
  nand g102 (n_151, B[16], n_148);
  nand g103 (n_153, n_149, n_150, n_151);
  xor g104 (n_152, A[16], B[16]);
  xor g105 (Z[16], n_148, n_152);
  nand g106 (n_154, A[17], B[17]);
  nand g107 (n_155, A[17], n_153);
  nand g108 (n_156, B[17], n_153);
  nand g109 (n_158, n_154, n_155, n_156);
  xor g110 (n_157, A[17], B[17]);
  xor g111 (Z[17], n_153, n_157);
  nand g112 (n_159, A[18], B[18]);
  nand g113 (n_160, A[18], n_158);
  nand g114 (n_161, B[18], n_158);
  nand g115 (n_163, n_159, n_160, n_161);
  xor g116 (n_162, A[18], B[18]);
  xor g117 (Z[18], n_158, n_162);
  nand g118 (n_164, A[19], B[19]);
  nand g119 (n_165, A[19], n_163);
  nand g120 (n_166, B[19], n_163);
  nand g121 (n_168, n_164, n_165, n_166);
  xor g122 (n_167, A[19], B[19]);
  xor g123 (Z[19], n_163, n_167);
  xor g129 (Z[20], n_168, n_172);
  xor g130 (n_172, A[20], B[20]);
endmodule

module add_signed_carry_GENERIC(A, B, CI, Z);
  input [20:0] A, B;
  input CI;
  output [20:0] Z;
  wire [20:0] A, B;
  wire CI;
  wire [20:0] Z;
  add_signed_carry_GENERIC_REAL g1(.A ({A[19], A[19:0]}), .B ({B[19],
       B[19:0]}), .CI (CI), .Z (Z));
endmodule

module add_signed_carry_3208_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_signed_carry
  input [21:0] A, B;
  input CI;
  output [21:0] Z;
  wire [21:0] A, B;
  wire CI;
  wire [21:0] Z;
  wire n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_180;
  nand g4 (n_72, A[0], B[0]);
  nand g5 (n_73, A[0], CI);
  nand g6 (n_74, B[0], CI);
  nand g7 (n_76, n_72, n_73, n_74);
  xor g8 (n_75, A[0], B[0]);
  xor g9 (Z[0], CI, n_75);
  nand g10 (n_77, A[1], B[1]);
  nand g11 (n_78, A[1], n_76);
  nand g12 (n_79, B[1], n_76);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  xor g15 (Z[1], n_76, n_80);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_117, A[9], B[9]);
  nand g59 (n_118, A[9], n_116);
  nand g60 (n_119, B[9], n_116);
  nand g61 (n_121, n_117, n_118, n_119);
  xor g62 (n_120, A[9], B[9]);
  xor g63 (Z[9], n_116, n_120);
  nand g64 (n_122, A[10], B[10]);
  nand g65 (n_123, A[10], n_121);
  nand g66 (n_124, B[10], n_121);
  nand g67 (n_126, n_122, n_123, n_124);
  xor g68 (n_125, A[10], B[10]);
  xor g69 (Z[10], n_121, n_125);
  nand g70 (n_127, A[11], B[11]);
  nand g71 (n_128, A[11], n_126);
  nand g72 (n_129, B[11], n_126);
  nand g73 (n_131, n_127, n_128, n_129);
  xor g74 (n_130, A[11], B[11]);
  xor g75 (Z[11], n_126, n_130);
  nand g76 (n_132, A[12], B[12]);
  nand g77 (n_133, A[12], n_131);
  nand g78 (n_134, B[12], n_131);
  nand g79 (n_136, n_132, n_133, n_134);
  xor g80 (n_135, A[12], B[12]);
  xor g81 (Z[12], n_131, n_135);
  nand g82 (n_137, A[13], B[13]);
  nand g83 (n_138, A[13], n_136);
  nand g84 (n_139, B[13], n_136);
  nand g85 (n_141, n_137, n_138, n_139);
  xor g86 (n_140, A[13], B[13]);
  xor g87 (Z[13], n_136, n_140);
  nand g88 (n_142, A[14], B[14]);
  nand g89 (n_143, A[14], n_141);
  nand g90 (n_144, B[14], n_141);
  nand g91 (n_146, n_142, n_143, n_144);
  xor g92 (n_145, A[14], B[14]);
  xor g93 (Z[14], n_141, n_145);
  nand g94 (n_147, A[15], B[15]);
  nand g95 (n_148, A[15], n_146);
  nand g96 (n_149, B[15], n_146);
  nand g97 (n_151, n_147, n_148, n_149);
  xor g98 (n_150, A[15], B[15]);
  xor g99 (Z[15], n_146, n_150);
  nand g100 (n_152, A[16], B[16]);
  nand g101 (n_153, A[16], n_151);
  nand g102 (n_154, B[16], n_151);
  nand g103 (n_156, n_152, n_153, n_154);
  xor g104 (n_155, A[16], B[16]);
  xor g105 (Z[16], n_151, n_155);
  nand g106 (n_157, A[17], B[17]);
  nand g107 (n_158, A[17], n_156);
  nand g108 (n_159, B[17], n_156);
  nand g109 (n_161, n_157, n_158, n_159);
  xor g110 (n_160, A[17], B[17]);
  xor g111 (Z[17], n_156, n_160);
  nand g112 (n_162, A[18], B[18]);
  nand g113 (n_163, A[18], n_161);
  nand g114 (n_164, B[18], n_161);
  nand g115 (n_166, n_162, n_163, n_164);
  xor g116 (n_165, A[18], B[18]);
  xor g117 (Z[18], n_161, n_165);
  nand g118 (n_167, A[19], B[19]);
  nand g119 (n_168, A[19], n_166);
  nand g120 (n_169, B[19], n_166);
  nand g121 (n_171, n_167, n_168, n_169);
  xor g122 (n_170, A[19], B[19]);
  xor g123 (Z[19], n_166, n_170);
  nand g124 (n_172, A[20], B[20]);
  nand g125 (n_173, A[20], n_171);
  nand g126 (n_174, B[20], n_171);
  nand g127 (n_176, n_172, n_173, n_174);
  xor g128 (n_175, A[20], B[20]);
  xor g129 (Z[20], n_171, n_175);
  xor g135 (Z[21], n_176, n_180);
  xor g136 (n_180, A[21], B[21]);
endmodule

module add_signed_carry_3208_GENERIC(A, B, CI, Z);
  input [21:0] A, B;
  input CI;
  output [21:0] Z;
  wire [21:0] A, B;
  wire CI;
  wire [21:0] Z;
  add_signed_carry_3208_GENERIC_REAL g1(.A ({A[20], A[20:0]}), .B
       ({B[20], B[20:0]}), .CI (CI), .Z (Z));
endmodule

module add_signed_carry_3208_1_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_signed_carry
  input [21:0] A, B;
  input CI;
  output [21:0] Z;
  wire [21:0] A, B;
  wire CI;
  wire [21:0] Z;
  wire n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_180;
  nand g4 (n_72, A[0], B[0]);
  nand g5 (n_73, A[0], CI);
  nand g6 (n_74, B[0], CI);
  nand g7 (n_76, n_72, n_73, n_74);
  xor g8 (n_75, A[0], B[0]);
  xor g9 (Z[0], CI, n_75);
  nand g10 (n_77, A[1], B[1]);
  nand g11 (n_78, A[1], n_76);
  nand g12 (n_79, B[1], n_76);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  xor g15 (Z[1], n_76, n_80);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_117, A[9], B[9]);
  nand g59 (n_118, A[9], n_116);
  nand g60 (n_119, B[9], n_116);
  nand g61 (n_121, n_117, n_118, n_119);
  xor g62 (n_120, A[9], B[9]);
  xor g63 (Z[9], n_116, n_120);
  nand g64 (n_122, A[10], B[10]);
  nand g65 (n_123, A[10], n_121);
  nand g66 (n_124, B[10], n_121);
  nand g67 (n_126, n_122, n_123, n_124);
  xor g68 (n_125, A[10], B[10]);
  xor g69 (Z[10], n_121, n_125);
  nand g70 (n_127, A[11], B[11]);
  nand g71 (n_128, A[11], n_126);
  nand g72 (n_129, B[11], n_126);
  nand g73 (n_131, n_127, n_128, n_129);
  xor g74 (n_130, A[11], B[11]);
  xor g75 (Z[11], n_126, n_130);
  nand g76 (n_132, A[12], B[12]);
  nand g77 (n_133, A[12], n_131);
  nand g78 (n_134, B[12], n_131);
  nand g79 (n_136, n_132, n_133, n_134);
  xor g80 (n_135, A[12], B[12]);
  xor g81 (Z[12], n_131, n_135);
  nand g82 (n_137, A[13], B[13]);
  nand g83 (n_138, A[13], n_136);
  nand g84 (n_139, B[13], n_136);
  nand g85 (n_141, n_137, n_138, n_139);
  xor g86 (n_140, A[13], B[13]);
  xor g87 (Z[13], n_136, n_140);
  nand g88 (n_142, A[14], B[14]);
  nand g89 (n_143, A[14], n_141);
  nand g90 (n_144, B[14], n_141);
  nand g91 (n_146, n_142, n_143, n_144);
  xor g92 (n_145, A[14], B[14]);
  xor g93 (Z[14], n_141, n_145);
  nand g94 (n_147, A[15], B[15]);
  nand g95 (n_148, A[15], n_146);
  nand g96 (n_149, B[15], n_146);
  nand g97 (n_151, n_147, n_148, n_149);
  xor g98 (n_150, A[15], B[15]);
  xor g99 (Z[15], n_146, n_150);
  nand g100 (n_152, A[16], B[16]);
  nand g101 (n_153, A[16], n_151);
  nand g102 (n_154, B[16], n_151);
  nand g103 (n_156, n_152, n_153, n_154);
  xor g104 (n_155, A[16], B[16]);
  xor g105 (Z[16], n_151, n_155);
  nand g106 (n_157, A[17], B[17]);
  nand g107 (n_158, A[17], n_156);
  nand g108 (n_159, B[17], n_156);
  nand g109 (n_161, n_157, n_158, n_159);
  xor g110 (n_160, A[17], B[17]);
  xor g111 (Z[17], n_156, n_160);
  nand g112 (n_162, A[18], B[18]);
  nand g113 (n_163, A[18], n_161);
  nand g114 (n_164, B[18], n_161);
  nand g115 (n_166, n_162, n_163, n_164);
  xor g116 (n_165, A[18], B[18]);
  xor g117 (Z[18], n_161, n_165);
  nand g118 (n_167, A[19], B[19]);
  nand g119 (n_168, A[19], n_166);
  nand g120 (n_169, B[19], n_166);
  nand g121 (n_171, n_167, n_168, n_169);
  xor g122 (n_170, A[19], B[19]);
  xor g123 (Z[19], n_166, n_170);
  nand g124 (n_172, A[20], B[20]);
  nand g125 (n_173, A[20], n_171);
  nand g126 (n_174, B[20], n_171);
  nand g127 (n_176, n_172, n_173, n_174);
  xor g128 (n_175, A[20], B[20]);
  xor g129 (Z[20], n_171, n_175);
  xor g135 (Z[21], n_176, n_180);
  xor g136 (n_180, A[21], B[21]);
endmodule

module add_signed_carry_3208_1_GENERIC(A, B, CI, Z);
  input [21:0] A, B;
  input CI;
  output [21:0] Z;
  wire [21:0] A, B;
  wire CI;
  wire [21:0] Z;
  add_signed_carry_3208_1_GENERIC_REAL g1(.A ({A[20], A[20:0]}), .B
       ({B[20], B[20:0]}), .CI (CI), .Z (Z));
endmodule

module add_signed_carry_6718_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_signed_carry
  input [22:0] A, B;
  input CI;
  output [22:0] Z;
  wire [22:0] A, B;
  wire CI;
  wire [22:0] Z;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_188;
  nand g4 (n_75, A[0], B[0]);
  nand g5 (n_76, A[0], CI);
  nand g6 (n_77, B[0], CI);
  nand g7 (n_79, n_75, n_76, n_77);
  xor g8 (n_78, A[0], B[0]);
  xor g9 (Z[0], CI, n_78);
  nand g10 (n_80, A[1], B[1]);
  nand g11 (n_81, A[1], n_79);
  nand g12 (n_82, B[1], n_79);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  xor g15 (Z[1], n_79, n_83);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_120, A[9], B[9]);
  nand g59 (n_121, A[9], n_119);
  nand g60 (n_122, B[9], n_119);
  nand g61 (n_124, n_120, n_121, n_122);
  xor g62 (n_123, A[9], B[9]);
  xor g63 (Z[9], n_119, n_123);
  nand g64 (n_125, A[10], B[10]);
  nand g65 (n_126, A[10], n_124);
  nand g66 (n_127, B[10], n_124);
  nand g67 (n_129, n_125, n_126, n_127);
  xor g68 (n_128, A[10], B[10]);
  xor g69 (Z[10], n_124, n_128);
  nand g70 (n_130, A[11], B[11]);
  nand g71 (n_131, A[11], n_129);
  nand g72 (n_132, B[11], n_129);
  nand g73 (n_134, n_130, n_131, n_132);
  xor g74 (n_133, A[11], B[11]);
  xor g75 (Z[11], n_129, n_133);
  nand g76 (n_135, A[12], B[12]);
  nand g77 (n_136, A[12], n_134);
  nand g78 (n_137, B[12], n_134);
  nand g79 (n_139, n_135, n_136, n_137);
  xor g80 (n_138, A[12], B[12]);
  xor g81 (Z[12], n_134, n_138);
  nand g82 (n_140, A[13], B[13]);
  nand g83 (n_141, A[13], n_139);
  nand g84 (n_142, B[13], n_139);
  nand g85 (n_144, n_140, n_141, n_142);
  xor g86 (n_143, A[13], B[13]);
  xor g87 (Z[13], n_139, n_143);
  nand g88 (n_145, A[14], B[14]);
  nand g89 (n_146, A[14], n_144);
  nand g90 (n_147, B[14], n_144);
  nand g91 (n_149, n_145, n_146, n_147);
  xor g92 (n_148, A[14], B[14]);
  xor g93 (Z[14], n_144, n_148);
  nand g94 (n_150, A[15], B[15]);
  nand g95 (n_151, A[15], n_149);
  nand g96 (n_152, B[15], n_149);
  nand g97 (n_154, n_150, n_151, n_152);
  xor g98 (n_153, A[15], B[15]);
  xor g99 (Z[15], n_149, n_153);
  nand g100 (n_155, A[16], B[16]);
  nand g101 (n_156, A[16], n_154);
  nand g102 (n_157, B[16], n_154);
  nand g103 (n_159, n_155, n_156, n_157);
  xor g104 (n_158, A[16], B[16]);
  xor g105 (Z[16], n_154, n_158);
  nand g106 (n_160, A[17], B[17]);
  nand g107 (n_161, A[17], n_159);
  nand g108 (n_162, B[17], n_159);
  nand g109 (n_164, n_160, n_161, n_162);
  xor g110 (n_163, A[17], B[17]);
  xor g111 (Z[17], n_159, n_163);
  nand g112 (n_165, A[18], B[18]);
  nand g113 (n_166, A[18], n_164);
  nand g114 (n_167, B[18], n_164);
  nand g115 (n_169, n_165, n_166, n_167);
  xor g116 (n_168, A[18], B[18]);
  xor g117 (Z[18], n_164, n_168);
  nand g118 (n_170, A[19], B[19]);
  nand g119 (n_171, A[19], n_169);
  nand g120 (n_172, B[19], n_169);
  nand g121 (n_174, n_170, n_171, n_172);
  xor g122 (n_173, A[19], B[19]);
  xor g123 (Z[19], n_169, n_173);
  nand g124 (n_175, A[20], B[20]);
  nand g125 (n_176, A[20], n_174);
  nand g126 (n_177, B[20], n_174);
  nand g127 (n_179, n_175, n_176, n_177);
  xor g128 (n_178, A[20], B[20]);
  xor g129 (Z[20], n_174, n_178);
  nand g130 (n_180, A[21], B[21]);
  nand g131 (n_181, A[21], n_179);
  nand g132 (n_182, B[21], n_179);
  nand g133 (n_184, n_180, n_181, n_182);
  xor g134 (n_183, A[21], B[21]);
  xor g135 (Z[21], n_179, n_183);
  xor g141 (Z[22], n_184, n_188);
  xor g142 (n_188, A[22], B[22]);
endmodule

module add_signed_carry_6718_GENERIC(A, B, CI, Z);
  input [22:0] A, B;
  input CI;
  output [22:0] Z;
  wire [22:0] A, B;
  wire CI;
  wire [22:0] Z;
  add_signed_carry_6718_GENERIC_REAL g1(.A ({A[21], A[21:0]}), .B
       ({B[21], B[21:0]}), .CI (CI), .Z (Z));
endmodule

module csa_tree_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 24'b0;"
  input [20:0] in_0, in_1, in_2;
  output [23:0] out_0, out_1;
  wire [20:0] in_0, in_1, in_2;
  wire [23:0] out_0, out_1;
  wire n_67, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_194;
  assign out_1[22] = 1'b0;
  assign out_1[23] = 1'b0;
  assign out_0[0] = in_1[0];
  assign out_0[22] = 1'b1;
  assign out_0[23] = 1'b1;
  xor g26 (out_1[0], in_0[0], in_2[0]);
  and g27 (out_0[1], in_0[0], in_2[0]);
  xor g28 (n_116, in_0[1], in_1[1]);
  xor g29 (out_1[1], n_116, in_2[1]);
  nand g30 (n_117, in_0[1], in_1[1]);
  nand g4 (n_118, in_2[1], in_1[1]);
  nand g5 (n_119, in_0[1], in_2[1]);
  nand g31 (out_0[2], n_117, n_118, n_119);
  xor g32 (n_120, in_0[2], in_1[2]);
  xor g33 (out_1[2], n_120, in_2[2]);
  nand g34 (n_121, in_0[2], in_1[2]);
  nand g35 (n_122, in_2[2], in_1[2]);
  nand g36 (n_123, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_121, n_122, n_123);
  xor g37 (n_124, in_0[3], in_1[3]);
  xor g38 (out_1[3], n_124, in_2[3]);
  nand g39 (n_125, in_0[3], in_1[3]);
  nand g40 (n_126, in_2[3], in_1[3]);
  nand g41 (n_127, in_0[3], in_2[3]);
  nand g42 (out_0[4], n_125, n_126, n_127);
  xor g43 (n_128, in_0[4], in_1[4]);
  xor g44 (out_1[4], n_128, in_2[4]);
  nand g45 (n_129, in_0[4], in_1[4]);
  nand g46 (n_130, in_2[4], in_1[4]);
  nand g47 (n_131, in_0[4], in_2[4]);
  nand g48 (out_0[5], n_129, n_130, n_131);
  xor g49 (n_132, in_0[5], in_1[5]);
  xor g50 (out_1[5], n_132, in_2[5]);
  nand g51 (n_133, in_0[5], in_1[5]);
  nand g52 (n_134, in_2[5], in_1[5]);
  nand g53 (n_135, in_0[5], in_2[5]);
  nand g54 (out_0[6], n_133, n_134, n_135);
  xor g55 (n_136, in_0[6], in_1[6]);
  xor g56 (out_1[6], n_136, in_2[6]);
  nand g57 (n_137, in_0[6], in_1[6]);
  nand g58 (n_138, in_2[6], in_1[6]);
  nand g59 (n_139, in_0[6], in_2[6]);
  nand g60 (out_0[7], n_137, n_138, n_139);
  xor g61 (n_140, in_0[7], in_1[7]);
  xor g62 (out_1[7], n_140, in_2[7]);
  nand g63 (n_141, in_0[7], in_1[7]);
  nand g64 (n_142, in_2[7], in_1[7]);
  nand g65 (n_143, in_0[7], in_2[7]);
  nand g66 (out_0[8], n_141, n_142, n_143);
  xor g67 (n_144, in_0[8], in_1[8]);
  xor g68 (out_1[8], n_144, in_2[8]);
  nand g69 (n_145, in_0[8], in_1[8]);
  nand g70 (n_146, in_2[8], in_1[8]);
  nand g71 (n_147, in_0[8], in_2[8]);
  nand g72 (out_0[9], n_145, n_146, n_147);
  xor g73 (n_148, in_0[9], in_1[9]);
  xor g74 (out_1[9], n_148, in_2[9]);
  nand g75 (n_149, in_0[9], in_1[9]);
  nand g76 (n_150, in_2[9], in_1[9]);
  nand g77 (n_151, in_0[9], in_2[9]);
  nand g78 (out_0[10], n_149, n_150, n_151);
  xor g79 (n_152, in_0[10], in_1[10]);
  xor g80 (out_1[10], n_152, in_2[10]);
  nand g81 (n_153, in_0[10], in_1[10]);
  nand g82 (n_154, in_2[10], in_1[10]);
  nand g83 (n_155, in_0[10], in_2[10]);
  nand g84 (out_0[11], n_153, n_154, n_155);
  xor g85 (n_156, in_0[11], in_1[11]);
  xor g86 (out_1[11], n_156, in_2[11]);
  nand g87 (n_157, in_0[11], in_1[11]);
  nand g88 (n_158, in_2[11], in_1[11]);
  nand g89 (n_159, in_0[11], in_2[11]);
  nand g90 (out_0[12], n_157, n_158, n_159);
  xor g91 (n_160, in_0[12], in_1[12]);
  xor g92 (out_1[12], n_160, in_2[12]);
  nand g93 (n_161, in_0[12], in_1[12]);
  nand g94 (n_162, in_2[12], in_1[12]);
  nand g95 (n_163, in_0[12], in_2[12]);
  nand g96 (out_0[13], n_161, n_162, n_163);
  xor g97 (n_164, in_0[13], in_1[13]);
  xor g98 (out_1[13], n_164, in_2[13]);
  nand g99 (n_165, in_0[13], in_1[13]);
  nand g100 (n_166, in_2[13], in_1[13]);
  nand g101 (n_167, in_0[13], in_2[13]);
  nand g102 (out_0[14], n_165, n_166, n_167);
  xor g103 (n_168, in_0[14], in_1[14]);
  xor g104 (out_1[14], n_168, in_2[14]);
  nand g105 (n_169, in_0[14], in_1[14]);
  nand g106 (n_170, in_2[14], in_1[14]);
  nand g107 (n_171, in_0[14], in_2[14]);
  nand g108 (out_0[15], n_169, n_170, n_171);
  xor g109 (n_172, in_0[15], in_1[15]);
  xor g110 (out_1[15], n_172, in_2[15]);
  nand g111 (n_173, in_0[15], in_1[15]);
  nand g112 (n_174, in_2[15], in_1[15]);
  nand g113 (n_175, in_0[15], in_2[15]);
  nand g114 (out_0[16], n_173, n_174, n_175);
  xor g115 (n_176, in_0[16], in_1[16]);
  xor g116 (out_1[16], n_176, in_2[16]);
  nand g117 (n_177, in_0[16], in_1[16]);
  nand g118 (n_178, in_2[16], in_1[16]);
  nand g119 (n_179, in_0[16], in_2[16]);
  nand g120 (out_0[17], n_177, n_178, n_179);
  xor g121 (n_180, in_0[17], in_1[17]);
  xor g122 (out_1[17], n_180, in_2[17]);
  nand g123 (n_181, in_0[17], in_1[17]);
  nand g124 (n_182, in_2[17], in_1[17]);
  nand g125 (n_183, in_0[17], in_2[17]);
  nand g126 (out_0[18], n_181, n_182, n_183);
  xor g127 (n_184, in_0[18], in_1[18]);
  xor g128 (out_1[18], n_184, in_2[18]);
  nand g129 (n_185, in_0[18], in_1[18]);
  nand g130 (n_186, in_2[18], in_1[18]);
  nand g131 (n_187, in_0[18], in_2[18]);
  nand g132 (out_0[19], n_185, n_186, n_187);
  xor g133 (n_188, in_0[19], in_1[19]);
  xor g134 (out_1[19], n_188, in_2[19]);
  nand g135 (n_189, in_0[19], in_1[19]);
  nand g136 (n_190, in_2[19], in_1[19]);
  nand g137 (n_191, in_0[19], in_2[19]);
  nand g138 (out_0[20], n_189, n_190, n_191);
  xor g142 (out_1[20], in_2[20], n_67);
  xor g147 (n_67, in_0[20], in_1[20]);
  nor g148 (out_0[21], in_0[20], in_1[20]);
  or g149 (n_194, in_2[20], wc);
  not gc (wc, n_67);
  or g151 (out_1[21], wc0, wc1, n_67);
  not gc1 (wc1, n_194);
  not gc0 (wc0, in_2[20]);
endmodule

module csa_tree_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [20:0] in_0, in_1, in_2;
  output [23:0] out_0, out_1;
  wire [20:0] in_0, in_1, in_2;
  wire [23:0] out_0, out_1;
  csa_tree_GENERIC_REAL g1(.in_0 ({in_0[19], in_0[19:0]}), .in_1
       ({in_1[19], in_1[19:0]}), .in_2 (in_2), .out_0 (out_0), .out_1
       (out_1));
endmodule

module csa_tree_3123_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 25'b0;"
  input [23:0] in_0, in_1;
  input [21:0] in_2;
  output [24:0] out_0, out_1;
  wire [23:0] in_0, in_1;
  wire [21:0] in_2;
  wire [24:0] out_0, out_1;
  wire n_70, n_74, n_75, n_79, n_80, n_131, n_132, n_133;
  wire n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_213, n_217, n_221;
  assign out_0[0] = in_1[0];
  xor g31 (out_1[0], in_0[0], in_2[0]);
  and g32 (out_0[1], in_0[0], in_2[0]);
  xor g33 (n_131, in_0[1], in_1[1]);
  xor g34 (out_1[1], n_131, in_2[1]);
  nand g35 (n_132, in_0[1], in_1[1]);
  nand g4 (n_133, in_2[1], in_1[1]);
  nand g5 (n_134, in_0[1], in_2[1]);
  nand g36 (out_0[2], n_132, n_133, n_134);
  xor g37 (n_135, in_0[2], in_1[2]);
  xor g38 (out_1[2], n_135, in_2[2]);
  nand g39 (n_136, in_0[2], in_1[2]);
  nand g40 (n_137, in_2[2], in_1[2]);
  nand g41 (n_138, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_136, n_137, n_138);
  xor g42 (n_139, in_0[3], in_1[3]);
  xor g43 (out_1[3], n_139, in_2[3]);
  nand g44 (n_140, in_0[3], in_1[3]);
  nand g45 (n_141, in_2[3], in_1[3]);
  nand g46 (n_142, in_0[3], in_2[3]);
  nand g47 (out_0[4], n_140, n_141, n_142);
  xor g48 (n_143, in_0[4], in_1[4]);
  xor g49 (out_1[4], n_143, in_2[4]);
  nand g50 (n_144, in_0[4], in_1[4]);
  nand g51 (n_145, in_2[4], in_1[4]);
  nand g52 (n_146, in_0[4], in_2[4]);
  nand g53 (out_0[5], n_144, n_145, n_146);
  xor g54 (n_147, in_0[5], in_1[5]);
  xor g55 (out_1[5], n_147, in_2[5]);
  nand g56 (n_148, in_0[5], in_1[5]);
  nand g57 (n_149, in_2[5], in_1[5]);
  nand g58 (n_150, in_0[5], in_2[5]);
  nand g59 (out_0[6], n_148, n_149, n_150);
  xor g60 (n_151, in_0[6], in_1[6]);
  xor g61 (out_1[6], n_151, in_2[6]);
  nand g62 (n_152, in_0[6], in_1[6]);
  nand g63 (n_153, in_2[6], in_1[6]);
  nand g64 (n_154, in_0[6], in_2[6]);
  nand g65 (out_0[7], n_152, n_153, n_154);
  xor g66 (n_155, in_0[7], in_1[7]);
  xor g67 (out_1[7], n_155, in_2[7]);
  nand g68 (n_156, in_0[7], in_1[7]);
  nand g69 (n_157, in_2[7], in_1[7]);
  nand g70 (n_158, in_0[7], in_2[7]);
  nand g71 (out_0[8], n_156, n_157, n_158);
  xor g72 (n_159, in_0[8], in_1[8]);
  xor g73 (out_1[8], n_159, in_2[8]);
  nand g74 (n_160, in_0[8], in_1[8]);
  nand g75 (n_161, in_2[8], in_1[8]);
  nand g76 (n_162, in_0[8], in_2[8]);
  nand g77 (out_0[9], n_160, n_161, n_162);
  xor g78 (n_163, in_0[9], in_1[9]);
  xor g79 (out_1[9], n_163, in_2[9]);
  nand g80 (n_164, in_0[9], in_1[9]);
  nand g81 (n_165, in_2[9], in_1[9]);
  nand g82 (n_166, in_0[9], in_2[9]);
  nand g83 (out_0[10], n_164, n_165, n_166);
  xor g84 (n_167, in_0[10], in_1[10]);
  xor g85 (out_1[10], n_167, in_2[10]);
  nand g86 (n_168, in_0[10], in_1[10]);
  nand g87 (n_169, in_2[10], in_1[10]);
  nand g88 (n_170, in_0[10], in_2[10]);
  nand g89 (out_0[11], n_168, n_169, n_170);
  xor g90 (n_171, in_0[11], in_1[11]);
  xor g91 (out_1[11], n_171, in_2[11]);
  nand g92 (n_172, in_0[11], in_1[11]);
  nand g93 (n_173, in_2[11], in_1[11]);
  nand g94 (n_174, in_0[11], in_2[11]);
  nand g95 (out_0[12], n_172, n_173, n_174);
  xor g96 (n_175, in_0[12], in_1[12]);
  xor g97 (out_1[12], n_175, in_2[12]);
  nand g98 (n_176, in_0[12], in_1[12]);
  nand g99 (n_177, in_2[12], in_1[12]);
  nand g100 (n_178, in_0[12], in_2[12]);
  nand g101 (out_0[13], n_176, n_177, n_178);
  xor g102 (n_179, in_0[13], in_1[13]);
  xor g103 (out_1[13], n_179, in_2[13]);
  nand g104 (n_180, in_0[13], in_1[13]);
  nand g105 (n_181, in_2[13], in_1[13]);
  nand g106 (n_182, in_0[13], in_2[13]);
  nand g107 (out_0[14], n_180, n_181, n_182);
  xor g108 (n_183, in_0[14], in_1[14]);
  xor g109 (out_1[14], n_183, in_2[14]);
  nand g110 (n_184, in_0[14], in_1[14]);
  nand g111 (n_185, in_2[14], in_1[14]);
  nand g112 (n_186, in_0[14], in_2[14]);
  nand g113 (out_0[15], n_184, n_185, n_186);
  xor g114 (n_187, in_0[15], in_1[15]);
  xor g115 (out_1[15], n_187, in_2[15]);
  nand g116 (n_188, in_0[15], in_1[15]);
  nand g117 (n_189, in_2[15], in_1[15]);
  nand g118 (n_190, in_0[15], in_2[15]);
  nand g119 (out_0[16], n_188, n_189, n_190);
  xor g120 (n_191, in_0[16], in_1[16]);
  xor g121 (out_1[16], n_191, in_2[16]);
  nand g122 (n_192, in_0[16], in_1[16]);
  nand g123 (n_193, in_2[16], in_1[16]);
  nand g124 (n_194, in_0[16], in_2[16]);
  nand g125 (out_0[17], n_192, n_193, n_194);
  xor g126 (n_195, in_0[17], in_1[17]);
  xor g127 (out_1[17], n_195, in_2[17]);
  nand g128 (n_196, in_0[17], in_1[17]);
  nand g129 (n_197, in_2[17], in_1[17]);
  nand g130 (n_198, in_0[17], in_2[17]);
  nand g131 (out_0[18], n_196, n_197, n_198);
  xor g132 (n_199, in_0[18], in_1[18]);
  xor g133 (out_1[18], n_199, in_2[18]);
  nand g134 (n_200, in_0[18], in_1[18]);
  nand g135 (n_201, in_2[18], in_1[18]);
  nand g136 (n_202, in_0[18], in_2[18]);
  nand g137 (out_0[19], n_200, n_201, n_202);
  xor g138 (n_203, in_0[19], in_1[19]);
  xor g139 (out_1[19], n_203, in_2[19]);
  nand g140 (n_204, in_0[19], in_1[19]);
  nand g141 (n_205, in_2[19], in_1[19]);
  nand g142 (n_206, in_0[19], in_2[19]);
  nand g143 (out_0[20], n_204, n_205, n_206);
  xor g144 (n_207, in_0[20], in_1[20]);
  xor g145 (out_1[20], n_207, in_2[20]);
  nand g146 (n_208, in_0[20], in_1[20]);
  nand g147 (n_209, in_2[20], in_1[20]);
  nand g148 (n_210, in_0[20], in_2[20]);
  nand g149 (out_0[21], n_208, n_209, n_210);
  xor g150 (n_70, in_0[21], in_1[21]);
  and g151 (n_75, in_0[21], in_1[21]);
  xor g153 (out_1[21], in_2[21], n_70);
  xor g158 (n_74, in_0[22], in_1[22]);
  and g159 (n_80, in_0[22], in_1[22]);
  nand g163 (n_217, n_75, n_74);
  nand g171 (n_221, n_80, n_79);
  or g174 (n_213, in_2[21], wc);
  not gc (wc, n_70);
  xor g178 (n_79, in_0[23], in_1[23]);
  nor g179 (out_0[24], in_0[23], in_1[23]);
  or g181 (out_0[22], wc0, wc1, n_70);
  not gc1 (wc1, n_213);
  not gc0 (wc0, in_2[21]);
  xnor g182 (out_1[22], n_75, n_74);
  or g183 (out_0[23], wc2, n_74, n_75);
  not gc2 (wc2, n_217);
  xnor g185 (out_1[23], n_80, n_79);
  or g186 (out_1[24], n_79, wc3, n_80);
  not gc3 (wc3, n_221);
endmodule

module csa_tree_3123_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [23:0] in_0, in_1;
  input [21:0] in_2;
  output [24:0] out_0, out_1;
  wire [23:0] in_0, in_1;
  wire [21:0] in_2;
  wire [24:0] out_0, out_1;
  csa_tree_3123_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_3151_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 26'b0;"
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  wire n_73, n_77, n_78, n_82, n_83, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_222, n_226, n_230;
  assign out_0[0] = in_1[0];
  xor g32 (out_1[0], in_0[0], in_2[0]);
  and g33 (out_0[1], in_0[0], in_2[0]);
  xor g34 (n_136, in_0[1], in_1[1]);
  xor g35 (out_1[1], n_136, in_2[1]);
  nand g36 (n_137, in_0[1], in_1[1]);
  nand g4 (n_138, in_2[1], in_1[1]);
  nand g5 (n_139, in_0[1], in_2[1]);
  nand g37 (out_0[2], n_137, n_138, n_139);
  xor g38 (n_140, in_0[2], in_1[2]);
  xor g39 (out_1[2], n_140, in_2[2]);
  nand g40 (n_141, in_0[2], in_1[2]);
  nand g41 (n_142, in_2[2], in_1[2]);
  nand g42 (n_143, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_141, n_142, n_143);
  xor g43 (n_144, in_0[3], in_1[3]);
  xor g44 (out_1[3], n_144, in_2[3]);
  nand g45 (n_145, in_0[3], in_1[3]);
  nand g46 (n_146, in_2[3], in_1[3]);
  nand g47 (n_147, in_0[3], in_2[3]);
  nand g48 (out_0[4], n_145, n_146, n_147);
  xor g49 (n_148, in_0[4], in_1[4]);
  xor g50 (out_1[4], n_148, in_2[4]);
  nand g51 (n_149, in_0[4], in_1[4]);
  nand g52 (n_150, in_2[4], in_1[4]);
  nand g53 (n_151, in_0[4], in_2[4]);
  nand g54 (out_0[5], n_149, n_150, n_151);
  xor g55 (n_152, in_0[5], in_1[5]);
  xor g56 (out_1[5], n_152, in_2[5]);
  nand g57 (n_153, in_0[5], in_1[5]);
  nand g58 (n_154, in_2[5], in_1[5]);
  nand g59 (n_155, in_0[5], in_2[5]);
  nand g60 (out_0[6], n_153, n_154, n_155);
  xor g61 (n_156, in_0[6], in_1[6]);
  xor g62 (out_1[6], n_156, in_2[6]);
  nand g63 (n_157, in_0[6], in_1[6]);
  nand g64 (n_158, in_2[6], in_1[6]);
  nand g65 (n_159, in_0[6], in_2[6]);
  nand g66 (out_0[7], n_157, n_158, n_159);
  xor g67 (n_160, in_0[7], in_1[7]);
  xor g68 (out_1[7], n_160, in_2[7]);
  nand g69 (n_161, in_0[7], in_1[7]);
  nand g70 (n_162, in_2[7], in_1[7]);
  nand g71 (n_163, in_0[7], in_2[7]);
  nand g72 (out_0[8], n_161, n_162, n_163);
  xor g73 (n_164, in_0[8], in_1[8]);
  xor g74 (out_1[8], n_164, in_2[8]);
  nand g75 (n_165, in_0[8], in_1[8]);
  nand g76 (n_166, in_2[8], in_1[8]);
  nand g77 (n_167, in_0[8], in_2[8]);
  nand g78 (out_0[9], n_165, n_166, n_167);
  xor g79 (n_168, in_0[9], in_1[9]);
  xor g80 (out_1[9], n_168, in_2[9]);
  nand g81 (n_169, in_0[9], in_1[9]);
  nand g82 (n_170, in_2[9], in_1[9]);
  nand g83 (n_171, in_0[9], in_2[9]);
  nand g84 (out_0[10], n_169, n_170, n_171);
  xor g85 (n_172, in_0[10], in_1[10]);
  xor g86 (out_1[10], n_172, in_2[10]);
  nand g87 (n_173, in_0[10], in_1[10]);
  nand g88 (n_174, in_2[10], in_1[10]);
  nand g89 (n_175, in_0[10], in_2[10]);
  nand g90 (out_0[11], n_173, n_174, n_175);
  xor g91 (n_176, in_0[11], in_1[11]);
  xor g92 (out_1[11], n_176, in_2[11]);
  nand g93 (n_177, in_0[11], in_1[11]);
  nand g94 (n_178, in_2[11], in_1[11]);
  nand g95 (n_179, in_0[11], in_2[11]);
  nand g96 (out_0[12], n_177, n_178, n_179);
  xor g97 (n_180, in_0[12], in_1[12]);
  xor g98 (out_1[12], n_180, in_2[12]);
  nand g99 (n_181, in_0[12], in_1[12]);
  nand g100 (n_182, in_2[12], in_1[12]);
  nand g101 (n_183, in_0[12], in_2[12]);
  nand g102 (out_0[13], n_181, n_182, n_183);
  xor g103 (n_184, in_0[13], in_1[13]);
  xor g104 (out_1[13], n_184, in_2[13]);
  nand g105 (n_185, in_0[13], in_1[13]);
  nand g106 (n_186, in_2[13], in_1[13]);
  nand g107 (n_187, in_0[13], in_2[13]);
  nand g108 (out_0[14], n_185, n_186, n_187);
  xor g109 (n_188, in_0[14], in_1[14]);
  xor g110 (out_1[14], n_188, in_2[14]);
  nand g111 (n_189, in_0[14], in_1[14]);
  nand g112 (n_190, in_2[14], in_1[14]);
  nand g113 (n_191, in_0[14], in_2[14]);
  nand g114 (out_0[15], n_189, n_190, n_191);
  xor g115 (n_192, in_0[15], in_1[15]);
  xor g116 (out_1[15], n_192, in_2[15]);
  nand g117 (n_193, in_0[15], in_1[15]);
  nand g118 (n_194, in_2[15], in_1[15]);
  nand g119 (n_195, in_0[15], in_2[15]);
  nand g120 (out_0[16], n_193, n_194, n_195);
  xor g121 (n_196, in_0[16], in_1[16]);
  xor g122 (out_1[16], n_196, in_2[16]);
  nand g123 (n_197, in_0[16], in_1[16]);
  nand g124 (n_198, in_2[16], in_1[16]);
  nand g125 (n_199, in_0[16], in_2[16]);
  nand g126 (out_0[17], n_197, n_198, n_199);
  xor g127 (n_200, in_0[17], in_1[17]);
  xor g128 (out_1[17], n_200, in_2[17]);
  nand g129 (n_201, in_0[17], in_1[17]);
  nand g130 (n_202, in_2[17], in_1[17]);
  nand g131 (n_203, in_0[17], in_2[17]);
  nand g132 (out_0[18], n_201, n_202, n_203);
  xor g133 (n_204, in_0[18], in_1[18]);
  xor g134 (out_1[18], n_204, in_2[18]);
  nand g135 (n_205, in_0[18], in_1[18]);
  nand g136 (n_206, in_2[18], in_1[18]);
  nand g137 (n_207, in_0[18], in_2[18]);
  nand g138 (out_0[19], n_205, n_206, n_207);
  xor g139 (n_208, in_0[19], in_1[19]);
  xor g140 (out_1[19], n_208, in_2[19]);
  nand g141 (n_209, in_0[19], in_1[19]);
  nand g142 (n_210, in_2[19], in_1[19]);
  nand g143 (n_211, in_0[19], in_2[19]);
  nand g144 (out_0[20], n_209, n_210, n_211);
  xor g145 (n_212, in_0[20], in_1[20]);
  xor g146 (out_1[20], n_212, in_2[20]);
  nand g147 (n_213, in_0[20], in_1[20]);
  nand g148 (n_214, in_2[20], in_1[20]);
  nand g149 (n_215, in_0[20], in_2[20]);
  nand g150 (out_0[21], n_213, n_214, n_215);
  xor g151 (n_216, in_0[21], in_1[21]);
  xor g152 (out_1[21], n_216, in_2[21]);
  nand g153 (n_217, in_0[21], in_1[21]);
  nand g154 (n_218, in_2[21], in_1[21]);
  nand g155 (n_219, in_0[21], in_2[21]);
  nand g156 (out_0[22], n_217, n_218, n_219);
  xor g157 (n_73, in_0[22], in_1[22]);
  and g158 (n_78, in_0[22], in_1[22]);
  xor g160 (out_1[22], in_2[22], n_73);
  xor g165 (n_77, in_0[23], in_1[23]);
  and g166 (n_83, in_0[23], in_1[23]);
  nand g170 (n_226, n_78, n_77);
  nand g178 (n_230, n_83, n_82);
  or g181 (n_222, in_2[22], wc);
  not gc (wc, n_73);
  xor g185 (n_82, in_0[24], in_1[24]);
  nor g186 (out_0[25], in_0[24], in_1[24]);
  or g188 (out_0[23], wc0, wc1, n_73);
  not gc1 (wc1, n_222);
  not gc0 (wc0, in_2[22]);
  xnor g189 (out_1[23], n_78, n_77);
  or g190 (out_0[24], wc2, n_77, n_78);
  not gc2 (wc2, n_226);
  xnor g192 (out_1[24], n_83, n_82);
  or g193 (out_1[25], n_82, wc3, n_83);
  not gc3 (wc3, n_230);
endmodule

module csa_tree_3151_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  csa_tree_3151_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_3151_1_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 26'b0;"
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  wire n_73, n_77, n_78, n_82, n_83, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_222, n_226, n_230;
  assign out_0[0] = in_1[0];
  xor g32 (out_1[0], in_0[0], in_2[0]);
  and g33 (out_0[1], in_0[0], in_2[0]);
  xor g34 (n_136, in_0[1], in_1[1]);
  xor g35 (out_1[1], n_136, in_2[1]);
  nand g36 (n_137, in_0[1], in_1[1]);
  nand g4 (n_138, in_2[1], in_1[1]);
  nand g5 (n_139, in_0[1], in_2[1]);
  nand g37 (out_0[2], n_137, n_138, n_139);
  xor g38 (n_140, in_0[2], in_1[2]);
  xor g39 (out_1[2], n_140, in_2[2]);
  nand g40 (n_141, in_0[2], in_1[2]);
  nand g41 (n_142, in_2[2], in_1[2]);
  nand g42 (n_143, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_141, n_142, n_143);
  xor g43 (n_144, in_0[3], in_1[3]);
  xor g44 (out_1[3], n_144, in_2[3]);
  nand g45 (n_145, in_0[3], in_1[3]);
  nand g46 (n_146, in_2[3], in_1[3]);
  nand g47 (n_147, in_0[3], in_2[3]);
  nand g48 (out_0[4], n_145, n_146, n_147);
  xor g49 (n_148, in_0[4], in_1[4]);
  xor g50 (out_1[4], n_148, in_2[4]);
  nand g51 (n_149, in_0[4], in_1[4]);
  nand g52 (n_150, in_2[4], in_1[4]);
  nand g53 (n_151, in_0[4], in_2[4]);
  nand g54 (out_0[5], n_149, n_150, n_151);
  xor g55 (n_152, in_0[5], in_1[5]);
  xor g56 (out_1[5], n_152, in_2[5]);
  nand g57 (n_153, in_0[5], in_1[5]);
  nand g58 (n_154, in_2[5], in_1[5]);
  nand g59 (n_155, in_0[5], in_2[5]);
  nand g60 (out_0[6], n_153, n_154, n_155);
  xor g61 (n_156, in_0[6], in_1[6]);
  xor g62 (out_1[6], n_156, in_2[6]);
  nand g63 (n_157, in_0[6], in_1[6]);
  nand g64 (n_158, in_2[6], in_1[6]);
  nand g65 (n_159, in_0[6], in_2[6]);
  nand g66 (out_0[7], n_157, n_158, n_159);
  xor g67 (n_160, in_0[7], in_1[7]);
  xor g68 (out_1[7], n_160, in_2[7]);
  nand g69 (n_161, in_0[7], in_1[7]);
  nand g70 (n_162, in_2[7], in_1[7]);
  nand g71 (n_163, in_0[7], in_2[7]);
  nand g72 (out_0[8], n_161, n_162, n_163);
  xor g73 (n_164, in_0[8], in_1[8]);
  xor g74 (out_1[8], n_164, in_2[8]);
  nand g75 (n_165, in_0[8], in_1[8]);
  nand g76 (n_166, in_2[8], in_1[8]);
  nand g77 (n_167, in_0[8], in_2[8]);
  nand g78 (out_0[9], n_165, n_166, n_167);
  xor g79 (n_168, in_0[9], in_1[9]);
  xor g80 (out_1[9], n_168, in_2[9]);
  nand g81 (n_169, in_0[9], in_1[9]);
  nand g82 (n_170, in_2[9], in_1[9]);
  nand g83 (n_171, in_0[9], in_2[9]);
  nand g84 (out_0[10], n_169, n_170, n_171);
  xor g85 (n_172, in_0[10], in_1[10]);
  xor g86 (out_1[10], n_172, in_2[10]);
  nand g87 (n_173, in_0[10], in_1[10]);
  nand g88 (n_174, in_2[10], in_1[10]);
  nand g89 (n_175, in_0[10], in_2[10]);
  nand g90 (out_0[11], n_173, n_174, n_175);
  xor g91 (n_176, in_0[11], in_1[11]);
  xor g92 (out_1[11], n_176, in_2[11]);
  nand g93 (n_177, in_0[11], in_1[11]);
  nand g94 (n_178, in_2[11], in_1[11]);
  nand g95 (n_179, in_0[11], in_2[11]);
  nand g96 (out_0[12], n_177, n_178, n_179);
  xor g97 (n_180, in_0[12], in_1[12]);
  xor g98 (out_1[12], n_180, in_2[12]);
  nand g99 (n_181, in_0[12], in_1[12]);
  nand g100 (n_182, in_2[12], in_1[12]);
  nand g101 (n_183, in_0[12], in_2[12]);
  nand g102 (out_0[13], n_181, n_182, n_183);
  xor g103 (n_184, in_0[13], in_1[13]);
  xor g104 (out_1[13], n_184, in_2[13]);
  nand g105 (n_185, in_0[13], in_1[13]);
  nand g106 (n_186, in_2[13], in_1[13]);
  nand g107 (n_187, in_0[13], in_2[13]);
  nand g108 (out_0[14], n_185, n_186, n_187);
  xor g109 (n_188, in_0[14], in_1[14]);
  xor g110 (out_1[14], n_188, in_2[14]);
  nand g111 (n_189, in_0[14], in_1[14]);
  nand g112 (n_190, in_2[14], in_1[14]);
  nand g113 (n_191, in_0[14], in_2[14]);
  nand g114 (out_0[15], n_189, n_190, n_191);
  xor g115 (n_192, in_0[15], in_1[15]);
  xor g116 (out_1[15], n_192, in_2[15]);
  nand g117 (n_193, in_0[15], in_1[15]);
  nand g118 (n_194, in_2[15], in_1[15]);
  nand g119 (n_195, in_0[15], in_2[15]);
  nand g120 (out_0[16], n_193, n_194, n_195);
  xor g121 (n_196, in_0[16], in_1[16]);
  xor g122 (out_1[16], n_196, in_2[16]);
  nand g123 (n_197, in_0[16], in_1[16]);
  nand g124 (n_198, in_2[16], in_1[16]);
  nand g125 (n_199, in_0[16], in_2[16]);
  nand g126 (out_0[17], n_197, n_198, n_199);
  xor g127 (n_200, in_0[17], in_1[17]);
  xor g128 (out_1[17], n_200, in_2[17]);
  nand g129 (n_201, in_0[17], in_1[17]);
  nand g130 (n_202, in_2[17], in_1[17]);
  nand g131 (n_203, in_0[17], in_2[17]);
  nand g132 (out_0[18], n_201, n_202, n_203);
  xor g133 (n_204, in_0[18], in_1[18]);
  xor g134 (out_1[18], n_204, in_2[18]);
  nand g135 (n_205, in_0[18], in_1[18]);
  nand g136 (n_206, in_2[18], in_1[18]);
  nand g137 (n_207, in_0[18], in_2[18]);
  nand g138 (out_0[19], n_205, n_206, n_207);
  xor g139 (n_208, in_0[19], in_1[19]);
  xor g140 (out_1[19], n_208, in_2[19]);
  nand g141 (n_209, in_0[19], in_1[19]);
  nand g142 (n_210, in_2[19], in_1[19]);
  nand g143 (n_211, in_0[19], in_2[19]);
  nand g144 (out_0[20], n_209, n_210, n_211);
  xor g145 (n_212, in_0[20], in_1[20]);
  xor g146 (out_1[20], n_212, in_2[20]);
  nand g147 (n_213, in_0[20], in_1[20]);
  nand g148 (n_214, in_2[20], in_1[20]);
  nand g149 (n_215, in_0[20], in_2[20]);
  nand g150 (out_0[21], n_213, n_214, n_215);
  xor g151 (n_216, in_0[21], in_1[21]);
  xor g152 (out_1[21], n_216, in_2[21]);
  nand g153 (n_217, in_0[21], in_1[21]);
  nand g154 (n_218, in_2[21], in_1[21]);
  nand g155 (n_219, in_0[21], in_2[21]);
  nand g156 (out_0[22], n_217, n_218, n_219);
  xor g157 (n_73, in_0[22], in_1[22]);
  and g158 (n_78, in_0[22], in_1[22]);
  xor g160 (out_1[22], in_2[22], n_73);
  xor g165 (n_77, in_0[23], in_1[23]);
  and g166 (n_83, in_0[23], in_1[23]);
  nand g170 (n_226, n_78, n_77);
  nand g178 (n_230, n_83, n_82);
  or g181 (n_222, in_2[22], wc);
  not gc (wc, n_73);
  xor g185 (n_82, in_0[24], in_1[24]);
  nor g186 (out_0[25], in_0[24], in_1[24]);
  or g188 (out_0[23], wc0, wc1, n_73);
  not gc1 (wc1, n_222);
  not gc0 (wc0, in_2[22]);
  xnor g189 (out_1[23], n_78, n_77);
  or g190 (out_0[24], wc2, n_77, n_78);
  not gc2 (wc2, n_226);
  xnor g192 (out_1[24], n_83, n_82);
  or g193 (out_1[25], n_82, wc3, n_83);
  not gc3 (wc3, n_230);
endmodule

module csa_tree_3151_1_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  csa_tree_3151_1_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_3151_2_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 26'b0;"
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  wire n_73, n_77, n_78, n_82, n_83, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_222, n_226, n_230;
  assign out_0[0] = in_1[0];
  xor g32 (out_1[0], in_0[0], in_2[0]);
  and g33 (out_0[1], in_0[0], in_2[0]);
  xor g34 (n_136, in_0[1], in_1[1]);
  xor g35 (out_1[1], n_136, in_2[1]);
  nand g36 (n_137, in_0[1], in_1[1]);
  nand g4 (n_138, in_2[1], in_1[1]);
  nand g5 (n_139, in_0[1], in_2[1]);
  nand g37 (out_0[2], n_137, n_138, n_139);
  xor g38 (n_140, in_0[2], in_1[2]);
  xor g39 (out_1[2], n_140, in_2[2]);
  nand g40 (n_141, in_0[2], in_1[2]);
  nand g41 (n_142, in_2[2], in_1[2]);
  nand g42 (n_143, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_141, n_142, n_143);
  xor g43 (n_144, in_0[3], in_1[3]);
  xor g44 (out_1[3], n_144, in_2[3]);
  nand g45 (n_145, in_0[3], in_1[3]);
  nand g46 (n_146, in_2[3], in_1[3]);
  nand g47 (n_147, in_0[3], in_2[3]);
  nand g48 (out_0[4], n_145, n_146, n_147);
  xor g49 (n_148, in_0[4], in_1[4]);
  xor g50 (out_1[4], n_148, in_2[4]);
  nand g51 (n_149, in_0[4], in_1[4]);
  nand g52 (n_150, in_2[4], in_1[4]);
  nand g53 (n_151, in_0[4], in_2[4]);
  nand g54 (out_0[5], n_149, n_150, n_151);
  xor g55 (n_152, in_0[5], in_1[5]);
  xor g56 (out_1[5], n_152, in_2[5]);
  nand g57 (n_153, in_0[5], in_1[5]);
  nand g58 (n_154, in_2[5], in_1[5]);
  nand g59 (n_155, in_0[5], in_2[5]);
  nand g60 (out_0[6], n_153, n_154, n_155);
  xor g61 (n_156, in_0[6], in_1[6]);
  xor g62 (out_1[6], n_156, in_2[6]);
  nand g63 (n_157, in_0[6], in_1[6]);
  nand g64 (n_158, in_2[6], in_1[6]);
  nand g65 (n_159, in_0[6], in_2[6]);
  nand g66 (out_0[7], n_157, n_158, n_159);
  xor g67 (n_160, in_0[7], in_1[7]);
  xor g68 (out_1[7], n_160, in_2[7]);
  nand g69 (n_161, in_0[7], in_1[7]);
  nand g70 (n_162, in_2[7], in_1[7]);
  nand g71 (n_163, in_0[7], in_2[7]);
  nand g72 (out_0[8], n_161, n_162, n_163);
  xor g73 (n_164, in_0[8], in_1[8]);
  xor g74 (out_1[8], n_164, in_2[8]);
  nand g75 (n_165, in_0[8], in_1[8]);
  nand g76 (n_166, in_2[8], in_1[8]);
  nand g77 (n_167, in_0[8], in_2[8]);
  nand g78 (out_0[9], n_165, n_166, n_167);
  xor g79 (n_168, in_0[9], in_1[9]);
  xor g80 (out_1[9], n_168, in_2[9]);
  nand g81 (n_169, in_0[9], in_1[9]);
  nand g82 (n_170, in_2[9], in_1[9]);
  nand g83 (n_171, in_0[9], in_2[9]);
  nand g84 (out_0[10], n_169, n_170, n_171);
  xor g85 (n_172, in_0[10], in_1[10]);
  xor g86 (out_1[10], n_172, in_2[10]);
  nand g87 (n_173, in_0[10], in_1[10]);
  nand g88 (n_174, in_2[10], in_1[10]);
  nand g89 (n_175, in_0[10], in_2[10]);
  nand g90 (out_0[11], n_173, n_174, n_175);
  xor g91 (n_176, in_0[11], in_1[11]);
  xor g92 (out_1[11], n_176, in_2[11]);
  nand g93 (n_177, in_0[11], in_1[11]);
  nand g94 (n_178, in_2[11], in_1[11]);
  nand g95 (n_179, in_0[11], in_2[11]);
  nand g96 (out_0[12], n_177, n_178, n_179);
  xor g97 (n_180, in_0[12], in_1[12]);
  xor g98 (out_1[12], n_180, in_2[12]);
  nand g99 (n_181, in_0[12], in_1[12]);
  nand g100 (n_182, in_2[12], in_1[12]);
  nand g101 (n_183, in_0[12], in_2[12]);
  nand g102 (out_0[13], n_181, n_182, n_183);
  xor g103 (n_184, in_0[13], in_1[13]);
  xor g104 (out_1[13], n_184, in_2[13]);
  nand g105 (n_185, in_0[13], in_1[13]);
  nand g106 (n_186, in_2[13], in_1[13]);
  nand g107 (n_187, in_0[13], in_2[13]);
  nand g108 (out_0[14], n_185, n_186, n_187);
  xor g109 (n_188, in_0[14], in_1[14]);
  xor g110 (out_1[14], n_188, in_2[14]);
  nand g111 (n_189, in_0[14], in_1[14]);
  nand g112 (n_190, in_2[14], in_1[14]);
  nand g113 (n_191, in_0[14], in_2[14]);
  nand g114 (out_0[15], n_189, n_190, n_191);
  xor g115 (n_192, in_0[15], in_1[15]);
  xor g116 (out_1[15], n_192, in_2[15]);
  nand g117 (n_193, in_0[15], in_1[15]);
  nand g118 (n_194, in_2[15], in_1[15]);
  nand g119 (n_195, in_0[15], in_2[15]);
  nand g120 (out_0[16], n_193, n_194, n_195);
  xor g121 (n_196, in_0[16], in_1[16]);
  xor g122 (out_1[16], n_196, in_2[16]);
  nand g123 (n_197, in_0[16], in_1[16]);
  nand g124 (n_198, in_2[16], in_1[16]);
  nand g125 (n_199, in_0[16], in_2[16]);
  nand g126 (out_0[17], n_197, n_198, n_199);
  xor g127 (n_200, in_0[17], in_1[17]);
  xor g128 (out_1[17], n_200, in_2[17]);
  nand g129 (n_201, in_0[17], in_1[17]);
  nand g130 (n_202, in_2[17], in_1[17]);
  nand g131 (n_203, in_0[17], in_2[17]);
  nand g132 (out_0[18], n_201, n_202, n_203);
  xor g133 (n_204, in_0[18], in_1[18]);
  xor g134 (out_1[18], n_204, in_2[18]);
  nand g135 (n_205, in_0[18], in_1[18]);
  nand g136 (n_206, in_2[18], in_1[18]);
  nand g137 (n_207, in_0[18], in_2[18]);
  nand g138 (out_0[19], n_205, n_206, n_207);
  xor g139 (n_208, in_0[19], in_1[19]);
  xor g140 (out_1[19], n_208, in_2[19]);
  nand g141 (n_209, in_0[19], in_1[19]);
  nand g142 (n_210, in_2[19], in_1[19]);
  nand g143 (n_211, in_0[19], in_2[19]);
  nand g144 (out_0[20], n_209, n_210, n_211);
  xor g145 (n_212, in_0[20], in_1[20]);
  xor g146 (out_1[20], n_212, in_2[20]);
  nand g147 (n_213, in_0[20], in_1[20]);
  nand g148 (n_214, in_2[20], in_1[20]);
  nand g149 (n_215, in_0[20], in_2[20]);
  nand g150 (out_0[21], n_213, n_214, n_215);
  xor g151 (n_216, in_0[21], in_1[21]);
  xor g152 (out_1[21], n_216, in_2[21]);
  nand g153 (n_217, in_0[21], in_1[21]);
  nand g154 (n_218, in_2[21], in_1[21]);
  nand g155 (n_219, in_0[21], in_2[21]);
  nand g156 (out_0[22], n_217, n_218, n_219);
  xor g157 (n_73, in_0[22], in_1[22]);
  and g158 (n_78, in_0[22], in_1[22]);
  xor g160 (out_1[22], in_2[22], n_73);
  xor g165 (n_77, in_0[23], in_1[23]);
  and g166 (n_83, in_0[23], in_1[23]);
  nand g170 (n_226, n_78, n_77);
  nand g178 (n_230, n_83, n_82);
  or g181 (n_222, in_2[22], wc);
  not gc (wc, n_73);
  xor g185 (n_82, in_0[24], in_1[24]);
  nor g186 (out_0[25], in_0[24], in_1[24]);
  or g188 (out_0[23], wc0, wc1, n_73);
  not gc1 (wc1, n_222);
  not gc0 (wc0, in_2[22]);
  xnor g189 (out_1[23], n_78, n_77);
  or g190 (out_0[24], wc2, n_77, n_78);
  not gc2 (wc2, n_226);
  xnor g192 (out_1[24], n_83, n_82);
  or g193 (out_1[25], n_82, wc3, n_83);
  not gc3 (wc3, n_230);
endmodule

module csa_tree_3151_2_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  csa_tree_3151_2_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_3209_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 25'b0;"
  input [21:0] in_0, in_1, in_2;
  output [24:0] out_0, out_1;
  wire [21:0] in_0, in_1, in_2;
  wire [24:0] out_0, out_1;
  wire n_70, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_203;
  assign out_1[23] = 1'b0;
  assign out_1[24] = 1'b0;
  assign out_0[0] = in_1[0];
  assign out_0[23] = 1'b1;
  assign out_0[24] = 1'b1;
  xor g27 (out_1[0], in_0[0], in_2[0]);
  and g28 (out_0[1], in_0[0], in_2[0]);
  xor g29 (n_121, in_0[1], in_1[1]);
  xor g30 (out_1[1], n_121, in_2[1]);
  nand g31 (n_122, in_0[1], in_1[1]);
  nand g4 (n_123, in_2[1], in_1[1]);
  nand g5 (n_124, in_0[1], in_2[1]);
  nand g32 (out_0[2], n_122, n_123, n_124);
  xor g33 (n_125, in_0[2], in_1[2]);
  xor g34 (out_1[2], n_125, in_2[2]);
  nand g35 (n_126, in_0[2], in_1[2]);
  nand g36 (n_127, in_2[2], in_1[2]);
  nand g37 (n_128, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_126, n_127, n_128);
  xor g38 (n_129, in_0[3], in_1[3]);
  xor g39 (out_1[3], n_129, in_2[3]);
  nand g40 (n_130, in_0[3], in_1[3]);
  nand g41 (n_131, in_2[3], in_1[3]);
  nand g42 (n_132, in_0[3], in_2[3]);
  nand g43 (out_0[4], n_130, n_131, n_132);
  xor g44 (n_133, in_0[4], in_1[4]);
  xor g45 (out_1[4], n_133, in_2[4]);
  nand g46 (n_134, in_0[4], in_1[4]);
  nand g47 (n_135, in_2[4], in_1[4]);
  nand g48 (n_136, in_0[4], in_2[4]);
  nand g49 (out_0[5], n_134, n_135, n_136);
  xor g50 (n_137, in_0[5], in_1[5]);
  xor g51 (out_1[5], n_137, in_2[5]);
  nand g52 (n_138, in_0[5], in_1[5]);
  nand g53 (n_139, in_2[5], in_1[5]);
  nand g54 (n_140, in_0[5], in_2[5]);
  nand g55 (out_0[6], n_138, n_139, n_140);
  xor g56 (n_141, in_0[6], in_1[6]);
  xor g57 (out_1[6], n_141, in_2[6]);
  nand g58 (n_142, in_0[6], in_1[6]);
  nand g59 (n_143, in_2[6], in_1[6]);
  nand g60 (n_144, in_0[6], in_2[6]);
  nand g61 (out_0[7], n_142, n_143, n_144);
  xor g62 (n_145, in_0[7], in_1[7]);
  xor g63 (out_1[7], n_145, in_2[7]);
  nand g64 (n_146, in_0[7], in_1[7]);
  nand g65 (n_147, in_2[7], in_1[7]);
  nand g66 (n_148, in_0[7], in_2[7]);
  nand g67 (out_0[8], n_146, n_147, n_148);
  xor g68 (n_149, in_0[8], in_1[8]);
  xor g69 (out_1[8], n_149, in_2[8]);
  nand g70 (n_150, in_0[8], in_1[8]);
  nand g71 (n_151, in_2[8], in_1[8]);
  nand g72 (n_152, in_0[8], in_2[8]);
  nand g73 (out_0[9], n_150, n_151, n_152);
  xor g74 (n_153, in_0[9], in_1[9]);
  xor g75 (out_1[9], n_153, in_2[9]);
  nand g76 (n_154, in_0[9], in_1[9]);
  nand g77 (n_155, in_2[9], in_1[9]);
  nand g78 (n_156, in_0[9], in_2[9]);
  nand g79 (out_0[10], n_154, n_155, n_156);
  xor g80 (n_157, in_0[10], in_1[10]);
  xor g81 (out_1[10], n_157, in_2[10]);
  nand g82 (n_158, in_0[10], in_1[10]);
  nand g83 (n_159, in_2[10], in_1[10]);
  nand g84 (n_160, in_0[10], in_2[10]);
  nand g85 (out_0[11], n_158, n_159, n_160);
  xor g86 (n_161, in_0[11], in_1[11]);
  xor g87 (out_1[11], n_161, in_2[11]);
  nand g88 (n_162, in_0[11], in_1[11]);
  nand g89 (n_163, in_2[11], in_1[11]);
  nand g90 (n_164, in_0[11], in_2[11]);
  nand g91 (out_0[12], n_162, n_163, n_164);
  xor g92 (n_165, in_0[12], in_1[12]);
  xor g93 (out_1[12], n_165, in_2[12]);
  nand g94 (n_166, in_0[12], in_1[12]);
  nand g95 (n_167, in_2[12], in_1[12]);
  nand g96 (n_168, in_0[12], in_2[12]);
  nand g97 (out_0[13], n_166, n_167, n_168);
  xor g98 (n_169, in_0[13], in_1[13]);
  xor g99 (out_1[13], n_169, in_2[13]);
  nand g100 (n_170, in_0[13], in_1[13]);
  nand g101 (n_171, in_2[13], in_1[13]);
  nand g102 (n_172, in_0[13], in_2[13]);
  nand g103 (out_0[14], n_170, n_171, n_172);
  xor g104 (n_173, in_0[14], in_1[14]);
  xor g105 (out_1[14], n_173, in_2[14]);
  nand g106 (n_174, in_0[14], in_1[14]);
  nand g107 (n_175, in_2[14], in_1[14]);
  nand g108 (n_176, in_0[14], in_2[14]);
  nand g109 (out_0[15], n_174, n_175, n_176);
  xor g110 (n_177, in_0[15], in_1[15]);
  xor g111 (out_1[15], n_177, in_2[15]);
  nand g112 (n_178, in_0[15], in_1[15]);
  nand g113 (n_179, in_2[15], in_1[15]);
  nand g114 (n_180, in_0[15], in_2[15]);
  nand g115 (out_0[16], n_178, n_179, n_180);
  xor g116 (n_181, in_0[16], in_1[16]);
  xor g117 (out_1[16], n_181, in_2[16]);
  nand g118 (n_182, in_0[16], in_1[16]);
  nand g119 (n_183, in_2[16], in_1[16]);
  nand g120 (n_184, in_0[16], in_2[16]);
  nand g121 (out_0[17], n_182, n_183, n_184);
  xor g122 (n_185, in_0[17], in_1[17]);
  xor g123 (out_1[17], n_185, in_2[17]);
  nand g124 (n_186, in_0[17], in_1[17]);
  nand g125 (n_187, in_2[17], in_1[17]);
  nand g126 (n_188, in_0[17], in_2[17]);
  nand g127 (out_0[18], n_186, n_187, n_188);
  xor g128 (n_189, in_0[18], in_1[18]);
  xor g129 (out_1[18], n_189, in_2[18]);
  nand g130 (n_190, in_0[18], in_1[18]);
  nand g131 (n_191, in_2[18], in_1[18]);
  nand g132 (n_192, in_0[18], in_2[18]);
  nand g133 (out_0[19], n_190, n_191, n_192);
  xor g134 (n_193, in_0[19], in_1[19]);
  xor g135 (out_1[19], n_193, in_2[19]);
  nand g136 (n_194, in_0[19], in_1[19]);
  nand g137 (n_195, in_2[19], in_1[19]);
  nand g138 (n_196, in_0[19], in_2[19]);
  nand g139 (out_0[20], n_194, n_195, n_196);
  xor g140 (n_197, in_0[20], in_1[20]);
  xor g141 (out_1[20], n_197, in_2[20]);
  nand g142 (n_198, in_0[20], in_1[20]);
  nand g143 (n_199, in_2[20], in_1[20]);
  nand g144 (n_200, in_0[20], in_2[20]);
  nand g145 (out_0[21], n_198, n_199, n_200);
  xor g149 (out_1[21], in_2[21], n_70);
  xor g154 (n_70, in_0[21], in_1[21]);
  nor g155 (out_0[22], in_0[21], in_1[21]);
  or g156 (n_203, in_2[21], wc);
  not gc (wc, n_70);
  or g158 (out_1[22], wc0, wc1, n_70);
  not gc1 (wc1, n_203);
  not gc0 (wc0, in_2[21]);
endmodule

module csa_tree_3209_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [21:0] in_0, in_1, in_2;
  output [24:0] out_0, out_1;
  wire [21:0] in_0, in_1, in_2;
  wire [24:0] out_0, out_1;
  csa_tree_3209_GENERIC_REAL g1(.in_0 ({in_0[20], in_0[20:0]}), .in_1
       ({in_1[20], in_1[20:0]}), .in_2 (in_2), .out_0 (out_0), .out_1
       (out_1));
endmodule

module csa_tree_3209_1_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 25'b0;"
  input [21:0] in_0, in_1, in_2;
  output [24:0] out_0, out_1;
  wire [21:0] in_0, in_1, in_2;
  wire [24:0] out_0, out_1;
  wire n_70, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_203;
  assign out_1[23] = 1'b0;
  assign out_1[24] = 1'b0;
  assign out_0[0] = in_1[0];
  assign out_0[23] = 1'b1;
  assign out_0[24] = 1'b1;
  xor g27 (out_1[0], in_0[0], in_2[0]);
  and g28 (out_0[1], in_0[0], in_2[0]);
  xor g29 (n_121, in_0[1], in_1[1]);
  xor g30 (out_1[1], n_121, in_2[1]);
  nand g31 (n_122, in_0[1], in_1[1]);
  nand g4 (n_123, in_2[1], in_1[1]);
  nand g5 (n_124, in_0[1], in_2[1]);
  nand g32 (out_0[2], n_122, n_123, n_124);
  xor g33 (n_125, in_0[2], in_1[2]);
  xor g34 (out_1[2], n_125, in_2[2]);
  nand g35 (n_126, in_0[2], in_1[2]);
  nand g36 (n_127, in_2[2], in_1[2]);
  nand g37 (n_128, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_126, n_127, n_128);
  xor g38 (n_129, in_0[3], in_1[3]);
  xor g39 (out_1[3], n_129, in_2[3]);
  nand g40 (n_130, in_0[3], in_1[3]);
  nand g41 (n_131, in_2[3], in_1[3]);
  nand g42 (n_132, in_0[3], in_2[3]);
  nand g43 (out_0[4], n_130, n_131, n_132);
  xor g44 (n_133, in_0[4], in_1[4]);
  xor g45 (out_1[4], n_133, in_2[4]);
  nand g46 (n_134, in_0[4], in_1[4]);
  nand g47 (n_135, in_2[4], in_1[4]);
  nand g48 (n_136, in_0[4], in_2[4]);
  nand g49 (out_0[5], n_134, n_135, n_136);
  xor g50 (n_137, in_0[5], in_1[5]);
  xor g51 (out_1[5], n_137, in_2[5]);
  nand g52 (n_138, in_0[5], in_1[5]);
  nand g53 (n_139, in_2[5], in_1[5]);
  nand g54 (n_140, in_0[5], in_2[5]);
  nand g55 (out_0[6], n_138, n_139, n_140);
  xor g56 (n_141, in_0[6], in_1[6]);
  xor g57 (out_1[6], n_141, in_2[6]);
  nand g58 (n_142, in_0[6], in_1[6]);
  nand g59 (n_143, in_2[6], in_1[6]);
  nand g60 (n_144, in_0[6], in_2[6]);
  nand g61 (out_0[7], n_142, n_143, n_144);
  xor g62 (n_145, in_0[7], in_1[7]);
  xor g63 (out_1[7], n_145, in_2[7]);
  nand g64 (n_146, in_0[7], in_1[7]);
  nand g65 (n_147, in_2[7], in_1[7]);
  nand g66 (n_148, in_0[7], in_2[7]);
  nand g67 (out_0[8], n_146, n_147, n_148);
  xor g68 (n_149, in_0[8], in_1[8]);
  xor g69 (out_1[8], n_149, in_2[8]);
  nand g70 (n_150, in_0[8], in_1[8]);
  nand g71 (n_151, in_2[8], in_1[8]);
  nand g72 (n_152, in_0[8], in_2[8]);
  nand g73 (out_0[9], n_150, n_151, n_152);
  xor g74 (n_153, in_0[9], in_1[9]);
  xor g75 (out_1[9], n_153, in_2[9]);
  nand g76 (n_154, in_0[9], in_1[9]);
  nand g77 (n_155, in_2[9], in_1[9]);
  nand g78 (n_156, in_0[9], in_2[9]);
  nand g79 (out_0[10], n_154, n_155, n_156);
  xor g80 (n_157, in_0[10], in_1[10]);
  xor g81 (out_1[10], n_157, in_2[10]);
  nand g82 (n_158, in_0[10], in_1[10]);
  nand g83 (n_159, in_2[10], in_1[10]);
  nand g84 (n_160, in_0[10], in_2[10]);
  nand g85 (out_0[11], n_158, n_159, n_160);
  xor g86 (n_161, in_0[11], in_1[11]);
  xor g87 (out_1[11], n_161, in_2[11]);
  nand g88 (n_162, in_0[11], in_1[11]);
  nand g89 (n_163, in_2[11], in_1[11]);
  nand g90 (n_164, in_0[11], in_2[11]);
  nand g91 (out_0[12], n_162, n_163, n_164);
  xor g92 (n_165, in_0[12], in_1[12]);
  xor g93 (out_1[12], n_165, in_2[12]);
  nand g94 (n_166, in_0[12], in_1[12]);
  nand g95 (n_167, in_2[12], in_1[12]);
  nand g96 (n_168, in_0[12], in_2[12]);
  nand g97 (out_0[13], n_166, n_167, n_168);
  xor g98 (n_169, in_0[13], in_1[13]);
  xor g99 (out_1[13], n_169, in_2[13]);
  nand g100 (n_170, in_0[13], in_1[13]);
  nand g101 (n_171, in_2[13], in_1[13]);
  nand g102 (n_172, in_0[13], in_2[13]);
  nand g103 (out_0[14], n_170, n_171, n_172);
  xor g104 (n_173, in_0[14], in_1[14]);
  xor g105 (out_1[14], n_173, in_2[14]);
  nand g106 (n_174, in_0[14], in_1[14]);
  nand g107 (n_175, in_2[14], in_1[14]);
  nand g108 (n_176, in_0[14], in_2[14]);
  nand g109 (out_0[15], n_174, n_175, n_176);
  xor g110 (n_177, in_0[15], in_1[15]);
  xor g111 (out_1[15], n_177, in_2[15]);
  nand g112 (n_178, in_0[15], in_1[15]);
  nand g113 (n_179, in_2[15], in_1[15]);
  nand g114 (n_180, in_0[15], in_2[15]);
  nand g115 (out_0[16], n_178, n_179, n_180);
  xor g116 (n_181, in_0[16], in_1[16]);
  xor g117 (out_1[16], n_181, in_2[16]);
  nand g118 (n_182, in_0[16], in_1[16]);
  nand g119 (n_183, in_2[16], in_1[16]);
  nand g120 (n_184, in_0[16], in_2[16]);
  nand g121 (out_0[17], n_182, n_183, n_184);
  xor g122 (n_185, in_0[17], in_1[17]);
  xor g123 (out_1[17], n_185, in_2[17]);
  nand g124 (n_186, in_0[17], in_1[17]);
  nand g125 (n_187, in_2[17], in_1[17]);
  nand g126 (n_188, in_0[17], in_2[17]);
  nand g127 (out_0[18], n_186, n_187, n_188);
  xor g128 (n_189, in_0[18], in_1[18]);
  xor g129 (out_1[18], n_189, in_2[18]);
  nand g130 (n_190, in_0[18], in_1[18]);
  nand g131 (n_191, in_2[18], in_1[18]);
  nand g132 (n_192, in_0[18], in_2[18]);
  nand g133 (out_0[19], n_190, n_191, n_192);
  xor g134 (n_193, in_0[19], in_1[19]);
  xor g135 (out_1[19], n_193, in_2[19]);
  nand g136 (n_194, in_0[19], in_1[19]);
  nand g137 (n_195, in_2[19], in_1[19]);
  nand g138 (n_196, in_0[19], in_2[19]);
  nand g139 (out_0[20], n_194, n_195, n_196);
  xor g140 (n_197, in_0[20], in_1[20]);
  xor g141 (out_1[20], n_197, in_2[20]);
  nand g142 (n_198, in_0[20], in_1[20]);
  nand g143 (n_199, in_2[20], in_1[20]);
  nand g144 (n_200, in_0[20], in_2[20]);
  nand g145 (out_0[21], n_198, n_199, n_200);
  xor g149 (out_1[21], in_2[21], n_70);
  xor g154 (n_70, in_0[21], in_1[21]);
  nor g155 (out_0[22], in_0[21], in_1[21]);
  or g156 (n_203, in_2[21], wc);
  not gc (wc, n_70);
  or g158 (out_1[22], wc0, wc1, n_70);
  not gc1 (wc1, n_203);
  not gc0 (wc0, in_2[21]);
endmodule

module csa_tree_3209_1_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [21:0] in_0, in_1, in_2;
  output [24:0] out_0, out_1;
  wire [21:0] in_0, in_1, in_2;
  wire [24:0] out_0, out_1;
  csa_tree_3209_1_GENERIC_REAL g1(.in_0 ({in_0[20], in_0[20:0]}), .in_1
       ({in_1[20], in_1[20:0]}), .in_2 (in_2), .out_0 (out_0), .out_1
       (out_1));
endmodule

module csa_tree_6719_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 26'b0;"
  input [22:0] in_0, in_1, in_2;
  output [25:0] out_0, out_1;
  wire [22:0] in_0, in_1, in_2;
  wire [25:0] out_0, out_1;
  wire n_73, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_212;
  assign out_1[24] = 1'b0;
  assign out_1[25] = 1'b0;
  assign out_0[0] = in_1[0];
  assign out_0[24] = 1'b1;
  assign out_0[25] = 1'b1;
  xor g28 (out_1[0], in_0[0], in_2[0]);
  and g29 (out_0[1], in_0[0], in_2[0]);
  xor g30 (n_126, in_0[1], in_1[1]);
  xor g31 (out_1[1], n_126, in_2[1]);
  nand g32 (n_127, in_0[1], in_1[1]);
  nand g4 (n_128, in_2[1], in_1[1]);
  nand g5 (n_129, in_0[1], in_2[1]);
  nand g33 (out_0[2], n_127, n_128, n_129);
  xor g34 (n_130, in_0[2], in_1[2]);
  xor g35 (out_1[2], n_130, in_2[2]);
  nand g36 (n_131, in_0[2], in_1[2]);
  nand g37 (n_132, in_2[2], in_1[2]);
  nand g38 (n_133, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_131, n_132, n_133);
  xor g39 (n_134, in_0[3], in_1[3]);
  xor g40 (out_1[3], n_134, in_2[3]);
  nand g41 (n_135, in_0[3], in_1[3]);
  nand g42 (n_136, in_2[3], in_1[3]);
  nand g43 (n_137, in_0[3], in_2[3]);
  nand g44 (out_0[4], n_135, n_136, n_137);
  xor g45 (n_138, in_0[4], in_1[4]);
  xor g46 (out_1[4], n_138, in_2[4]);
  nand g47 (n_139, in_0[4], in_1[4]);
  nand g48 (n_140, in_2[4], in_1[4]);
  nand g49 (n_141, in_0[4], in_2[4]);
  nand g50 (out_0[5], n_139, n_140, n_141);
  xor g51 (n_142, in_0[5], in_1[5]);
  xor g52 (out_1[5], n_142, in_2[5]);
  nand g53 (n_143, in_0[5], in_1[5]);
  nand g54 (n_144, in_2[5], in_1[5]);
  nand g55 (n_145, in_0[5], in_2[5]);
  nand g56 (out_0[6], n_143, n_144, n_145);
  xor g57 (n_146, in_0[6], in_1[6]);
  xor g58 (out_1[6], n_146, in_2[6]);
  nand g59 (n_147, in_0[6], in_1[6]);
  nand g60 (n_148, in_2[6], in_1[6]);
  nand g61 (n_149, in_0[6], in_2[6]);
  nand g62 (out_0[7], n_147, n_148, n_149);
  xor g63 (n_150, in_0[7], in_1[7]);
  xor g64 (out_1[7], n_150, in_2[7]);
  nand g65 (n_151, in_0[7], in_1[7]);
  nand g66 (n_152, in_2[7], in_1[7]);
  nand g67 (n_153, in_0[7], in_2[7]);
  nand g68 (out_0[8], n_151, n_152, n_153);
  xor g69 (n_154, in_0[8], in_1[8]);
  xor g70 (out_1[8], n_154, in_2[8]);
  nand g71 (n_155, in_0[8], in_1[8]);
  nand g72 (n_156, in_2[8], in_1[8]);
  nand g73 (n_157, in_0[8], in_2[8]);
  nand g74 (out_0[9], n_155, n_156, n_157);
  xor g75 (n_158, in_0[9], in_1[9]);
  xor g76 (out_1[9], n_158, in_2[9]);
  nand g77 (n_159, in_0[9], in_1[9]);
  nand g78 (n_160, in_2[9], in_1[9]);
  nand g79 (n_161, in_0[9], in_2[9]);
  nand g80 (out_0[10], n_159, n_160, n_161);
  xor g81 (n_162, in_0[10], in_1[10]);
  xor g82 (out_1[10], n_162, in_2[10]);
  nand g83 (n_163, in_0[10], in_1[10]);
  nand g84 (n_164, in_2[10], in_1[10]);
  nand g85 (n_165, in_0[10], in_2[10]);
  nand g86 (out_0[11], n_163, n_164, n_165);
  xor g87 (n_166, in_0[11], in_1[11]);
  xor g88 (out_1[11], n_166, in_2[11]);
  nand g89 (n_167, in_0[11], in_1[11]);
  nand g90 (n_168, in_2[11], in_1[11]);
  nand g91 (n_169, in_0[11], in_2[11]);
  nand g92 (out_0[12], n_167, n_168, n_169);
  xor g93 (n_170, in_0[12], in_1[12]);
  xor g94 (out_1[12], n_170, in_2[12]);
  nand g95 (n_171, in_0[12], in_1[12]);
  nand g96 (n_172, in_2[12], in_1[12]);
  nand g97 (n_173, in_0[12], in_2[12]);
  nand g98 (out_0[13], n_171, n_172, n_173);
  xor g99 (n_174, in_0[13], in_1[13]);
  xor g100 (out_1[13], n_174, in_2[13]);
  nand g101 (n_175, in_0[13], in_1[13]);
  nand g102 (n_176, in_2[13], in_1[13]);
  nand g103 (n_177, in_0[13], in_2[13]);
  nand g104 (out_0[14], n_175, n_176, n_177);
  xor g105 (n_178, in_0[14], in_1[14]);
  xor g106 (out_1[14], n_178, in_2[14]);
  nand g107 (n_179, in_0[14], in_1[14]);
  nand g108 (n_180, in_2[14], in_1[14]);
  nand g109 (n_181, in_0[14], in_2[14]);
  nand g110 (out_0[15], n_179, n_180, n_181);
  xor g111 (n_182, in_0[15], in_1[15]);
  xor g112 (out_1[15], n_182, in_2[15]);
  nand g113 (n_183, in_0[15], in_1[15]);
  nand g114 (n_184, in_2[15], in_1[15]);
  nand g115 (n_185, in_0[15], in_2[15]);
  nand g116 (out_0[16], n_183, n_184, n_185);
  xor g117 (n_186, in_0[16], in_1[16]);
  xor g118 (out_1[16], n_186, in_2[16]);
  nand g119 (n_187, in_0[16], in_1[16]);
  nand g120 (n_188, in_2[16], in_1[16]);
  nand g121 (n_189, in_0[16], in_2[16]);
  nand g122 (out_0[17], n_187, n_188, n_189);
  xor g123 (n_190, in_0[17], in_1[17]);
  xor g124 (out_1[17], n_190, in_2[17]);
  nand g125 (n_191, in_0[17], in_1[17]);
  nand g126 (n_192, in_2[17], in_1[17]);
  nand g127 (n_193, in_0[17], in_2[17]);
  nand g128 (out_0[18], n_191, n_192, n_193);
  xor g129 (n_194, in_0[18], in_1[18]);
  xor g130 (out_1[18], n_194, in_2[18]);
  nand g131 (n_195, in_0[18], in_1[18]);
  nand g132 (n_196, in_2[18], in_1[18]);
  nand g133 (n_197, in_0[18], in_2[18]);
  nand g134 (out_0[19], n_195, n_196, n_197);
  xor g135 (n_198, in_0[19], in_1[19]);
  xor g136 (out_1[19], n_198, in_2[19]);
  nand g137 (n_199, in_0[19], in_1[19]);
  nand g138 (n_200, in_2[19], in_1[19]);
  nand g139 (n_201, in_0[19], in_2[19]);
  nand g140 (out_0[20], n_199, n_200, n_201);
  xor g141 (n_202, in_0[20], in_1[20]);
  xor g142 (out_1[20], n_202, in_2[20]);
  nand g143 (n_203, in_0[20], in_1[20]);
  nand g144 (n_204, in_2[20], in_1[20]);
  nand g145 (n_205, in_0[20], in_2[20]);
  nand g146 (out_0[21], n_203, n_204, n_205);
  xor g147 (n_206, in_0[21], in_1[21]);
  xor g148 (out_1[21], n_206, in_2[21]);
  nand g149 (n_207, in_0[21], in_1[21]);
  nand g150 (n_208, in_2[21], in_1[21]);
  nand g151 (n_209, in_0[21], in_2[21]);
  nand g152 (out_0[22], n_207, n_208, n_209);
  xor g156 (out_1[22], in_2[22], n_73);
  xor g161 (n_73, in_0[22], in_1[22]);
  nor g162 (out_0[23], in_0[22], in_1[22]);
  or g163 (n_212, in_2[22], wc);
  not gc (wc, n_73);
  or g165 (out_1[23], wc0, wc1, n_73);
  not gc1 (wc1, n_212);
  not gc0 (wc0, in_2[22]);
endmodule

module csa_tree_6719_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [22:0] in_0, in_1, in_2;
  output [25:0] out_0, out_1;
  wire [22:0] in_0, in_1, in_2;
  wire [25:0] out_0, out_1;
  csa_tree_6719_GENERIC_REAL g1(.in_0 ({in_0[21], in_0[21:0]}), .in_1
       ({in_1[21], in_1[21:0]}), .in_2 (in_2), .out_0 (out_0), .out_1
       (out_1));
endmodule

module csa_tree_6744_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 27'b0;"
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [26:0] out_0, out_1;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [26:0] out_0, out_1;
  wire n_76, n_80, n_81, n_85, n_86, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_231, n_235, n_239;
  assign out_0[0] = in_1[0];
  xor g33 (out_1[0], in_0[0], in_2[0]);
  and g34 (out_0[1], in_0[0], in_2[0]);
  xor g35 (n_141, in_0[1], in_1[1]);
  xor g36 (out_1[1], n_141, in_2[1]);
  nand g37 (n_142, in_0[1], in_1[1]);
  nand g4 (n_143, in_2[1], in_1[1]);
  nand g5 (n_144, in_0[1], in_2[1]);
  nand g38 (out_0[2], n_142, n_143, n_144);
  xor g39 (n_145, in_0[2], in_1[2]);
  xor g40 (out_1[2], n_145, in_2[2]);
  nand g41 (n_146, in_0[2], in_1[2]);
  nand g42 (n_147, in_2[2], in_1[2]);
  nand g43 (n_148, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_146, n_147, n_148);
  xor g44 (n_149, in_0[3], in_1[3]);
  xor g45 (out_1[3], n_149, in_2[3]);
  nand g46 (n_150, in_0[3], in_1[3]);
  nand g47 (n_151, in_2[3], in_1[3]);
  nand g48 (n_152, in_0[3], in_2[3]);
  nand g49 (out_0[4], n_150, n_151, n_152);
  xor g50 (n_153, in_0[4], in_1[4]);
  xor g51 (out_1[4], n_153, in_2[4]);
  nand g52 (n_154, in_0[4], in_1[4]);
  nand g53 (n_155, in_2[4], in_1[4]);
  nand g54 (n_156, in_0[4], in_2[4]);
  nand g55 (out_0[5], n_154, n_155, n_156);
  xor g56 (n_157, in_0[5], in_1[5]);
  xor g57 (out_1[5], n_157, in_2[5]);
  nand g58 (n_158, in_0[5], in_1[5]);
  nand g59 (n_159, in_2[5], in_1[5]);
  nand g60 (n_160, in_0[5], in_2[5]);
  nand g61 (out_0[6], n_158, n_159, n_160);
  xor g62 (n_161, in_0[6], in_1[6]);
  xor g63 (out_1[6], n_161, in_2[6]);
  nand g64 (n_162, in_0[6], in_1[6]);
  nand g65 (n_163, in_2[6], in_1[6]);
  nand g66 (n_164, in_0[6], in_2[6]);
  nand g67 (out_0[7], n_162, n_163, n_164);
  xor g68 (n_165, in_0[7], in_1[7]);
  xor g69 (out_1[7], n_165, in_2[7]);
  nand g70 (n_166, in_0[7], in_1[7]);
  nand g71 (n_167, in_2[7], in_1[7]);
  nand g72 (n_168, in_0[7], in_2[7]);
  nand g73 (out_0[8], n_166, n_167, n_168);
  xor g74 (n_169, in_0[8], in_1[8]);
  xor g75 (out_1[8], n_169, in_2[8]);
  nand g76 (n_170, in_0[8], in_1[8]);
  nand g77 (n_171, in_2[8], in_1[8]);
  nand g78 (n_172, in_0[8], in_2[8]);
  nand g79 (out_0[9], n_170, n_171, n_172);
  xor g80 (n_173, in_0[9], in_1[9]);
  xor g81 (out_1[9], n_173, in_2[9]);
  nand g82 (n_174, in_0[9], in_1[9]);
  nand g83 (n_175, in_2[9], in_1[9]);
  nand g84 (n_176, in_0[9], in_2[9]);
  nand g85 (out_0[10], n_174, n_175, n_176);
  xor g86 (n_177, in_0[10], in_1[10]);
  xor g87 (out_1[10], n_177, in_2[10]);
  nand g88 (n_178, in_0[10], in_1[10]);
  nand g89 (n_179, in_2[10], in_1[10]);
  nand g90 (n_180, in_0[10], in_2[10]);
  nand g91 (out_0[11], n_178, n_179, n_180);
  xor g92 (n_181, in_0[11], in_1[11]);
  xor g93 (out_1[11], n_181, in_2[11]);
  nand g94 (n_182, in_0[11], in_1[11]);
  nand g95 (n_183, in_2[11], in_1[11]);
  nand g96 (n_184, in_0[11], in_2[11]);
  nand g97 (out_0[12], n_182, n_183, n_184);
  xor g98 (n_185, in_0[12], in_1[12]);
  xor g99 (out_1[12], n_185, in_2[12]);
  nand g100 (n_186, in_0[12], in_1[12]);
  nand g101 (n_187, in_2[12], in_1[12]);
  nand g102 (n_188, in_0[12], in_2[12]);
  nand g103 (out_0[13], n_186, n_187, n_188);
  xor g104 (n_189, in_0[13], in_1[13]);
  xor g105 (out_1[13], n_189, in_2[13]);
  nand g106 (n_190, in_0[13], in_1[13]);
  nand g107 (n_191, in_2[13], in_1[13]);
  nand g108 (n_192, in_0[13], in_2[13]);
  nand g109 (out_0[14], n_190, n_191, n_192);
  xor g110 (n_193, in_0[14], in_1[14]);
  xor g111 (out_1[14], n_193, in_2[14]);
  nand g112 (n_194, in_0[14], in_1[14]);
  nand g113 (n_195, in_2[14], in_1[14]);
  nand g114 (n_196, in_0[14], in_2[14]);
  nand g115 (out_0[15], n_194, n_195, n_196);
  xor g116 (n_197, in_0[15], in_1[15]);
  xor g117 (out_1[15], n_197, in_2[15]);
  nand g118 (n_198, in_0[15], in_1[15]);
  nand g119 (n_199, in_2[15], in_1[15]);
  nand g120 (n_200, in_0[15], in_2[15]);
  nand g121 (out_0[16], n_198, n_199, n_200);
  xor g122 (n_201, in_0[16], in_1[16]);
  xor g123 (out_1[16], n_201, in_2[16]);
  nand g124 (n_202, in_0[16], in_1[16]);
  nand g125 (n_203, in_2[16], in_1[16]);
  nand g126 (n_204, in_0[16], in_2[16]);
  nand g127 (out_0[17], n_202, n_203, n_204);
  xor g128 (n_205, in_0[17], in_1[17]);
  xor g129 (out_1[17], n_205, in_2[17]);
  nand g130 (n_206, in_0[17], in_1[17]);
  nand g131 (n_207, in_2[17], in_1[17]);
  nand g132 (n_208, in_0[17], in_2[17]);
  nand g133 (out_0[18], n_206, n_207, n_208);
  xor g134 (n_209, in_0[18], in_1[18]);
  xor g135 (out_1[18], n_209, in_2[18]);
  nand g136 (n_210, in_0[18], in_1[18]);
  nand g137 (n_211, in_2[18], in_1[18]);
  nand g138 (n_212, in_0[18], in_2[18]);
  nand g139 (out_0[19], n_210, n_211, n_212);
  xor g140 (n_213, in_0[19], in_1[19]);
  xor g141 (out_1[19], n_213, in_2[19]);
  nand g142 (n_214, in_0[19], in_1[19]);
  nand g143 (n_215, in_2[19], in_1[19]);
  nand g144 (n_216, in_0[19], in_2[19]);
  nand g145 (out_0[20], n_214, n_215, n_216);
  xor g146 (n_217, in_0[20], in_1[20]);
  xor g147 (out_1[20], n_217, in_2[20]);
  nand g148 (n_218, in_0[20], in_1[20]);
  nand g149 (n_219, in_2[20], in_1[20]);
  nand g150 (n_220, in_0[20], in_2[20]);
  nand g151 (out_0[21], n_218, n_219, n_220);
  xor g152 (n_221, in_0[21], in_1[21]);
  xor g153 (out_1[21], n_221, in_2[21]);
  nand g154 (n_222, in_0[21], in_1[21]);
  nand g155 (n_223, in_2[21], in_1[21]);
  nand g156 (n_224, in_0[21], in_2[21]);
  nand g157 (out_0[22], n_222, n_223, n_224);
  xor g158 (n_225, in_0[22], in_1[22]);
  xor g159 (out_1[22], n_225, in_2[22]);
  nand g160 (n_226, in_0[22], in_1[22]);
  nand g161 (n_227, in_2[22], in_1[22]);
  nand g162 (n_228, in_0[22], in_2[22]);
  nand g163 (out_0[23], n_226, n_227, n_228);
  xor g164 (n_76, in_0[23], in_1[23]);
  and g165 (n_81, in_0[23], in_1[23]);
  xor g167 (out_1[23], in_2[23], n_76);
  xor g172 (n_80, in_0[24], in_1[24]);
  and g173 (n_86, in_0[24], in_1[24]);
  nand g177 (n_235, n_81, n_80);
  nand g185 (n_239, n_86, n_85);
  or g188 (n_231, in_2[23], wc);
  not gc (wc, n_76);
  xor g192 (n_85, in_0[25], in_1[25]);
  nor g193 (out_0[26], in_0[25], in_1[25]);
  or g195 (out_0[24], wc0, wc1, n_76);
  not gc1 (wc1, n_231);
  not gc0 (wc0, in_2[23]);
  xnor g196 (out_1[24], n_81, n_80);
  or g197 (out_0[25], wc2, n_80, n_81);
  not gc2 (wc2, n_235);
  xnor g199 (out_1[25], n_86, n_85);
  or g200 (out_1[26], n_85, wc3, n_86);
  not gc3 (wc3, n_239);
endmodule

module csa_tree_6744_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [26:0] out_0, out_1;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [26:0] out_0, out_1;
  csa_tree_6744_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_add_178_36_group_6829_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_242, n_243;
  wire n_244, n_245, n_246, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_255, n_256, n_257, n_258, n_259, n_261, n_262;
  wire n_263, n_264, n_265, n_267, n_268, n_269, n_270, n_271;
  wire n_273, n_274, n_275, n_276, n_277, n_279, n_280, n_281;
  wire n_282, n_283, n_285, n_286, n_287, n_288, n_289, n_291;
  wire n_292, n_293, n_294, n_295, n_297, n_298, n_299, n_300;
  wire n_301, n_303, n_304, n_305, n_306, n_307, n_309, n_310;
  wire n_311, n_312, n_313, n_315, n_316, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_325, n_327, n_329, n_330, n_332;
  wire n_333, n_335, n_337, n_339, n_340, n_342, n_343, n_345;
  wire n_347, n_349, n_350, n_352, n_353, n_355, n_357, n_359;
  wire n_360, n_362, n_363, n_365, n_367, n_369, n_370, n_372;
  wire n_374, n_375, n_376, n_378, n_379, n_380, n_382, n_383;
  wire n_384, n_385, n_387, n_389, n_391, n_392, n_393, n_395;
  wire n_396, n_397, n_399, n_400, n_402, n_404, n_406, n_407;
  wire n_408, n_410, n_411, n_412, n_414, n_416, n_417, n_418;
  wire n_420, n_421, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_441, n_443, n_444, n_445, n_447;
  wire n_448, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_464, n_465;
  wire n_466, n_468, n_469, n_470, n_471, n_473, n_474, n_475;
  wire n_477, n_478, n_479, n_480, n_482, n_483, n_485, n_486;
  wire n_488, n_489, n_490, n_491, n_493, n_494, n_495, n_497;
  wire n_498, n_499, n_500, n_502, n_503, n_505, n_506, n_508;
  wire n_509, n_510, n_511, n_513, n_514, n_515, n_516, n_517;
  xor g26 (n_125, in_2[1], in_0[1]);
  and g2 (n_153, in_2[1], in_0[1]);
  xor g27 (n_157, in_2[2], n_153);
  xor g28 (n_149, n_157, in_0[2]);
  nand g3 (n_124, in_2[2], n_153);
  nand g29 (n_158, in_0[2], n_153);
  nand g30 (n_126, in_2[2], in_0[2]);
  nand g31 (n_123, n_124, n_158, n_126);
  xor g32 (n_159, in_2[3], in_0[3]);
  xor g33 (n_148, n_159, in_1[3]);
  nand g34 (n_160, in_2[3], in_0[3]);
  nand g4 (n_161, in_1[3], in_0[3]);
  nand g35 (n_162, in_2[3], in_1[3]);
  nand g36 (n_122, n_160, n_161, n_162);
  xor g37 (n_163, in_2[4], in_0[4]);
  xor g38 (n_147, n_163, in_1[4]);
  nand g39 (n_164, in_2[4], in_0[4]);
  nand g40 (n_165, in_1[4], in_0[4]);
  nand g5 (n_166, in_2[4], in_1[4]);
  nand g41 (n_121, n_164, n_165, n_166);
  xor g42 (n_167, in_2[5], in_0[5]);
  xor g43 (n_146, n_167, in_1[5]);
  nand g44 (n_168, in_2[5], in_0[5]);
  nand g45 (n_169, in_1[5], in_0[5]);
  nand g46 (n_170, in_2[5], in_1[5]);
  nand g6 (n_120, n_168, n_169, n_170);
  xor g47 (n_171, in_2[6], in_0[6]);
  xor g48 (n_145, n_171, in_1[6]);
  nand g49 (n_172, in_2[6], in_0[6]);
  nand g50 (n_173, in_1[6], in_0[6]);
  nand g51 (n_174, in_2[6], in_1[6]);
  nand g52 (n_119, n_172, n_173, n_174);
  xor g53 (n_175, in_2[7], in_0[7]);
  xor g54 (n_144, n_175, in_1[7]);
  nand g55 (n_176, in_2[7], in_0[7]);
  nand g56 (n_177, in_1[7], in_0[7]);
  nand g57 (n_178, in_2[7], in_1[7]);
  nand g58 (n_118, n_176, n_177, n_178);
  xor g59 (n_179, in_2[8], in_0[8]);
  xor g60 (n_143, n_179, in_1[8]);
  nand g61 (n_180, in_2[8], in_0[8]);
  nand g62 (n_181, in_1[8], in_0[8]);
  nand g63 (n_150, in_2[8], in_1[8]);
  nand g64 (n_117, n_180, n_181, n_150);
  xor g65 (n_151, in_2[9], in_0[9]);
  xor g66 (n_142, n_151, in_1[9]);
  nand g67 (n_152, in_2[9], in_0[9]);
  nand g68 (n_182, in_1[9], in_0[9]);
  nand g69 (n_183, in_2[9], in_1[9]);
  nand g70 (n_116, n_152, n_182, n_183);
  xor g71 (n_184, in_2[10], in_0[10]);
  xor g72 (n_141, n_184, in_1[10]);
  nand g73 (n_185, in_2[10], in_0[10]);
  nand g74 (n_186, in_1[10], in_0[10]);
  nand g75 (n_187, in_2[10], in_1[10]);
  nand g76 (n_115, n_185, n_186, n_187);
  xor g77 (n_188, in_2[11], in_0[11]);
  xor g78 (n_140, n_188, in_1[11]);
  nand g79 (n_189, in_2[11], in_0[11]);
  nand g80 (n_190, in_1[11], in_0[11]);
  nand g81 (n_191, in_2[11], in_1[11]);
  nand g82 (n_114, n_189, n_190, n_191);
  xor g83 (n_192, in_2[12], in_0[12]);
  xor g84 (n_139, n_192, in_1[12]);
  nand g85 (n_193, in_2[12], in_0[12]);
  nand g86 (n_194, in_1[12], in_0[12]);
  nand g87 (n_195, in_2[12], in_1[12]);
  nand g88 (n_113, n_193, n_194, n_195);
  xor g89 (n_196, in_2[13], in_0[13]);
  xor g90 (n_138, n_196, in_1[13]);
  nand g91 (n_197, in_2[13], in_0[13]);
  nand g92 (n_198, in_1[13], in_0[13]);
  nand g93 (n_199, in_2[13], in_1[13]);
  nand g94 (n_112, n_197, n_198, n_199);
  xor g95 (n_200, in_2[14], in_0[14]);
  xor g96 (n_137, n_200, in_1[14]);
  nand g97 (n_201, in_2[14], in_0[14]);
  nand g98 (n_202, in_1[14], in_0[14]);
  nand g99 (n_203, in_2[14], in_1[14]);
  nand g100 (n_111, n_201, n_202, n_203);
  xor g101 (n_204, in_2[15], in_0[15]);
  xor g102 (n_136, n_204, in_1[15]);
  nand g103 (n_205, in_2[15], in_0[15]);
  nand g104 (n_206, in_1[15], in_0[15]);
  nand g105 (n_207, in_2[15], in_1[15]);
  nand g106 (n_110, n_205, n_206, n_207);
  xor g107 (n_208, in_2[16], in_0[16]);
  xor g108 (n_135, n_208, in_1[16]);
  nand g109 (n_209, in_2[16], in_0[16]);
  nand g110 (n_210, in_1[16], in_0[16]);
  nand g111 (n_211, in_2[16], in_1[16]);
  nand g112 (n_109, n_209, n_210, n_211);
  xor g113 (n_212, in_2[17], in_0[17]);
  xor g114 (n_134, n_212, in_1[17]);
  nand g115 (n_213, in_2[17], in_0[17]);
  nand g116 (n_214, in_1[17], in_0[17]);
  nand g117 (n_215, in_2[17], in_1[17]);
  nand g118 (n_108, n_213, n_214, n_215);
  xor g119 (n_216, in_2[18], in_0[18]);
  xor g120 (n_133, n_216, in_1[18]);
  nand g121 (n_217, in_2[18], in_0[18]);
  nand g122 (n_218, in_1[18], in_0[18]);
  nand g123 (n_219, in_2[18], in_1[18]);
  nand g124 (n_107, n_217, n_218, n_219);
  xor g125 (n_220, in_2[19], in_0[19]);
  xor g126 (n_132, n_220, in_1[19]);
  nand g127 (n_221, in_2[19], in_0[19]);
  nand g128 (n_222, in_1[19], in_0[19]);
  nand g129 (n_223, in_2[19], in_1[19]);
  nand g130 (n_106, n_221, n_222, n_223);
  xor g131 (n_224, in_2[20], in_0[20]);
  xor g132 (n_131, n_224, in_1[20]);
  nand g133 (n_225, in_2[20], in_0[20]);
  nand g134 (n_226, in_1[20], in_0[20]);
  nand g135 (n_227, in_2[20], in_1[20]);
  nand g136 (n_105, n_225, n_226, n_227);
  xor g137 (n_228, in_2[21], in_0[21]);
  xor g138 (n_130, n_228, in_1[21]);
  nand g139 (n_229, in_2[21], in_0[21]);
  nand g140 (n_230, in_1[21], in_0[21]);
  nand g141 (n_231, in_2[21], in_1[21]);
  nand g142 (n_129, n_229, n_230, n_231);
  xor g143 (n_232, in_2[22], in_0[22]);
  xor g144 (n_104, n_232, in_1[22]);
  nand g145 (n_233, in_2[22], in_0[22]);
  nand g146 (n_234, in_1[22], in_0[22]);
  nand g147 (n_235, in_2[22], in_1[22]);
  nand g148 (n_103, n_233, n_234, n_235);
  xor g151 (n_236, in_2[23], in_1[23]);
  xor g152 (n_128, n_236, in_0[23]);
  nand g153 (n_237, in_2[23], in_1[23]);
  nand g154 (n_238, in_0[23], in_1[23]);
  nand g155 (n_239, in_2[23], in_0[23]);
  nand g156 (n_127, n_237, n_238, n_239);
  xor g159 (n_517, in_0[0], in_1[0]);
  nand g160 (n_242, in_0[0], in_1[0]);
  nand g161 (n_243, in_0[0], in_2[0]);
  nand g7 (n_244, in_1[0], in_2[0]);
  nand g8 (n_246, n_242, n_243, n_244);
  nor g9 (n_245, n_125, in_1[1]);
  nand g10 (n_248, n_125, in_1[1]);
  nor g11 (n_255, in_1[2], n_149);
  nand g12 (n_250, in_1[2], n_149);
  nor g13 (n_251, n_123, n_148);
  nand g14 (n_252, n_123, n_148);
  nor g15 (n_261, n_122, n_147);
  nand g16 (n_256, n_122, n_147);
  nor g17 (n_257, n_121, n_146);
  nand g18 (n_258, n_121, n_146);
  nor g19 (n_267, n_120, n_145);
  nand g20 (n_262, n_120, n_145);
  nor g21 (n_263, n_119, n_144);
  nand g22 (n_264, n_119, n_144);
  nor g23 (n_273, n_118, n_143);
  nand g24 (n_268, n_118, n_143);
  nor g25 (n_269, n_117, n_142);
  nand g162 (n_270, n_117, n_142);
  nor g163 (n_279, n_116, n_141);
  nand g164 (n_274, n_116, n_141);
  nor g165 (n_275, n_115, n_140);
  nand g166 (n_276, n_115, n_140);
  nor g167 (n_285, n_114, n_139);
  nand g168 (n_280, n_114, n_139);
  nor g169 (n_281, n_113, n_138);
  nand g170 (n_282, n_113, n_138);
  nor g171 (n_291, n_112, n_137);
  nand g172 (n_286, n_112, n_137);
  nor g173 (n_287, n_111, n_136);
  nand g174 (n_288, n_111, n_136);
  nor g175 (n_297, n_110, n_135);
  nand g176 (n_292, n_110, n_135);
  nor g177 (n_293, n_109, n_134);
  nand g178 (n_294, n_109, n_134);
  nor g179 (n_303, n_108, n_133);
  nand g180 (n_298, n_108, n_133);
  nor g181 (n_299, n_107, n_132);
  nand g182 (n_300, n_107, n_132);
  nor g183 (n_309, n_106, n_131);
  nand g184 (n_304, n_106, n_131);
  nor g185 (n_305, n_105, n_130);
  nand g186 (n_306, n_105, n_130);
  nor g187 (n_315, n_104, n_129);
  nand g188 (n_310, n_104, n_129);
  nor g189 (n_311, n_103, n_128);
  nand g190 (n_312, n_103, n_128);
  nand g195 (n_316, n_248, n_249);
  nor g196 (n_253, n_250, n_251);
  nor g199 (n_319, n_255, n_251);
  nor g200 (n_259, n_256, n_257);
  nor g203 (n_325, n_261, n_257);
  nor g204 (n_265, n_262, n_263);
  nor g207 (n_327, n_267, n_263);
  nor g208 (n_271, n_268, n_269);
  nor g211 (n_335, n_273, n_269);
  nor g212 (n_277, n_274, n_275);
  nor g215 (n_337, n_279, n_275);
  nor g216 (n_283, n_280, n_281);
  nor g219 (n_345, n_285, n_281);
  nor g220 (n_289, n_286, n_287);
  nor g223 (n_347, n_291, n_287);
  nor g224 (n_295, n_292, n_293);
  nor g227 (n_355, n_297, n_293);
  nor g228 (n_301, n_298, n_299);
  nor g231 (n_357, n_303, n_299);
  nor g232 (n_307, n_304, n_305);
  nor g235 (n_365, n_309, n_305);
  nor g236 (n_313, n_310, n_311);
  nor g239 (n_367, n_315, n_311);
  nand g242 (n_464, n_250, n_318);
  nand g243 (n_321, n_319, n_316);
  nand g244 (n_372, n_320, n_321);
  nor g245 (n_323, n_267, n_322);
  nand g254 (n_380, n_325, n_327);
  nor g255 (n_333, n_279, n_332);
  nand g264 (n_387, n_335, n_337);
  nor g265 (n_343, n_291, n_342);
  nand g274 (n_395, n_345, n_347);
  nor g275 (n_353, n_303, n_352);
  nand g284 (n_402, n_355, n_357);
  nor g285 (n_363, n_315, n_362);
  nand g294 (n_410, n_365, n_367);
  nand g297 (n_468, n_256, n_374);
  nand g298 (n_375, n_325, n_372);
  nand g299 (n_470, n_322, n_375);
  nand g302 (n_473, n_378, n_379);
  nand g305 (n_414, n_382, n_383);
  nor g306 (n_385, n_285, n_384);
  nor g309 (n_424, n_285, n_387);
  nor g315 (n_393, n_391, n_384);
  nor g318 (n_430, n_387, n_391);
  nor g319 (n_397, n_395, n_384);
  nor g322 (n_433, n_387, n_395);
  nor g323 (n_400, n_309, n_399);
  nor g326 (n_451, n_309, n_402);
  nor g332 (n_408, n_406, n_399);
  nor g335 (n_457, n_402, n_406);
  nor g336 (n_412, n_410, n_399);
  nor g339 (n_439, n_402, n_410);
  nand g342 (n_477, n_268, n_416);
  nand g343 (n_417, n_335, n_414);
  nand g344 (n_479, n_332, n_417);
  nand g347 (n_482, n_420, n_421);
  nand g350 (n_485, n_384, n_423);
  nand g351 (n_426, n_424, n_414);
  nand g352 (n_488, n_425, n_426);
  nand g353 (n_429, n_427, n_414);
  nand g354 (n_490, n_428, n_429);
  nand g355 (n_432, n_430, n_414);
  nand g356 (n_493, n_431, n_432);
  nand g357 (n_435, n_433, n_414);
  nand g358 (n_441, n_434, n_435);
  nand g362 (n_497, n_292, n_443);
  nand g363 (n_444, n_355, n_441);
  nand g364 (n_499, n_352, n_444);
  nand g367 (n_502, n_447, n_448);
  nand g370 (n_505, n_399, n_450);
  nand g371 (n_453, n_451, n_441);
  nand g372 (n_508, n_452, n_453);
  nand g373 (n_456, n_454, n_441);
  nand g374 (n_510, n_455, n_456);
  nand g375 (n_459, n_457, n_441);
  nand g376 (n_513, n_458, n_459);
  nand g377 (n_460, n_439, n_441);
  nand g378 (n_515, n_437, n_460);
  xnor g380 (out_0[1], n_246, n_461);
  xnor g382 (out_0[2], n_316, n_462);
  xnor g385 (out_0[3], n_464, n_465);
  xnor g387 (out_0[4], n_372, n_466);
  xnor g390 (out_0[5], n_468, n_469);
  xnor g392 (out_0[6], n_470, n_471);
  xnor g395 (out_0[7], n_473, n_474);
  xnor g397 (out_0[8], n_414, n_475);
  xnor g400 (out_0[9], n_477, n_478);
  xnor g402 (out_0[10], n_479, n_480);
  xnor g405 (out_0[11], n_482, n_483);
  xnor g408 (out_0[12], n_485, n_486);
  xnor g411 (out_0[13], n_488, n_489);
  xnor g413 (out_0[14], n_490, n_491);
  xnor g416 (out_0[15], n_493, n_494);
  xnor g418 (out_0[16], n_441, n_495);
  xnor g421 (out_0[17], n_497, n_498);
  xnor g423 (out_0[18], n_499, n_500);
  xnor g426 (out_0[19], n_502, n_503);
  xnor g429 (out_0[20], n_505, n_506);
  xnor g432 (out_0[21], n_508, n_509);
  xnor g434 (out_0[22], n_510, n_511);
  xnor g437 (out_0[23], n_513, n_514);
  xnor g439 (out_0[24], n_515, n_516);
  xor g440 (out_0[0], in_2[0], n_517);
  or g441 (n_249, n_245, wc);
  not gc (wc, n_246);
  or g442 (n_461, wc0, n_245);
  not gc0 (wc0, n_248);
  and g443 (n_322, wc1, n_258);
  not gc1 (wc1, n_259);
  and g444 (n_329, wc2, n_264);
  not gc2 (wc2, n_265);
  and g445 (n_332, wc3, n_270);
  not gc3 (wc3, n_271);
  and g446 (n_339, wc4, n_276);
  not gc4 (wc4, n_277);
  and g447 (n_342, wc5, n_282);
  not gc5 (wc5, n_283);
  and g448 (n_349, wc6, n_288);
  not gc6 (wc6, n_289);
  and g449 (n_352, wc7, n_294);
  not gc7 (wc7, n_295);
  and g450 (n_359, wc8, n_300);
  not gc8 (wc8, n_301);
  and g451 (n_362, wc9, n_306);
  not gc9 (wc9, n_307);
  or g452 (n_376, wc10, n_267);
  not gc10 (wc10, n_325);
  or g453 (n_418, wc11, n_279);
  not gc11 (wc11, n_335);
  or g454 (n_391, wc12, n_291);
  not gc12 (wc12, n_345);
  or g455 (n_445, wc13, n_303);
  not gc13 (wc13, n_355);
  or g456 (n_406, wc14, n_315);
  not gc14 (wc14, n_365);
  or g457 (n_466, wc15, n_261);
  not gc15 (wc15, n_256);
  or g458 (n_469, wc16, n_257);
  not gc16 (wc16, n_258);
  or g459 (n_471, wc17, n_267);
  not gc17 (wc17, n_262);
  or g460 (n_474, wc18, n_263);
  not gc18 (wc18, n_264);
  or g461 (n_475, wc19, n_273);
  not gc19 (wc19, n_268);
  or g462 (n_478, wc20, n_269);
  not gc20 (wc20, n_270);
  or g463 (n_480, wc21, n_279);
  not gc21 (wc21, n_274);
  or g464 (n_483, wc22, n_275);
  not gc22 (wc22, n_276);
  or g465 (n_486, wc23, n_285);
  not gc23 (wc23, n_280);
  or g466 (n_489, wc24, n_281);
  not gc24 (wc24, n_282);
  or g467 (n_491, wc25, n_291);
  not gc25 (wc25, n_286);
  or g468 (n_494, wc26, n_287);
  not gc26 (wc26, n_288);
  or g469 (n_495, wc27, n_297);
  not gc27 (wc27, n_292);
  or g470 (n_498, wc28, n_293);
  not gc28 (wc28, n_294);
  or g471 (n_500, wc29, n_303);
  not gc29 (wc29, n_298);
  or g472 (n_503, wc30, n_299);
  not gc30 (wc30, n_300);
  or g473 (n_506, wc31, n_309);
  not gc31 (wc31, n_304);
  or g474 (n_509, wc32, n_305);
  not gc32 (wc32, n_306);
  or g475 (n_511, wc33, n_315);
  not gc33 (wc33, n_310);
  and g476 (n_436, wc34, n_127);
  not gc34 (wc34, in_2[23]);
  or g477 (n_438, wc35, n_127);
  not gc35 (wc35, in_2[23]);
  and g478 (n_320, wc36, n_252);
  not gc36 (wc36, n_253);
  or g479 (n_318, wc37, n_255);
  not gc37 (wc37, n_316);
  and g480 (n_330, wc38, n_327);
  not gc38 (wc38, n_322);
  and g481 (n_340, wc39, n_337);
  not gc39 (wc39, n_332);
  and g482 (n_350, wc40, n_347);
  not gc40 (wc40, n_342);
  and g483 (n_360, wc41, n_357);
  not gc41 (wc41, n_352);
  and g484 (n_427, wc42, n_345);
  not gc42 (wc42, n_387);
  and g485 (n_454, wc43, n_365);
  not gc43 (wc43, n_402);
  or g486 (n_462, wc44, n_255);
  not gc44 (wc44, n_250);
  or g487 (n_465, wc45, n_251);
  not gc45 (wc45, n_252);
  and g488 (n_369, wc46, n_312);
  not gc46 (wc46, n_313);
  and g489 (n_378, wc47, n_262);
  not gc47 (wc47, n_323);
  and g490 (n_382, wc48, n_329);
  not gc48 (wc48, n_330);
  and g491 (n_420, wc49, n_274);
  not gc49 (wc49, n_333);
  and g492 (n_384, wc50, n_339);
  not gc50 (wc50, n_340);
  and g493 (n_392, wc51, n_286);
  not gc51 (wc51, n_343);
  and g494 (n_396, wc52, n_349);
  not gc52 (wc52, n_350);
  and g495 (n_447, wc53, n_298);
  not gc53 (wc53, n_353);
  and g496 (n_399, wc54, n_359);
  not gc54 (wc54, n_360);
  and g497 (n_407, wc55, n_310);
  not gc55 (wc55, n_363);
  or g498 (n_514, wc56, n_311);
  not gc56 (wc56, n_312);
  and g499 (n_370, wc57, n_367);
  not gc57 (wc57, n_362);
  or g500 (n_374, wc58, n_261);
  not gc58 (wc58, n_372);
  or g501 (n_379, n_376, wc59);
  not gc59 (wc59, n_372);
  or g502 (n_383, n_380, wc60);
  not gc60 (wc60, n_372);
  and g503 (n_389, wc61, n_345);
  not gc61 (wc61, n_384);
  and g504 (n_404, wc62, n_365);
  not gc62 (wc62, n_399);
  or g505 (n_516, wc63, n_436);
  not gc63 (wc63, n_438);
  and g506 (n_411, wc64, n_369);
  not gc64 (wc64, n_370);
  and g507 (n_425, wc65, n_280);
  not gc65 (wc65, n_385);
  and g508 (n_428, wc66, n_342);
  not gc66 (wc66, n_389);
  and g509 (n_431, n_392, wc67);
  not gc67 (wc67, n_393);
  and g510 (n_434, n_396, wc68);
  not gc68 (wc68, n_397);
  and g511 (n_452, wc69, n_304);
  not gc69 (wc69, n_400);
  and g512 (n_455, wc70, n_362);
  not gc70 (wc70, n_404);
  and g513 (n_458, n_407, wc71);
  not gc71 (wc71, n_408);
  or g514 (n_416, wc72, n_273);
  not gc72 (wc72, n_414);
  or g515 (n_421, n_418, wc73);
  not gc73 (wc73, n_414);
  or g516 (n_423, wc74, n_387);
  not gc74 (wc74, n_414);
  and g517 (n_437, n_411, wc75);
  not gc75 (wc75, n_412);
  or g518 (n_443, wc76, n_297);
  not gc76 (wc76, n_441);
  or g519 (n_448, n_445, wc77);
  not gc77 (wc77, n_441);
  or g520 (n_450, wc78, n_402);
  not gc78 (wc78, n_441);
endmodule

module csa_tree_add_178_36_group_6829_GENERIC(in_0, in_1, in_2, out_0);
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  csa_tree_add_178_36_group_6829_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_181_36_group_6825_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_242, n_243;
  wire n_244, n_245, n_246, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_255, n_256, n_257, n_258, n_259, n_261, n_262;
  wire n_263, n_264, n_265, n_267, n_268, n_269, n_270, n_271;
  wire n_273, n_274, n_275, n_276, n_277, n_279, n_280, n_281;
  wire n_282, n_283, n_285, n_286, n_287, n_288, n_289, n_291;
  wire n_292, n_293, n_294, n_295, n_297, n_298, n_299, n_300;
  wire n_301, n_303, n_304, n_305, n_306, n_307, n_309, n_310;
  wire n_311, n_312, n_313, n_315, n_316, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_325, n_327, n_329, n_330, n_332;
  wire n_333, n_335, n_337, n_339, n_340, n_342, n_343, n_345;
  wire n_347, n_349, n_350, n_352, n_353, n_355, n_357, n_359;
  wire n_360, n_362, n_363, n_365, n_367, n_369, n_370, n_372;
  wire n_374, n_375, n_376, n_378, n_379, n_380, n_382, n_383;
  wire n_384, n_385, n_387, n_389, n_391, n_392, n_393, n_395;
  wire n_396, n_397, n_399, n_400, n_402, n_404, n_406, n_407;
  wire n_408, n_410, n_411, n_412, n_414, n_416, n_417, n_418;
  wire n_420, n_421, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_441, n_443, n_444, n_445, n_447;
  wire n_448, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_464, n_465;
  wire n_466, n_468, n_469, n_470, n_471, n_473, n_474, n_475;
  wire n_477, n_478, n_479, n_480, n_482, n_483, n_485, n_486;
  wire n_488, n_489, n_490, n_491, n_493, n_494, n_495, n_497;
  wire n_498, n_499, n_500, n_502, n_503, n_505, n_506, n_508;
  wire n_509, n_510, n_511, n_513, n_514, n_515, n_516, n_517;
  xor g26 (n_125, in_2[1], in_0[1]);
  and g2 (n_153, in_2[1], in_0[1]);
  xor g27 (n_157, in_2[2], n_153);
  xor g28 (n_149, n_157, in_0[2]);
  nand g3 (n_124, in_2[2], n_153);
  nand g29 (n_158, in_0[2], n_153);
  nand g30 (n_126, in_2[2], in_0[2]);
  nand g31 (n_123, n_124, n_158, n_126);
  xor g32 (n_159, in_2[3], in_0[3]);
  xor g33 (n_148, n_159, in_1[3]);
  nand g34 (n_160, in_2[3], in_0[3]);
  nand g4 (n_161, in_1[3], in_0[3]);
  nand g35 (n_162, in_2[3], in_1[3]);
  nand g36 (n_122, n_160, n_161, n_162);
  xor g37 (n_163, in_2[4], in_0[4]);
  xor g38 (n_147, n_163, in_1[4]);
  nand g39 (n_164, in_2[4], in_0[4]);
  nand g40 (n_165, in_1[4], in_0[4]);
  nand g5 (n_166, in_2[4], in_1[4]);
  nand g41 (n_121, n_164, n_165, n_166);
  xor g42 (n_167, in_2[5], in_0[5]);
  xor g43 (n_146, n_167, in_1[5]);
  nand g44 (n_168, in_2[5], in_0[5]);
  nand g45 (n_169, in_1[5], in_0[5]);
  nand g46 (n_170, in_2[5], in_1[5]);
  nand g6 (n_120, n_168, n_169, n_170);
  xor g47 (n_171, in_2[6], in_0[6]);
  xor g48 (n_145, n_171, in_1[6]);
  nand g49 (n_172, in_2[6], in_0[6]);
  nand g50 (n_173, in_1[6], in_0[6]);
  nand g51 (n_174, in_2[6], in_1[6]);
  nand g52 (n_119, n_172, n_173, n_174);
  xor g53 (n_175, in_2[7], in_0[7]);
  xor g54 (n_144, n_175, in_1[7]);
  nand g55 (n_176, in_2[7], in_0[7]);
  nand g56 (n_177, in_1[7], in_0[7]);
  nand g57 (n_178, in_2[7], in_1[7]);
  nand g58 (n_118, n_176, n_177, n_178);
  xor g59 (n_179, in_2[8], in_0[8]);
  xor g60 (n_143, n_179, in_1[8]);
  nand g61 (n_180, in_2[8], in_0[8]);
  nand g62 (n_181, in_1[8], in_0[8]);
  nand g63 (n_150, in_2[8], in_1[8]);
  nand g64 (n_117, n_180, n_181, n_150);
  xor g65 (n_151, in_2[9], in_0[9]);
  xor g66 (n_142, n_151, in_1[9]);
  nand g67 (n_152, in_2[9], in_0[9]);
  nand g68 (n_182, in_1[9], in_0[9]);
  nand g69 (n_183, in_2[9], in_1[9]);
  nand g70 (n_116, n_152, n_182, n_183);
  xor g71 (n_184, in_2[10], in_0[10]);
  xor g72 (n_141, n_184, in_1[10]);
  nand g73 (n_185, in_2[10], in_0[10]);
  nand g74 (n_186, in_1[10], in_0[10]);
  nand g75 (n_187, in_2[10], in_1[10]);
  nand g76 (n_115, n_185, n_186, n_187);
  xor g77 (n_188, in_2[11], in_0[11]);
  xor g78 (n_140, n_188, in_1[11]);
  nand g79 (n_189, in_2[11], in_0[11]);
  nand g80 (n_190, in_1[11], in_0[11]);
  nand g81 (n_191, in_2[11], in_1[11]);
  nand g82 (n_114, n_189, n_190, n_191);
  xor g83 (n_192, in_2[12], in_0[12]);
  xor g84 (n_139, n_192, in_1[12]);
  nand g85 (n_193, in_2[12], in_0[12]);
  nand g86 (n_194, in_1[12], in_0[12]);
  nand g87 (n_195, in_2[12], in_1[12]);
  nand g88 (n_113, n_193, n_194, n_195);
  xor g89 (n_196, in_2[13], in_0[13]);
  xor g90 (n_138, n_196, in_1[13]);
  nand g91 (n_197, in_2[13], in_0[13]);
  nand g92 (n_198, in_1[13], in_0[13]);
  nand g93 (n_199, in_2[13], in_1[13]);
  nand g94 (n_112, n_197, n_198, n_199);
  xor g95 (n_200, in_2[14], in_0[14]);
  xor g96 (n_137, n_200, in_1[14]);
  nand g97 (n_201, in_2[14], in_0[14]);
  nand g98 (n_202, in_1[14], in_0[14]);
  nand g99 (n_203, in_2[14], in_1[14]);
  nand g100 (n_111, n_201, n_202, n_203);
  xor g101 (n_204, in_2[15], in_0[15]);
  xor g102 (n_136, n_204, in_1[15]);
  nand g103 (n_205, in_2[15], in_0[15]);
  nand g104 (n_206, in_1[15], in_0[15]);
  nand g105 (n_207, in_2[15], in_1[15]);
  nand g106 (n_110, n_205, n_206, n_207);
  xor g107 (n_208, in_2[16], in_0[16]);
  xor g108 (n_135, n_208, in_1[16]);
  nand g109 (n_209, in_2[16], in_0[16]);
  nand g110 (n_210, in_1[16], in_0[16]);
  nand g111 (n_211, in_2[16], in_1[16]);
  nand g112 (n_109, n_209, n_210, n_211);
  xor g113 (n_212, in_2[17], in_0[17]);
  xor g114 (n_134, n_212, in_1[17]);
  nand g115 (n_213, in_2[17], in_0[17]);
  nand g116 (n_214, in_1[17], in_0[17]);
  nand g117 (n_215, in_2[17], in_1[17]);
  nand g118 (n_108, n_213, n_214, n_215);
  xor g119 (n_216, in_2[18], in_0[18]);
  xor g120 (n_133, n_216, in_1[18]);
  nand g121 (n_217, in_2[18], in_0[18]);
  nand g122 (n_218, in_1[18], in_0[18]);
  nand g123 (n_219, in_2[18], in_1[18]);
  nand g124 (n_107, n_217, n_218, n_219);
  xor g125 (n_220, in_2[19], in_0[19]);
  xor g126 (n_132, n_220, in_1[19]);
  nand g127 (n_221, in_2[19], in_0[19]);
  nand g128 (n_222, in_1[19], in_0[19]);
  nand g129 (n_223, in_2[19], in_1[19]);
  nand g130 (n_106, n_221, n_222, n_223);
  xor g131 (n_224, in_2[20], in_0[20]);
  xor g132 (n_131, n_224, in_1[20]);
  nand g133 (n_225, in_2[20], in_0[20]);
  nand g134 (n_226, in_1[20], in_0[20]);
  nand g135 (n_227, in_2[20], in_1[20]);
  nand g136 (n_105, n_225, n_226, n_227);
  xor g137 (n_228, in_2[21], in_0[21]);
  xor g138 (n_130, n_228, in_1[21]);
  nand g139 (n_229, in_2[21], in_0[21]);
  nand g140 (n_230, in_1[21], in_0[21]);
  nand g141 (n_231, in_2[21], in_1[21]);
  nand g142 (n_104, n_229, n_230, n_231);
  xor g143 (n_232, in_2[22], in_0[22]);
  xor g144 (n_129, n_232, in_1[22]);
  nand g145 (n_233, in_2[22], in_0[22]);
  nand g146 (n_234, in_1[22], in_0[22]);
  nand g147 (n_235, in_2[22], in_1[22]);
  nand g148 (n_103, n_233, n_234, n_235);
  xor g151 (n_236, in_2[23], in_1[23]);
  xor g152 (n_128, n_236, in_0[23]);
  nand g153 (n_237, in_2[23], in_1[23]);
  nand g154 (n_238, in_0[23], in_1[23]);
  nand g155 (n_239, in_2[23], in_0[23]);
  nand g156 (n_127, n_237, n_238, n_239);
  xor g159 (n_517, in_1[0], in_0[0]);
  nand g160 (n_242, in_1[0], in_0[0]);
  nand g161 (n_243, in_1[0], in_2[0]);
  nand g7 (n_244, in_0[0], in_2[0]);
  nand g8 (n_246, n_242, n_243, n_244);
  nor g9 (n_245, n_125, in_1[1]);
  nand g10 (n_248, n_125, in_1[1]);
  nor g11 (n_255, in_1[2], n_149);
  nand g12 (n_250, in_1[2], n_149);
  nor g13 (n_251, n_123, n_148);
  nand g14 (n_252, n_123, n_148);
  nor g15 (n_261, n_122, n_147);
  nand g16 (n_256, n_122, n_147);
  nor g17 (n_257, n_121, n_146);
  nand g18 (n_258, n_121, n_146);
  nor g19 (n_267, n_120, n_145);
  nand g20 (n_262, n_120, n_145);
  nor g21 (n_263, n_119, n_144);
  nand g22 (n_264, n_119, n_144);
  nor g23 (n_273, n_118, n_143);
  nand g24 (n_268, n_118, n_143);
  nor g25 (n_269, n_117, n_142);
  nand g162 (n_270, n_117, n_142);
  nor g163 (n_279, n_116, n_141);
  nand g164 (n_274, n_116, n_141);
  nor g165 (n_275, n_115, n_140);
  nand g166 (n_276, n_115, n_140);
  nor g167 (n_285, n_114, n_139);
  nand g168 (n_280, n_114, n_139);
  nor g169 (n_281, n_113, n_138);
  nand g170 (n_282, n_113, n_138);
  nor g171 (n_291, n_112, n_137);
  nand g172 (n_286, n_112, n_137);
  nor g173 (n_287, n_111, n_136);
  nand g174 (n_288, n_111, n_136);
  nor g175 (n_297, n_110, n_135);
  nand g176 (n_292, n_110, n_135);
  nor g177 (n_293, n_109, n_134);
  nand g178 (n_294, n_109, n_134);
  nor g179 (n_303, n_108, n_133);
  nand g180 (n_298, n_108, n_133);
  nor g181 (n_299, n_107, n_132);
  nand g182 (n_300, n_107, n_132);
  nor g183 (n_309, n_106, n_131);
  nand g184 (n_304, n_106, n_131);
  nor g185 (n_305, n_105, n_130);
  nand g186 (n_306, n_105, n_130);
  nor g187 (n_315, n_104, n_129);
  nand g188 (n_310, n_104, n_129);
  nor g189 (n_311, n_103, n_128);
  nand g190 (n_312, n_103, n_128);
  nand g195 (n_316, n_248, n_249);
  nor g196 (n_253, n_250, n_251);
  nor g199 (n_319, n_255, n_251);
  nor g200 (n_259, n_256, n_257);
  nor g203 (n_325, n_261, n_257);
  nor g204 (n_265, n_262, n_263);
  nor g207 (n_327, n_267, n_263);
  nor g208 (n_271, n_268, n_269);
  nor g211 (n_335, n_273, n_269);
  nor g212 (n_277, n_274, n_275);
  nor g215 (n_337, n_279, n_275);
  nor g216 (n_283, n_280, n_281);
  nor g219 (n_345, n_285, n_281);
  nor g220 (n_289, n_286, n_287);
  nor g223 (n_347, n_291, n_287);
  nor g224 (n_295, n_292, n_293);
  nor g227 (n_355, n_297, n_293);
  nor g228 (n_301, n_298, n_299);
  nor g231 (n_357, n_303, n_299);
  nor g232 (n_307, n_304, n_305);
  nor g235 (n_365, n_309, n_305);
  nor g236 (n_313, n_310, n_311);
  nor g239 (n_367, n_315, n_311);
  nand g242 (n_464, n_250, n_318);
  nand g243 (n_321, n_319, n_316);
  nand g244 (n_372, n_320, n_321);
  nor g245 (n_323, n_267, n_322);
  nand g254 (n_380, n_325, n_327);
  nor g255 (n_333, n_279, n_332);
  nand g264 (n_387, n_335, n_337);
  nor g265 (n_343, n_291, n_342);
  nand g274 (n_395, n_345, n_347);
  nor g275 (n_353, n_303, n_352);
  nand g284 (n_402, n_355, n_357);
  nor g285 (n_363, n_315, n_362);
  nand g294 (n_410, n_365, n_367);
  nand g297 (n_468, n_256, n_374);
  nand g298 (n_375, n_325, n_372);
  nand g299 (n_470, n_322, n_375);
  nand g302 (n_473, n_378, n_379);
  nand g305 (n_414, n_382, n_383);
  nor g306 (n_385, n_285, n_384);
  nor g309 (n_424, n_285, n_387);
  nor g315 (n_393, n_391, n_384);
  nor g318 (n_430, n_387, n_391);
  nor g319 (n_397, n_395, n_384);
  nor g322 (n_433, n_387, n_395);
  nor g323 (n_400, n_309, n_399);
  nor g326 (n_451, n_309, n_402);
  nor g332 (n_408, n_406, n_399);
  nor g335 (n_457, n_402, n_406);
  nor g336 (n_412, n_410, n_399);
  nor g339 (n_439, n_402, n_410);
  nand g342 (n_477, n_268, n_416);
  nand g343 (n_417, n_335, n_414);
  nand g344 (n_479, n_332, n_417);
  nand g347 (n_482, n_420, n_421);
  nand g350 (n_485, n_384, n_423);
  nand g351 (n_426, n_424, n_414);
  nand g352 (n_488, n_425, n_426);
  nand g353 (n_429, n_427, n_414);
  nand g354 (n_490, n_428, n_429);
  nand g355 (n_432, n_430, n_414);
  nand g356 (n_493, n_431, n_432);
  nand g357 (n_435, n_433, n_414);
  nand g358 (n_441, n_434, n_435);
  nand g362 (n_497, n_292, n_443);
  nand g363 (n_444, n_355, n_441);
  nand g364 (n_499, n_352, n_444);
  nand g367 (n_502, n_447, n_448);
  nand g370 (n_505, n_399, n_450);
  nand g371 (n_453, n_451, n_441);
  nand g372 (n_508, n_452, n_453);
  nand g373 (n_456, n_454, n_441);
  nand g374 (n_510, n_455, n_456);
  nand g375 (n_459, n_457, n_441);
  nand g376 (n_513, n_458, n_459);
  nand g377 (n_460, n_439, n_441);
  nand g378 (n_515, n_437, n_460);
  xnor g380 (out_0[1], n_246, n_461);
  xnor g382 (out_0[2], n_316, n_462);
  xnor g385 (out_0[3], n_464, n_465);
  xnor g387 (out_0[4], n_372, n_466);
  xnor g390 (out_0[5], n_468, n_469);
  xnor g392 (out_0[6], n_470, n_471);
  xnor g395 (out_0[7], n_473, n_474);
  xnor g397 (out_0[8], n_414, n_475);
  xnor g400 (out_0[9], n_477, n_478);
  xnor g402 (out_0[10], n_479, n_480);
  xnor g405 (out_0[11], n_482, n_483);
  xnor g408 (out_0[12], n_485, n_486);
  xnor g411 (out_0[13], n_488, n_489);
  xnor g413 (out_0[14], n_490, n_491);
  xnor g416 (out_0[15], n_493, n_494);
  xnor g418 (out_0[16], n_441, n_495);
  xnor g421 (out_0[17], n_497, n_498);
  xnor g423 (out_0[18], n_499, n_500);
  xnor g426 (out_0[19], n_502, n_503);
  xnor g429 (out_0[20], n_505, n_506);
  xnor g432 (out_0[21], n_508, n_509);
  xnor g434 (out_0[22], n_510, n_511);
  xnor g437 (out_0[23], n_513, n_514);
  xnor g439 (out_0[24], n_515, n_516);
  xor g440 (out_0[0], in_2[0], n_517);
  or g441 (n_249, n_245, wc);
  not gc (wc, n_246);
  or g442 (n_461, wc0, n_245);
  not gc0 (wc0, n_248);
  and g443 (n_322, wc1, n_258);
  not gc1 (wc1, n_259);
  and g444 (n_329, wc2, n_264);
  not gc2 (wc2, n_265);
  and g445 (n_332, wc3, n_270);
  not gc3 (wc3, n_271);
  and g446 (n_339, wc4, n_276);
  not gc4 (wc4, n_277);
  and g447 (n_342, wc5, n_282);
  not gc5 (wc5, n_283);
  and g448 (n_349, wc6, n_288);
  not gc6 (wc6, n_289);
  and g449 (n_352, wc7, n_294);
  not gc7 (wc7, n_295);
  and g450 (n_359, wc8, n_300);
  not gc8 (wc8, n_301);
  and g451 (n_362, wc9, n_306);
  not gc9 (wc9, n_307);
  or g452 (n_376, wc10, n_267);
  not gc10 (wc10, n_325);
  or g453 (n_418, wc11, n_279);
  not gc11 (wc11, n_335);
  or g454 (n_391, wc12, n_291);
  not gc12 (wc12, n_345);
  or g455 (n_445, wc13, n_303);
  not gc13 (wc13, n_355);
  or g456 (n_406, wc14, n_315);
  not gc14 (wc14, n_365);
  or g457 (n_466, wc15, n_261);
  not gc15 (wc15, n_256);
  or g458 (n_469, wc16, n_257);
  not gc16 (wc16, n_258);
  or g459 (n_471, wc17, n_267);
  not gc17 (wc17, n_262);
  or g460 (n_474, wc18, n_263);
  not gc18 (wc18, n_264);
  or g461 (n_475, wc19, n_273);
  not gc19 (wc19, n_268);
  or g462 (n_478, wc20, n_269);
  not gc20 (wc20, n_270);
  or g463 (n_480, wc21, n_279);
  not gc21 (wc21, n_274);
  or g464 (n_483, wc22, n_275);
  not gc22 (wc22, n_276);
  or g465 (n_486, wc23, n_285);
  not gc23 (wc23, n_280);
  or g466 (n_489, wc24, n_281);
  not gc24 (wc24, n_282);
  or g467 (n_491, wc25, n_291);
  not gc25 (wc25, n_286);
  or g468 (n_494, wc26, n_287);
  not gc26 (wc26, n_288);
  or g469 (n_495, wc27, n_297);
  not gc27 (wc27, n_292);
  or g470 (n_498, wc28, n_293);
  not gc28 (wc28, n_294);
  or g471 (n_500, wc29, n_303);
  not gc29 (wc29, n_298);
  or g472 (n_503, wc30, n_299);
  not gc30 (wc30, n_300);
  or g473 (n_506, wc31, n_309);
  not gc31 (wc31, n_304);
  or g474 (n_509, wc32, n_305);
  not gc32 (wc32, n_306);
  or g475 (n_511, wc33, n_315);
  not gc33 (wc33, n_310);
  and g476 (n_436, wc34, n_127);
  not gc34 (wc34, in_2[23]);
  or g477 (n_438, wc35, n_127);
  not gc35 (wc35, in_2[23]);
  and g478 (n_320, wc36, n_252);
  not gc36 (wc36, n_253);
  or g479 (n_318, wc37, n_255);
  not gc37 (wc37, n_316);
  and g480 (n_330, wc38, n_327);
  not gc38 (wc38, n_322);
  and g481 (n_340, wc39, n_337);
  not gc39 (wc39, n_332);
  and g482 (n_350, wc40, n_347);
  not gc40 (wc40, n_342);
  and g483 (n_360, wc41, n_357);
  not gc41 (wc41, n_352);
  and g484 (n_427, wc42, n_345);
  not gc42 (wc42, n_387);
  and g485 (n_454, wc43, n_365);
  not gc43 (wc43, n_402);
  or g486 (n_462, wc44, n_255);
  not gc44 (wc44, n_250);
  or g487 (n_465, wc45, n_251);
  not gc45 (wc45, n_252);
  and g488 (n_369, wc46, n_312);
  not gc46 (wc46, n_313);
  and g489 (n_378, wc47, n_262);
  not gc47 (wc47, n_323);
  and g490 (n_382, wc48, n_329);
  not gc48 (wc48, n_330);
  and g491 (n_420, wc49, n_274);
  not gc49 (wc49, n_333);
  and g492 (n_384, wc50, n_339);
  not gc50 (wc50, n_340);
  and g493 (n_392, wc51, n_286);
  not gc51 (wc51, n_343);
  and g494 (n_396, wc52, n_349);
  not gc52 (wc52, n_350);
  and g495 (n_447, wc53, n_298);
  not gc53 (wc53, n_353);
  and g496 (n_399, wc54, n_359);
  not gc54 (wc54, n_360);
  and g497 (n_407, wc55, n_310);
  not gc55 (wc55, n_363);
  or g498 (n_514, wc56, n_311);
  not gc56 (wc56, n_312);
  and g499 (n_370, wc57, n_367);
  not gc57 (wc57, n_362);
  or g500 (n_374, wc58, n_261);
  not gc58 (wc58, n_372);
  or g501 (n_379, n_376, wc59);
  not gc59 (wc59, n_372);
  or g502 (n_383, n_380, wc60);
  not gc60 (wc60, n_372);
  and g503 (n_389, wc61, n_345);
  not gc61 (wc61, n_384);
  and g504 (n_404, wc62, n_365);
  not gc62 (wc62, n_399);
  or g505 (n_516, wc63, n_436);
  not gc63 (wc63, n_438);
  and g506 (n_411, wc64, n_369);
  not gc64 (wc64, n_370);
  and g507 (n_425, wc65, n_280);
  not gc65 (wc65, n_385);
  and g508 (n_428, wc66, n_342);
  not gc66 (wc66, n_389);
  and g509 (n_431, n_392, wc67);
  not gc67 (wc67, n_393);
  and g510 (n_434, n_396, wc68);
  not gc68 (wc68, n_397);
  and g511 (n_452, wc69, n_304);
  not gc69 (wc69, n_400);
  and g512 (n_455, wc70, n_362);
  not gc70 (wc70, n_404);
  and g513 (n_458, n_407, wc71);
  not gc71 (wc71, n_408);
  or g514 (n_416, wc72, n_273);
  not gc72 (wc72, n_414);
  or g515 (n_421, n_418, wc73);
  not gc73 (wc73, n_414);
  or g516 (n_423, wc74, n_387);
  not gc74 (wc74, n_414);
  and g517 (n_437, n_411, wc75);
  not gc75 (wc75, n_412);
  or g518 (n_443, wc76, n_297);
  not gc76 (wc76, n_441);
  or g519 (n_448, n_445, wc77);
  not gc77 (wc77, n_441);
  or g520 (n_450, wc78, n_402);
  not gc78 (wc78, n_441);
endmodule

module csa_tree_add_181_36_group_6825_GENERIC(in_0, in_1, in_2, out_0);
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  csa_tree_add_181_36_group_6825_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_237_42_group_6823_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [20:0] in_0, in_1, in_2, in_3, in_4;
  output [23:0] out_0;
  wire [20:0] in_0, in_1, in_2, in_3, in_4;
  wire [23:0] out_0;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213;
  wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_256, n_257, n_258;
  wire n_259, n_260, n_263, n_265, n_266, n_267, n_268, n_269;
  wire n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285;
  wire n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381;
  wire n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389;
  wire n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397;
  wire n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405;
  wire n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413;
  wire n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421;
  wire n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429;
  wire n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437;
  wire n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445;
  wire n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453;
  wire n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461;
  wire n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477;
  wire n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485;
  wire n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_496, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_508, n_509, n_510, n_511, n_512, n_514, n_515;
  wire n_516, n_517, n_518, n_519, n_521, n_522, n_523, n_524;
  wire n_525, n_527, n_528, n_529, n_530, n_531, n_533, n_534;
  wire n_535, n_536, n_537, n_539, n_540, n_541, n_542, n_543;
  wire n_545, n_546, n_547, n_548, n_549, n_551, n_552, n_553;
  wire n_554, n_555, n_557, n_558, n_559, n_560, n_561, n_563;
  wire n_564, n_565, n_566, n_567, n_569, n_570, n_571, n_572;
  wire n_573, n_575, n_576, n_579, n_580, n_581, n_582, n_583;
  wire n_584, n_585, n_586, n_588, n_590, n_592, n_593, n_595;
  wire n_596, n_598, n_600, n_602, n_603, n_605, n_606, n_608;
  wire n_610, n_612, n_613, n_615, n_616, n_618, n_620, n_622;
  wire n_623, n_625, n_626, n_628, n_630, n_632, n_633, n_634;
  wire n_636, n_637, n_638, n_640, n_641, n_642, n_643, n_645;
  wire n_647, n_649, n_650, n_651, n_653, n_654, n_655, n_657;
  wire n_658, n_660, n_662, n_664, n_665, n_666, n_668, n_670;
  wire n_671, n_672, n_674, n_675, n_677, n_678, n_679, n_680;
  wire n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_692, n_693, n_694, n_696, n_697, n_699;
  wire n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_712, n_713, n_714, n_716, n_717;
  wire n_718, n_719, n_721, n_722, n_723, n_725, n_726, n_727;
  wire n_728, n_730, n_731, n_733, n_734, n_736, n_737, n_738;
  wire n_739, n_741, n_742, n_743, n_745, n_746, n_747, n_748;
  wire n_750, n_751, n_753, n_754, n_756, n_757, n_758, n_759;
  wire n_761, n_763;
  xor g69 (n_266, in_0[0], in_4[0]);
  xor g70 (n_177, n_266, in_3[0]);
  nand g71 (n_267, in_0[0], in_4[0]);
  nand g72 (n_268, in_3[0], in_4[0]);
  nand g73 (n_269, in_0[0], in_3[0]);
  nand g6 (n_179, n_267, n_268, n_269);
  xor g74 (n_270, in_0[1], in_1[1]);
  xor g75 (n_152, n_270, in_4[1]);
  nand g76 (n_271, in_0[1], in_1[1]);
  nand g77 (n_272, in_4[1], in_1[1]);
  nand g78 (n_273, in_0[1], in_4[1]);
  nand g79 (n_181, n_271, n_272, n_273);
  xor g80 (n_274, in_3[1], in_2[1]);
  xor g81 (n_176, n_274, n_179);
  nand g82 (n_275, in_3[1], in_2[1]);
  nand g83 (n_276, n_179, in_2[1]);
  nand g84 (n_277, in_3[1], n_179);
  nand g85 (n_151, n_275, n_276, n_277);
  xor g86 (n_180, in_0[2], in_1[2]);
  and g87 (n_183, in_0[2], in_1[2]);
  xor g88 (n_278, in_3[2], in_4[2]);
  xor g89 (n_182, n_278, in_2[2]);
  nand g90 (n_279, in_3[2], in_4[2]);
  nand g91 (n_280, in_2[2], in_4[2]);
  nand g92 (n_281, in_3[2], in_2[2]);
  nand g93 (n_184, n_279, n_280, n_281);
  xor g94 (n_282, n_180, n_181);
  xor g95 (n_175, n_282, n_182);
  nand g96 (n_283, n_180, n_181);
  nand g97 (n_284, n_182, n_181);
  nand g98 (n_285, n_180, n_182);
  nand g99 (n_150, n_283, n_284, n_285);
  xor g100 (n_286, in_0[3], in_1[3]);
  xor g101 (n_185, n_286, in_3[3]);
  nand g102 (n_287, in_0[3], in_1[3]);
  nand g103 (n_288, in_3[3], in_1[3]);
  nand g104 (n_289, in_0[3], in_3[3]);
  nand g105 (n_187, n_287, n_288, n_289);
  xor g106 (n_290, in_4[3], in_2[3]);
  xor g107 (n_186, n_290, n_183);
  nand g108 (n_291, in_4[3], in_2[3]);
  nand g109 (n_292, n_183, in_2[3]);
  nand g110 (n_293, in_4[3], n_183);
  nand g111 (n_189, n_291, n_292, n_293);
  xor g112 (n_294, n_184, n_185);
  xor g113 (n_174, n_294, n_186);
  nand g114 (n_295, n_184, n_185);
  nand g115 (n_296, n_186, n_185);
  nand g116 (n_297, n_184, n_186);
  nand g117 (n_149, n_295, n_296, n_297);
  xor g118 (n_298, in_0[4], in_1[4]);
  xor g119 (n_188, n_298, in_3[4]);
  nand g120 (n_299, in_0[4], in_1[4]);
  nand g121 (n_300, in_3[4], in_1[4]);
  nand g122 (n_301, in_0[4], in_3[4]);
  nand g123 (n_191, n_299, n_300, n_301);
  xor g124 (n_302, in_4[4], in_2[4]);
  xor g125 (n_190, n_302, n_187);
  nand g126 (n_303, in_4[4], in_2[4]);
  nand g127 (n_304, n_187, in_2[4]);
  nand g128 (n_305, in_4[4], n_187);
  nand g129 (n_194, n_303, n_304, n_305);
  xor g130 (n_306, n_188, n_189);
  xor g131 (n_173, n_306, n_190);
  nand g132 (n_307, n_188, n_189);
  nand g133 (n_308, n_190, n_189);
  nand g134 (n_309, n_188, n_190);
  nand g135 (n_148, n_307, n_308, n_309);
  xor g136 (n_310, in_0[5], in_1[5]);
  xor g137 (n_192, n_310, in_3[5]);
  nand g138 (n_311, in_0[5], in_1[5]);
  nand g139 (n_312, in_3[5], in_1[5]);
  nand g140 (n_313, in_0[5], in_3[5]);
  nand g141 (n_195, n_311, n_312, n_313);
  xor g142 (n_314, in_4[5], in_2[5]);
  xor g143 (n_193, n_314, n_191);
  nand g144 (n_315, in_4[5], in_2[5]);
  nand g145 (n_316, n_191, in_2[5]);
  nand g146 (n_317, in_4[5], n_191);
  nand g147 (n_198, n_315, n_316, n_317);
  xor g148 (n_318, n_192, n_193);
  xor g149 (n_172, n_318, n_194);
  nand g150 (n_319, n_192, n_193);
  nand g151 (n_320, n_194, n_193);
  nand g152 (n_321, n_192, n_194);
  nand g153 (n_147, n_319, n_320, n_321);
  xor g154 (n_322, in_0[6], in_1[6]);
  xor g155 (n_196, n_322, in_3[6]);
  nand g156 (n_323, in_0[6], in_1[6]);
  nand g157 (n_324, in_3[6], in_1[6]);
  nand g158 (n_325, in_0[6], in_3[6]);
  nand g159 (n_199, n_323, n_324, n_325);
  xor g160 (n_326, in_4[6], in_2[6]);
  xor g161 (n_197, n_326, n_195);
  nand g162 (n_327, in_4[6], in_2[6]);
  nand g163 (n_328, n_195, in_2[6]);
  nand g164 (n_329, in_4[6], n_195);
  nand g165 (n_202, n_327, n_328, n_329);
  xor g166 (n_330, n_196, n_197);
  xor g167 (n_171, n_330, n_198);
  nand g168 (n_331, n_196, n_197);
  nand g169 (n_332, n_198, n_197);
  nand g170 (n_333, n_196, n_198);
  nand g171 (n_146, n_331, n_332, n_333);
  xor g172 (n_334, in_0[7], in_1[7]);
  xor g173 (n_200, n_334, in_3[7]);
  nand g174 (n_335, in_0[7], in_1[7]);
  nand g175 (n_336, in_3[7], in_1[7]);
  nand g176 (n_337, in_0[7], in_3[7]);
  nand g177 (n_203, n_335, n_336, n_337);
  xor g178 (n_338, in_4[7], in_2[7]);
  xor g179 (n_201, n_338, n_199);
  nand g180 (n_339, in_4[7], in_2[7]);
  nand g181 (n_340, n_199, in_2[7]);
  nand g182 (n_341, in_4[7], n_199);
  nand g183 (n_206, n_339, n_340, n_341);
  xor g184 (n_342, n_200, n_201);
  xor g185 (n_170, n_342, n_202);
  nand g186 (n_343, n_200, n_201);
  nand g187 (n_344, n_202, n_201);
  nand g188 (n_345, n_200, n_202);
  nand g189 (n_145, n_343, n_344, n_345);
  xor g190 (n_346, in_0[8], in_1[8]);
  xor g191 (n_204, n_346, in_3[8]);
  nand g192 (n_347, in_0[8], in_1[8]);
  nand g193 (n_348, in_3[8], in_1[8]);
  nand g194 (n_349, in_0[8], in_3[8]);
  nand g195 (n_207, n_347, n_348, n_349);
  xor g196 (n_350, in_4[8], in_2[8]);
  xor g197 (n_205, n_350, n_203);
  nand g198 (n_351, in_4[8], in_2[8]);
  nand g199 (n_352, n_203, in_2[8]);
  nand g200 (n_353, in_4[8], n_203);
  nand g201 (n_210, n_351, n_352, n_353);
  xor g202 (n_354, n_204, n_205);
  xor g203 (n_169, n_354, n_206);
  nand g204 (n_355, n_204, n_205);
  nand g205 (n_356, n_206, n_205);
  nand g206 (n_357, n_204, n_206);
  nand g207 (n_144, n_355, n_356, n_357);
  xor g208 (n_358, in_0[9], in_1[9]);
  xor g209 (n_208, n_358, in_3[9]);
  nand g210 (n_359, in_0[9], in_1[9]);
  nand g211 (n_360, in_3[9], in_1[9]);
  nand g212 (n_361, in_0[9], in_3[9]);
  nand g213 (n_211, n_359, n_360, n_361);
  xor g214 (n_362, in_4[9], in_2[9]);
  xor g215 (n_209, n_362, n_207);
  nand g216 (n_363, in_4[9], in_2[9]);
  nand g217 (n_364, n_207, in_2[9]);
  nand g218 (n_365, in_4[9], n_207);
  nand g219 (n_214, n_363, n_364, n_365);
  xor g220 (n_366, n_208, n_209);
  xor g221 (n_168, n_366, n_210);
  nand g222 (n_367, n_208, n_209);
  nand g223 (n_368, n_210, n_209);
  nand g224 (n_369, n_208, n_210);
  nand g225 (n_143, n_367, n_368, n_369);
  xor g226 (n_370, in_0[10], in_1[10]);
  xor g227 (n_212, n_370, in_3[10]);
  nand g228 (n_371, in_0[10], in_1[10]);
  nand g229 (n_372, in_3[10], in_1[10]);
  nand g230 (n_373, in_0[10], in_3[10]);
  nand g231 (n_215, n_371, n_372, n_373);
  xor g232 (n_374, in_4[10], in_2[10]);
  xor g233 (n_213, n_374, n_211);
  nand g234 (n_375, in_4[10], in_2[10]);
  nand g235 (n_376, n_211, in_2[10]);
  nand g236 (n_377, in_4[10], n_211);
  nand g237 (n_218, n_375, n_376, n_377);
  xor g238 (n_378, n_212, n_213);
  xor g239 (n_167, n_378, n_214);
  nand g240 (n_379, n_212, n_213);
  nand g241 (n_380, n_214, n_213);
  nand g242 (n_381, n_212, n_214);
  nand g243 (n_142, n_379, n_380, n_381);
  xor g244 (n_382, in_0[11], in_1[11]);
  xor g245 (n_216, n_382, in_3[11]);
  nand g246 (n_383, in_0[11], in_1[11]);
  nand g247 (n_384, in_3[11], in_1[11]);
  nand g248 (n_385, in_0[11], in_3[11]);
  nand g249 (n_219, n_383, n_384, n_385);
  xor g250 (n_386, in_4[11], in_2[11]);
  xor g251 (n_217, n_386, n_215);
  nand g252 (n_387, in_4[11], in_2[11]);
  nand g253 (n_388, n_215, in_2[11]);
  nand g254 (n_389, in_4[11], n_215);
  nand g255 (n_222, n_387, n_388, n_389);
  xor g256 (n_390, n_216, n_217);
  xor g257 (n_166, n_390, n_218);
  nand g258 (n_391, n_216, n_217);
  nand g259 (n_392, n_218, n_217);
  nand g260 (n_393, n_216, n_218);
  nand g261 (n_141, n_391, n_392, n_393);
  xor g262 (n_394, in_0[12], in_1[12]);
  xor g263 (n_220, n_394, in_3[12]);
  nand g264 (n_395, in_0[12], in_1[12]);
  nand g265 (n_396, in_3[12], in_1[12]);
  nand g266 (n_397, in_0[12], in_3[12]);
  nand g267 (n_223, n_395, n_396, n_397);
  xor g268 (n_398, in_4[12], in_2[12]);
  xor g269 (n_221, n_398, n_219);
  nand g270 (n_399, in_4[12], in_2[12]);
  nand g271 (n_400, n_219, in_2[12]);
  nand g272 (n_401, in_4[12], n_219);
  nand g273 (n_226, n_399, n_400, n_401);
  xor g274 (n_402, n_220, n_221);
  xor g275 (n_165, n_402, n_222);
  nand g276 (n_403, n_220, n_221);
  nand g277 (n_404, n_222, n_221);
  nand g278 (n_405, n_220, n_222);
  nand g279 (n_140, n_403, n_404, n_405);
  xor g280 (n_406, in_0[13], in_1[13]);
  xor g281 (n_224, n_406, in_3[13]);
  nand g282 (n_407, in_0[13], in_1[13]);
  nand g283 (n_408, in_3[13], in_1[13]);
  nand g284 (n_409, in_0[13], in_3[13]);
  nand g285 (n_227, n_407, n_408, n_409);
  xor g286 (n_410, in_4[13], in_2[13]);
  xor g287 (n_225, n_410, n_223);
  nand g288 (n_411, in_4[13], in_2[13]);
  nand g289 (n_412, n_223, in_2[13]);
  nand g290 (n_413, in_4[13], n_223);
  nand g291 (n_230, n_411, n_412, n_413);
  xor g292 (n_414, n_224, n_225);
  xor g293 (n_164, n_414, n_226);
  nand g294 (n_415, n_224, n_225);
  nand g295 (n_416, n_226, n_225);
  nand g296 (n_417, n_224, n_226);
  nand g297 (n_139, n_415, n_416, n_417);
  xor g298 (n_418, in_0[14], in_1[14]);
  xor g299 (n_228, n_418, in_3[14]);
  nand g300 (n_419, in_0[14], in_1[14]);
  nand g301 (n_420, in_3[14], in_1[14]);
  nand g302 (n_421, in_0[14], in_3[14]);
  nand g303 (n_231, n_419, n_420, n_421);
  xor g304 (n_422, in_4[14], in_2[14]);
  xor g305 (n_229, n_422, n_227);
  nand g306 (n_423, in_4[14], in_2[14]);
  nand g307 (n_424, n_227, in_2[14]);
  nand g308 (n_425, in_4[14], n_227);
  nand g309 (n_234, n_423, n_424, n_425);
  xor g310 (n_426, n_228, n_229);
  xor g311 (n_163, n_426, n_230);
  nand g312 (n_427, n_228, n_229);
  nand g313 (n_428, n_230, n_229);
  nand g314 (n_429, n_228, n_230);
  nand g315 (n_138, n_427, n_428, n_429);
  xor g316 (n_430, in_0[15], in_1[15]);
  xor g317 (n_232, n_430, in_3[15]);
  nand g318 (n_431, in_0[15], in_1[15]);
  nand g319 (n_432, in_3[15], in_1[15]);
  nand g320 (n_433, in_0[15], in_3[15]);
  nand g321 (n_235, n_431, n_432, n_433);
  xor g322 (n_434, in_4[15], in_2[15]);
  xor g323 (n_233, n_434, n_231);
  nand g324 (n_435, in_4[15], in_2[15]);
  nand g325 (n_436, n_231, in_2[15]);
  nand g326 (n_437, in_4[15], n_231);
  nand g327 (n_238, n_435, n_436, n_437);
  xor g328 (n_438, n_232, n_233);
  xor g329 (n_162, n_438, n_234);
  nand g330 (n_439, n_232, n_233);
  nand g331 (n_440, n_234, n_233);
  nand g332 (n_441, n_232, n_234);
  nand g333 (n_137, n_439, n_440, n_441);
  xor g334 (n_442, in_0[16], in_1[16]);
  xor g335 (n_236, n_442, in_3[16]);
  nand g336 (n_443, in_0[16], in_1[16]);
  nand g337 (n_444, in_3[16], in_1[16]);
  nand g338 (n_445, in_0[16], in_3[16]);
  nand g339 (n_239, n_443, n_444, n_445);
  xor g340 (n_446, in_4[16], in_2[16]);
  xor g341 (n_237, n_446, n_235);
  nand g342 (n_447, in_4[16], in_2[16]);
  nand g343 (n_448, n_235, in_2[16]);
  nand g344 (n_449, in_4[16], n_235);
  nand g345 (n_242, n_447, n_448, n_449);
  xor g346 (n_450, n_236, n_237);
  xor g347 (n_161, n_450, n_238);
  nand g348 (n_451, n_236, n_237);
  nand g349 (n_452, n_238, n_237);
  nand g350 (n_453, n_236, n_238);
  nand g351 (n_136, n_451, n_452, n_453);
  xor g352 (n_454, in_0[17], in_1[17]);
  xor g353 (n_240, n_454, in_3[17]);
  nand g354 (n_455, in_0[17], in_1[17]);
  nand g355 (n_456, in_3[17], in_1[17]);
  nand g356 (n_457, in_0[17], in_3[17]);
  nand g357 (n_243, n_455, n_456, n_457);
  xor g358 (n_458, in_4[17], in_2[17]);
  xor g359 (n_241, n_458, n_239);
  nand g360 (n_459, in_4[17], in_2[17]);
  nand g361 (n_460, n_239, in_2[17]);
  nand g362 (n_461, in_4[17], n_239);
  nand g363 (n_246, n_459, n_460, n_461);
  xor g364 (n_462, n_240, n_241);
  xor g365 (n_160, n_462, n_242);
  nand g366 (n_463, n_240, n_241);
  nand g367 (n_464, n_242, n_241);
  nand g368 (n_465, n_240, n_242);
  nand g369 (n_135, n_463, n_464, n_465);
  xor g370 (n_466, in_0[18], in_1[18]);
  xor g371 (n_244, n_466, in_3[18]);
  nand g372 (n_467, in_0[18], in_1[18]);
  nand g373 (n_468, in_3[18], in_1[18]);
  nand g374 (n_469, in_0[18], in_3[18]);
  nand g375 (n_247, n_467, n_468, n_469);
  xor g376 (n_470, in_4[18], in_2[18]);
  xor g377 (n_245, n_470, n_243);
  nand g378 (n_471, in_4[18], in_2[18]);
  nand g379 (n_472, n_243, in_2[18]);
  nand g380 (n_473, in_4[18], n_243);
  nand g381 (n_250, n_471, n_472, n_473);
  xor g382 (n_474, n_244, n_245);
  xor g383 (n_159, n_474, n_246);
  nand g384 (n_475, n_244, n_245);
  nand g385 (n_476, n_246, n_245);
  nand g386 (n_477, n_244, n_246);
  nand g387 (n_134, n_475, n_476, n_477);
  xor g388 (n_478, in_0[19], in_1[19]);
  xor g389 (n_248, n_478, in_3[19]);
  nand g390 (n_479, in_0[19], in_1[19]);
  nand g391 (n_480, in_3[19], in_1[19]);
  nand g392 (n_481, in_0[19], in_3[19]);
  nand g393 (n_257, n_479, n_480, n_481);
  xor g394 (n_482, in_4[19], in_2[19]);
  xor g395 (n_249, n_482, n_247);
  nand g396 (n_483, in_4[19], in_2[19]);
  nand g397 (n_484, n_247, in_2[19]);
  nand g398 (n_485, in_4[19], n_247);
  nand g399 (n_260, n_483, n_484, n_485);
  xor g400 (n_486, n_248, n_249);
  xor g401 (n_158, n_486, n_250);
  nand g402 (n_487, n_248, n_249);
  nand g403 (n_488, n_250, n_249);
  nand g404 (n_489, n_248, n_250);
  nand g405 (n_133, n_487, n_488, n_489);
  nand g413 (n_263, n_491, n_492, n_493);
  nand g417 (n_496, n_257, n_256);
  xor g420 (n_498, n_258, n_259);
  xor g421 (n_157, n_498, n_260);
  nand g422 (n_499, n_258, n_259);
  nand g423 (n_500, n_260, n_259);
  nand g424 (n_501, n_258, n_260);
  nand g425 (n_132, n_499, n_500, n_501);
  xor g429 (n_156, n_502, n_265);
  nand g432 (n_505, n_263, n_265);
  nand g433 (n_155, n_503, n_504, n_505);
  xor g436 (n_763, in_1[0], n_177);
  nand g437 (n_508, in_1[0], n_177);
  nand g438 (n_509, in_1[0], in_2[0]);
  nand g7 (n_510, n_177, in_2[0]);
  nand g8 (n_512, n_508, n_509, n_510);
  nor g9 (n_511, n_152, n_176);
  nand g10 (n_514, n_152, n_176);
  nor g11 (n_521, n_151, n_175);
  nand g12 (n_516, n_151, n_175);
  nor g13 (n_517, n_150, n_174);
  nand g14 (n_518, n_150, n_174);
  nor g15 (n_527, n_149, n_173);
  nand g16 (n_522, n_149, n_173);
  nor g17 (n_523, n_148, n_172);
  nand g18 (n_524, n_148, n_172);
  nor g19 (n_533, n_147, n_171);
  nand g20 (n_528, n_147, n_171);
  nor g21 (n_529, n_146, n_170);
  nand g22 (n_530, n_146, n_170);
  nor g23 (n_539, n_145, n_169);
  nand g24 (n_534, n_145, n_169);
  nor g25 (n_535, n_144, n_168);
  nand g26 (n_536, n_144, n_168);
  nor g27 (n_545, n_143, n_167);
  nand g28 (n_540, n_143, n_167);
  nor g29 (n_541, n_142, n_166);
  nand g30 (n_542, n_142, n_166);
  nor g31 (n_551, n_141, n_165);
  nand g32 (n_546, n_141, n_165);
  nor g33 (n_547, n_140, n_164);
  nand g34 (n_548, n_140, n_164);
  nor g35 (n_557, n_139, n_163);
  nand g36 (n_552, n_139, n_163);
  nor g37 (n_553, n_138, n_162);
  nand g38 (n_554, n_138, n_162);
  nor g39 (n_563, n_137, n_161);
  nand g40 (n_558, n_137, n_161);
  nor g41 (n_559, n_136, n_160);
  nand g42 (n_560, n_136, n_160);
  nor g43 (n_569, n_135, n_159);
  nand g44 (n_564, n_135, n_159);
  nor g45 (n_565, n_134, n_158);
  nand g46 (n_566, n_134, n_158);
  nor g47 (n_575, n_133, n_157);
  nand g48 (n_570, n_133, n_157);
  nor g49 (n_571, n_132, n_156);
  nand g50 (n_572, n_132, n_156);
  nor g51 (n_579, n_131, n_155);
  nand g52 (n_576, n_131, n_155);
  nand g57 (n_580, n_514, n_515);
  nor g58 (n_519, n_516, n_517);
  nor g61 (n_582, n_521, n_517);
  nor g62 (n_525, n_522, n_523);
  nor g65 (n_588, n_527, n_523);
  nor g66 (n_531, n_528, n_529);
  nor g439 (n_590, n_533, n_529);
  nor g440 (n_537, n_534, n_535);
  nor g443 (n_598, n_539, n_535);
  nor g444 (n_543, n_540, n_541);
  nor g447 (n_600, n_545, n_541);
  nor g448 (n_549, n_546, n_547);
  nor g451 (n_608, n_551, n_547);
  nor g452 (n_555, n_552, n_553);
  nor g455 (n_610, n_557, n_553);
  nor g456 (n_561, n_558, n_559);
  nor g459 (n_618, n_563, n_559);
  nor g460 (n_567, n_564, n_565);
  nor g463 (n_620, n_569, n_565);
  nor g464 (n_573, n_570, n_571);
  nor g467 (n_628, n_575, n_571);
  nand g470 (n_712, n_516, n_581);
  nand g471 (n_584, n_582, n_580);
  nand g472 (n_630, n_583, n_584);
  nor g473 (n_586, n_533, n_585);
  nand g482 (n_638, n_588, n_590);
  nor g483 (n_596, n_545, n_595);
  nand g492 (n_645, n_598, n_600);
  nor g493 (n_606, n_557, n_605);
  nand g502 (n_653, n_608, n_610);
  nor g503 (n_616, n_569, n_615);
  nand g512 (n_660, n_618, n_620);
  nor g513 (n_626, n_579, n_625);
  nand g520 (n_716, n_522, n_632);
  nand g521 (n_633, n_588, n_630);
  nand g522 (n_718, n_585, n_633);
  nand g525 (n_721, n_636, n_637);
  nand g528 (n_668, n_640, n_641);
  nor g529 (n_643, n_551, n_642);
  nor g532 (n_678, n_551, n_645);
  nor g538 (n_651, n_649, n_642);
  nor g541 (n_684, n_645, n_649);
  nor g542 (n_655, n_653, n_642);
  nor g545 (n_687, n_645, n_653);
  nor g546 (n_658, n_575, n_657);
  nor g549 (n_700, n_575, n_660);
  nor g555 (n_666, n_664, n_657);
  nor g558 (n_706, n_660, n_664);
  nand g561 (n_725, n_534, n_670);
  nand g562 (n_671, n_598, n_668);
  nand g563 (n_727, n_595, n_671);
  nand g566 (n_730, n_674, n_675);
  nand g569 (n_733, n_642, n_677);
  nand g570 (n_680, n_678, n_668);
  nand g571 (n_736, n_679, n_680);
  nand g572 (n_683, n_681, n_668);
  nand g573 (n_738, n_682, n_683);
  nand g574 (n_686, n_684, n_668);
  nand g575 (n_741, n_685, n_686);
  nand g576 (n_689, n_687, n_668);
  nand g577 (n_690, n_688, n_689);
  nand g580 (n_745, n_558, n_692);
  nand g581 (n_693, n_618, n_690);
  nand g582 (n_747, n_615, n_693);
  nand g585 (n_750, n_696, n_697);
  nand g588 (n_753, n_657, n_699);
  nand g589 (n_702, n_700, n_690);
  nand g590 (n_756, n_701, n_702);
  nand g591 (n_705, n_703, n_690);
  nand g592 (n_758, n_704, n_705);
  nand g593 (n_708, n_706, n_690);
  nand g594 (n_761, n_707, n_708);
  xnor g596 (out_0[1], n_512, n_709);
  xnor g598 (out_0[2], n_580, n_710);
  xnor g601 (out_0[3], n_712, n_713);
  xnor g603 (out_0[4], n_630, n_714);
  xnor g606 (out_0[5], n_716, n_717);
  xnor g608 (out_0[6], n_718, n_719);
  xnor g611 (out_0[7], n_721, n_722);
  xnor g613 (out_0[8], n_668, n_723);
  xnor g616 (out_0[9], n_725, n_726);
  xnor g618 (out_0[10], n_727, n_728);
  xnor g621 (out_0[11], n_730, n_731);
  xnor g624 (out_0[12], n_733, n_734);
  xnor g627 (out_0[13], n_736, n_737);
  xnor g629 (out_0[14], n_738, n_739);
  xnor g632 (out_0[15], n_741, n_742);
  xnor g634 (out_0[16], n_690, n_743);
  xnor g637 (out_0[17], n_745, n_746);
  xnor g639 (out_0[18], n_747, n_748);
  xnor g642 (out_0[19], n_750, n_751);
  xnor g645 (out_0[20], n_753, n_754);
  xnor g648 (out_0[21], n_756, n_757);
  xnor g650 (out_0[22], n_758, n_759);
  xor g654 (out_0[0], in_2[0], n_763);
  xor g655 (n_256, in_0[20], in_1[20]);
  nor g656 (n_131, in_0[20], in_1[20]);
  xor g657 (n_490, in_3[20], in_4[20]);
  or g658 (n_491, in_3[20], in_4[20]);
  or g659 (n_492, in_2[20], in_4[20]);
  or g660 (n_493, in_2[20], in_3[20]);
  xnor g661 (n_258, n_490, in_2[20]);
  xnor g665 (n_259, n_257, n_256);
  or g666 (n_265, n_256, wc, n_257);
  not gc (wc, n_496);
  xnor g667 (n_502, n_263, n_131);
  or g668 (n_503, n_131, wc0);
  not gc0 (wc0, n_263);
  or g669 (n_504, wc1, n_131);
  not gc1 (wc1, n_265);
  or g670 (n_515, n_511, wc2);
  not gc2 (wc2, n_512);
  or g671 (n_709, wc3, n_511);
  not gc3 (wc3, n_514);
  and g672 (n_583, wc4, n_518);
  not gc4 (wc4, n_519);
  or g673 (n_710, wc5, n_521);
  not gc5 (wc5, n_516);
  or g674 (n_713, wc6, n_517);
  not gc6 (wc6, n_518);
  and g675 (n_585, wc7, n_524);
  not gc7 (wc7, n_525);
  or g676 (n_581, wc8, n_521);
  not gc8 (wc8, n_580);
  or g677 (n_714, wc9, n_527);
  not gc9 (wc9, n_522);
  or g678 (n_717, wc10, n_523);
  not gc10 (wc10, n_524);
  and g679 (n_592, wc11, n_530);
  not gc11 (wc11, n_531);
  and g680 (n_595, wc12, n_536);
  not gc12 (wc12, n_537);
  and g681 (n_602, wc13, n_542);
  not gc13 (wc13, n_543);
  and g682 (n_605, wc14, n_548);
  not gc14 (wc14, n_549);
  and g683 (n_612, wc15, n_554);
  not gc15 (wc15, n_555);
  and g684 (n_615, wc16, n_560);
  not gc16 (wc16, n_561);
  and g685 (n_622, wc17, n_566);
  not gc17 (wc17, n_567);
  and g686 (n_625, wc18, n_572);
  not gc18 (wc18, n_573);
  or g687 (n_634, wc19, n_533);
  not gc19 (wc19, n_588);
  or g688 (n_672, wc20, n_545);
  not gc20 (wc20, n_598);
  or g689 (n_649, wc21, n_557);
  not gc21 (wc21, n_608);
  or g690 (n_694, wc22, n_569);
  not gc22 (wc22, n_618);
  or g691 (n_664, wc23, n_579);
  not gc23 (wc23, n_628);
  or g692 (n_719, wc24, n_533);
  not gc24 (wc24, n_528);
  or g693 (n_722, wc25, n_529);
  not gc25 (wc25, n_530);
  or g694 (n_723, wc26, n_539);
  not gc26 (wc26, n_534);
  or g695 (n_726, wc27, n_535);
  not gc27 (wc27, n_536);
  or g696 (n_728, wc28, n_545);
  not gc28 (wc28, n_540);
  or g697 (n_731, wc29, n_541);
  not gc29 (wc29, n_542);
  or g698 (n_734, wc30, n_551);
  not gc30 (wc30, n_546);
  or g699 (n_737, wc31, n_547);
  not gc31 (wc31, n_548);
  or g700 (n_739, wc32, n_557);
  not gc32 (wc32, n_552);
  or g701 (n_742, wc33, n_553);
  not gc33 (wc33, n_554);
  or g702 (n_743, wc34, n_563);
  not gc34 (wc34, n_558);
  or g703 (n_746, wc35, n_559);
  not gc35 (wc35, n_560);
  or g704 (n_748, wc36, n_569);
  not gc36 (wc36, n_564);
  or g705 (n_751, wc37, n_565);
  not gc37 (wc37, n_566);
  or g706 (n_754, wc38, n_575);
  not gc38 (wc38, n_570);
  or g707 (n_757, wc39, n_571);
  not gc39 (wc39, n_572);
  or g708 (n_759, wc40, n_579);
  not gc40 (wc40, n_576);
  and g709 (n_636, wc41, n_528);
  not gc41 (wc41, n_586);
  and g710 (n_593, wc42, n_590);
  not gc42 (wc42, n_585);
  and g711 (n_603, wc43, n_600);
  not gc43 (wc43, n_595);
  and g712 (n_613, wc44, n_610);
  not gc44 (wc44, n_605);
  and g713 (n_623, wc45, n_620);
  not gc45 (wc45, n_615);
  or g714 (n_632, wc46, n_527);
  not gc46 (wc46, n_630);
  and g715 (n_681, wc47, n_608);
  not gc47 (wc47, n_645);
  and g716 (n_703, wc48, n_628);
  not gc48 (wc48, n_660);
  and g717 (n_640, wc49, n_592);
  not gc49 (wc49, n_593);
  and g718 (n_674, wc50, n_540);
  not gc50 (wc50, n_596);
  and g719 (n_642, wc51, n_602);
  not gc51 (wc51, n_603);
  and g720 (n_650, wc52, n_552);
  not gc52 (wc52, n_606);
  and g721 (n_654, wc53, n_612);
  not gc53 (wc53, n_613);
  and g722 (n_696, wc54, n_564);
  not gc54 (wc54, n_616);
  and g723 (n_657, wc55, n_622);
  not gc55 (wc55, n_623);
  and g724 (n_665, wc56, n_576);
  not gc56 (wc56, n_626);
  or g725 (n_637, n_634, wc57);
  not gc57 (wc57, n_630);
  or g726 (n_641, n_638, wc58);
  not gc58 (wc58, n_630);
  and g727 (n_647, wc59, n_608);
  not gc59 (wc59, n_642);
  and g728 (n_662, wc60, n_628);
  not gc60 (wc60, n_657);
  and g729 (n_679, wc61, n_546);
  not gc61 (wc61, n_643);
  and g730 (n_682, wc62, n_605);
  not gc62 (wc62, n_647);
  and g731 (n_685, n_650, wc63);
  not gc63 (wc63, n_651);
  and g732 (n_688, n_654, wc64);
  not gc64 (wc64, n_655);
  and g733 (n_701, wc65, n_570);
  not gc65 (wc65, n_658);
  and g734 (n_704, wc66, n_625);
  not gc66 (wc66, n_662);
  and g735 (n_707, n_665, wc67);
  not gc67 (wc67, n_666);
  or g736 (n_670, wc68, n_539);
  not gc68 (wc68, n_668);
  or g737 (n_675, n_672, wc69);
  not gc69 (wc69, n_668);
  or g738 (n_677, wc70, n_645);
  not gc70 (wc70, n_668);
  or g739 (n_692, wc71, n_563);
  not gc71 (wc71, n_690);
  or g740 (n_697, n_694, wc72);
  not gc72 (wc72, n_690);
  or g741 (n_699, wc73, n_660);
  not gc73 (wc73, n_690);
  not g742 (out_0[23], n_761);
endmodule

module csa_tree_add_237_42_group_6823_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [20:0] in_0, in_1, in_2, in_3, in_4;
  output [23:0] out_0;
  wire [20:0] in_0, in_1, in_2, in_3, in_4;
  wire [23:0] out_0;
  csa_tree_add_237_42_group_6823_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_284_36_group_6827_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_242, n_243;
  wire n_244, n_245, n_246, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_255, n_256, n_257, n_258, n_259, n_261, n_262;
  wire n_263, n_264, n_265, n_267, n_268, n_269, n_270, n_271;
  wire n_273, n_274, n_275, n_276, n_277, n_279, n_280, n_281;
  wire n_282, n_283, n_285, n_286, n_287, n_288, n_289, n_291;
  wire n_292, n_293, n_294, n_295, n_297, n_298, n_299, n_300;
  wire n_301, n_303, n_304, n_305, n_306, n_307, n_309, n_310;
  wire n_311, n_312, n_313, n_315, n_316, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_325, n_327, n_329, n_330, n_332;
  wire n_333, n_335, n_337, n_339, n_340, n_342, n_343, n_345;
  wire n_347, n_349, n_350, n_352, n_353, n_355, n_357, n_359;
  wire n_360, n_362, n_363, n_365, n_367, n_369, n_370, n_372;
  wire n_374, n_375, n_376, n_378, n_379, n_380, n_382, n_383;
  wire n_384, n_385, n_387, n_389, n_391, n_392, n_393, n_395;
  wire n_396, n_397, n_399, n_400, n_402, n_404, n_406, n_407;
  wire n_408, n_410, n_411, n_412, n_414, n_416, n_417, n_418;
  wire n_420, n_421, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_441, n_443, n_444, n_445, n_447;
  wire n_448, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_464, n_465;
  wire n_466, n_468, n_469, n_470, n_471, n_473, n_474, n_475;
  wire n_477, n_478, n_479, n_480, n_482, n_483, n_485, n_486;
  wire n_488, n_489, n_490, n_491, n_493, n_494, n_495, n_497;
  wire n_498, n_499, n_500, n_502, n_503, n_505, n_506, n_508;
  wire n_509, n_510, n_511, n_513, n_514, n_515, n_516, n_517;
  xor g26 (n_125, in_2[1], in_0[1]);
  and g2 (n_153, in_2[1], in_0[1]);
  xor g27 (n_123, in_2[2], n_153);
  xor g28 (n_149, n_123, in_0[2]);
  nand g3 (n_124, in_2[2], n_153);
  nand g29 (n_158, in_0[2], n_153);
  nand g30 (n_126, in_2[2], in_0[2]);
  nand g31 (n_154, n_124, n_158, n_126);
  xor g32 (n_159, in_2[3], in_0[3]);
  xor g33 (n_148, n_159, n_154);
  nand g34 (n_160, in_2[3], in_0[3]);
  nand g4 (n_161, n_154, in_0[3]);
  nand g35 (n_162, in_2[3], n_154);
  nand g36 (n_122, n_160, n_161, n_162);
  xor g37 (n_163, in_2[4], in_0[4]);
  xor g38 (n_147, n_163, in_1[4]);
  nand g39 (n_164, in_2[4], in_0[4]);
  nand g40 (n_165, in_1[4], in_0[4]);
  nand g5 (n_166, in_2[4], in_1[4]);
  nand g41 (n_121, n_164, n_165, n_166);
  xor g42 (n_167, in_2[5], in_0[5]);
  xor g43 (n_146, n_167, in_1[5]);
  nand g44 (n_168, in_2[5], in_0[5]);
  nand g45 (n_169, in_1[5], in_0[5]);
  nand g46 (n_170, in_2[5], in_1[5]);
  nand g6 (n_120, n_168, n_169, n_170);
  xor g47 (n_171, in_2[6], in_0[6]);
  xor g48 (n_145, n_171, in_1[6]);
  nand g49 (n_172, in_2[6], in_0[6]);
  nand g50 (n_173, in_1[6], in_0[6]);
  nand g51 (n_174, in_2[6], in_1[6]);
  nand g52 (n_119, n_172, n_173, n_174);
  xor g53 (n_175, in_2[7], in_0[7]);
  xor g54 (n_144, n_175, in_1[7]);
  nand g55 (n_176, in_2[7], in_0[7]);
  nand g56 (n_177, in_1[7], in_0[7]);
  nand g57 (n_178, in_2[7], in_1[7]);
  nand g58 (n_118, n_176, n_177, n_178);
  xor g59 (n_179, in_2[8], in_0[8]);
  xor g60 (n_143, n_179, in_1[8]);
  nand g61 (n_180, in_2[8], in_0[8]);
  nand g62 (n_181, in_1[8], in_0[8]);
  nand g63 (n_150, in_2[8], in_1[8]);
  nand g64 (n_117, n_180, n_181, n_150);
  xor g65 (n_151, in_2[9], in_0[9]);
  xor g66 (n_142, n_151, in_1[9]);
  nand g67 (n_152, in_2[9], in_0[9]);
  nand g68 (n_182, in_1[9], in_0[9]);
  nand g69 (n_183, in_2[9], in_1[9]);
  nand g70 (n_116, n_152, n_182, n_183);
  xor g71 (n_184, in_2[10], in_0[10]);
  xor g72 (n_141, n_184, in_1[10]);
  nand g73 (n_185, in_2[10], in_0[10]);
  nand g74 (n_186, in_1[10], in_0[10]);
  nand g75 (n_187, in_2[10], in_1[10]);
  nand g76 (n_115, n_185, n_186, n_187);
  xor g77 (n_188, in_2[11], in_0[11]);
  xor g78 (n_140, n_188, in_1[11]);
  nand g79 (n_189, in_2[11], in_0[11]);
  nand g80 (n_190, in_1[11], in_0[11]);
  nand g81 (n_191, in_2[11], in_1[11]);
  nand g82 (n_114, n_189, n_190, n_191);
  xor g83 (n_192, in_2[12], in_0[12]);
  xor g84 (n_139, n_192, in_1[12]);
  nand g85 (n_193, in_2[12], in_0[12]);
  nand g86 (n_194, in_1[12], in_0[12]);
  nand g87 (n_195, in_2[12], in_1[12]);
  nand g88 (n_113, n_193, n_194, n_195);
  xor g89 (n_196, in_2[13], in_0[13]);
  xor g90 (n_138, n_196, in_1[13]);
  nand g91 (n_197, in_2[13], in_0[13]);
  nand g92 (n_198, in_1[13], in_0[13]);
  nand g93 (n_199, in_2[13], in_1[13]);
  nand g94 (n_112, n_197, n_198, n_199);
  xor g95 (n_200, in_2[14], in_0[14]);
  xor g96 (n_137, n_200, in_1[14]);
  nand g97 (n_201, in_2[14], in_0[14]);
  nand g98 (n_202, in_1[14], in_0[14]);
  nand g99 (n_203, in_2[14], in_1[14]);
  nand g100 (n_111, n_201, n_202, n_203);
  xor g101 (n_204, in_2[15], in_0[15]);
  xor g102 (n_136, n_204, in_1[15]);
  nand g103 (n_205, in_2[15], in_0[15]);
  nand g104 (n_206, in_1[15], in_0[15]);
  nand g105 (n_207, in_2[15], in_1[15]);
  nand g106 (n_110, n_205, n_206, n_207);
  xor g107 (n_208, in_2[16], in_0[16]);
  xor g108 (n_135, n_208, in_1[16]);
  nand g109 (n_209, in_2[16], in_0[16]);
  nand g110 (n_210, in_1[16], in_0[16]);
  nand g111 (n_211, in_2[16], in_1[16]);
  nand g112 (n_109, n_209, n_210, n_211);
  xor g113 (n_212, in_2[17], in_0[17]);
  xor g114 (n_134, n_212, in_1[17]);
  nand g115 (n_213, in_2[17], in_0[17]);
  nand g116 (n_214, in_1[17], in_0[17]);
  nand g117 (n_215, in_2[17], in_1[17]);
  nand g118 (n_108, n_213, n_214, n_215);
  xor g119 (n_216, in_2[18], in_0[18]);
  xor g120 (n_133, n_216, in_1[18]);
  nand g121 (n_217, in_2[18], in_0[18]);
  nand g122 (n_218, in_1[18], in_0[18]);
  nand g123 (n_219, in_2[18], in_1[18]);
  nand g124 (n_107, n_217, n_218, n_219);
  xor g125 (n_220, in_2[19], in_0[19]);
  xor g126 (n_132, n_220, in_1[19]);
  nand g127 (n_221, in_2[19], in_0[19]);
  nand g128 (n_222, in_1[19], in_0[19]);
  nand g129 (n_223, in_2[19], in_1[19]);
  nand g130 (n_131, n_221, n_222, n_223);
  xor g131 (n_224, in_2[20], in_0[20]);
  xor g132 (n_106, n_224, in_1[20]);
  nand g133 (n_225, in_2[20], in_0[20]);
  nand g134 (n_226, in_1[20], in_0[20]);
  nand g135 (n_227, in_2[20], in_1[20]);
  nand g136 (n_105, n_225, n_226, n_227);
  xor g137 (n_228, in_2[21], in_0[21]);
  xor g138 (n_130, n_228, in_1[21]);
  nand g139 (n_229, in_2[21], in_0[21]);
  nand g140 (n_230, in_1[21], in_0[21]);
  nand g141 (n_231, in_2[21], in_1[21]);
  nand g142 (n_104, n_229, n_230, n_231);
  xor g143 (n_232, in_2[22], in_0[22]);
  xor g144 (n_129, n_232, in_1[22]);
  nand g145 (n_233, in_2[22], in_0[22]);
  nand g146 (n_234, in_1[22], in_0[22]);
  nand g147 (n_235, in_2[22], in_1[22]);
  nand g148 (n_128, n_233, n_234, n_235);
  xor g151 (n_236, in_2[23], in_1[23]);
  xor g152 (n_103, n_236, in_0[23]);
  nand g153 (n_237, in_2[23], in_1[23]);
  nand g154 (n_238, in_0[23], in_1[23]);
  nand g155 (n_239, in_2[23], in_0[23]);
  nand g156 (n_127, n_237, n_238, n_239);
  xor g159 (n_517, in_1[0], in_0[0]);
  nand g160 (n_242, in_1[0], in_0[0]);
  nand g161 (n_243, in_1[0], in_2[0]);
  nand g7 (n_244, in_0[0], in_2[0]);
  nand g8 (n_246, n_242, n_243, n_244);
  nor g9 (n_245, n_125, in_1[1]);
  nand g10 (n_248, n_125, in_1[1]);
  nor g11 (n_255, in_1[2], n_149);
  nand g12 (n_250, in_1[2], n_149);
  nor g13 (n_251, in_1[3], n_148);
  nand g14 (n_252, in_1[3], n_148);
  nor g15 (n_261, n_122, n_147);
  nand g16 (n_256, n_122, n_147);
  nor g17 (n_257, n_121, n_146);
  nand g18 (n_258, n_121, n_146);
  nor g19 (n_267, n_120, n_145);
  nand g20 (n_262, n_120, n_145);
  nor g21 (n_263, n_119, n_144);
  nand g22 (n_264, n_119, n_144);
  nor g23 (n_273, n_118, n_143);
  nand g24 (n_268, n_118, n_143);
  nor g25 (n_269, n_117, n_142);
  nand g162 (n_270, n_117, n_142);
  nor g163 (n_279, n_116, n_141);
  nand g164 (n_274, n_116, n_141);
  nor g165 (n_275, n_115, n_140);
  nand g166 (n_276, n_115, n_140);
  nor g167 (n_285, n_114, n_139);
  nand g168 (n_280, n_114, n_139);
  nor g169 (n_281, n_113, n_138);
  nand g170 (n_282, n_113, n_138);
  nor g171 (n_291, n_112, n_137);
  nand g172 (n_286, n_112, n_137);
  nor g173 (n_287, n_111, n_136);
  nand g174 (n_288, n_111, n_136);
  nor g175 (n_297, n_110, n_135);
  nand g176 (n_292, n_110, n_135);
  nor g177 (n_293, n_109, n_134);
  nand g178 (n_294, n_109, n_134);
  nor g179 (n_303, n_108, n_133);
  nand g180 (n_298, n_108, n_133);
  nor g181 (n_299, n_107, n_132);
  nand g182 (n_300, n_107, n_132);
  nor g183 (n_309, n_106, n_131);
  nand g184 (n_304, n_106, n_131);
  nor g185 (n_305, n_105, n_130);
  nand g186 (n_306, n_105, n_130);
  nor g187 (n_315, n_104, n_129);
  nand g188 (n_310, n_104, n_129);
  nor g189 (n_311, n_103, n_128);
  nand g190 (n_312, n_103, n_128);
  nand g195 (n_316, n_248, n_249);
  nor g196 (n_253, n_250, n_251);
  nor g199 (n_319, n_255, n_251);
  nor g200 (n_259, n_256, n_257);
  nor g203 (n_325, n_261, n_257);
  nor g204 (n_265, n_262, n_263);
  nor g207 (n_327, n_267, n_263);
  nor g208 (n_271, n_268, n_269);
  nor g211 (n_335, n_273, n_269);
  nor g212 (n_277, n_274, n_275);
  nor g215 (n_337, n_279, n_275);
  nor g216 (n_283, n_280, n_281);
  nor g219 (n_345, n_285, n_281);
  nor g220 (n_289, n_286, n_287);
  nor g223 (n_347, n_291, n_287);
  nor g224 (n_295, n_292, n_293);
  nor g227 (n_355, n_297, n_293);
  nor g228 (n_301, n_298, n_299);
  nor g231 (n_357, n_303, n_299);
  nor g232 (n_307, n_304, n_305);
  nor g235 (n_365, n_309, n_305);
  nor g236 (n_313, n_310, n_311);
  nor g239 (n_367, n_315, n_311);
  nand g242 (n_464, n_250, n_318);
  nand g243 (n_321, n_319, n_316);
  nand g244 (n_372, n_320, n_321);
  nor g245 (n_323, n_267, n_322);
  nand g254 (n_380, n_325, n_327);
  nor g255 (n_333, n_279, n_332);
  nand g264 (n_387, n_335, n_337);
  nor g265 (n_343, n_291, n_342);
  nand g274 (n_395, n_345, n_347);
  nor g275 (n_353, n_303, n_352);
  nand g284 (n_402, n_355, n_357);
  nor g285 (n_363, n_315, n_362);
  nand g294 (n_410, n_365, n_367);
  nand g297 (n_468, n_256, n_374);
  nand g298 (n_375, n_325, n_372);
  nand g299 (n_470, n_322, n_375);
  nand g302 (n_473, n_378, n_379);
  nand g305 (n_414, n_382, n_383);
  nor g306 (n_385, n_285, n_384);
  nor g309 (n_424, n_285, n_387);
  nor g315 (n_393, n_391, n_384);
  nor g318 (n_430, n_387, n_391);
  nor g319 (n_397, n_395, n_384);
  nor g322 (n_433, n_387, n_395);
  nor g323 (n_400, n_309, n_399);
  nor g326 (n_451, n_309, n_402);
  nor g332 (n_408, n_406, n_399);
  nor g335 (n_457, n_402, n_406);
  nor g336 (n_412, n_410, n_399);
  nor g339 (n_439, n_402, n_410);
  nand g342 (n_477, n_268, n_416);
  nand g343 (n_417, n_335, n_414);
  nand g344 (n_479, n_332, n_417);
  nand g347 (n_482, n_420, n_421);
  nand g350 (n_485, n_384, n_423);
  nand g351 (n_426, n_424, n_414);
  nand g352 (n_488, n_425, n_426);
  nand g353 (n_429, n_427, n_414);
  nand g354 (n_490, n_428, n_429);
  nand g355 (n_432, n_430, n_414);
  nand g356 (n_493, n_431, n_432);
  nand g357 (n_435, n_433, n_414);
  nand g358 (n_441, n_434, n_435);
  nand g362 (n_497, n_292, n_443);
  nand g363 (n_444, n_355, n_441);
  nand g364 (n_499, n_352, n_444);
  nand g367 (n_502, n_447, n_448);
  nand g370 (n_505, n_399, n_450);
  nand g371 (n_453, n_451, n_441);
  nand g372 (n_508, n_452, n_453);
  nand g373 (n_456, n_454, n_441);
  nand g374 (n_510, n_455, n_456);
  nand g375 (n_459, n_457, n_441);
  nand g376 (n_513, n_458, n_459);
  nand g377 (n_460, n_439, n_441);
  nand g378 (n_515, n_437, n_460);
  xnor g380 (out_0[1], n_246, n_461);
  xnor g382 (out_0[2], n_316, n_462);
  xnor g385 (out_0[3], n_464, n_465);
  xnor g387 (out_0[4], n_372, n_466);
  xnor g390 (out_0[5], n_468, n_469);
  xnor g392 (out_0[6], n_470, n_471);
  xnor g395 (out_0[7], n_473, n_474);
  xnor g397 (out_0[8], n_414, n_475);
  xnor g400 (out_0[9], n_477, n_478);
  xnor g402 (out_0[10], n_479, n_480);
  xnor g405 (out_0[11], n_482, n_483);
  xnor g408 (out_0[12], n_485, n_486);
  xnor g411 (out_0[13], n_488, n_489);
  xnor g413 (out_0[14], n_490, n_491);
  xnor g416 (out_0[15], n_493, n_494);
  xnor g418 (out_0[16], n_441, n_495);
  xnor g421 (out_0[17], n_497, n_498);
  xnor g423 (out_0[18], n_499, n_500);
  xnor g426 (out_0[19], n_502, n_503);
  xnor g429 (out_0[20], n_505, n_506);
  xnor g432 (out_0[21], n_508, n_509);
  xnor g434 (out_0[22], n_510, n_511);
  xnor g437 (out_0[23], n_513, n_514);
  xnor g439 (out_0[24], n_515, n_516);
  xor g440 (out_0[0], in_2[0], n_517);
  or g441 (n_249, n_245, wc);
  not gc (wc, n_246);
  or g442 (n_461, wc0, n_245);
  not gc0 (wc0, n_248);
  and g443 (n_329, wc1, n_264);
  not gc1 (wc1, n_265);
  and g444 (n_332, wc2, n_270);
  not gc2 (wc2, n_271);
  and g445 (n_339, wc3, n_276);
  not gc3 (wc3, n_277);
  and g446 (n_342, wc4, n_282);
  not gc4 (wc4, n_283);
  and g447 (n_349, wc5, n_288);
  not gc5 (wc5, n_289);
  and g448 (n_352, wc6, n_294);
  not gc6 (wc6, n_295);
  and g449 (n_359, wc7, n_300);
  not gc7 (wc7, n_301);
  and g450 (n_362, wc8, n_306);
  not gc8 (wc8, n_307);
  or g451 (n_418, wc9, n_279);
  not gc9 (wc9, n_335);
  or g452 (n_391, wc10, n_291);
  not gc10 (wc10, n_345);
  or g453 (n_445, wc11, n_303);
  not gc11 (wc11, n_355);
  or g454 (n_406, wc12, n_315);
  not gc12 (wc12, n_365);
  or g455 (n_469, wc13, n_257);
  not gc13 (wc13, n_258);
  or g456 (n_471, wc14, n_267);
  not gc14 (wc14, n_262);
  or g457 (n_474, wc15, n_263);
  not gc15 (wc15, n_264);
  or g458 (n_475, wc16, n_273);
  not gc16 (wc16, n_268);
  or g459 (n_478, wc17, n_269);
  not gc17 (wc17, n_270);
  or g460 (n_480, wc18, n_279);
  not gc18 (wc18, n_274);
  or g461 (n_483, wc19, n_275);
  not gc19 (wc19, n_276);
  or g462 (n_486, wc20, n_285);
  not gc20 (wc20, n_280);
  or g463 (n_489, wc21, n_281);
  not gc21 (wc21, n_282);
  or g464 (n_491, wc22, n_291);
  not gc22 (wc22, n_286);
  or g465 (n_494, wc23, n_287);
  not gc23 (wc23, n_288);
  or g466 (n_495, wc24, n_297);
  not gc24 (wc24, n_292);
  or g467 (n_498, wc25, n_293);
  not gc25 (wc25, n_294);
  or g468 (n_500, wc26, n_303);
  not gc26 (wc26, n_298);
  or g469 (n_503, wc27, n_299);
  not gc27 (wc27, n_300);
  or g470 (n_506, wc28, n_309);
  not gc28 (wc28, n_304);
  or g471 (n_509, wc29, n_305);
  not gc29 (wc29, n_306);
  or g472 (n_511, wc30, n_315);
  not gc30 (wc30, n_310);
  and g473 (n_436, wc31, n_127);
  not gc31 (wc31, in_2[23]);
  or g474 (n_438, wc32, n_127);
  not gc32 (wc32, in_2[23]);
  or g475 (n_318, wc33, n_255);
  not gc33 (wc33, n_316);
  and g476 (n_340, wc34, n_337);
  not gc34 (wc34, n_332);
  and g477 (n_350, wc35, n_347);
  not gc35 (wc35, n_342);
  and g478 (n_360, wc36, n_357);
  not gc36 (wc36, n_352);
  and g479 (n_427, wc37, n_345);
  not gc37 (wc37, n_387);
  and g480 (n_454, wc38, n_365);
  not gc38 (wc38, n_402);
  or g481 (n_462, wc39, n_255);
  not gc39 (wc39, n_250);
  and g482 (n_320, wc40, n_252);
  not gc40 (wc40, n_253);
  and g483 (n_369, wc41, n_312);
  not gc41 (wc41, n_313);
  and g484 (n_420, wc42, n_274);
  not gc42 (wc42, n_333);
  and g485 (n_384, wc43, n_339);
  not gc43 (wc43, n_340);
  and g486 (n_392, wc44, n_286);
  not gc44 (wc44, n_343);
  and g487 (n_396, wc45, n_349);
  not gc45 (wc45, n_350);
  and g488 (n_447, wc46, n_298);
  not gc46 (wc46, n_353);
  and g489 (n_399, wc47, n_359);
  not gc47 (wc47, n_360);
  and g490 (n_407, wc48, n_310);
  not gc48 (wc48, n_363);
  or g491 (n_465, wc49, n_251);
  not gc49 (wc49, n_252);
  or g492 (n_514, wc50, n_311);
  not gc50 (wc50, n_312);
  and g493 (n_322, wc51, n_258);
  not gc51 (wc51, n_259);
  or g494 (n_376, wc52, n_267);
  not gc52 (wc52, n_325);
  and g495 (n_370, wc53, n_367);
  not gc53 (wc53, n_362);
  and g496 (n_389, wc54, n_345);
  not gc54 (wc54, n_384);
  and g497 (n_404, wc55, n_365);
  not gc55 (wc55, n_399);
  or g498 (n_466, wc56, n_261);
  not gc56 (wc56, n_256);
  or g499 (n_516, wc57, n_436);
  not gc57 (wc57, n_438);
  and g500 (n_330, wc58, n_327);
  not gc58 (wc58, n_322);
  and g501 (n_411, wc59, n_369);
  not gc59 (wc59, n_370);
  or g502 (n_374, wc60, n_261);
  not gc60 (wc60, n_372);
  and g503 (n_425, wc61, n_280);
  not gc61 (wc61, n_385);
  and g504 (n_428, wc62, n_342);
  not gc62 (wc62, n_389);
  and g505 (n_431, n_392, wc63);
  not gc63 (wc63, n_393);
  and g506 (n_434, n_396, wc64);
  not gc64 (wc64, n_397);
  and g507 (n_452, wc65, n_304);
  not gc65 (wc65, n_400);
  and g508 (n_455, wc66, n_362);
  not gc66 (wc66, n_404);
  and g509 (n_458, n_407, wc67);
  not gc67 (wc67, n_408);
  and g510 (n_378, wc68, n_262);
  not gc68 (wc68, n_323);
  and g511 (n_382, wc69, n_329);
  not gc69 (wc69, n_330);
  or g512 (n_379, n_376, wc70);
  not gc70 (wc70, n_372);
  or g513 (n_383, n_380, wc71);
  not gc71 (wc71, n_372);
  and g514 (n_437, n_411, wc72);
  not gc72 (wc72, n_412);
  or g515 (n_416, wc73, n_273);
  not gc73 (wc73, n_414);
  or g516 (n_421, n_418, wc74);
  not gc74 (wc74, n_414);
  or g517 (n_423, wc75, n_387);
  not gc75 (wc75, n_414);
  or g518 (n_443, wc76, n_297);
  not gc76 (wc76, n_441);
  or g519 (n_448, n_445, wc77);
  not gc77 (wc77, n_441);
  or g520 (n_450, wc78, n_402);
  not gc78 (wc78, n_441);
endmodule

module csa_tree_add_284_36_group_6827_GENERIC(in_0, in_1, in_2, out_0);
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  csa_tree_add_284_36_group_6827_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_287_40_group_6803_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [26:0] in_0, in_1;
  input [24:0] in_2;
  output [25:0] out_0;
  wire [26:0] in_0, in_1;
  wire [24:0] in_2;
  wire [25:0] out_0;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_163, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213;
  wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_252, n_253, n_254, n_255;
  wire n_256, n_258, n_259, n_260, n_261, n_262, n_263, n_265;
  wire n_266, n_267, n_268, n_269, n_271, n_272, n_273, n_274;
  wire n_275, n_277, n_278, n_279, n_280, n_281, n_283, n_284;
  wire n_285, n_286, n_287, n_289, n_290, n_291, n_292, n_293;
  wire n_295, n_296, n_297, n_298, n_299, n_301, n_302, n_303;
  wire n_304, n_305, n_307, n_308, n_309, n_310, n_311, n_313;
  wire n_314, n_315, n_316, n_317, n_319, n_320, n_321, n_322;
  wire n_323, n_325, n_326, n_327, n_328, n_329, n_330, n_332;
  wire n_333, n_334, n_335, n_336, n_337, n_339, n_341, n_343;
  wire n_344, n_346, n_347, n_349, n_351, n_353, n_354, n_356;
  wire n_357, n_359, n_361, n_363, n_364, n_366, n_367, n_369;
  wire n_371, n_373, n_374, n_376, n_377, n_379, n_381, n_383;
  wire n_384, n_386, n_388, n_389, n_390, n_392, n_393, n_394;
  wire n_396, n_397, n_398, n_399, n_401, n_403, n_405, n_406;
  wire n_407, n_409, n_410, n_411, n_413, n_414, n_416, n_418;
  wire n_420, n_421, n_422, n_424, n_425, n_426, n_428, n_430;
  wire n_431, n_432, n_434, n_435, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_453, n_455, n_457, n_458, n_459;
  wire n_461, n_462, n_464, n_465, n_466, n_467, n_468, n_469;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_477, n_478;
  wire n_479, n_480, n_482, n_483, n_484, n_486, n_487, n_488;
  wire n_489, n_491, n_492, n_493, n_495, n_496, n_497, n_498;
  wire n_500, n_501, n_503, n_504, n_506, n_507, n_508, n_509;
  wire n_511, n_512, n_513, n_515, n_516, n_517, n_518, n_520;
  wire n_521, n_523, n_524, n_526, n_527, n_528, n_529, n_531;
  wire n_532, n_533, n_534, n_536, n_537, n_538;
  xor g27 (n_130, in_2[1], in_0[1]);
  and g2 (n_159, in_2[1], in_0[1]);
  xor g28 (n_163, in_2[2], n_159);
  xor g29 (n_155, n_163, in_0[2]);
  nand g3 (n_129, in_2[2], n_159);
  nand g30 (n_164, in_0[2], n_159);
  nand g31 (n_131, in_2[2], in_0[2]);
  nand g32 (n_128, n_129, n_164, n_131);
  xor g33 (n_165, in_2[3], in_0[3]);
  xor g34 (n_154, n_165, in_1[3]);
  nand g35 (n_166, in_2[3], in_0[3]);
  nand g4 (n_167, in_1[3], in_0[3]);
  nand g36 (n_168, in_2[3], in_1[3]);
  nand g37 (n_127, n_166, n_167, n_168);
  xor g38 (n_169, in_2[4], in_0[4]);
  xor g39 (n_153, n_169, in_1[4]);
  nand g40 (n_170, in_2[4], in_0[4]);
  nand g41 (n_171, in_1[4], in_0[4]);
  nand g5 (n_172, in_2[4], in_1[4]);
  nand g42 (n_126, n_170, n_171, n_172);
  xor g43 (n_173, in_2[5], in_0[5]);
  xor g44 (n_152, n_173, in_1[5]);
  nand g45 (n_174, in_2[5], in_0[5]);
  nand g46 (n_175, in_1[5], in_0[5]);
  nand g47 (n_176, in_2[5], in_1[5]);
  nand g6 (n_125, n_174, n_175, n_176);
  xor g48 (n_177, in_2[6], in_0[6]);
  xor g49 (n_151, n_177, in_1[6]);
  nand g50 (n_178, in_2[6], in_0[6]);
  nand g51 (n_179, in_1[6], in_0[6]);
  nand g52 (n_180, in_2[6], in_1[6]);
  nand g53 (n_124, n_178, n_179, n_180);
  xor g54 (n_181, in_2[7], in_0[7]);
  xor g55 (n_150, n_181, in_1[7]);
  nand g56 (n_182, in_2[7], in_0[7]);
  nand g57 (n_183, in_1[7], in_0[7]);
  nand g58 (n_184, in_2[7], in_1[7]);
  nand g59 (n_123, n_182, n_183, n_184);
  xor g60 (n_185, in_2[8], in_0[8]);
  xor g61 (n_149, n_185, in_1[8]);
  nand g62 (n_186, in_2[8], in_0[8]);
  nand g63 (n_187, in_1[8], in_0[8]);
  nand g64 (n_188, in_2[8], in_1[8]);
  nand g65 (n_122, n_186, n_187, n_188);
  xor g66 (n_156, in_2[9], in_0[9]);
  xor g67 (n_148, n_156, in_1[9]);
  nand g68 (n_157, in_2[9], in_0[9]);
  nand g69 (n_158, in_1[9], in_0[9]);
  nand g70 (n_189, in_2[9], in_1[9]);
  nand g71 (n_121, n_157, n_158, n_189);
  xor g72 (n_190, in_2[10], in_0[10]);
  xor g73 (n_147, n_190, in_1[10]);
  nand g74 (n_191, in_2[10], in_0[10]);
  nand g75 (n_192, in_1[10], in_0[10]);
  nand g76 (n_193, in_2[10], in_1[10]);
  nand g77 (n_120, n_191, n_192, n_193);
  xor g78 (n_194, in_2[11], in_0[11]);
  xor g79 (n_146, n_194, in_1[11]);
  nand g80 (n_195, in_2[11], in_0[11]);
  nand g81 (n_196, in_1[11], in_0[11]);
  nand g82 (n_197, in_2[11], in_1[11]);
  nand g83 (n_119, n_195, n_196, n_197);
  xor g84 (n_198, in_2[12], in_0[12]);
  xor g85 (n_145, n_198, in_1[12]);
  nand g86 (n_199, in_2[12], in_0[12]);
  nand g87 (n_200, in_1[12], in_0[12]);
  nand g88 (n_201, in_2[12], in_1[12]);
  nand g89 (n_118, n_199, n_200, n_201);
  xor g90 (n_202, in_2[13], in_0[13]);
  xor g91 (n_144, n_202, in_1[13]);
  nand g92 (n_203, in_2[13], in_0[13]);
  nand g93 (n_204, in_1[13], in_0[13]);
  nand g94 (n_205, in_2[13], in_1[13]);
  nand g95 (n_117, n_203, n_204, n_205);
  xor g96 (n_206, in_2[14], in_0[14]);
  xor g97 (n_143, n_206, in_1[14]);
  nand g98 (n_207, in_2[14], in_0[14]);
  nand g99 (n_208, in_1[14], in_0[14]);
  nand g100 (n_209, in_2[14], in_1[14]);
  nand g101 (n_116, n_207, n_208, n_209);
  xor g102 (n_210, in_2[15], in_0[15]);
  xor g103 (n_142, n_210, in_1[15]);
  nand g104 (n_211, in_2[15], in_0[15]);
  nand g105 (n_212, in_1[15], in_0[15]);
  nand g106 (n_213, in_2[15], in_1[15]);
  nand g107 (n_115, n_211, n_212, n_213);
  xor g108 (n_214, in_2[16], in_0[16]);
  xor g109 (n_141, n_214, in_1[16]);
  nand g110 (n_215, in_2[16], in_0[16]);
  nand g111 (n_216, in_1[16], in_0[16]);
  nand g112 (n_217, in_2[16], in_1[16]);
  nand g113 (n_114, n_215, n_216, n_217);
  xor g114 (n_218, in_2[17], in_0[17]);
  xor g115 (n_140, n_218, in_1[17]);
  nand g116 (n_219, in_2[17], in_0[17]);
  nand g117 (n_220, in_1[17], in_0[17]);
  nand g118 (n_221, in_2[17], in_1[17]);
  nand g119 (n_113, n_219, n_220, n_221);
  xor g120 (n_222, in_2[18], in_0[18]);
  xor g121 (n_139, n_222, in_1[18]);
  nand g122 (n_223, in_2[18], in_0[18]);
  nand g123 (n_224, in_1[18], in_0[18]);
  nand g124 (n_225, in_2[18], in_1[18]);
  nand g125 (n_112, n_223, n_224, n_225);
  xor g126 (n_226, in_2[19], in_0[19]);
  xor g127 (n_138, n_226, in_1[19]);
  nand g128 (n_227, in_2[19], in_0[19]);
  nand g129 (n_228, in_1[19], in_0[19]);
  nand g130 (n_229, in_2[19], in_1[19]);
  nand g131 (n_111, n_227, n_228, n_229);
  xor g132 (n_230, in_2[20], in_0[20]);
  xor g133 (n_137, n_230, in_1[20]);
  nand g134 (n_231, in_2[20], in_0[20]);
  nand g135 (n_232, in_1[20], in_0[20]);
  nand g136 (n_233, in_2[20], in_1[20]);
  nand g137 (n_110, n_231, n_232, n_233);
  xor g138 (n_234, in_2[21], in_0[21]);
  xor g139 (n_136, n_234, in_1[21]);
  nand g140 (n_235, in_2[21], in_0[21]);
  nand g141 (n_236, in_1[21], in_0[21]);
  nand g142 (n_237, in_2[21], in_1[21]);
  nand g143 (n_109, n_235, n_236, n_237);
  xor g144 (n_238, in_2[22], in_0[22]);
  xor g145 (n_135, n_238, in_1[22]);
  nand g146 (n_239, in_2[22], in_0[22]);
  nand g147 (n_240, in_1[22], in_0[22]);
  nand g148 (n_241, in_2[22], in_1[22]);
  nand g149 (n_108, n_239, n_240, n_241);
  xor g150 (n_242, in_2[23], in_0[23]);
  xor g151 (n_134, n_242, in_1[23]);
  nand g152 (n_243, in_2[23], in_0[23]);
  nand g153 (n_244, in_1[23], in_0[23]);
  nand g154 (n_245, in_2[23], in_1[23]);
  nand g155 (n_107, n_243, n_244, n_245);
  xor g158 (n_246, in_2[24], in_1[24]);
  xor g159 (n_133, n_246, in_0[24]);
  nand g160 (n_247, in_2[24], in_1[24]);
  nand g161 (n_248, in_0[24], in_1[24]);
  nand g162 (n_249, in_2[24], in_0[24]);
  nand g163 (n_132, n_247, n_248, n_249);
  xor g166 (n_538, in_1[0], in_0[0]);
  nand g167 (n_252, in_1[0], in_0[0]);
  nand g168 (n_253, in_1[0], in_2[0]);
  nand g7 (n_254, in_0[0], in_2[0]);
  nand g8 (n_256, n_252, n_253, n_254);
  nor g9 (n_255, n_130, in_1[1]);
  nand g10 (n_258, n_130, in_1[1]);
  nor g11 (n_265, in_1[2], n_155);
  nand g12 (n_260, in_1[2], n_155);
  nor g13 (n_261, n_128, n_154);
  nand g14 (n_262, n_128, n_154);
  nor g15 (n_271, n_127, n_153);
  nand g16 (n_266, n_127, n_153);
  nor g17 (n_267, n_126, n_152);
  nand g18 (n_268, n_126, n_152);
  nor g19 (n_277, n_125, n_151);
  nand g20 (n_272, n_125, n_151);
  nor g21 (n_273, n_124, n_150);
  nand g22 (n_274, n_124, n_150);
  nor g23 (n_283, n_123, n_149);
  nand g24 (n_278, n_123, n_149);
  nor g25 (n_279, n_122, n_148);
  nand g26 (n_280, n_122, n_148);
  nor g169 (n_289, n_121, n_147);
  nand g170 (n_284, n_121, n_147);
  nor g171 (n_285, n_120, n_146);
  nand g172 (n_286, n_120, n_146);
  nor g173 (n_295, n_119, n_145);
  nand g174 (n_290, n_119, n_145);
  nor g175 (n_291, n_118, n_144);
  nand g176 (n_292, n_118, n_144);
  nor g177 (n_301, n_117, n_143);
  nand g178 (n_296, n_117, n_143);
  nor g179 (n_297, n_116, n_142);
  nand g180 (n_298, n_116, n_142);
  nor g181 (n_307, n_115, n_141);
  nand g182 (n_302, n_115, n_141);
  nor g183 (n_303, n_114, n_140);
  nand g184 (n_304, n_114, n_140);
  nor g185 (n_313, n_113, n_139);
  nand g186 (n_308, n_113, n_139);
  nor g187 (n_309, n_112, n_138);
  nand g188 (n_310, n_112, n_138);
  nor g189 (n_319, n_111, n_137);
  nand g190 (n_314, n_111, n_137);
  nor g191 (n_315, n_110, n_136);
  nand g192 (n_316, n_110, n_136);
  nor g193 (n_325, n_109, n_135);
  nand g194 (n_320, n_109, n_135);
  nor g195 (n_321, n_108, n_134);
  nand g196 (n_322, n_108, n_134);
  nor g197 (n_329, n_107, n_133);
  nand g198 (n_326, n_107, n_133);
  nand g203 (n_330, n_258, n_259);
  nor g204 (n_263, n_260, n_261);
  nor g207 (n_333, n_265, n_261);
  nor g208 (n_269, n_266, n_267);
  nor g211 (n_339, n_271, n_267);
  nor g212 (n_275, n_272, n_273);
  nor g215 (n_341, n_277, n_273);
  nor g216 (n_281, n_278, n_279);
  nor g219 (n_349, n_283, n_279);
  nor g220 (n_287, n_284, n_285);
  nor g223 (n_351, n_289, n_285);
  nor g224 (n_293, n_290, n_291);
  nor g227 (n_359, n_295, n_291);
  nor g228 (n_299, n_296, n_297);
  nor g231 (n_361, n_301, n_297);
  nor g232 (n_305, n_302, n_303);
  nor g235 (n_369, n_307, n_303);
  nor g236 (n_311, n_308, n_309);
  nor g239 (n_371, n_313, n_309);
  nor g240 (n_317, n_314, n_315);
  nor g243 (n_379, n_319, n_315);
  nor g244 (n_323, n_320, n_321);
  nor g247 (n_381, n_325, n_321);
  nand g250 (n_482, n_260, n_332);
  nand g251 (n_335, n_333, n_330);
  nand g252 (n_386, n_334, n_335);
  nor g253 (n_337, n_277, n_336);
  nand g262 (n_394, n_339, n_341);
  nor g263 (n_347, n_289, n_346);
  nand g272 (n_401, n_349, n_351);
  nor g273 (n_357, n_301, n_356);
  nand g282 (n_409, n_359, n_361);
  nor g283 (n_367, n_313, n_366);
  nand g292 (n_416, n_369, n_371);
  nor g293 (n_377, n_325, n_376);
  nand g302 (n_424, n_379, n_381);
  nand g305 (n_486, n_266, n_388);
  nand g306 (n_389, n_339, n_386);
  nand g307 (n_488, n_336, n_389);
  nand g310 (n_491, n_392, n_393);
  nand g313 (n_428, n_396, n_397);
  nor g314 (n_399, n_295, n_398);
  nor g317 (n_438, n_295, n_401);
  nor g323 (n_407, n_405, n_398);
  nor g326 (n_444, n_401, n_405);
  nor g327 (n_411, n_409, n_398);
  nor g330 (n_447, n_401, n_409);
  nor g331 (n_414, n_319, n_413);
  nor g334 (n_465, n_319, n_416);
  nor g340 (n_422, n_420, n_413);
  nor g343 (n_471, n_416, n_420);
  nor g344 (n_426, n_424, n_413);
  nor g347 (n_453, n_416, n_424);
  nand g350 (n_495, n_278, n_430);
  nand g351 (n_431, n_349, n_428);
  nand g352 (n_497, n_346, n_431);
  nand g355 (n_500, n_434, n_435);
  nand g358 (n_503, n_398, n_437);
  nand g359 (n_440, n_438, n_428);
  nand g360 (n_506, n_439, n_440);
  nand g361 (n_443, n_441, n_428);
  nand g362 (n_508, n_442, n_443);
  nand g363 (n_446, n_444, n_428);
  nand g364 (n_511, n_445, n_446);
  nand g365 (n_449, n_447, n_428);
  nand g366 (n_455, n_448, n_449);
  nor g367 (n_451, n_329, n_450);
  nand g374 (n_515, n_302, n_457);
  nand g375 (n_458, n_369, n_455);
  nand g376 (n_517, n_366, n_458);
  nand g379 (n_520, n_461, n_462);
  nand g382 (n_523, n_413, n_464);
  nand g383 (n_467, n_465, n_455);
  nand g384 (n_526, n_466, n_467);
  nand g385 (n_470, n_468, n_455);
  nand g386 (n_528, n_469, n_470);
  nand g387 (n_473, n_471, n_455);
  nand g388 (n_531, n_472, n_473);
  nand g389 (n_474, n_453, n_455);
  nand g390 (n_533, n_450, n_474);
  nand g393 (n_536, n_477, n_478);
  xnor g395 (out_0[1], n_256, n_479);
  xnor g397 (out_0[2], n_330, n_480);
  xnor g400 (out_0[3], n_482, n_483);
  xnor g402 (out_0[4], n_386, n_484);
  xnor g405 (out_0[5], n_486, n_487);
  xnor g407 (out_0[6], n_488, n_489);
  xnor g410 (out_0[7], n_491, n_492);
  xnor g412 (out_0[8], n_428, n_493);
  xnor g415 (out_0[9], n_495, n_496);
  xnor g417 (out_0[10], n_497, n_498);
  xnor g420 (out_0[11], n_500, n_501);
  xnor g423 (out_0[12], n_503, n_504);
  xnor g426 (out_0[13], n_506, n_507);
  xnor g428 (out_0[14], n_508, n_509);
  xnor g431 (out_0[15], n_511, n_512);
  xnor g433 (out_0[16], n_455, n_513);
  xnor g436 (out_0[17], n_515, n_516);
  xnor g438 (out_0[18], n_517, n_518);
  xnor g441 (out_0[19], n_520, n_521);
  xnor g444 (out_0[20], n_523, n_524);
  xnor g447 (out_0[21], n_526, n_527);
  xnor g449 (out_0[22], n_528, n_529);
  xnor g452 (out_0[23], n_531, n_532);
  xnor g454 (out_0[24], n_533, n_534);
  xnor g457 (out_0[25], n_536, n_537);
  xor g458 (out_0[0], in_2[0], n_538);
  or g459 (n_259, n_255, wc);
  not gc (wc, n_256);
  or g460 (n_479, wc0, n_255);
  not gc0 (wc0, n_258);
  and g461 (n_336, wc1, n_268);
  not gc1 (wc1, n_269);
  and g462 (n_343, wc2, n_274);
  not gc2 (wc2, n_275);
  and g463 (n_346, wc3, n_280);
  not gc3 (wc3, n_281);
  and g464 (n_353, wc4, n_286);
  not gc4 (wc4, n_287);
  and g465 (n_356, wc5, n_292);
  not gc5 (wc5, n_293);
  and g466 (n_363, wc6, n_298);
  not gc6 (wc6, n_299);
  and g467 (n_366, wc7, n_304);
  not gc7 (wc7, n_305);
  and g468 (n_373, wc8, n_310);
  not gc8 (wc8, n_311);
  and g469 (n_376, wc9, n_316);
  not gc9 (wc9, n_317);
  and g470 (n_383, wc10, n_322);
  not gc10 (wc10, n_323);
  or g471 (n_390, wc11, n_277);
  not gc11 (wc11, n_339);
  or g472 (n_432, wc12, n_289);
  not gc12 (wc12, n_349);
  or g473 (n_405, wc13, n_301);
  not gc13 (wc13, n_359);
  or g474 (n_459, wc14, n_313);
  not gc14 (wc14, n_369);
  or g475 (n_420, wc15, n_325);
  not gc15 (wc15, n_379);
  or g476 (n_484, wc16, n_271);
  not gc16 (wc16, n_266);
  or g477 (n_487, wc17, n_267);
  not gc17 (wc17, n_268);
  or g478 (n_489, wc18, n_277);
  not gc18 (wc18, n_272);
  or g479 (n_492, wc19, n_273);
  not gc19 (wc19, n_274);
  or g480 (n_493, wc20, n_283);
  not gc20 (wc20, n_278);
  or g481 (n_496, wc21, n_279);
  not gc21 (wc21, n_280);
  or g482 (n_498, wc22, n_289);
  not gc22 (wc22, n_284);
  or g483 (n_501, wc23, n_285);
  not gc23 (wc23, n_286);
  or g484 (n_504, wc24, n_295);
  not gc24 (wc24, n_290);
  or g485 (n_507, wc25, n_291);
  not gc25 (wc25, n_292);
  or g486 (n_509, wc26, n_301);
  not gc26 (wc26, n_296);
  or g487 (n_512, wc27, n_297);
  not gc27 (wc27, n_298);
  or g488 (n_513, wc28, n_307);
  not gc28 (wc28, n_302);
  or g489 (n_516, wc29, n_303);
  not gc29 (wc29, n_304);
  or g490 (n_518, wc30, n_313);
  not gc30 (wc30, n_308);
  or g491 (n_521, wc31, n_309);
  not gc31 (wc31, n_310);
  or g492 (n_524, wc32, n_319);
  not gc32 (wc32, n_314);
  or g493 (n_527, wc33, n_315);
  not gc33 (wc33, n_316);
  or g494 (n_529, wc34, n_325);
  not gc34 (wc34, n_320);
  or g495 (n_532, wc35, n_321);
  not gc35 (wc35, n_322);
  and g496 (n_327, wc36, n_132);
  not gc36 (wc36, in_2[24]);
  or g497 (n_328, wc37, n_132);
  not gc37 (wc37, in_2[24]);
  and g498 (n_334, wc38, n_262);
  not gc38 (wc38, n_263);
  or g499 (n_332, wc39, n_265);
  not gc39 (wc39, n_330);
  and g500 (n_344, wc40, n_341);
  not gc40 (wc40, n_336);
  and g501 (n_354, wc41, n_351);
  not gc41 (wc41, n_346);
  and g502 (n_364, wc42, n_361);
  not gc42 (wc42, n_356);
  and g503 (n_374, wc43, n_371);
  not gc43 (wc43, n_366);
  and g504 (n_384, wc44, n_381);
  not gc44 (wc44, n_376);
  and g505 (n_441, wc45, n_359);
  not gc45 (wc45, n_401);
  and g506 (n_468, wc46, n_379);
  not gc46 (wc46, n_416);
  or g507 (n_480, wc47, n_265);
  not gc47 (wc47, n_260);
  or g508 (n_483, wc48, n_261);
  not gc48 (wc48, n_262);
  and g509 (n_392, wc49, n_272);
  not gc49 (wc49, n_337);
  and g510 (n_396, wc50, n_343);
  not gc50 (wc50, n_344);
  and g511 (n_434, wc51, n_284);
  not gc51 (wc51, n_347);
  and g512 (n_398, wc52, n_353);
  not gc52 (wc52, n_354);
  and g513 (n_406, wc53, n_296);
  not gc53 (wc53, n_357);
  and g514 (n_410, wc54, n_363);
  not gc54 (wc54, n_364);
  and g515 (n_461, wc55, n_308);
  not gc55 (wc55, n_367);
  and g516 (n_413, wc56, n_373);
  not gc56 (wc56, n_374);
  and g517 (n_421, wc57, n_320);
  not gc57 (wc57, n_377);
  and g518 (n_425, wc58, n_383);
  not gc58 (wc58, n_384);
  or g519 (n_475, wc59, n_329);
  not gc59 (wc59, n_453);
  or g520 (n_534, wc60, n_329);
  not gc60 (wc60, n_326);
  or g521 (n_388, wc61, n_271);
  not gc61 (wc61, n_386);
  or g522 (n_393, n_390, wc62);
  not gc62 (wc62, n_386);
  or g523 (n_397, n_394, wc63);
  not gc63 (wc63, n_386);
  and g524 (n_403, wc64, n_359);
  not gc64 (wc64, n_398);
  and g525 (n_418, wc65, n_379);
  not gc65 (wc65, n_413);
  or g526 (n_537, wc66, n_327);
  not gc66 (wc66, n_328);
  and g527 (n_439, wc67, n_290);
  not gc67 (wc67, n_399);
  and g528 (n_442, wc68, n_356);
  not gc68 (wc68, n_403);
  and g529 (n_445, n_406, wc69);
  not gc69 (wc69, n_407);
  and g530 (n_448, n_410, wc70);
  not gc70 (wc70, n_411);
  and g531 (n_466, wc71, n_314);
  not gc71 (wc71, n_414);
  and g532 (n_469, wc72, n_376);
  not gc72 (wc72, n_418);
  and g533 (n_472, n_421, wc73);
  not gc73 (wc73, n_422);
  and g534 (n_450, n_425, wc74);
  not gc74 (wc74, n_426);
  or g535 (n_430, wc75, n_283);
  not gc75 (wc75, n_428);
  or g536 (n_435, n_432, wc76);
  not gc76 (wc76, n_428);
  or g537 (n_437, wc77, n_401);
  not gc77 (wc77, n_428);
  and g538 (n_477, wc78, n_326);
  not gc78 (wc78, n_451);
  or g539 (n_457, wc79, n_307);
  not gc79 (wc79, n_455);
  or g540 (n_462, n_459, wc80);
  not gc80 (wc80, n_455);
  or g541 (n_464, wc81, n_416);
  not gc81 (wc81, n_455);
  or g542 (n_478, n_475, wc82);
  not gc82 (wc82, n_455);
endmodule

module csa_tree_add_287_40_group_6803_GENERIC(in_0, in_1, in_2, out_0);
  input [26:0] in_0, in_1;
  input [24:0] in_2;
  output [25:0] out_0;
  wire [26:0] in_0, in_1;
  wire [24:0] in_2;
  wire [25:0] out_0;
  csa_tree_add_287_40_group_6803_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_311_38_group_6821_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_311_38_group_6821_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_311_38_group_6821_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_384_38_group_6813_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_384_38_group_6813_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_384_38_group_6813_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_457_38_group_6815_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_457_38_group_6815_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_457_38_group_6815_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_530_38_group_6817_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_530_38_group_6817_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_530_38_group_6817_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_603_38_group_6819_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_603_38_group_6819_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_603_38_group_6819_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_676_38_group_6811_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_676_38_group_6811_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_676_38_group_6811_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_749_44_group_6809_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_280, n_281, n_282, n_283, n_284, n_287;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_544, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_556, n_557;
  wire n_558, n_559, n_560, n_562, n_563, n_564, n_565, n_566;
  wire n_567, n_569, n_570, n_571, n_572, n_573, n_575, n_576;
  wire n_577, n_578, n_579, n_581, n_582, n_583, n_584, n_585;
  wire n_587, n_588, n_589, n_590, n_591, n_593, n_594, n_595;
  wire n_596, n_597, n_599, n_600, n_601, n_602, n_603, n_605;
  wire n_606, n_607, n_608, n_609, n_611, n_612, n_613, n_614;
  wire n_615, n_617, n_618, n_619, n_620, n_621, n_623, n_624;
  wire n_625, n_626, n_627, n_629, n_630, n_633, n_634, n_636;
  wire n_637, n_638, n_639, n_640, n_642, n_644, n_646, n_647;
  wire n_649, n_650, n_652, n_654, n_656, n_657, n_659, n_660;
  wire n_662, n_664, n_666, n_667, n_669, n_670, n_672, n_674;
  wire n_676, n_677, n_679, n_680, n_682, n_684, n_686, n_687;
  wire n_689, n_691, n_692, n_693, n_695, n_696, n_697, n_699;
  wire n_700, n_701, n_702, n_704, n_706, n_708, n_709, n_710;
  wire n_712, n_713, n_714, n_716, n_717, n_719, n_721, n_723;
  wire n_724, n_725, n_727, n_728, n_729, n_731, n_733, n_734;
  wire n_735, n_737, n_738, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_756, n_758, n_760, n_761, n_762, n_764;
  wire n_765, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_780, n_781, n_782;
  wire n_783, n_785, n_786, n_787, n_789, n_790, n_791, n_792;
  wire n_794, n_795, n_796, n_798, n_799, n_800, n_801, n_803;
  wire n_804, n_806, n_807, n_809, n_810, n_811, n_812, n_814;
  wire n_815, n_816, n_818, n_819, n_820, n_821, n_823, n_824;
  wire n_826, n_827, n_829, n_830, n_831, n_832, n_834, n_835;
  wire n_836, n_837, n_839, n_841;
  xor g75 (n_290, in_0[0], in_4[0]);
  xor g76 (n_193, n_290, in_3[0]);
  nand g77 (n_291, in_0[0], in_4[0]);
  nand g78 (n_292, in_3[0], in_4[0]);
  nand g79 (n_293, in_0[0], in_3[0]);
  nand g6 (n_195, n_291, n_292, n_293);
  xor g80 (n_294, in_0[1], in_1[1]);
  xor g81 (n_166, n_294, in_4[1]);
  nand g82 (n_295, in_0[1], in_1[1]);
  nand g83 (n_296, in_4[1], in_1[1]);
  nand g84 (n_297, in_0[1], in_4[1]);
  nand g85 (n_197, n_295, n_296, n_297);
  xor g86 (n_298, in_3[1], in_2[1]);
  xor g87 (n_192, n_298, n_195);
  nand g88 (n_299, in_3[1], in_2[1]);
  nand g89 (n_300, n_195, in_2[1]);
  nand g90 (n_301, in_3[1], n_195);
  nand g91 (n_165, n_299, n_300, n_301);
  xor g92 (n_196, in_0[2], in_1[2]);
  and g93 (n_199, in_0[2], in_1[2]);
  xor g94 (n_302, in_3[2], in_4[2]);
  xor g95 (n_198, n_302, in_2[2]);
  nand g96 (n_303, in_3[2], in_4[2]);
  nand g97 (n_304, in_2[2], in_4[2]);
  nand g98 (n_305, in_3[2], in_2[2]);
  nand g99 (n_200, n_303, n_304, n_305);
  xor g100 (n_306, n_196, n_197);
  xor g101 (n_191, n_306, n_198);
  nand g102 (n_307, n_196, n_197);
  nand g103 (n_308, n_198, n_197);
  nand g104 (n_309, n_196, n_198);
  nand g105 (n_164, n_307, n_308, n_309);
  xor g106 (n_310, in_0[3], in_1[3]);
  xor g107 (n_201, n_310, in_3[3]);
  nand g108 (n_311, in_0[3], in_1[3]);
  nand g109 (n_312, in_3[3], in_1[3]);
  nand g110 (n_313, in_0[3], in_3[3]);
  nand g111 (n_203, n_311, n_312, n_313);
  xor g112 (n_314, in_4[3], in_2[3]);
  xor g113 (n_202, n_314, n_199);
  nand g114 (n_315, in_4[3], in_2[3]);
  nand g115 (n_316, n_199, in_2[3]);
  nand g116 (n_317, in_4[3], n_199);
  nand g117 (n_205, n_315, n_316, n_317);
  xor g118 (n_318, n_200, n_201);
  xor g119 (n_190, n_318, n_202);
  nand g120 (n_319, n_200, n_201);
  nand g121 (n_320, n_202, n_201);
  nand g122 (n_321, n_200, n_202);
  nand g123 (n_163, n_319, n_320, n_321);
  xor g124 (n_322, in_0[4], in_1[4]);
  xor g125 (n_204, n_322, in_3[4]);
  nand g126 (n_323, in_0[4], in_1[4]);
  nand g127 (n_324, in_3[4], in_1[4]);
  nand g128 (n_325, in_0[4], in_3[4]);
  nand g129 (n_207, n_323, n_324, n_325);
  xor g130 (n_326, in_4[4], in_2[4]);
  xor g131 (n_206, n_326, n_203);
  nand g132 (n_327, in_4[4], in_2[4]);
  nand g133 (n_328, n_203, in_2[4]);
  nand g134 (n_329, in_4[4], n_203);
  nand g135 (n_210, n_327, n_328, n_329);
  xor g136 (n_330, n_204, n_205);
  xor g137 (n_189, n_330, n_206);
  nand g138 (n_331, n_204, n_205);
  nand g139 (n_332, n_206, n_205);
  nand g140 (n_333, n_204, n_206);
  nand g141 (n_162, n_331, n_332, n_333);
  xor g142 (n_334, in_0[5], in_1[5]);
  xor g143 (n_208, n_334, in_3[5]);
  nand g144 (n_335, in_0[5], in_1[5]);
  nand g145 (n_336, in_3[5], in_1[5]);
  nand g146 (n_337, in_0[5], in_3[5]);
  nand g147 (n_211, n_335, n_336, n_337);
  xor g148 (n_338, in_4[5], in_2[5]);
  xor g149 (n_209, n_338, n_207);
  nand g150 (n_339, in_4[5], in_2[5]);
  nand g151 (n_340, n_207, in_2[5]);
  nand g152 (n_341, in_4[5], n_207);
  nand g153 (n_214, n_339, n_340, n_341);
  xor g154 (n_342, n_208, n_209);
  xor g155 (n_188, n_342, n_210);
  nand g156 (n_343, n_208, n_209);
  nand g157 (n_344, n_210, n_209);
  nand g158 (n_345, n_208, n_210);
  nand g159 (n_161, n_343, n_344, n_345);
  xor g160 (n_346, in_0[6], in_1[6]);
  xor g161 (n_212, n_346, in_3[6]);
  nand g162 (n_347, in_0[6], in_1[6]);
  nand g163 (n_348, in_3[6], in_1[6]);
  nand g164 (n_349, in_0[6], in_3[6]);
  nand g165 (n_215, n_347, n_348, n_349);
  xor g166 (n_350, in_4[6], in_2[6]);
  xor g167 (n_213, n_350, n_211);
  nand g168 (n_351, in_4[6], in_2[6]);
  nand g169 (n_352, n_211, in_2[6]);
  nand g170 (n_353, in_4[6], n_211);
  nand g171 (n_218, n_351, n_352, n_353);
  xor g172 (n_354, n_212, n_213);
  xor g173 (n_187, n_354, n_214);
  nand g174 (n_355, n_212, n_213);
  nand g175 (n_356, n_214, n_213);
  nand g176 (n_357, n_212, n_214);
  nand g177 (n_160, n_355, n_356, n_357);
  xor g178 (n_358, in_0[7], in_1[7]);
  xor g179 (n_216, n_358, in_3[7]);
  nand g180 (n_359, in_0[7], in_1[7]);
  nand g181 (n_360, in_3[7], in_1[7]);
  nand g182 (n_361, in_0[7], in_3[7]);
  nand g183 (n_219, n_359, n_360, n_361);
  xor g184 (n_362, in_4[7], in_2[7]);
  xor g185 (n_217, n_362, n_215);
  nand g186 (n_363, in_4[7], in_2[7]);
  nand g187 (n_364, n_215, in_2[7]);
  nand g188 (n_365, in_4[7], n_215);
  nand g189 (n_222, n_363, n_364, n_365);
  xor g190 (n_366, n_216, n_217);
  xor g191 (n_186, n_366, n_218);
  nand g192 (n_367, n_216, n_217);
  nand g193 (n_368, n_218, n_217);
  nand g194 (n_369, n_216, n_218);
  nand g195 (n_159, n_367, n_368, n_369);
  xor g196 (n_370, in_0[8], in_1[8]);
  xor g197 (n_220, n_370, in_3[8]);
  nand g198 (n_371, in_0[8], in_1[8]);
  nand g199 (n_372, in_3[8], in_1[8]);
  nand g200 (n_373, in_0[8], in_3[8]);
  nand g201 (n_223, n_371, n_372, n_373);
  xor g202 (n_374, in_4[8], in_2[8]);
  xor g203 (n_221, n_374, n_219);
  nand g204 (n_375, in_4[8], in_2[8]);
  nand g205 (n_376, n_219, in_2[8]);
  nand g206 (n_377, in_4[8], n_219);
  nand g207 (n_226, n_375, n_376, n_377);
  xor g208 (n_378, n_220, n_221);
  xor g209 (n_185, n_378, n_222);
  nand g210 (n_379, n_220, n_221);
  nand g211 (n_380, n_222, n_221);
  nand g212 (n_381, n_220, n_222);
  nand g213 (n_158, n_379, n_380, n_381);
  xor g214 (n_382, in_0[9], in_1[9]);
  xor g215 (n_224, n_382, in_3[9]);
  nand g216 (n_383, in_0[9], in_1[9]);
  nand g217 (n_384, in_3[9], in_1[9]);
  nand g218 (n_385, in_0[9], in_3[9]);
  nand g219 (n_227, n_383, n_384, n_385);
  xor g220 (n_386, in_4[9], in_2[9]);
  xor g221 (n_225, n_386, n_223);
  nand g222 (n_387, in_4[9], in_2[9]);
  nand g223 (n_388, n_223, in_2[9]);
  nand g224 (n_389, in_4[9], n_223);
  nand g225 (n_230, n_387, n_388, n_389);
  xor g226 (n_390, n_224, n_225);
  xor g227 (n_184, n_390, n_226);
  nand g228 (n_391, n_224, n_225);
  nand g229 (n_392, n_226, n_225);
  nand g230 (n_393, n_224, n_226);
  nand g231 (n_157, n_391, n_392, n_393);
  xor g232 (n_394, in_0[10], in_1[10]);
  xor g233 (n_228, n_394, in_3[10]);
  nand g234 (n_395, in_0[10], in_1[10]);
  nand g235 (n_396, in_3[10], in_1[10]);
  nand g236 (n_397, in_0[10], in_3[10]);
  nand g237 (n_231, n_395, n_396, n_397);
  xor g238 (n_398, in_4[10], in_2[10]);
  xor g239 (n_229, n_398, n_227);
  nand g240 (n_399, in_4[10], in_2[10]);
  nand g241 (n_400, n_227, in_2[10]);
  nand g242 (n_401, in_4[10], n_227);
  nand g243 (n_234, n_399, n_400, n_401);
  xor g244 (n_402, n_228, n_229);
  xor g245 (n_183, n_402, n_230);
  nand g246 (n_403, n_228, n_229);
  nand g247 (n_404, n_230, n_229);
  nand g248 (n_405, n_228, n_230);
  nand g249 (n_156, n_403, n_404, n_405);
  xor g250 (n_406, in_0[11], in_1[11]);
  xor g251 (n_232, n_406, in_3[11]);
  nand g252 (n_407, in_0[11], in_1[11]);
  nand g253 (n_408, in_3[11], in_1[11]);
  nand g254 (n_409, in_0[11], in_3[11]);
  nand g255 (n_235, n_407, n_408, n_409);
  xor g256 (n_410, in_4[11], in_2[11]);
  xor g257 (n_233, n_410, n_231);
  nand g258 (n_411, in_4[11], in_2[11]);
  nand g259 (n_412, n_231, in_2[11]);
  nand g260 (n_413, in_4[11], n_231);
  nand g261 (n_238, n_411, n_412, n_413);
  xor g262 (n_414, n_232, n_233);
  xor g263 (n_182, n_414, n_234);
  nand g264 (n_415, n_232, n_233);
  nand g265 (n_416, n_234, n_233);
  nand g266 (n_417, n_232, n_234);
  nand g267 (n_155, n_415, n_416, n_417);
  xor g268 (n_418, in_0[12], in_1[12]);
  xor g269 (n_236, n_418, in_3[12]);
  nand g270 (n_419, in_0[12], in_1[12]);
  nand g271 (n_420, in_3[12], in_1[12]);
  nand g272 (n_421, in_0[12], in_3[12]);
  nand g273 (n_239, n_419, n_420, n_421);
  xor g274 (n_422, in_4[12], in_2[12]);
  xor g275 (n_237, n_422, n_235);
  nand g276 (n_423, in_4[12], in_2[12]);
  nand g277 (n_424, n_235, in_2[12]);
  nand g278 (n_425, in_4[12], n_235);
  nand g279 (n_242, n_423, n_424, n_425);
  xor g280 (n_426, n_236, n_237);
  xor g281 (n_181, n_426, n_238);
  nand g282 (n_427, n_236, n_237);
  nand g283 (n_428, n_238, n_237);
  nand g284 (n_429, n_236, n_238);
  nand g285 (n_154, n_427, n_428, n_429);
  xor g286 (n_430, in_0[13], in_1[13]);
  xor g287 (n_240, n_430, in_3[13]);
  nand g288 (n_431, in_0[13], in_1[13]);
  nand g289 (n_432, in_3[13], in_1[13]);
  nand g290 (n_433, in_0[13], in_3[13]);
  nand g291 (n_243, n_431, n_432, n_433);
  xor g292 (n_434, in_4[13], in_2[13]);
  xor g293 (n_241, n_434, n_239);
  nand g294 (n_435, in_4[13], in_2[13]);
  nand g295 (n_436, n_239, in_2[13]);
  nand g296 (n_437, in_4[13], n_239);
  nand g297 (n_246, n_435, n_436, n_437);
  xor g298 (n_438, n_240, n_241);
  xor g299 (n_180, n_438, n_242);
  nand g300 (n_439, n_240, n_241);
  nand g301 (n_440, n_242, n_241);
  nand g302 (n_441, n_240, n_242);
  nand g303 (n_153, n_439, n_440, n_441);
  xor g304 (n_442, in_0[14], in_1[14]);
  xor g305 (n_244, n_442, in_3[14]);
  nand g306 (n_443, in_0[14], in_1[14]);
  nand g307 (n_444, in_3[14], in_1[14]);
  nand g308 (n_445, in_0[14], in_3[14]);
  nand g309 (n_247, n_443, n_444, n_445);
  xor g310 (n_446, in_4[14], in_2[14]);
  xor g311 (n_245, n_446, n_243);
  nand g312 (n_447, in_4[14], in_2[14]);
  nand g313 (n_448, n_243, in_2[14]);
  nand g314 (n_449, in_4[14], n_243);
  nand g315 (n_250, n_447, n_448, n_449);
  xor g316 (n_450, n_244, n_245);
  xor g317 (n_179, n_450, n_246);
  nand g318 (n_451, n_244, n_245);
  nand g319 (n_452, n_246, n_245);
  nand g320 (n_453, n_244, n_246);
  nand g321 (n_152, n_451, n_452, n_453);
  xor g322 (n_454, in_0[15], in_1[15]);
  xor g323 (n_248, n_454, in_3[15]);
  nand g324 (n_455, in_0[15], in_1[15]);
  nand g325 (n_456, in_3[15], in_1[15]);
  nand g326 (n_457, in_0[15], in_3[15]);
  nand g327 (n_251, n_455, n_456, n_457);
  xor g328 (n_458, in_4[15], in_2[15]);
  xor g329 (n_249, n_458, n_247);
  nand g330 (n_459, in_4[15], in_2[15]);
  nand g331 (n_460, n_247, in_2[15]);
  nand g332 (n_461, in_4[15], n_247);
  nand g333 (n_254, n_459, n_460, n_461);
  xor g334 (n_462, n_248, n_249);
  xor g335 (n_178, n_462, n_250);
  nand g336 (n_463, n_248, n_249);
  nand g337 (n_464, n_250, n_249);
  nand g338 (n_465, n_248, n_250);
  nand g339 (n_151, n_463, n_464, n_465);
  xor g340 (n_466, in_0[16], in_1[16]);
  xor g341 (n_252, n_466, in_3[16]);
  nand g342 (n_467, in_0[16], in_1[16]);
  nand g343 (n_468, in_3[16], in_1[16]);
  nand g344 (n_469, in_0[16], in_3[16]);
  nand g345 (n_255, n_467, n_468, n_469);
  xor g346 (n_470, in_4[16], in_2[16]);
  xor g347 (n_253, n_470, n_251);
  nand g348 (n_471, in_4[16], in_2[16]);
  nand g349 (n_472, n_251, in_2[16]);
  nand g350 (n_473, in_4[16], n_251);
  nand g351 (n_258, n_471, n_472, n_473);
  xor g352 (n_474, n_252, n_253);
  xor g353 (n_177, n_474, n_254);
  nand g354 (n_475, n_252, n_253);
  nand g355 (n_476, n_254, n_253);
  nand g356 (n_477, n_252, n_254);
  nand g357 (n_150, n_475, n_476, n_477);
  xor g358 (n_478, in_0[17], in_1[17]);
  xor g359 (n_256, n_478, in_3[17]);
  nand g360 (n_479, in_0[17], in_1[17]);
  nand g361 (n_480, in_3[17], in_1[17]);
  nand g362 (n_481, in_0[17], in_3[17]);
  nand g363 (n_259, n_479, n_480, n_481);
  xor g364 (n_482, in_4[17], in_2[17]);
  xor g365 (n_257, n_482, n_255);
  nand g366 (n_483, in_4[17], in_2[17]);
  nand g367 (n_484, n_255, in_2[17]);
  nand g368 (n_485, in_4[17], n_255);
  nand g369 (n_262, n_483, n_484, n_485);
  xor g370 (n_486, n_256, n_257);
  xor g371 (n_176, n_486, n_258);
  nand g372 (n_487, n_256, n_257);
  nand g373 (n_488, n_258, n_257);
  nand g374 (n_489, n_256, n_258);
  nand g375 (n_149, n_487, n_488, n_489);
  xor g376 (n_490, in_0[18], in_1[18]);
  xor g377 (n_260, n_490, in_3[18]);
  nand g378 (n_491, in_0[18], in_1[18]);
  nand g379 (n_492, in_3[18], in_1[18]);
  nand g380 (n_493, in_0[18], in_3[18]);
  nand g381 (n_263, n_491, n_492, n_493);
  xor g382 (n_494, in_4[18], in_2[18]);
  xor g383 (n_261, n_494, n_259);
  nand g384 (n_495, in_4[18], in_2[18]);
  nand g385 (n_496, n_259, in_2[18]);
  nand g386 (n_497, in_4[18], n_259);
  nand g387 (n_266, n_495, n_496, n_497);
  xor g388 (n_498, n_260, n_261);
  xor g389 (n_175, n_498, n_262);
  nand g390 (n_499, n_260, n_261);
  nand g391 (n_500, n_262, n_261);
  nand g392 (n_501, n_260, n_262);
  nand g393 (n_148, n_499, n_500, n_501);
  xor g394 (n_502, in_0[19], in_1[19]);
  xor g395 (n_264, n_502, in_3[19]);
  nand g396 (n_503, in_0[19], in_1[19]);
  nand g397 (n_504, in_3[19], in_1[19]);
  nand g398 (n_505, in_0[19], in_3[19]);
  nand g399 (n_267, n_503, n_504, n_505);
  xor g400 (n_506, in_4[19], in_2[19]);
  xor g401 (n_265, n_506, n_263);
  nand g402 (n_507, in_4[19], in_2[19]);
  nand g403 (n_508, n_263, in_2[19]);
  nand g404 (n_509, in_4[19], n_263);
  nand g405 (n_270, n_507, n_508, n_509);
  xor g406 (n_510, n_264, n_265);
  xor g407 (n_174, n_510, n_266);
  nand g408 (n_511, n_264, n_265);
  nand g409 (n_512, n_266, n_265);
  nand g410 (n_513, n_264, n_266);
  nand g411 (n_147, n_511, n_512, n_513);
  xor g412 (n_514, in_0[20], in_1[20]);
  xor g413 (n_268, n_514, in_3[20]);
  nand g414 (n_515, in_0[20], in_1[20]);
  nand g415 (n_516, in_3[20], in_1[20]);
  nand g416 (n_517, in_0[20], in_3[20]);
  nand g417 (n_271, n_515, n_516, n_517);
  xor g418 (n_518, in_4[20], in_2[20]);
  xor g419 (n_269, n_518, n_267);
  nand g420 (n_519, in_4[20], in_2[20]);
  nand g421 (n_520, n_267, in_2[20]);
  nand g422 (n_521, in_4[20], n_267);
  nand g423 (n_274, n_519, n_520, n_521);
  xor g424 (n_522, n_268, n_269);
  xor g425 (n_173, n_522, n_270);
  nand g426 (n_523, n_268, n_269);
  nand g427 (n_524, n_270, n_269);
  nand g428 (n_525, n_268, n_270);
  nand g429 (n_146, n_523, n_524, n_525);
  xor g430 (n_526, in_0[21], in_1[21]);
  xor g431 (n_272, n_526, in_3[21]);
  nand g432 (n_527, in_0[21], in_1[21]);
  nand g433 (n_528, in_3[21], in_1[21]);
  nand g434 (n_529, in_0[21], in_3[21]);
  nand g435 (n_281, n_527, n_528, n_529);
  xor g436 (n_530, in_4[21], in_2[21]);
  xor g437 (n_273, n_530, n_271);
  nand g438 (n_531, in_4[21], in_2[21]);
  nand g439 (n_532, n_271, in_2[21]);
  nand g440 (n_533, in_4[21], n_271);
  nand g441 (n_284, n_531, n_532, n_533);
  xor g442 (n_534, n_272, n_273);
  xor g443 (n_172, n_534, n_274);
  nand g444 (n_535, n_272, n_273);
  nand g445 (n_536, n_274, n_273);
  nand g446 (n_537, n_272, n_274);
  nand g447 (n_145, n_535, n_536, n_537);
  nand g455 (n_287, n_539, n_540, n_541);
  nand g459 (n_544, n_281, n_280);
  xor g462 (n_546, n_282, n_283);
  xor g463 (n_171, n_546, n_284);
  nand g464 (n_547, n_282, n_283);
  nand g465 (n_548, n_284, n_283);
  nand g466 (n_549, n_282, n_284);
  nand g467 (n_144, n_547, n_548, n_549);
  xor g471 (n_170, n_550, n_289);
  nand g474 (n_553, n_287, n_289);
  nand g475 (n_169, n_551, n_552, n_553);
  xor g478 (n_841, in_1[0], n_193);
  nand g479 (n_556, in_1[0], n_193);
  nand g480 (n_557, in_1[0], in_2[0]);
  nand g7 (n_558, n_193, in_2[0]);
  nand g8 (n_560, n_556, n_557, n_558);
  nor g9 (n_559, n_166, n_192);
  nand g10 (n_562, n_166, n_192);
  nor g11 (n_569, n_165, n_191);
  nand g12 (n_564, n_165, n_191);
  nor g13 (n_565, n_164, n_190);
  nand g14 (n_566, n_164, n_190);
  nor g15 (n_575, n_163, n_189);
  nand g16 (n_570, n_163, n_189);
  nor g17 (n_571, n_162, n_188);
  nand g18 (n_572, n_162, n_188);
  nor g19 (n_581, n_161, n_187);
  nand g20 (n_576, n_161, n_187);
  nor g21 (n_577, n_160, n_186);
  nand g22 (n_578, n_160, n_186);
  nor g23 (n_587, n_159, n_185);
  nand g24 (n_582, n_159, n_185);
  nor g25 (n_583, n_158, n_184);
  nand g26 (n_584, n_158, n_184);
  nor g27 (n_593, n_157, n_183);
  nand g28 (n_588, n_157, n_183);
  nor g29 (n_589, n_156, n_182);
  nand g30 (n_590, n_156, n_182);
  nor g31 (n_599, n_155, n_181);
  nand g32 (n_594, n_155, n_181);
  nor g33 (n_595, n_154, n_180);
  nand g34 (n_596, n_154, n_180);
  nor g35 (n_605, n_153, n_179);
  nand g36 (n_600, n_153, n_179);
  nor g37 (n_601, n_152, n_178);
  nand g38 (n_602, n_152, n_178);
  nor g39 (n_611, n_151, n_177);
  nand g40 (n_606, n_151, n_177);
  nor g41 (n_607, n_150, n_176);
  nand g42 (n_608, n_150, n_176);
  nor g43 (n_617, n_149, n_175);
  nand g44 (n_612, n_149, n_175);
  nor g45 (n_613, n_148, n_174);
  nand g46 (n_614, n_148, n_174);
  nor g47 (n_623, n_147, n_173);
  nand g48 (n_618, n_147, n_173);
  nor g49 (n_619, n_146, n_172);
  nand g50 (n_620, n_146, n_172);
  nor g51 (n_629, n_145, n_171);
  nand g52 (n_624, n_145, n_171);
  nor g53 (n_625, n_144, n_170);
  nand g54 (n_626, n_144, n_170);
  nor g55 (n_633, n_143, n_169);
  nand g56 (n_630, n_143, n_169);
  nand g61 (n_634, n_562, n_563);
  nor g62 (n_567, n_564, n_565);
  nor g65 (n_167, n_569, n_565);
  nor g66 (n_573, n_570, n_571);
  nor g69 (n_642, n_575, n_571);
  nor g70 (n_579, n_576, n_577);
  nor g73 (n_644, n_581, n_577);
  nor g74 (n_585, n_582, n_583);
  nor g483 (n_652, n_587, n_583);
  nor g484 (n_591, n_588, n_589);
  nor g487 (n_654, n_593, n_589);
  nor g488 (n_597, n_594, n_595);
  nor g491 (n_662, n_599, n_595);
  nor g492 (n_603, n_600, n_601);
  nor g495 (n_664, n_605, n_601);
  nor g496 (n_609, n_606, n_607);
  nor g499 (n_672, n_611, n_607);
  nor g500 (n_615, n_612, n_613);
  nor g503 (n_674, n_617, n_613);
  nor g504 (n_621, n_618, n_619);
  nor g507 (n_682, n_623, n_619);
  nor g508 (n_627, n_624, n_625);
  nor g511 (n_684, n_629, n_625);
  nand g514 (n_785, n_564, n_636);
  nand g515 (n_638, n_167, n_634);
  nand g516 (n_689, n_637, n_638);
  nor g517 (n_640, n_581, n_639);
  nand g526 (n_697, n_642, n_644);
  nor g527 (n_650, n_593, n_649);
  nand g536 (n_704, n_652, n_654);
  nor g537 (n_660, n_605, n_659);
  nand g546 (n_712, n_662, n_664);
  nor g547 (n_670, n_617, n_669);
  nand g556 (n_719, n_672, n_674);
  nor g557 (n_680, n_629, n_679);
  nand g566 (n_727, n_682, n_684);
  nand g569 (n_789, n_570, n_691);
  nand g570 (n_692, n_642, n_689);
  nand g571 (n_791, n_639, n_692);
  nand g574 (n_794, n_695, n_696);
  nand g577 (n_731, n_699, n_700);
  nor g578 (n_702, n_599, n_701);
  nor g581 (n_741, n_599, n_704);
  nor g587 (n_710, n_708, n_701);
  nor g590 (n_747, n_704, n_708);
  nor g591 (n_714, n_712, n_701);
  nor g594 (n_750, n_704, n_712);
  nor g595 (n_717, n_623, n_716);
  nor g598 (n_768, n_623, n_719);
  nor g604 (n_725, n_723, n_716);
  nor g607 (n_774, n_719, n_723);
  nor g608 (n_729, n_727, n_716);
  nor g611 (n_756, n_719, n_727);
  nand g614 (n_798, n_582, n_733);
  nand g615 (n_734, n_652, n_731);
  nand g616 (n_800, n_649, n_734);
  nand g619 (n_803, n_737, n_738);
  nand g622 (n_806, n_701, n_740);
  nand g623 (n_743, n_741, n_731);
  nand g624 (n_809, n_742, n_743);
  nand g625 (n_746, n_744, n_731);
  nand g626 (n_811, n_745, n_746);
  nand g627 (n_749, n_747, n_731);
  nand g628 (n_814, n_748, n_749);
  nand g629 (n_752, n_750, n_731);
  nand g630 (n_758, n_751, n_752);
  nor g631 (n_754, n_633, n_753);
  nand g638 (n_818, n_606, n_760);
  nand g639 (n_761, n_672, n_758);
  nand g640 (n_820, n_669, n_761);
  nand g643 (n_823, n_764, n_765);
  nand g646 (n_826, n_716, n_767);
  nand g647 (n_770, n_768, n_758);
  nand g648 (n_829, n_769, n_770);
  nand g649 (n_773, n_771, n_758);
  nand g650 (n_831, n_772, n_773);
  nand g651 (n_776, n_774, n_758);
  nand g652 (n_834, n_775, n_776);
  nand g653 (n_777, n_756, n_758);
  nand g654 (n_836, n_753, n_777);
  nand g657 (n_839, n_780, n_781);
  xnor g659 (out_0[1], n_560, n_782);
  xnor g661 (out_0[2], n_634, n_783);
  xnor g664 (out_0[3], n_785, n_786);
  xnor g666 (out_0[4], n_689, n_787);
  xnor g669 (out_0[5], n_789, n_790);
  xnor g671 (out_0[6], n_791, n_792);
  xnor g674 (out_0[7], n_794, n_795);
  xnor g676 (out_0[8], n_731, n_796);
  xnor g679 (out_0[9], n_798, n_799);
  xnor g681 (out_0[10], n_800, n_801);
  xnor g684 (out_0[11], n_803, n_804);
  xnor g687 (out_0[12], n_806, n_807);
  xnor g690 (out_0[13], n_809, n_810);
  xnor g692 (out_0[14], n_811, n_812);
  xnor g695 (out_0[15], n_814, n_815);
  xnor g697 (out_0[16], n_758, n_816);
  xnor g700 (out_0[17], n_818, n_819);
  xnor g702 (out_0[18], n_820, n_821);
  xnor g705 (out_0[19], n_823, n_824);
  xnor g708 (out_0[20], n_826, n_827);
  xnor g711 (out_0[21], n_829, n_830);
  xnor g713 (out_0[22], n_831, n_832);
  xnor g716 (out_0[23], n_834, n_835);
  xnor g718 (out_0[24], n_836, n_837);
  xor g722 (out_0[0], in_2[0], n_841);
  xor g723 (n_280, in_0[22], in_1[22]);
  nor g724 (n_143, in_0[22], in_1[22]);
  xor g725 (n_538, in_3[22], in_4[22]);
  or g726 (n_539, in_3[22], in_4[22]);
  or g727 (n_540, in_2[22], in_4[22]);
  or g728 (n_541, in_2[22], in_3[22]);
  xnor g729 (n_282, n_538, in_2[22]);
  xnor g733 (n_283, n_281, n_280);
  or g734 (n_289, n_280, wc, n_281);
  not gc (wc, n_544);
  xnor g735 (n_550, n_287, n_143);
  or g736 (n_551, n_143, wc0);
  not gc0 (wc0, n_287);
  or g737 (n_552, wc1, n_143);
  not gc1 (wc1, n_289);
  or g738 (n_563, n_559, wc2);
  not gc2 (wc2, n_560);
  or g739 (n_782, wc3, n_559);
  not gc3 (wc3, n_562);
  and g740 (n_637, wc4, n_566);
  not gc4 (wc4, n_567);
  or g741 (n_783, wc5, n_569);
  not gc5 (wc5, n_564);
  or g742 (n_786, wc6, n_565);
  not gc6 (wc6, n_566);
  and g743 (n_639, wc7, n_572);
  not gc7 (wc7, n_573);
  or g744 (n_636, wc8, n_569);
  not gc8 (wc8, n_634);
  or g745 (n_787, wc9, n_575);
  not gc9 (wc9, n_570);
  or g746 (n_790, wc10, n_571);
  not gc10 (wc10, n_572);
  and g747 (n_646, wc11, n_578);
  not gc11 (wc11, n_579);
  and g748 (n_649, wc12, n_584);
  not gc12 (wc12, n_585);
  and g749 (n_656, wc13, n_590);
  not gc13 (wc13, n_591);
  and g750 (n_659, wc14, n_596);
  not gc14 (wc14, n_597);
  and g751 (n_666, wc15, n_602);
  not gc15 (wc15, n_603);
  and g752 (n_669, wc16, n_608);
  not gc16 (wc16, n_609);
  and g753 (n_676, wc17, n_614);
  not gc17 (wc17, n_615);
  and g754 (n_679, wc18, n_620);
  not gc18 (wc18, n_621);
  and g755 (n_686, wc19, n_626);
  not gc19 (wc19, n_627);
  or g756 (n_693, wc20, n_581);
  not gc20 (wc20, n_642);
  or g757 (n_735, wc21, n_593);
  not gc21 (wc21, n_652);
  or g758 (n_708, wc22, n_605);
  not gc22 (wc22, n_662);
  or g759 (n_762, wc23, n_617);
  not gc23 (wc23, n_672);
  or g760 (n_723, wc24, n_629);
  not gc24 (wc24, n_682);
  or g761 (n_792, wc25, n_581);
  not gc25 (wc25, n_576);
  or g762 (n_795, wc26, n_577);
  not gc26 (wc26, n_578);
  or g763 (n_796, wc27, n_587);
  not gc27 (wc27, n_582);
  or g764 (n_799, wc28, n_583);
  not gc28 (wc28, n_584);
  or g765 (n_801, wc29, n_593);
  not gc29 (wc29, n_588);
  or g766 (n_804, wc30, n_589);
  not gc30 (wc30, n_590);
  or g767 (n_807, wc31, n_599);
  not gc31 (wc31, n_594);
  or g768 (n_810, wc32, n_595);
  not gc32 (wc32, n_596);
  or g769 (n_812, wc33, n_605);
  not gc33 (wc33, n_600);
  or g770 (n_815, wc34, n_601);
  not gc34 (wc34, n_602);
  or g771 (n_816, wc35, n_611);
  not gc35 (wc35, n_606);
  or g772 (n_819, wc36, n_607);
  not gc36 (wc36, n_608);
  or g773 (n_821, wc37, n_617);
  not gc37 (wc37, n_612);
  or g774 (n_824, wc38, n_613);
  not gc38 (wc38, n_614);
  or g775 (n_827, wc39, n_623);
  not gc39 (wc39, n_618);
  or g776 (n_830, wc40, n_619);
  not gc40 (wc40, n_620);
  or g777 (n_832, wc41, n_629);
  not gc41 (wc41, n_624);
  or g778 (n_835, wc42, n_625);
  not gc42 (wc42, n_626);
  or g779 (n_837, wc43, n_633);
  not gc43 (wc43, n_630);
  and g780 (n_695, wc44, n_576);
  not gc44 (wc44, n_640);
  and g781 (n_647, wc45, n_644);
  not gc45 (wc45, n_639);
  and g782 (n_657, wc46, n_654);
  not gc46 (wc46, n_649);
  and g783 (n_667, wc47, n_664);
  not gc47 (wc47, n_659);
  and g784 (n_677, wc48, n_674);
  not gc48 (wc48, n_669);
  and g785 (n_687, wc49, n_684);
  not gc49 (wc49, n_679);
  or g786 (n_691, wc50, n_575);
  not gc50 (wc50, n_689);
  and g787 (n_744, wc51, n_662);
  not gc51 (wc51, n_704);
  and g788 (n_771, wc52, n_682);
  not gc52 (wc52, n_719);
  and g789 (n_699, wc53, n_646);
  not gc53 (wc53, n_647);
  and g790 (n_737, wc54, n_588);
  not gc54 (wc54, n_650);
  and g791 (n_701, wc55, n_656);
  not gc55 (wc55, n_657);
  and g792 (n_709, wc56, n_600);
  not gc56 (wc56, n_660);
  and g793 (n_713, wc57, n_666);
  not gc57 (wc57, n_667);
  and g794 (n_764, wc58, n_612);
  not gc58 (wc58, n_670);
  and g795 (n_716, wc59, n_676);
  not gc59 (wc59, n_677);
  and g796 (n_724, wc60, n_624);
  not gc60 (wc60, n_680);
  and g797 (n_728, wc61, n_686);
  not gc61 (wc61, n_687);
  or g798 (n_696, n_693, wc62);
  not gc62 (wc62, n_689);
  or g799 (n_700, n_697, wc63);
  not gc63 (wc63, n_689);
  or g800 (n_778, wc64, n_633);
  not gc64 (wc64, n_756);
  and g801 (n_706, wc65, n_662);
  not gc65 (wc65, n_701);
  and g802 (n_721, wc66, n_682);
  not gc66 (wc66, n_716);
  and g803 (n_742, wc67, n_594);
  not gc67 (wc67, n_702);
  and g804 (n_745, wc68, n_659);
  not gc68 (wc68, n_706);
  and g805 (n_748, n_709, wc69);
  not gc69 (wc69, n_710);
  and g806 (n_751, n_713, wc70);
  not gc70 (wc70, n_714);
  and g807 (n_769, wc71, n_618);
  not gc71 (wc71, n_717);
  and g808 (n_772, wc72, n_679);
  not gc72 (wc72, n_721);
  and g809 (n_775, n_724, wc73);
  not gc73 (wc73, n_725);
  and g810 (n_753, n_728, wc74);
  not gc74 (wc74, n_729);
  or g811 (n_733, wc75, n_587);
  not gc75 (wc75, n_731);
  or g812 (n_738, n_735, wc76);
  not gc76 (wc76, n_731);
  or g813 (n_740, wc77, n_704);
  not gc77 (wc77, n_731);
  and g814 (n_780, wc78, n_630);
  not gc78 (wc78, n_754);
  or g815 (n_760, wc79, n_611);
  not gc79 (wc79, n_758);
  or g816 (n_765, n_762, wc80);
  not gc80 (wc80, n_758);
  or g817 (n_767, wc81, n_719);
  not gc81 (wc81, n_758);
  or g818 (n_781, n_778, wc82);
  not gc82 (wc82, n_758);
  not g819 (out_0[25], n_839);
endmodule

module csa_tree_add_749_44_group_6809_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  csa_tree_add_749_44_group_6809_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_823_44_group_6807_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_280, n_281, n_282, n_283, n_284, n_287;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_544, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_556, n_557;
  wire n_558, n_559, n_560, n_562, n_563, n_564, n_565, n_566;
  wire n_567, n_569, n_570, n_571, n_572, n_573, n_575, n_576;
  wire n_577, n_578, n_579, n_581, n_582, n_583, n_584, n_585;
  wire n_587, n_588, n_589, n_590, n_591, n_593, n_594, n_595;
  wire n_596, n_597, n_599, n_600, n_601, n_602, n_603, n_605;
  wire n_606, n_607, n_608, n_609, n_611, n_612, n_613, n_614;
  wire n_615, n_617, n_618, n_619, n_620, n_621, n_623, n_624;
  wire n_625, n_626, n_627, n_629, n_630, n_633, n_634, n_636;
  wire n_637, n_638, n_639, n_640, n_642, n_644, n_646, n_647;
  wire n_649, n_650, n_652, n_654, n_656, n_657, n_659, n_660;
  wire n_662, n_664, n_666, n_667, n_669, n_670, n_672, n_674;
  wire n_676, n_677, n_679, n_680, n_682, n_684, n_686, n_687;
  wire n_689, n_691, n_692, n_693, n_695, n_696, n_697, n_699;
  wire n_700, n_701, n_702, n_704, n_706, n_708, n_709, n_710;
  wire n_712, n_713, n_714, n_716, n_717, n_719, n_721, n_723;
  wire n_724, n_725, n_727, n_728, n_729, n_731, n_733, n_734;
  wire n_735, n_737, n_738, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_756, n_758, n_760, n_761, n_762, n_764;
  wire n_765, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_780, n_781, n_782;
  wire n_783, n_785, n_786, n_787, n_789, n_790, n_791, n_792;
  wire n_794, n_795, n_796, n_798, n_799, n_800, n_801, n_803;
  wire n_804, n_806, n_807, n_809, n_810, n_811, n_812, n_814;
  wire n_815, n_816, n_818, n_819, n_820, n_821, n_823, n_824;
  wire n_826, n_827, n_829, n_830, n_831, n_832, n_834, n_835;
  wire n_836, n_837, n_839, n_841;
  xor g75 (n_290, in_0[0], in_4[0]);
  xor g76 (n_193, n_290, in_3[0]);
  nand g77 (n_291, in_0[0], in_4[0]);
  nand g78 (n_292, in_3[0], in_4[0]);
  nand g79 (n_293, in_0[0], in_3[0]);
  nand g6 (n_195, n_291, n_292, n_293);
  xor g80 (n_294, in_0[1], in_1[1]);
  xor g81 (n_166, n_294, in_4[1]);
  nand g82 (n_295, in_0[1], in_1[1]);
  nand g83 (n_296, in_4[1], in_1[1]);
  nand g84 (n_297, in_0[1], in_4[1]);
  nand g85 (n_197, n_295, n_296, n_297);
  xor g86 (n_298, in_3[1], in_2[1]);
  xor g87 (n_192, n_298, n_195);
  nand g88 (n_299, in_3[1], in_2[1]);
  nand g89 (n_300, n_195, in_2[1]);
  nand g90 (n_301, in_3[1], n_195);
  nand g91 (n_165, n_299, n_300, n_301);
  xor g92 (n_196, in_0[2], in_1[2]);
  and g93 (n_199, in_0[2], in_1[2]);
  xor g94 (n_302, in_3[2], in_4[2]);
  xor g95 (n_198, n_302, in_2[2]);
  nand g96 (n_303, in_3[2], in_4[2]);
  nand g97 (n_304, in_2[2], in_4[2]);
  nand g98 (n_305, in_3[2], in_2[2]);
  nand g99 (n_200, n_303, n_304, n_305);
  xor g100 (n_306, n_196, n_197);
  xor g101 (n_191, n_306, n_198);
  nand g102 (n_307, n_196, n_197);
  nand g103 (n_308, n_198, n_197);
  nand g104 (n_309, n_196, n_198);
  nand g105 (n_164, n_307, n_308, n_309);
  xor g106 (n_310, in_0[3], in_1[3]);
  xor g107 (n_201, n_310, in_3[3]);
  nand g108 (n_311, in_0[3], in_1[3]);
  nand g109 (n_312, in_3[3], in_1[3]);
  nand g110 (n_313, in_0[3], in_3[3]);
  nand g111 (n_203, n_311, n_312, n_313);
  xor g112 (n_314, in_4[3], in_2[3]);
  xor g113 (n_202, n_314, n_199);
  nand g114 (n_315, in_4[3], in_2[3]);
  nand g115 (n_316, n_199, in_2[3]);
  nand g116 (n_317, in_4[3], n_199);
  nand g117 (n_205, n_315, n_316, n_317);
  xor g118 (n_318, n_200, n_201);
  xor g119 (n_190, n_318, n_202);
  nand g120 (n_319, n_200, n_201);
  nand g121 (n_320, n_202, n_201);
  nand g122 (n_321, n_200, n_202);
  nand g123 (n_163, n_319, n_320, n_321);
  xor g124 (n_322, in_0[4], in_1[4]);
  xor g125 (n_204, n_322, in_3[4]);
  nand g126 (n_323, in_0[4], in_1[4]);
  nand g127 (n_324, in_3[4], in_1[4]);
  nand g128 (n_325, in_0[4], in_3[4]);
  nand g129 (n_207, n_323, n_324, n_325);
  xor g130 (n_326, in_4[4], in_2[4]);
  xor g131 (n_206, n_326, n_203);
  nand g132 (n_327, in_4[4], in_2[4]);
  nand g133 (n_328, n_203, in_2[4]);
  nand g134 (n_329, in_4[4], n_203);
  nand g135 (n_210, n_327, n_328, n_329);
  xor g136 (n_330, n_204, n_205);
  xor g137 (n_189, n_330, n_206);
  nand g138 (n_331, n_204, n_205);
  nand g139 (n_332, n_206, n_205);
  nand g140 (n_333, n_204, n_206);
  nand g141 (n_162, n_331, n_332, n_333);
  xor g142 (n_334, in_0[5], in_1[5]);
  xor g143 (n_208, n_334, in_3[5]);
  nand g144 (n_335, in_0[5], in_1[5]);
  nand g145 (n_336, in_3[5], in_1[5]);
  nand g146 (n_337, in_0[5], in_3[5]);
  nand g147 (n_211, n_335, n_336, n_337);
  xor g148 (n_338, in_4[5], in_2[5]);
  xor g149 (n_209, n_338, n_207);
  nand g150 (n_339, in_4[5], in_2[5]);
  nand g151 (n_340, n_207, in_2[5]);
  nand g152 (n_341, in_4[5], n_207);
  nand g153 (n_214, n_339, n_340, n_341);
  xor g154 (n_342, n_208, n_209);
  xor g155 (n_188, n_342, n_210);
  nand g156 (n_343, n_208, n_209);
  nand g157 (n_344, n_210, n_209);
  nand g158 (n_345, n_208, n_210);
  nand g159 (n_161, n_343, n_344, n_345);
  xor g160 (n_346, in_0[6], in_1[6]);
  xor g161 (n_212, n_346, in_3[6]);
  nand g162 (n_347, in_0[6], in_1[6]);
  nand g163 (n_348, in_3[6], in_1[6]);
  nand g164 (n_349, in_0[6], in_3[6]);
  nand g165 (n_215, n_347, n_348, n_349);
  xor g166 (n_350, in_4[6], in_2[6]);
  xor g167 (n_213, n_350, n_211);
  nand g168 (n_351, in_4[6], in_2[6]);
  nand g169 (n_352, n_211, in_2[6]);
  nand g170 (n_353, in_4[6], n_211);
  nand g171 (n_218, n_351, n_352, n_353);
  xor g172 (n_354, n_212, n_213);
  xor g173 (n_187, n_354, n_214);
  nand g174 (n_355, n_212, n_213);
  nand g175 (n_356, n_214, n_213);
  nand g176 (n_357, n_212, n_214);
  nand g177 (n_160, n_355, n_356, n_357);
  xor g178 (n_358, in_0[7], in_1[7]);
  xor g179 (n_216, n_358, in_3[7]);
  nand g180 (n_359, in_0[7], in_1[7]);
  nand g181 (n_360, in_3[7], in_1[7]);
  nand g182 (n_361, in_0[7], in_3[7]);
  nand g183 (n_219, n_359, n_360, n_361);
  xor g184 (n_362, in_4[7], in_2[7]);
  xor g185 (n_217, n_362, n_215);
  nand g186 (n_363, in_4[7], in_2[7]);
  nand g187 (n_364, n_215, in_2[7]);
  nand g188 (n_365, in_4[7], n_215);
  nand g189 (n_222, n_363, n_364, n_365);
  xor g190 (n_366, n_216, n_217);
  xor g191 (n_186, n_366, n_218);
  nand g192 (n_367, n_216, n_217);
  nand g193 (n_368, n_218, n_217);
  nand g194 (n_369, n_216, n_218);
  nand g195 (n_159, n_367, n_368, n_369);
  xor g196 (n_370, in_0[8], in_1[8]);
  xor g197 (n_220, n_370, in_3[8]);
  nand g198 (n_371, in_0[8], in_1[8]);
  nand g199 (n_372, in_3[8], in_1[8]);
  nand g200 (n_373, in_0[8], in_3[8]);
  nand g201 (n_223, n_371, n_372, n_373);
  xor g202 (n_374, in_4[8], in_2[8]);
  xor g203 (n_221, n_374, n_219);
  nand g204 (n_375, in_4[8], in_2[8]);
  nand g205 (n_376, n_219, in_2[8]);
  nand g206 (n_377, in_4[8], n_219);
  nand g207 (n_226, n_375, n_376, n_377);
  xor g208 (n_378, n_220, n_221);
  xor g209 (n_185, n_378, n_222);
  nand g210 (n_379, n_220, n_221);
  nand g211 (n_380, n_222, n_221);
  nand g212 (n_381, n_220, n_222);
  nand g213 (n_158, n_379, n_380, n_381);
  xor g214 (n_382, in_0[9], in_1[9]);
  xor g215 (n_224, n_382, in_3[9]);
  nand g216 (n_383, in_0[9], in_1[9]);
  nand g217 (n_384, in_3[9], in_1[9]);
  nand g218 (n_385, in_0[9], in_3[9]);
  nand g219 (n_227, n_383, n_384, n_385);
  xor g220 (n_386, in_4[9], in_2[9]);
  xor g221 (n_225, n_386, n_223);
  nand g222 (n_387, in_4[9], in_2[9]);
  nand g223 (n_388, n_223, in_2[9]);
  nand g224 (n_389, in_4[9], n_223);
  nand g225 (n_230, n_387, n_388, n_389);
  xor g226 (n_390, n_224, n_225);
  xor g227 (n_184, n_390, n_226);
  nand g228 (n_391, n_224, n_225);
  nand g229 (n_392, n_226, n_225);
  nand g230 (n_393, n_224, n_226);
  nand g231 (n_157, n_391, n_392, n_393);
  xor g232 (n_394, in_0[10], in_1[10]);
  xor g233 (n_228, n_394, in_3[10]);
  nand g234 (n_395, in_0[10], in_1[10]);
  nand g235 (n_396, in_3[10], in_1[10]);
  nand g236 (n_397, in_0[10], in_3[10]);
  nand g237 (n_231, n_395, n_396, n_397);
  xor g238 (n_398, in_4[10], in_2[10]);
  xor g239 (n_229, n_398, n_227);
  nand g240 (n_399, in_4[10], in_2[10]);
  nand g241 (n_400, n_227, in_2[10]);
  nand g242 (n_401, in_4[10], n_227);
  nand g243 (n_234, n_399, n_400, n_401);
  xor g244 (n_402, n_228, n_229);
  xor g245 (n_183, n_402, n_230);
  nand g246 (n_403, n_228, n_229);
  nand g247 (n_404, n_230, n_229);
  nand g248 (n_405, n_228, n_230);
  nand g249 (n_156, n_403, n_404, n_405);
  xor g250 (n_406, in_0[11], in_1[11]);
  xor g251 (n_232, n_406, in_3[11]);
  nand g252 (n_407, in_0[11], in_1[11]);
  nand g253 (n_408, in_3[11], in_1[11]);
  nand g254 (n_409, in_0[11], in_3[11]);
  nand g255 (n_235, n_407, n_408, n_409);
  xor g256 (n_410, in_4[11], in_2[11]);
  xor g257 (n_233, n_410, n_231);
  nand g258 (n_411, in_4[11], in_2[11]);
  nand g259 (n_412, n_231, in_2[11]);
  nand g260 (n_413, in_4[11], n_231);
  nand g261 (n_238, n_411, n_412, n_413);
  xor g262 (n_414, n_232, n_233);
  xor g263 (n_182, n_414, n_234);
  nand g264 (n_415, n_232, n_233);
  nand g265 (n_416, n_234, n_233);
  nand g266 (n_417, n_232, n_234);
  nand g267 (n_155, n_415, n_416, n_417);
  xor g268 (n_418, in_0[12], in_1[12]);
  xor g269 (n_236, n_418, in_3[12]);
  nand g270 (n_419, in_0[12], in_1[12]);
  nand g271 (n_420, in_3[12], in_1[12]);
  nand g272 (n_421, in_0[12], in_3[12]);
  nand g273 (n_239, n_419, n_420, n_421);
  xor g274 (n_422, in_4[12], in_2[12]);
  xor g275 (n_237, n_422, n_235);
  nand g276 (n_423, in_4[12], in_2[12]);
  nand g277 (n_424, n_235, in_2[12]);
  nand g278 (n_425, in_4[12], n_235);
  nand g279 (n_242, n_423, n_424, n_425);
  xor g280 (n_426, n_236, n_237);
  xor g281 (n_181, n_426, n_238);
  nand g282 (n_427, n_236, n_237);
  nand g283 (n_428, n_238, n_237);
  nand g284 (n_429, n_236, n_238);
  nand g285 (n_154, n_427, n_428, n_429);
  xor g286 (n_430, in_0[13], in_1[13]);
  xor g287 (n_240, n_430, in_3[13]);
  nand g288 (n_431, in_0[13], in_1[13]);
  nand g289 (n_432, in_3[13], in_1[13]);
  nand g290 (n_433, in_0[13], in_3[13]);
  nand g291 (n_243, n_431, n_432, n_433);
  xor g292 (n_434, in_4[13], in_2[13]);
  xor g293 (n_241, n_434, n_239);
  nand g294 (n_435, in_4[13], in_2[13]);
  nand g295 (n_436, n_239, in_2[13]);
  nand g296 (n_437, in_4[13], n_239);
  nand g297 (n_246, n_435, n_436, n_437);
  xor g298 (n_438, n_240, n_241);
  xor g299 (n_180, n_438, n_242);
  nand g300 (n_439, n_240, n_241);
  nand g301 (n_440, n_242, n_241);
  nand g302 (n_441, n_240, n_242);
  nand g303 (n_153, n_439, n_440, n_441);
  xor g304 (n_442, in_0[14], in_1[14]);
  xor g305 (n_244, n_442, in_3[14]);
  nand g306 (n_443, in_0[14], in_1[14]);
  nand g307 (n_444, in_3[14], in_1[14]);
  nand g308 (n_445, in_0[14], in_3[14]);
  nand g309 (n_247, n_443, n_444, n_445);
  xor g310 (n_446, in_4[14], in_2[14]);
  xor g311 (n_245, n_446, n_243);
  nand g312 (n_447, in_4[14], in_2[14]);
  nand g313 (n_448, n_243, in_2[14]);
  nand g314 (n_449, in_4[14], n_243);
  nand g315 (n_250, n_447, n_448, n_449);
  xor g316 (n_450, n_244, n_245);
  xor g317 (n_179, n_450, n_246);
  nand g318 (n_451, n_244, n_245);
  nand g319 (n_452, n_246, n_245);
  nand g320 (n_453, n_244, n_246);
  nand g321 (n_152, n_451, n_452, n_453);
  xor g322 (n_454, in_0[15], in_1[15]);
  xor g323 (n_248, n_454, in_3[15]);
  nand g324 (n_455, in_0[15], in_1[15]);
  nand g325 (n_456, in_3[15], in_1[15]);
  nand g326 (n_457, in_0[15], in_3[15]);
  nand g327 (n_251, n_455, n_456, n_457);
  xor g328 (n_458, in_4[15], in_2[15]);
  xor g329 (n_249, n_458, n_247);
  nand g330 (n_459, in_4[15], in_2[15]);
  nand g331 (n_460, n_247, in_2[15]);
  nand g332 (n_461, in_4[15], n_247);
  nand g333 (n_254, n_459, n_460, n_461);
  xor g334 (n_462, n_248, n_249);
  xor g335 (n_178, n_462, n_250);
  nand g336 (n_463, n_248, n_249);
  nand g337 (n_464, n_250, n_249);
  nand g338 (n_465, n_248, n_250);
  nand g339 (n_151, n_463, n_464, n_465);
  xor g340 (n_466, in_0[16], in_1[16]);
  xor g341 (n_252, n_466, in_3[16]);
  nand g342 (n_467, in_0[16], in_1[16]);
  nand g343 (n_468, in_3[16], in_1[16]);
  nand g344 (n_469, in_0[16], in_3[16]);
  nand g345 (n_255, n_467, n_468, n_469);
  xor g346 (n_470, in_4[16], in_2[16]);
  xor g347 (n_253, n_470, n_251);
  nand g348 (n_471, in_4[16], in_2[16]);
  nand g349 (n_472, n_251, in_2[16]);
  nand g350 (n_473, in_4[16], n_251);
  nand g351 (n_258, n_471, n_472, n_473);
  xor g352 (n_474, n_252, n_253);
  xor g353 (n_177, n_474, n_254);
  nand g354 (n_475, n_252, n_253);
  nand g355 (n_476, n_254, n_253);
  nand g356 (n_477, n_252, n_254);
  nand g357 (n_150, n_475, n_476, n_477);
  xor g358 (n_478, in_0[17], in_1[17]);
  xor g359 (n_256, n_478, in_3[17]);
  nand g360 (n_479, in_0[17], in_1[17]);
  nand g361 (n_480, in_3[17], in_1[17]);
  nand g362 (n_481, in_0[17], in_3[17]);
  nand g363 (n_259, n_479, n_480, n_481);
  xor g364 (n_482, in_4[17], in_2[17]);
  xor g365 (n_257, n_482, n_255);
  nand g366 (n_483, in_4[17], in_2[17]);
  nand g367 (n_484, n_255, in_2[17]);
  nand g368 (n_485, in_4[17], n_255);
  nand g369 (n_262, n_483, n_484, n_485);
  xor g370 (n_486, n_256, n_257);
  xor g371 (n_176, n_486, n_258);
  nand g372 (n_487, n_256, n_257);
  nand g373 (n_488, n_258, n_257);
  nand g374 (n_489, n_256, n_258);
  nand g375 (n_149, n_487, n_488, n_489);
  xor g376 (n_490, in_0[18], in_1[18]);
  xor g377 (n_260, n_490, in_3[18]);
  nand g378 (n_491, in_0[18], in_1[18]);
  nand g379 (n_492, in_3[18], in_1[18]);
  nand g380 (n_493, in_0[18], in_3[18]);
  nand g381 (n_263, n_491, n_492, n_493);
  xor g382 (n_494, in_4[18], in_2[18]);
  xor g383 (n_261, n_494, n_259);
  nand g384 (n_495, in_4[18], in_2[18]);
  nand g385 (n_496, n_259, in_2[18]);
  nand g386 (n_497, in_4[18], n_259);
  nand g387 (n_266, n_495, n_496, n_497);
  xor g388 (n_498, n_260, n_261);
  xor g389 (n_175, n_498, n_262);
  nand g390 (n_499, n_260, n_261);
  nand g391 (n_500, n_262, n_261);
  nand g392 (n_501, n_260, n_262);
  nand g393 (n_148, n_499, n_500, n_501);
  xor g394 (n_502, in_0[19], in_1[19]);
  xor g395 (n_264, n_502, in_3[19]);
  nand g396 (n_503, in_0[19], in_1[19]);
  nand g397 (n_504, in_3[19], in_1[19]);
  nand g398 (n_505, in_0[19], in_3[19]);
  nand g399 (n_267, n_503, n_504, n_505);
  xor g400 (n_506, in_4[19], in_2[19]);
  xor g401 (n_265, n_506, n_263);
  nand g402 (n_507, in_4[19], in_2[19]);
  nand g403 (n_508, n_263, in_2[19]);
  nand g404 (n_509, in_4[19], n_263);
  nand g405 (n_270, n_507, n_508, n_509);
  xor g406 (n_510, n_264, n_265);
  xor g407 (n_174, n_510, n_266);
  nand g408 (n_511, n_264, n_265);
  nand g409 (n_512, n_266, n_265);
  nand g410 (n_513, n_264, n_266);
  nand g411 (n_147, n_511, n_512, n_513);
  xor g412 (n_514, in_0[20], in_1[20]);
  xor g413 (n_268, n_514, in_3[20]);
  nand g414 (n_515, in_0[20], in_1[20]);
  nand g415 (n_516, in_3[20], in_1[20]);
  nand g416 (n_517, in_0[20], in_3[20]);
  nand g417 (n_271, n_515, n_516, n_517);
  xor g418 (n_518, in_4[20], in_2[20]);
  xor g419 (n_269, n_518, n_267);
  nand g420 (n_519, in_4[20], in_2[20]);
  nand g421 (n_520, n_267, in_2[20]);
  nand g422 (n_521, in_4[20], n_267);
  nand g423 (n_274, n_519, n_520, n_521);
  xor g424 (n_522, n_268, n_269);
  xor g425 (n_173, n_522, n_270);
  nand g426 (n_523, n_268, n_269);
  nand g427 (n_524, n_270, n_269);
  nand g428 (n_525, n_268, n_270);
  nand g429 (n_146, n_523, n_524, n_525);
  xor g430 (n_526, in_0[21], in_1[21]);
  xor g431 (n_272, n_526, in_3[21]);
  nand g432 (n_527, in_0[21], in_1[21]);
  nand g433 (n_528, in_3[21], in_1[21]);
  nand g434 (n_529, in_0[21], in_3[21]);
  nand g435 (n_281, n_527, n_528, n_529);
  xor g436 (n_530, in_4[21], in_2[21]);
  xor g437 (n_273, n_530, n_271);
  nand g438 (n_531, in_4[21], in_2[21]);
  nand g439 (n_532, n_271, in_2[21]);
  nand g440 (n_533, in_4[21], n_271);
  nand g441 (n_284, n_531, n_532, n_533);
  xor g442 (n_534, n_272, n_273);
  xor g443 (n_172, n_534, n_274);
  nand g444 (n_535, n_272, n_273);
  nand g445 (n_536, n_274, n_273);
  nand g446 (n_537, n_272, n_274);
  nand g447 (n_145, n_535, n_536, n_537);
  nand g455 (n_287, n_539, n_540, n_541);
  nand g459 (n_544, n_281, n_280);
  xor g462 (n_546, n_282, n_283);
  xor g463 (n_171, n_546, n_284);
  nand g464 (n_547, n_282, n_283);
  nand g465 (n_548, n_284, n_283);
  nand g466 (n_549, n_282, n_284);
  nand g467 (n_144, n_547, n_548, n_549);
  xor g471 (n_170, n_550, n_289);
  nand g474 (n_553, n_287, n_289);
  nand g475 (n_169, n_551, n_552, n_553);
  xor g478 (n_841, in_1[0], n_193);
  nand g479 (n_556, in_1[0], n_193);
  nand g480 (n_557, in_1[0], in_2[0]);
  nand g7 (n_558, n_193, in_2[0]);
  nand g8 (n_560, n_556, n_557, n_558);
  nor g9 (n_559, n_166, n_192);
  nand g10 (n_562, n_166, n_192);
  nor g11 (n_569, n_165, n_191);
  nand g12 (n_564, n_165, n_191);
  nor g13 (n_565, n_164, n_190);
  nand g14 (n_566, n_164, n_190);
  nor g15 (n_575, n_163, n_189);
  nand g16 (n_570, n_163, n_189);
  nor g17 (n_571, n_162, n_188);
  nand g18 (n_572, n_162, n_188);
  nor g19 (n_581, n_161, n_187);
  nand g20 (n_576, n_161, n_187);
  nor g21 (n_577, n_160, n_186);
  nand g22 (n_578, n_160, n_186);
  nor g23 (n_587, n_159, n_185);
  nand g24 (n_582, n_159, n_185);
  nor g25 (n_583, n_158, n_184);
  nand g26 (n_584, n_158, n_184);
  nor g27 (n_593, n_157, n_183);
  nand g28 (n_588, n_157, n_183);
  nor g29 (n_589, n_156, n_182);
  nand g30 (n_590, n_156, n_182);
  nor g31 (n_599, n_155, n_181);
  nand g32 (n_594, n_155, n_181);
  nor g33 (n_595, n_154, n_180);
  nand g34 (n_596, n_154, n_180);
  nor g35 (n_605, n_153, n_179);
  nand g36 (n_600, n_153, n_179);
  nor g37 (n_601, n_152, n_178);
  nand g38 (n_602, n_152, n_178);
  nor g39 (n_611, n_151, n_177);
  nand g40 (n_606, n_151, n_177);
  nor g41 (n_607, n_150, n_176);
  nand g42 (n_608, n_150, n_176);
  nor g43 (n_617, n_149, n_175);
  nand g44 (n_612, n_149, n_175);
  nor g45 (n_613, n_148, n_174);
  nand g46 (n_614, n_148, n_174);
  nor g47 (n_623, n_147, n_173);
  nand g48 (n_618, n_147, n_173);
  nor g49 (n_619, n_146, n_172);
  nand g50 (n_620, n_146, n_172);
  nor g51 (n_629, n_145, n_171);
  nand g52 (n_624, n_145, n_171);
  nor g53 (n_625, n_144, n_170);
  nand g54 (n_626, n_144, n_170);
  nor g55 (n_633, n_143, n_169);
  nand g56 (n_630, n_143, n_169);
  nand g61 (n_634, n_562, n_563);
  nor g62 (n_567, n_564, n_565);
  nor g65 (n_167, n_569, n_565);
  nor g66 (n_573, n_570, n_571);
  nor g69 (n_642, n_575, n_571);
  nor g70 (n_579, n_576, n_577);
  nor g73 (n_644, n_581, n_577);
  nor g74 (n_585, n_582, n_583);
  nor g483 (n_652, n_587, n_583);
  nor g484 (n_591, n_588, n_589);
  nor g487 (n_654, n_593, n_589);
  nor g488 (n_597, n_594, n_595);
  nor g491 (n_662, n_599, n_595);
  nor g492 (n_603, n_600, n_601);
  nor g495 (n_664, n_605, n_601);
  nor g496 (n_609, n_606, n_607);
  nor g499 (n_672, n_611, n_607);
  nor g500 (n_615, n_612, n_613);
  nor g503 (n_674, n_617, n_613);
  nor g504 (n_621, n_618, n_619);
  nor g507 (n_682, n_623, n_619);
  nor g508 (n_627, n_624, n_625);
  nor g511 (n_684, n_629, n_625);
  nand g514 (n_785, n_564, n_636);
  nand g515 (n_638, n_167, n_634);
  nand g516 (n_689, n_637, n_638);
  nor g517 (n_640, n_581, n_639);
  nand g526 (n_697, n_642, n_644);
  nor g527 (n_650, n_593, n_649);
  nand g536 (n_704, n_652, n_654);
  nor g537 (n_660, n_605, n_659);
  nand g546 (n_712, n_662, n_664);
  nor g547 (n_670, n_617, n_669);
  nand g556 (n_719, n_672, n_674);
  nor g557 (n_680, n_629, n_679);
  nand g566 (n_727, n_682, n_684);
  nand g569 (n_789, n_570, n_691);
  nand g570 (n_692, n_642, n_689);
  nand g571 (n_791, n_639, n_692);
  nand g574 (n_794, n_695, n_696);
  nand g577 (n_731, n_699, n_700);
  nor g578 (n_702, n_599, n_701);
  nor g581 (n_741, n_599, n_704);
  nor g587 (n_710, n_708, n_701);
  nor g590 (n_747, n_704, n_708);
  nor g591 (n_714, n_712, n_701);
  nor g594 (n_750, n_704, n_712);
  nor g595 (n_717, n_623, n_716);
  nor g598 (n_768, n_623, n_719);
  nor g604 (n_725, n_723, n_716);
  nor g607 (n_774, n_719, n_723);
  nor g608 (n_729, n_727, n_716);
  nor g611 (n_756, n_719, n_727);
  nand g614 (n_798, n_582, n_733);
  nand g615 (n_734, n_652, n_731);
  nand g616 (n_800, n_649, n_734);
  nand g619 (n_803, n_737, n_738);
  nand g622 (n_806, n_701, n_740);
  nand g623 (n_743, n_741, n_731);
  nand g624 (n_809, n_742, n_743);
  nand g625 (n_746, n_744, n_731);
  nand g626 (n_811, n_745, n_746);
  nand g627 (n_749, n_747, n_731);
  nand g628 (n_814, n_748, n_749);
  nand g629 (n_752, n_750, n_731);
  nand g630 (n_758, n_751, n_752);
  nor g631 (n_754, n_633, n_753);
  nand g638 (n_818, n_606, n_760);
  nand g639 (n_761, n_672, n_758);
  nand g640 (n_820, n_669, n_761);
  nand g643 (n_823, n_764, n_765);
  nand g646 (n_826, n_716, n_767);
  nand g647 (n_770, n_768, n_758);
  nand g648 (n_829, n_769, n_770);
  nand g649 (n_773, n_771, n_758);
  nand g650 (n_831, n_772, n_773);
  nand g651 (n_776, n_774, n_758);
  nand g652 (n_834, n_775, n_776);
  nand g653 (n_777, n_756, n_758);
  nand g654 (n_836, n_753, n_777);
  nand g657 (n_839, n_780, n_781);
  xnor g659 (out_0[1], n_560, n_782);
  xnor g661 (out_0[2], n_634, n_783);
  xnor g664 (out_0[3], n_785, n_786);
  xnor g666 (out_0[4], n_689, n_787);
  xnor g669 (out_0[5], n_789, n_790);
  xnor g671 (out_0[6], n_791, n_792);
  xnor g674 (out_0[7], n_794, n_795);
  xnor g676 (out_0[8], n_731, n_796);
  xnor g679 (out_0[9], n_798, n_799);
  xnor g681 (out_0[10], n_800, n_801);
  xnor g684 (out_0[11], n_803, n_804);
  xnor g687 (out_0[12], n_806, n_807);
  xnor g690 (out_0[13], n_809, n_810);
  xnor g692 (out_0[14], n_811, n_812);
  xnor g695 (out_0[15], n_814, n_815);
  xnor g697 (out_0[16], n_758, n_816);
  xnor g700 (out_0[17], n_818, n_819);
  xnor g702 (out_0[18], n_820, n_821);
  xnor g705 (out_0[19], n_823, n_824);
  xnor g708 (out_0[20], n_826, n_827);
  xnor g711 (out_0[21], n_829, n_830);
  xnor g713 (out_0[22], n_831, n_832);
  xnor g716 (out_0[23], n_834, n_835);
  xnor g718 (out_0[24], n_836, n_837);
  xor g722 (out_0[0], in_2[0], n_841);
  xor g723 (n_280, in_0[22], in_1[22]);
  nor g724 (n_143, in_0[22], in_1[22]);
  xor g725 (n_538, in_3[22], in_4[22]);
  or g726 (n_539, in_3[22], in_4[22]);
  or g727 (n_540, in_2[22], in_4[22]);
  or g728 (n_541, in_2[22], in_3[22]);
  xnor g729 (n_282, n_538, in_2[22]);
  xnor g733 (n_283, n_281, n_280);
  or g734 (n_289, n_280, wc, n_281);
  not gc (wc, n_544);
  xnor g735 (n_550, n_287, n_143);
  or g736 (n_551, n_143, wc0);
  not gc0 (wc0, n_287);
  or g737 (n_552, wc1, n_143);
  not gc1 (wc1, n_289);
  or g738 (n_563, n_559, wc2);
  not gc2 (wc2, n_560);
  or g739 (n_782, wc3, n_559);
  not gc3 (wc3, n_562);
  and g740 (n_637, wc4, n_566);
  not gc4 (wc4, n_567);
  or g741 (n_783, wc5, n_569);
  not gc5 (wc5, n_564);
  or g742 (n_786, wc6, n_565);
  not gc6 (wc6, n_566);
  and g743 (n_639, wc7, n_572);
  not gc7 (wc7, n_573);
  or g744 (n_636, wc8, n_569);
  not gc8 (wc8, n_634);
  or g745 (n_787, wc9, n_575);
  not gc9 (wc9, n_570);
  or g746 (n_790, wc10, n_571);
  not gc10 (wc10, n_572);
  and g747 (n_646, wc11, n_578);
  not gc11 (wc11, n_579);
  and g748 (n_649, wc12, n_584);
  not gc12 (wc12, n_585);
  and g749 (n_656, wc13, n_590);
  not gc13 (wc13, n_591);
  and g750 (n_659, wc14, n_596);
  not gc14 (wc14, n_597);
  and g751 (n_666, wc15, n_602);
  not gc15 (wc15, n_603);
  and g752 (n_669, wc16, n_608);
  not gc16 (wc16, n_609);
  and g753 (n_676, wc17, n_614);
  not gc17 (wc17, n_615);
  and g754 (n_679, wc18, n_620);
  not gc18 (wc18, n_621);
  and g755 (n_686, wc19, n_626);
  not gc19 (wc19, n_627);
  or g756 (n_693, wc20, n_581);
  not gc20 (wc20, n_642);
  or g757 (n_735, wc21, n_593);
  not gc21 (wc21, n_652);
  or g758 (n_708, wc22, n_605);
  not gc22 (wc22, n_662);
  or g759 (n_762, wc23, n_617);
  not gc23 (wc23, n_672);
  or g760 (n_723, wc24, n_629);
  not gc24 (wc24, n_682);
  or g761 (n_792, wc25, n_581);
  not gc25 (wc25, n_576);
  or g762 (n_795, wc26, n_577);
  not gc26 (wc26, n_578);
  or g763 (n_796, wc27, n_587);
  not gc27 (wc27, n_582);
  or g764 (n_799, wc28, n_583);
  not gc28 (wc28, n_584);
  or g765 (n_801, wc29, n_593);
  not gc29 (wc29, n_588);
  or g766 (n_804, wc30, n_589);
  not gc30 (wc30, n_590);
  or g767 (n_807, wc31, n_599);
  not gc31 (wc31, n_594);
  or g768 (n_810, wc32, n_595);
  not gc32 (wc32, n_596);
  or g769 (n_812, wc33, n_605);
  not gc33 (wc33, n_600);
  or g770 (n_815, wc34, n_601);
  not gc34 (wc34, n_602);
  or g771 (n_816, wc35, n_611);
  not gc35 (wc35, n_606);
  or g772 (n_819, wc36, n_607);
  not gc36 (wc36, n_608);
  or g773 (n_821, wc37, n_617);
  not gc37 (wc37, n_612);
  or g774 (n_824, wc38, n_613);
  not gc38 (wc38, n_614);
  or g775 (n_827, wc39, n_623);
  not gc39 (wc39, n_618);
  or g776 (n_830, wc40, n_619);
  not gc40 (wc40, n_620);
  or g777 (n_832, wc41, n_629);
  not gc41 (wc41, n_624);
  or g778 (n_835, wc42, n_625);
  not gc42 (wc42, n_626);
  or g779 (n_837, wc43, n_633);
  not gc43 (wc43, n_630);
  and g780 (n_695, wc44, n_576);
  not gc44 (wc44, n_640);
  and g781 (n_647, wc45, n_644);
  not gc45 (wc45, n_639);
  and g782 (n_657, wc46, n_654);
  not gc46 (wc46, n_649);
  and g783 (n_667, wc47, n_664);
  not gc47 (wc47, n_659);
  and g784 (n_677, wc48, n_674);
  not gc48 (wc48, n_669);
  and g785 (n_687, wc49, n_684);
  not gc49 (wc49, n_679);
  or g786 (n_691, wc50, n_575);
  not gc50 (wc50, n_689);
  and g787 (n_744, wc51, n_662);
  not gc51 (wc51, n_704);
  and g788 (n_771, wc52, n_682);
  not gc52 (wc52, n_719);
  and g789 (n_699, wc53, n_646);
  not gc53 (wc53, n_647);
  and g790 (n_737, wc54, n_588);
  not gc54 (wc54, n_650);
  and g791 (n_701, wc55, n_656);
  not gc55 (wc55, n_657);
  and g792 (n_709, wc56, n_600);
  not gc56 (wc56, n_660);
  and g793 (n_713, wc57, n_666);
  not gc57 (wc57, n_667);
  and g794 (n_764, wc58, n_612);
  not gc58 (wc58, n_670);
  and g795 (n_716, wc59, n_676);
  not gc59 (wc59, n_677);
  and g796 (n_724, wc60, n_624);
  not gc60 (wc60, n_680);
  and g797 (n_728, wc61, n_686);
  not gc61 (wc61, n_687);
  or g798 (n_696, n_693, wc62);
  not gc62 (wc62, n_689);
  or g799 (n_700, n_697, wc63);
  not gc63 (wc63, n_689);
  or g800 (n_778, wc64, n_633);
  not gc64 (wc64, n_756);
  and g801 (n_706, wc65, n_662);
  not gc65 (wc65, n_701);
  and g802 (n_721, wc66, n_682);
  not gc66 (wc66, n_716);
  and g803 (n_742, wc67, n_594);
  not gc67 (wc67, n_702);
  and g804 (n_745, wc68, n_659);
  not gc68 (wc68, n_706);
  and g805 (n_748, n_709, wc69);
  not gc69 (wc69, n_710);
  and g806 (n_751, n_713, wc70);
  not gc70 (wc70, n_714);
  and g807 (n_769, wc71, n_618);
  not gc71 (wc71, n_717);
  and g808 (n_772, wc72, n_679);
  not gc72 (wc72, n_721);
  and g809 (n_775, n_724, wc73);
  not gc73 (wc73, n_725);
  and g810 (n_753, n_728, wc74);
  not gc74 (wc74, n_729);
  or g811 (n_733, wc75, n_587);
  not gc75 (wc75, n_731);
  or g812 (n_738, n_735, wc76);
  not gc76 (wc76, n_731);
  or g813 (n_740, wc77, n_704);
  not gc77 (wc77, n_731);
  and g814 (n_780, wc78, n_630);
  not gc78 (wc78, n_754);
  or g815 (n_760, wc79, n_611);
  not gc79 (wc79, n_758);
  or g816 (n_765, n_762, wc80);
  not gc80 (wc80, n_758);
  or g817 (n_767, wc81, n_719);
  not gc81 (wc81, n_758);
  or g818 (n_781, n_778, wc82);
  not gc82 (wc82, n_758);
  not g819 (out_0[25], n_839);
endmodule

module csa_tree_add_823_44_group_6807_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  csa_tree_add_823_44_group_6807_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_897_44_group_6805_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_280, n_281, n_282, n_283, n_284, n_287;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_544, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_556, n_557;
  wire n_558, n_559, n_560, n_562, n_563, n_564, n_565, n_566;
  wire n_567, n_569, n_570, n_571, n_572, n_573, n_575, n_576;
  wire n_577, n_578, n_579, n_581, n_582, n_583, n_584, n_585;
  wire n_587, n_588, n_589, n_590, n_591, n_593, n_594, n_595;
  wire n_596, n_597, n_599, n_600, n_601, n_602, n_603, n_605;
  wire n_606, n_607, n_608, n_609, n_611, n_612, n_613, n_614;
  wire n_615, n_617, n_618, n_619, n_620, n_621, n_623, n_624;
  wire n_625, n_626, n_627, n_629, n_630, n_633, n_634, n_636;
  wire n_637, n_638, n_639, n_640, n_642, n_644, n_646, n_647;
  wire n_649, n_650, n_652, n_654, n_656, n_657, n_659, n_660;
  wire n_662, n_664, n_666, n_667, n_669, n_670, n_672, n_674;
  wire n_676, n_677, n_679, n_680, n_682, n_684, n_686, n_687;
  wire n_689, n_691, n_692, n_693, n_695, n_696, n_697, n_699;
  wire n_700, n_701, n_702, n_704, n_706, n_708, n_709, n_710;
  wire n_712, n_713, n_714, n_716, n_717, n_719, n_721, n_723;
  wire n_724, n_725, n_727, n_728, n_729, n_731, n_733, n_734;
  wire n_735, n_737, n_738, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_756, n_758, n_760, n_761, n_762, n_764;
  wire n_765, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_780, n_781, n_782;
  wire n_783, n_785, n_786, n_787, n_789, n_790, n_791, n_792;
  wire n_794, n_795, n_796, n_798, n_799, n_800, n_801, n_803;
  wire n_804, n_806, n_807, n_809, n_810, n_811, n_812, n_814;
  wire n_815, n_816, n_818, n_819, n_820, n_821, n_823, n_824;
  wire n_826, n_827, n_829, n_830, n_831, n_832, n_834, n_835;
  wire n_836, n_837, n_839, n_841;
  xor g75 (n_290, in_0[0], in_4[0]);
  xor g76 (n_193, n_290, in_3[0]);
  nand g77 (n_291, in_0[0], in_4[0]);
  nand g78 (n_292, in_3[0], in_4[0]);
  nand g79 (n_293, in_0[0], in_3[0]);
  nand g6 (n_195, n_291, n_292, n_293);
  xor g80 (n_294, in_0[1], in_1[1]);
  xor g81 (n_166, n_294, in_4[1]);
  nand g82 (n_295, in_0[1], in_1[1]);
  nand g83 (n_296, in_4[1], in_1[1]);
  nand g84 (n_297, in_0[1], in_4[1]);
  nand g85 (n_197, n_295, n_296, n_297);
  xor g86 (n_298, in_3[1], in_2[1]);
  xor g87 (n_192, n_298, n_195);
  nand g88 (n_299, in_3[1], in_2[1]);
  nand g89 (n_300, n_195, in_2[1]);
  nand g90 (n_301, in_3[1], n_195);
  nand g91 (n_165, n_299, n_300, n_301);
  xor g92 (n_196, in_0[2], in_1[2]);
  and g93 (n_199, in_0[2], in_1[2]);
  xor g94 (n_302, in_3[2], in_4[2]);
  xor g95 (n_198, n_302, in_2[2]);
  nand g96 (n_303, in_3[2], in_4[2]);
  nand g97 (n_304, in_2[2], in_4[2]);
  nand g98 (n_305, in_3[2], in_2[2]);
  nand g99 (n_200, n_303, n_304, n_305);
  xor g100 (n_306, n_196, n_197);
  xor g101 (n_191, n_306, n_198);
  nand g102 (n_307, n_196, n_197);
  nand g103 (n_308, n_198, n_197);
  nand g104 (n_309, n_196, n_198);
  nand g105 (n_164, n_307, n_308, n_309);
  xor g106 (n_310, in_0[3], in_1[3]);
  xor g107 (n_201, n_310, in_3[3]);
  nand g108 (n_311, in_0[3], in_1[3]);
  nand g109 (n_312, in_3[3], in_1[3]);
  nand g110 (n_313, in_0[3], in_3[3]);
  nand g111 (n_203, n_311, n_312, n_313);
  xor g112 (n_314, in_4[3], in_2[3]);
  xor g113 (n_202, n_314, n_199);
  nand g114 (n_315, in_4[3], in_2[3]);
  nand g115 (n_316, n_199, in_2[3]);
  nand g116 (n_317, in_4[3], n_199);
  nand g117 (n_205, n_315, n_316, n_317);
  xor g118 (n_318, n_200, n_201);
  xor g119 (n_190, n_318, n_202);
  nand g120 (n_319, n_200, n_201);
  nand g121 (n_320, n_202, n_201);
  nand g122 (n_321, n_200, n_202);
  nand g123 (n_163, n_319, n_320, n_321);
  xor g124 (n_322, in_0[4], in_1[4]);
  xor g125 (n_204, n_322, in_3[4]);
  nand g126 (n_323, in_0[4], in_1[4]);
  nand g127 (n_324, in_3[4], in_1[4]);
  nand g128 (n_325, in_0[4], in_3[4]);
  nand g129 (n_207, n_323, n_324, n_325);
  xor g130 (n_326, in_4[4], in_2[4]);
  xor g131 (n_206, n_326, n_203);
  nand g132 (n_327, in_4[4], in_2[4]);
  nand g133 (n_328, n_203, in_2[4]);
  nand g134 (n_329, in_4[4], n_203);
  nand g135 (n_210, n_327, n_328, n_329);
  xor g136 (n_330, n_204, n_205);
  xor g137 (n_189, n_330, n_206);
  nand g138 (n_331, n_204, n_205);
  nand g139 (n_332, n_206, n_205);
  nand g140 (n_333, n_204, n_206);
  nand g141 (n_162, n_331, n_332, n_333);
  xor g142 (n_334, in_0[5], in_1[5]);
  xor g143 (n_208, n_334, in_3[5]);
  nand g144 (n_335, in_0[5], in_1[5]);
  nand g145 (n_336, in_3[5], in_1[5]);
  nand g146 (n_337, in_0[5], in_3[5]);
  nand g147 (n_211, n_335, n_336, n_337);
  xor g148 (n_338, in_4[5], in_2[5]);
  xor g149 (n_209, n_338, n_207);
  nand g150 (n_339, in_4[5], in_2[5]);
  nand g151 (n_340, n_207, in_2[5]);
  nand g152 (n_341, in_4[5], n_207);
  nand g153 (n_214, n_339, n_340, n_341);
  xor g154 (n_342, n_208, n_209);
  xor g155 (n_188, n_342, n_210);
  nand g156 (n_343, n_208, n_209);
  nand g157 (n_344, n_210, n_209);
  nand g158 (n_345, n_208, n_210);
  nand g159 (n_161, n_343, n_344, n_345);
  xor g160 (n_346, in_0[6], in_1[6]);
  xor g161 (n_212, n_346, in_3[6]);
  nand g162 (n_347, in_0[6], in_1[6]);
  nand g163 (n_348, in_3[6], in_1[6]);
  nand g164 (n_349, in_0[6], in_3[6]);
  nand g165 (n_215, n_347, n_348, n_349);
  xor g166 (n_350, in_4[6], in_2[6]);
  xor g167 (n_213, n_350, n_211);
  nand g168 (n_351, in_4[6], in_2[6]);
  nand g169 (n_352, n_211, in_2[6]);
  nand g170 (n_353, in_4[6], n_211);
  nand g171 (n_218, n_351, n_352, n_353);
  xor g172 (n_354, n_212, n_213);
  xor g173 (n_187, n_354, n_214);
  nand g174 (n_355, n_212, n_213);
  nand g175 (n_356, n_214, n_213);
  nand g176 (n_357, n_212, n_214);
  nand g177 (n_160, n_355, n_356, n_357);
  xor g178 (n_358, in_0[7], in_1[7]);
  xor g179 (n_216, n_358, in_3[7]);
  nand g180 (n_359, in_0[7], in_1[7]);
  nand g181 (n_360, in_3[7], in_1[7]);
  nand g182 (n_361, in_0[7], in_3[7]);
  nand g183 (n_219, n_359, n_360, n_361);
  xor g184 (n_362, in_4[7], in_2[7]);
  xor g185 (n_217, n_362, n_215);
  nand g186 (n_363, in_4[7], in_2[7]);
  nand g187 (n_364, n_215, in_2[7]);
  nand g188 (n_365, in_4[7], n_215);
  nand g189 (n_222, n_363, n_364, n_365);
  xor g190 (n_366, n_216, n_217);
  xor g191 (n_186, n_366, n_218);
  nand g192 (n_367, n_216, n_217);
  nand g193 (n_368, n_218, n_217);
  nand g194 (n_369, n_216, n_218);
  nand g195 (n_159, n_367, n_368, n_369);
  xor g196 (n_370, in_0[8], in_1[8]);
  xor g197 (n_220, n_370, in_3[8]);
  nand g198 (n_371, in_0[8], in_1[8]);
  nand g199 (n_372, in_3[8], in_1[8]);
  nand g200 (n_373, in_0[8], in_3[8]);
  nand g201 (n_223, n_371, n_372, n_373);
  xor g202 (n_374, in_4[8], in_2[8]);
  xor g203 (n_221, n_374, n_219);
  nand g204 (n_375, in_4[8], in_2[8]);
  nand g205 (n_376, n_219, in_2[8]);
  nand g206 (n_377, in_4[8], n_219);
  nand g207 (n_226, n_375, n_376, n_377);
  xor g208 (n_378, n_220, n_221);
  xor g209 (n_185, n_378, n_222);
  nand g210 (n_379, n_220, n_221);
  nand g211 (n_380, n_222, n_221);
  nand g212 (n_381, n_220, n_222);
  nand g213 (n_158, n_379, n_380, n_381);
  xor g214 (n_382, in_0[9], in_1[9]);
  xor g215 (n_224, n_382, in_3[9]);
  nand g216 (n_383, in_0[9], in_1[9]);
  nand g217 (n_384, in_3[9], in_1[9]);
  nand g218 (n_385, in_0[9], in_3[9]);
  nand g219 (n_227, n_383, n_384, n_385);
  xor g220 (n_386, in_4[9], in_2[9]);
  xor g221 (n_225, n_386, n_223);
  nand g222 (n_387, in_4[9], in_2[9]);
  nand g223 (n_388, n_223, in_2[9]);
  nand g224 (n_389, in_4[9], n_223);
  nand g225 (n_230, n_387, n_388, n_389);
  xor g226 (n_390, n_224, n_225);
  xor g227 (n_184, n_390, n_226);
  nand g228 (n_391, n_224, n_225);
  nand g229 (n_392, n_226, n_225);
  nand g230 (n_393, n_224, n_226);
  nand g231 (n_157, n_391, n_392, n_393);
  xor g232 (n_394, in_0[10], in_1[10]);
  xor g233 (n_228, n_394, in_3[10]);
  nand g234 (n_395, in_0[10], in_1[10]);
  nand g235 (n_396, in_3[10], in_1[10]);
  nand g236 (n_397, in_0[10], in_3[10]);
  nand g237 (n_231, n_395, n_396, n_397);
  xor g238 (n_398, in_4[10], in_2[10]);
  xor g239 (n_229, n_398, n_227);
  nand g240 (n_399, in_4[10], in_2[10]);
  nand g241 (n_400, n_227, in_2[10]);
  nand g242 (n_401, in_4[10], n_227);
  nand g243 (n_234, n_399, n_400, n_401);
  xor g244 (n_402, n_228, n_229);
  xor g245 (n_183, n_402, n_230);
  nand g246 (n_403, n_228, n_229);
  nand g247 (n_404, n_230, n_229);
  nand g248 (n_405, n_228, n_230);
  nand g249 (n_156, n_403, n_404, n_405);
  xor g250 (n_406, in_0[11], in_1[11]);
  xor g251 (n_232, n_406, in_3[11]);
  nand g252 (n_407, in_0[11], in_1[11]);
  nand g253 (n_408, in_3[11], in_1[11]);
  nand g254 (n_409, in_0[11], in_3[11]);
  nand g255 (n_235, n_407, n_408, n_409);
  xor g256 (n_410, in_4[11], in_2[11]);
  xor g257 (n_233, n_410, n_231);
  nand g258 (n_411, in_4[11], in_2[11]);
  nand g259 (n_412, n_231, in_2[11]);
  nand g260 (n_413, in_4[11], n_231);
  nand g261 (n_238, n_411, n_412, n_413);
  xor g262 (n_414, n_232, n_233);
  xor g263 (n_182, n_414, n_234);
  nand g264 (n_415, n_232, n_233);
  nand g265 (n_416, n_234, n_233);
  nand g266 (n_417, n_232, n_234);
  nand g267 (n_155, n_415, n_416, n_417);
  xor g268 (n_418, in_0[12], in_1[12]);
  xor g269 (n_236, n_418, in_3[12]);
  nand g270 (n_419, in_0[12], in_1[12]);
  nand g271 (n_420, in_3[12], in_1[12]);
  nand g272 (n_421, in_0[12], in_3[12]);
  nand g273 (n_239, n_419, n_420, n_421);
  xor g274 (n_422, in_4[12], in_2[12]);
  xor g275 (n_237, n_422, n_235);
  nand g276 (n_423, in_4[12], in_2[12]);
  nand g277 (n_424, n_235, in_2[12]);
  nand g278 (n_425, in_4[12], n_235);
  nand g279 (n_242, n_423, n_424, n_425);
  xor g280 (n_426, n_236, n_237);
  xor g281 (n_181, n_426, n_238);
  nand g282 (n_427, n_236, n_237);
  nand g283 (n_428, n_238, n_237);
  nand g284 (n_429, n_236, n_238);
  nand g285 (n_154, n_427, n_428, n_429);
  xor g286 (n_430, in_0[13], in_1[13]);
  xor g287 (n_240, n_430, in_3[13]);
  nand g288 (n_431, in_0[13], in_1[13]);
  nand g289 (n_432, in_3[13], in_1[13]);
  nand g290 (n_433, in_0[13], in_3[13]);
  nand g291 (n_243, n_431, n_432, n_433);
  xor g292 (n_434, in_4[13], in_2[13]);
  xor g293 (n_241, n_434, n_239);
  nand g294 (n_435, in_4[13], in_2[13]);
  nand g295 (n_436, n_239, in_2[13]);
  nand g296 (n_437, in_4[13], n_239);
  nand g297 (n_246, n_435, n_436, n_437);
  xor g298 (n_438, n_240, n_241);
  xor g299 (n_180, n_438, n_242);
  nand g300 (n_439, n_240, n_241);
  nand g301 (n_440, n_242, n_241);
  nand g302 (n_441, n_240, n_242);
  nand g303 (n_153, n_439, n_440, n_441);
  xor g304 (n_442, in_0[14], in_1[14]);
  xor g305 (n_244, n_442, in_3[14]);
  nand g306 (n_443, in_0[14], in_1[14]);
  nand g307 (n_444, in_3[14], in_1[14]);
  nand g308 (n_445, in_0[14], in_3[14]);
  nand g309 (n_247, n_443, n_444, n_445);
  xor g310 (n_446, in_4[14], in_2[14]);
  xor g311 (n_245, n_446, n_243);
  nand g312 (n_447, in_4[14], in_2[14]);
  nand g313 (n_448, n_243, in_2[14]);
  nand g314 (n_449, in_4[14], n_243);
  nand g315 (n_250, n_447, n_448, n_449);
  xor g316 (n_450, n_244, n_245);
  xor g317 (n_179, n_450, n_246);
  nand g318 (n_451, n_244, n_245);
  nand g319 (n_452, n_246, n_245);
  nand g320 (n_453, n_244, n_246);
  nand g321 (n_152, n_451, n_452, n_453);
  xor g322 (n_454, in_0[15], in_1[15]);
  xor g323 (n_248, n_454, in_3[15]);
  nand g324 (n_455, in_0[15], in_1[15]);
  nand g325 (n_456, in_3[15], in_1[15]);
  nand g326 (n_457, in_0[15], in_3[15]);
  nand g327 (n_251, n_455, n_456, n_457);
  xor g328 (n_458, in_4[15], in_2[15]);
  xor g329 (n_249, n_458, n_247);
  nand g330 (n_459, in_4[15], in_2[15]);
  nand g331 (n_460, n_247, in_2[15]);
  nand g332 (n_461, in_4[15], n_247);
  nand g333 (n_254, n_459, n_460, n_461);
  xor g334 (n_462, n_248, n_249);
  xor g335 (n_178, n_462, n_250);
  nand g336 (n_463, n_248, n_249);
  nand g337 (n_464, n_250, n_249);
  nand g338 (n_465, n_248, n_250);
  nand g339 (n_151, n_463, n_464, n_465);
  xor g340 (n_466, in_0[16], in_1[16]);
  xor g341 (n_252, n_466, in_3[16]);
  nand g342 (n_467, in_0[16], in_1[16]);
  nand g343 (n_468, in_3[16], in_1[16]);
  nand g344 (n_469, in_0[16], in_3[16]);
  nand g345 (n_255, n_467, n_468, n_469);
  xor g346 (n_470, in_4[16], in_2[16]);
  xor g347 (n_253, n_470, n_251);
  nand g348 (n_471, in_4[16], in_2[16]);
  nand g349 (n_472, n_251, in_2[16]);
  nand g350 (n_473, in_4[16], n_251);
  nand g351 (n_258, n_471, n_472, n_473);
  xor g352 (n_474, n_252, n_253);
  xor g353 (n_177, n_474, n_254);
  nand g354 (n_475, n_252, n_253);
  nand g355 (n_476, n_254, n_253);
  nand g356 (n_477, n_252, n_254);
  nand g357 (n_150, n_475, n_476, n_477);
  xor g358 (n_478, in_0[17], in_1[17]);
  xor g359 (n_256, n_478, in_3[17]);
  nand g360 (n_479, in_0[17], in_1[17]);
  nand g361 (n_480, in_3[17], in_1[17]);
  nand g362 (n_481, in_0[17], in_3[17]);
  nand g363 (n_259, n_479, n_480, n_481);
  xor g364 (n_482, in_4[17], in_2[17]);
  xor g365 (n_257, n_482, n_255);
  nand g366 (n_483, in_4[17], in_2[17]);
  nand g367 (n_484, n_255, in_2[17]);
  nand g368 (n_485, in_4[17], n_255);
  nand g369 (n_262, n_483, n_484, n_485);
  xor g370 (n_486, n_256, n_257);
  xor g371 (n_176, n_486, n_258);
  nand g372 (n_487, n_256, n_257);
  nand g373 (n_488, n_258, n_257);
  nand g374 (n_489, n_256, n_258);
  nand g375 (n_149, n_487, n_488, n_489);
  xor g376 (n_490, in_0[18], in_1[18]);
  xor g377 (n_260, n_490, in_3[18]);
  nand g378 (n_491, in_0[18], in_1[18]);
  nand g379 (n_492, in_3[18], in_1[18]);
  nand g380 (n_493, in_0[18], in_3[18]);
  nand g381 (n_263, n_491, n_492, n_493);
  xor g382 (n_494, in_4[18], in_2[18]);
  xor g383 (n_261, n_494, n_259);
  nand g384 (n_495, in_4[18], in_2[18]);
  nand g385 (n_496, n_259, in_2[18]);
  nand g386 (n_497, in_4[18], n_259);
  nand g387 (n_266, n_495, n_496, n_497);
  xor g388 (n_498, n_260, n_261);
  xor g389 (n_175, n_498, n_262);
  nand g390 (n_499, n_260, n_261);
  nand g391 (n_500, n_262, n_261);
  nand g392 (n_501, n_260, n_262);
  nand g393 (n_148, n_499, n_500, n_501);
  xor g394 (n_502, in_0[19], in_1[19]);
  xor g395 (n_264, n_502, in_3[19]);
  nand g396 (n_503, in_0[19], in_1[19]);
  nand g397 (n_504, in_3[19], in_1[19]);
  nand g398 (n_505, in_0[19], in_3[19]);
  nand g399 (n_267, n_503, n_504, n_505);
  xor g400 (n_506, in_4[19], in_2[19]);
  xor g401 (n_265, n_506, n_263);
  nand g402 (n_507, in_4[19], in_2[19]);
  nand g403 (n_508, n_263, in_2[19]);
  nand g404 (n_509, in_4[19], n_263);
  nand g405 (n_270, n_507, n_508, n_509);
  xor g406 (n_510, n_264, n_265);
  xor g407 (n_174, n_510, n_266);
  nand g408 (n_511, n_264, n_265);
  nand g409 (n_512, n_266, n_265);
  nand g410 (n_513, n_264, n_266);
  nand g411 (n_147, n_511, n_512, n_513);
  xor g412 (n_514, in_0[20], in_1[20]);
  xor g413 (n_268, n_514, in_3[20]);
  nand g414 (n_515, in_0[20], in_1[20]);
  nand g415 (n_516, in_3[20], in_1[20]);
  nand g416 (n_517, in_0[20], in_3[20]);
  nand g417 (n_271, n_515, n_516, n_517);
  xor g418 (n_518, in_4[20], in_2[20]);
  xor g419 (n_269, n_518, n_267);
  nand g420 (n_519, in_4[20], in_2[20]);
  nand g421 (n_520, n_267, in_2[20]);
  nand g422 (n_521, in_4[20], n_267);
  nand g423 (n_274, n_519, n_520, n_521);
  xor g424 (n_522, n_268, n_269);
  xor g425 (n_173, n_522, n_270);
  nand g426 (n_523, n_268, n_269);
  nand g427 (n_524, n_270, n_269);
  nand g428 (n_525, n_268, n_270);
  nand g429 (n_146, n_523, n_524, n_525);
  xor g430 (n_526, in_0[21], in_1[21]);
  xor g431 (n_272, n_526, in_3[21]);
  nand g432 (n_527, in_0[21], in_1[21]);
  nand g433 (n_528, in_3[21], in_1[21]);
  nand g434 (n_529, in_0[21], in_3[21]);
  nand g435 (n_281, n_527, n_528, n_529);
  xor g436 (n_530, in_4[21], in_2[21]);
  xor g437 (n_273, n_530, n_271);
  nand g438 (n_531, in_4[21], in_2[21]);
  nand g439 (n_532, n_271, in_2[21]);
  nand g440 (n_533, in_4[21], n_271);
  nand g441 (n_284, n_531, n_532, n_533);
  xor g442 (n_534, n_272, n_273);
  xor g443 (n_172, n_534, n_274);
  nand g444 (n_535, n_272, n_273);
  nand g445 (n_536, n_274, n_273);
  nand g446 (n_537, n_272, n_274);
  nand g447 (n_145, n_535, n_536, n_537);
  nand g455 (n_287, n_539, n_540, n_541);
  nand g459 (n_544, n_281, n_280);
  xor g462 (n_546, n_282, n_283);
  xor g463 (n_171, n_546, n_284);
  nand g464 (n_547, n_282, n_283);
  nand g465 (n_548, n_284, n_283);
  nand g466 (n_549, n_282, n_284);
  nand g467 (n_144, n_547, n_548, n_549);
  xor g471 (n_170, n_550, n_289);
  nand g474 (n_553, n_287, n_289);
  nand g475 (n_169, n_551, n_552, n_553);
  xor g478 (n_841, in_1[0], n_193);
  nand g479 (n_556, in_1[0], n_193);
  nand g480 (n_557, in_1[0], in_2[0]);
  nand g7 (n_558, n_193, in_2[0]);
  nand g8 (n_560, n_556, n_557, n_558);
  nor g9 (n_559, n_166, n_192);
  nand g10 (n_562, n_166, n_192);
  nor g11 (n_569, n_165, n_191);
  nand g12 (n_564, n_165, n_191);
  nor g13 (n_565, n_164, n_190);
  nand g14 (n_566, n_164, n_190);
  nor g15 (n_575, n_163, n_189);
  nand g16 (n_570, n_163, n_189);
  nor g17 (n_571, n_162, n_188);
  nand g18 (n_572, n_162, n_188);
  nor g19 (n_581, n_161, n_187);
  nand g20 (n_576, n_161, n_187);
  nor g21 (n_577, n_160, n_186);
  nand g22 (n_578, n_160, n_186);
  nor g23 (n_587, n_159, n_185);
  nand g24 (n_582, n_159, n_185);
  nor g25 (n_583, n_158, n_184);
  nand g26 (n_584, n_158, n_184);
  nor g27 (n_593, n_157, n_183);
  nand g28 (n_588, n_157, n_183);
  nor g29 (n_589, n_156, n_182);
  nand g30 (n_590, n_156, n_182);
  nor g31 (n_599, n_155, n_181);
  nand g32 (n_594, n_155, n_181);
  nor g33 (n_595, n_154, n_180);
  nand g34 (n_596, n_154, n_180);
  nor g35 (n_605, n_153, n_179);
  nand g36 (n_600, n_153, n_179);
  nor g37 (n_601, n_152, n_178);
  nand g38 (n_602, n_152, n_178);
  nor g39 (n_611, n_151, n_177);
  nand g40 (n_606, n_151, n_177);
  nor g41 (n_607, n_150, n_176);
  nand g42 (n_608, n_150, n_176);
  nor g43 (n_617, n_149, n_175);
  nand g44 (n_612, n_149, n_175);
  nor g45 (n_613, n_148, n_174);
  nand g46 (n_614, n_148, n_174);
  nor g47 (n_623, n_147, n_173);
  nand g48 (n_618, n_147, n_173);
  nor g49 (n_619, n_146, n_172);
  nand g50 (n_620, n_146, n_172);
  nor g51 (n_629, n_145, n_171);
  nand g52 (n_624, n_145, n_171);
  nor g53 (n_625, n_144, n_170);
  nand g54 (n_626, n_144, n_170);
  nor g55 (n_633, n_143, n_169);
  nand g56 (n_630, n_143, n_169);
  nand g61 (n_634, n_562, n_563);
  nor g62 (n_567, n_564, n_565);
  nor g65 (n_167, n_569, n_565);
  nor g66 (n_573, n_570, n_571);
  nor g69 (n_642, n_575, n_571);
  nor g70 (n_579, n_576, n_577);
  nor g73 (n_644, n_581, n_577);
  nor g74 (n_585, n_582, n_583);
  nor g483 (n_652, n_587, n_583);
  nor g484 (n_591, n_588, n_589);
  nor g487 (n_654, n_593, n_589);
  nor g488 (n_597, n_594, n_595);
  nor g491 (n_662, n_599, n_595);
  nor g492 (n_603, n_600, n_601);
  nor g495 (n_664, n_605, n_601);
  nor g496 (n_609, n_606, n_607);
  nor g499 (n_672, n_611, n_607);
  nor g500 (n_615, n_612, n_613);
  nor g503 (n_674, n_617, n_613);
  nor g504 (n_621, n_618, n_619);
  nor g507 (n_682, n_623, n_619);
  nor g508 (n_627, n_624, n_625);
  nor g511 (n_684, n_629, n_625);
  nand g514 (n_785, n_564, n_636);
  nand g515 (n_638, n_167, n_634);
  nand g516 (n_689, n_637, n_638);
  nor g517 (n_640, n_581, n_639);
  nand g526 (n_697, n_642, n_644);
  nor g527 (n_650, n_593, n_649);
  nand g536 (n_704, n_652, n_654);
  nor g537 (n_660, n_605, n_659);
  nand g546 (n_712, n_662, n_664);
  nor g547 (n_670, n_617, n_669);
  nand g556 (n_719, n_672, n_674);
  nor g557 (n_680, n_629, n_679);
  nand g566 (n_727, n_682, n_684);
  nand g569 (n_789, n_570, n_691);
  nand g570 (n_692, n_642, n_689);
  nand g571 (n_791, n_639, n_692);
  nand g574 (n_794, n_695, n_696);
  nand g577 (n_731, n_699, n_700);
  nor g578 (n_702, n_599, n_701);
  nor g581 (n_741, n_599, n_704);
  nor g587 (n_710, n_708, n_701);
  nor g590 (n_747, n_704, n_708);
  nor g591 (n_714, n_712, n_701);
  nor g594 (n_750, n_704, n_712);
  nor g595 (n_717, n_623, n_716);
  nor g598 (n_768, n_623, n_719);
  nor g604 (n_725, n_723, n_716);
  nor g607 (n_774, n_719, n_723);
  nor g608 (n_729, n_727, n_716);
  nor g611 (n_756, n_719, n_727);
  nand g614 (n_798, n_582, n_733);
  nand g615 (n_734, n_652, n_731);
  nand g616 (n_800, n_649, n_734);
  nand g619 (n_803, n_737, n_738);
  nand g622 (n_806, n_701, n_740);
  nand g623 (n_743, n_741, n_731);
  nand g624 (n_809, n_742, n_743);
  nand g625 (n_746, n_744, n_731);
  nand g626 (n_811, n_745, n_746);
  nand g627 (n_749, n_747, n_731);
  nand g628 (n_814, n_748, n_749);
  nand g629 (n_752, n_750, n_731);
  nand g630 (n_758, n_751, n_752);
  nor g631 (n_754, n_633, n_753);
  nand g638 (n_818, n_606, n_760);
  nand g639 (n_761, n_672, n_758);
  nand g640 (n_820, n_669, n_761);
  nand g643 (n_823, n_764, n_765);
  nand g646 (n_826, n_716, n_767);
  nand g647 (n_770, n_768, n_758);
  nand g648 (n_829, n_769, n_770);
  nand g649 (n_773, n_771, n_758);
  nand g650 (n_831, n_772, n_773);
  nand g651 (n_776, n_774, n_758);
  nand g652 (n_834, n_775, n_776);
  nand g653 (n_777, n_756, n_758);
  nand g654 (n_836, n_753, n_777);
  nand g657 (n_839, n_780, n_781);
  xnor g659 (out_0[1], n_560, n_782);
  xnor g661 (out_0[2], n_634, n_783);
  xnor g664 (out_0[3], n_785, n_786);
  xnor g666 (out_0[4], n_689, n_787);
  xnor g669 (out_0[5], n_789, n_790);
  xnor g671 (out_0[6], n_791, n_792);
  xnor g674 (out_0[7], n_794, n_795);
  xnor g676 (out_0[8], n_731, n_796);
  xnor g679 (out_0[9], n_798, n_799);
  xnor g681 (out_0[10], n_800, n_801);
  xnor g684 (out_0[11], n_803, n_804);
  xnor g687 (out_0[12], n_806, n_807);
  xnor g690 (out_0[13], n_809, n_810);
  xnor g692 (out_0[14], n_811, n_812);
  xnor g695 (out_0[15], n_814, n_815);
  xnor g697 (out_0[16], n_758, n_816);
  xnor g700 (out_0[17], n_818, n_819);
  xnor g702 (out_0[18], n_820, n_821);
  xnor g705 (out_0[19], n_823, n_824);
  xnor g708 (out_0[20], n_826, n_827);
  xnor g711 (out_0[21], n_829, n_830);
  xnor g713 (out_0[22], n_831, n_832);
  xnor g716 (out_0[23], n_834, n_835);
  xnor g718 (out_0[24], n_836, n_837);
  xor g722 (out_0[0], in_2[0], n_841);
  xor g723 (n_280, in_0[22], in_1[22]);
  nor g724 (n_143, in_0[22], in_1[22]);
  xor g725 (n_538, in_3[22], in_4[22]);
  or g726 (n_539, in_3[22], in_4[22]);
  or g727 (n_540, in_2[22], in_4[22]);
  or g728 (n_541, in_2[22], in_3[22]);
  xnor g729 (n_282, n_538, in_2[22]);
  xnor g733 (n_283, n_281, n_280);
  or g734 (n_289, n_280, wc, n_281);
  not gc (wc, n_544);
  xnor g735 (n_550, n_287, n_143);
  or g736 (n_551, n_143, wc0);
  not gc0 (wc0, n_287);
  or g737 (n_552, wc1, n_143);
  not gc1 (wc1, n_289);
  or g738 (n_563, n_559, wc2);
  not gc2 (wc2, n_560);
  or g739 (n_782, wc3, n_559);
  not gc3 (wc3, n_562);
  and g740 (n_637, wc4, n_566);
  not gc4 (wc4, n_567);
  or g741 (n_783, wc5, n_569);
  not gc5 (wc5, n_564);
  or g742 (n_786, wc6, n_565);
  not gc6 (wc6, n_566);
  and g743 (n_639, wc7, n_572);
  not gc7 (wc7, n_573);
  or g744 (n_636, wc8, n_569);
  not gc8 (wc8, n_634);
  or g745 (n_787, wc9, n_575);
  not gc9 (wc9, n_570);
  or g746 (n_790, wc10, n_571);
  not gc10 (wc10, n_572);
  and g747 (n_646, wc11, n_578);
  not gc11 (wc11, n_579);
  and g748 (n_649, wc12, n_584);
  not gc12 (wc12, n_585);
  and g749 (n_656, wc13, n_590);
  not gc13 (wc13, n_591);
  and g750 (n_659, wc14, n_596);
  not gc14 (wc14, n_597);
  and g751 (n_666, wc15, n_602);
  not gc15 (wc15, n_603);
  and g752 (n_669, wc16, n_608);
  not gc16 (wc16, n_609);
  and g753 (n_676, wc17, n_614);
  not gc17 (wc17, n_615);
  and g754 (n_679, wc18, n_620);
  not gc18 (wc18, n_621);
  and g755 (n_686, wc19, n_626);
  not gc19 (wc19, n_627);
  or g756 (n_693, wc20, n_581);
  not gc20 (wc20, n_642);
  or g757 (n_735, wc21, n_593);
  not gc21 (wc21, n_652);
  or g758 (n_708, wc22, n_605);
  not gc22 (wc22, n_662);
  or g759 (n_762, wc23, n_617);
  not gc23 (wc23, n_672);
  or g760 (n_723, wc24, n_629);
  not gc24 (wc24, n_682);
  or g761 (n_792, wc25, n_581);
  not gc25 (wc25, n_576);
  or g762 (n_795, wc26, n_577);
  not gc26 (wc26, n_578);
  or g763 (n_796, wc27, n_587);
  not gc27 (wc27, n_582);
  or g764 (n_799, wc28, n_583);
  not gc28 (wc28, n_584);
  or g765 (n_801, wc29, n_593);
  not gc29 (wc29, n_588);
  or g766 (n_804, wc30, n_589);
  not gc30 (wc30, n_590);
  or g767 (n_807, wc31, n_599);
  not gc31 (wc31, n_594);
  or g768 (n_810, wc32, n_595);
  not gc32 (wc32, n_596);
  or g769 (n_812, wc33, n_605);
  not gc33 (wc33, n_600);
  or g770 (n_815, wc34, n_601);
  not gc34 (wc34, n_602);
  or g771 (n_816, wc35, n_611);
  not gc35 (wc35, n_606);
  or g772 (n_819, wc36, n_607);
  not gc36 (wc36, n_608);
  or g773 (n_821, wc37, n_617);
  not gc37 (wc37, n_612);
  or g774 (n_824, wc38, n_613);
  not gc38 (wc38, n_614);
  or g775 (n_827, wc39, n_623);
  not gc39 (wc39, n_618);
  or g776 (n_830, wc40, n_619);
  not gc40 (wc40, n_620);
  or g777 (n_832, wc41, n_629);
  not gc41 (wc41, n_624);
  or g778 (n_835, wc42, n_625);
  not gc42 (wc42, n_626);
  or g779 (n_837, wc43, n_633);
  not gc43 (wc43, n_630);
  and g780 (n_695, wc44, n_576);
  not gc44 (wc44, n_640);
  and g781 (n_647, wc45, n_644);
  not gc45 (wc45, n_639);
  and g782 (n_657, wc46, n_654);
  not gc46 (wc46, n_649);
  and g783 (n_667, wc47, n_664);
  not gc47 (wc47, n_659);
  and g784 (n_677, wc48, n_674);
  not gc48 (wc48, n_669);
  and g785 (n_687, wc49, n_684);
  not gc49 (wc49, n_679);
  or g786 (n_691, wc50, n_575);
  not gc50 (wc50, n_689);
  and g787 (n_744, wc51, n_662);
  not gc51 (wc51, n_704);
  and g788 (n_771, wc52, n_682);
  not gc52 (wc52, n_719);
  and g789 (n_699, wc53, n_646);
  not gc53 (wc53, n_647);
  and g790 (n_737, wc54, n_588);
  not gc54 (wc54, n_650);
  and g791 (n_701, wc55, n_656);
  not gc55 (wc55, n_657);
  and g792 (n_709, wc56, n_600);
  not gc56 (wc56, n_660);
  and g793 (n_713, wc57, n_666);
  not gc57 (wc57, n_667);
  and g794 (n_764, wc58, n_612);
  not gc58 (wc58, n_670);
  and g795 (n_716, wc59, n_676);
  not gc59 (wc59, n_677);
  and g796 (n_724, wc60, n_624);
  not gc60 (wc60, n_680);
  and g797 (n_728, wc61, n_686);
  not gc61 (wc61, n_687);
  or g798 (n_696, n_693, wc62);
  not gc62 (wc62, n_689);
  or g799 (n_700, n_697, wc63);
  not gc63 (wc63, n_689);
  or g800 (n_778, wc64, n_633);
  not gc64 (wc64, n_756);
  and g801 (n_706, wc65, n_662);
  not gc65 (wc65, n_701);
  and g802 (n_721, wc66, n_682);
  not gc66 (wc66, n_716);
  and g803 (n_742, wc67, n_594);
  not gc67 (wc67, n_702);
  and g804 (n_745, wc68, n_659);
  not gc68 (wc68, n_706);
  and g805 (n_748, n_709, wc69);
  not gc69 (wc69, n_710);
  and g806 (n_751, n_713, wc70);
  not gc70 (wc70, n_714);
  and g807 (n_769, wc71, n_618);
  not gc71 (wc71, n_717);
  and g808 (n_772, wc72, n_679);
  not gc72 (wc72, n_721);
  and g809 (n_775, n_724, wc73);
  not gc73 (wc73, n_725);
  and g810 (n_753, n_728, wc74);
  not gc74 (wc74, n_729);
  or g811 (n_733, wc75, n_587);
  not gc75 (wc75, n_731);
  or g812 (n_738, n_735, wc76);
  not gc76 (wc76, n_731);
  or g813 (n_740, wc77, n_704);
  not gc77 (wc77, n_731);
  and g814 (n_780, wc78, n_630);
  not gc78 (wc78, n_754);
  or g815 (n_760, wc79, n_611);
  not gc79 (wc79, n_758);
  or g816 (n_765, n_762, wc80);
  not gc80 (wc80, n_758);
  or g817 (n_767, wc81, n_719);
  not gc81 (wc81, n_758);
  or g818 (n_781, n_778, wc82);
  not gc82 (wc82, n_758);
  not g819 (out_0[25], n_839);
endmodule

module csa_tree_add_897_44_group_6805_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  csa_tree_add_897_44_group_6805_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module mult_signed_const_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_67;
  wire n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_174;
  wire n_181, n_182, n_184, n_185, n_186, n_190, n_191, n_197;
  wire n_198, n_204, n_205, n_206, n_210, n_211, n_212, n_213;
  wire n_214, n_218, n_220, n_221, n_226, n_227, n_228, n_229;
  wire n_237, n_238, n_239, n_240, n_241, n_247, n_248, n_249;
  wire n_250, n_251, n_252, n_253, n_259, n_260, n_261, n_262;
  wire n_263, n_271, n_273, n_274, n_275, n_276, n_277, n_278;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_327, n_335, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_358, n_359, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_372, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_391, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_450, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_469, n_471, n_472, n_473, n_474, n_475, n_476, n_477;
  wire n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485;
  wire n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_516, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_531, n_533, n_534, n_535, n_536, n_537, n_538, n_539;
  wire n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_555;
  wire n_558, n_560, n_561, n_562, n_563, n_564, n_565, n_566;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_577;
  wire n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586;
  wire n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_596;
  wire n_597, n_598, n_599, n_600, n_604, n_605, n_606, n_607;
  wire n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_618;
  wire n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630;
  wire n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638;
  wire n_639, n_640, n_641, n_642, n_647, n_648, n_649, n_650;
  wire n_651, n_652, n_653, n_654, n_655, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_666, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_678, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_694, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_719;
  wire n_720, n_721, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_767, n_768, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_793, n_794, n_795;
  wire n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803;
  wire n_804, n_805, n_806, n_817, n_821, n_823, n_824, n_825;
  wire n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833;
  wire n_834, n_843, n_844, n_845, n_846, n_847, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_917, n_918, n_919;
  wire n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_927;
  wire n_928, n_929, n_930, n_945, n_946, n_947, n_948, n_950;
  wire n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958;
  wire n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966;
  wire n_975, n_979, n_980, n_981, n_982, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1019;
  wire n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027;
  wire n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035;
  wire n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1044;
  wire n_1045, n_1048, n_1050, n_1052, n_1053, n_1057, n_1058, n_1059;
  wire n_1064, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072;
  wire n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080;
  wire n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1089;
  wire n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098;
  wire n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106;
  wire n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114;
  wire n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122;
  wire n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130;
  wire n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138;
  wire n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1146, n_1147;
  wire n_1148, n_1149, n_1150, n_1153, n_1154, n_1155, n_1156, n_1157;
  wire n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165;
  wire n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173;
  wire n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181;
  wire n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190;
  wire n_1191, n_1192, n_1194, n_1195, n_1196, n_1197, n_1198, n_1201;
  wire n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209;
  wire n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217;
  wire n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225;
  wire n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233;
  wire n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241;
  wire n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249;
  wire n_1250, n_1251, n_1252, n_1253, n_1254, n_1257, n_1258, n_1259;
  wire n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1269;
  wire n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
  wire n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285;
  wire n_1286, n_1287, n_1289, n_1291, n_1292, n_1293, n_1294, n_1295;
  wire n_1296, n_1297, n_1298, n_1301, n_1302, n_1303, n_1304, n_1305;
  wire n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313;
  wire n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321;
  wire n_1322, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331;
  wire n_1335, n_1336, n_1337, n_1338, n_1339, n_1341, n_1342, n_1343;
  wire n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351;
  wire n_1352, n_1353, n_1354, n_1356, n_1357, n_1358, n_1359, n_1362;
  wire n_1363, n_1364, n_1365, n_1366, n_1367, n_1369, n_1370, n_1371;
  wire n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379;
  wire n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387;
  wire n_1389, n_1390, n_1391, n_1392, n_1394, n_1395, n_1396, n_1397;
  wire n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405;
  wire n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1415, n_1416;
  wire n_1417, n_1418, n_1419, n_1421, n_1422, n_1425, n_1426, n_1427;
  wire n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435;
  wire n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1445;
  wire n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453;
  wire n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461;
  wire n_1462, n_1464, n_1465, n_1467, n_1468, n_1470, n_1471, n_1472;
  wire n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480;
  wire n_1481, n_1482, n_1486, n_1489, n_1490, n_1491, n_1492, n_1493;
  wire n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501;
  wire n_1502, n_1505, n_1507, n_1508, n_1509, n_1511, n_1513, n_1514;
  wire n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522;
  wire n_1525, n_1526, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534;
  wire n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1543;
  wire n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1552;
  wire n_1553, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561;
  wire n_1562, n_1563, n_1566, n_1568, n_1569, n_1570, n_1571, n_1572;
  wire n_1573, n_1574, n_1575, n_1579, n_1580, n_1581, n_1582, n_1584;
  wire n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592;
  wire n_1593, n_1594, n_1605, n_1606, n_1607, n_1608, n_1610, n_1611;
  wire n_1612, n_1613, n_1614, n_1616, n_1617, n_1618, n_1619, n_1620;
  wire n_1622, n_1623, n_1624, n_1625, n_1626, n_1628, n_1629, n_1630;
  wire n_1631, n_1632, n_1634, n_1635, n_1636, n_1637, n_1638, n_1640;
  wire n_1641, n_1642, n_1643, n_1644, n_1646, n_1647, n_1648, n_1649;
  wire n_1650, n_1652, n_1653, n_1654, n_1655, n_1656, n_1658, n_1659;
  wire n_1660, n_1661, n_1662, n_1664, n_1665, n_1666, n_1667, n_1668;
  wire n_1670, n_1671, n_1672, n_1673, n_1674, n_1676, n_1677, n_1678;
  wire n_1679, n_1680, n_1682, n_1683, n_1684, n_1685, n_1686, n_1688;
  wire n_1689, n_1690, n_1691, n_1692, n_1694, n_1695, n_1696, n_1697;
  wire n_1698, n_1700, n_1701, n_1702, n_1703, n_1704, n_1706, n_1707;
  wire n_1708, n_1709, n_1710, n_1712, n_1713, n_1714, n_1715, n_1716;
  wire n_1718, n_1719, n_1720, n_1721, n_1722, n_1724, n_1725, n_1726;
  wire n_1727, n_1728, n_1730, n_1731, n_1732, n_1733, n_1734, n_1736;
  wire n_1737, n_1738, n_1739, n_1740, n_1745, n_1747, n_1748, n_1750;
  wire n_1752, n_1754, n_1755, n_1757, n_1758, n_1760, n_1762, n_1764;
  wire n_1765, n_1767, n_1768, n_1770, n_1772, n_1774, n_1775, n_1777;
  wire n_1778, n_1780, n_1782, n_1784, n_1785, n_1787, n_1788, n_1790;
  wire n_1792, n_1794, n_1795, n_1797, n_1798, n_1800, n_1802, n_1804;
  wire n_1805, n_1807, n_1808, n_1810, n_1812, n_1814, n_1815, n_1817;
  wire n_1818, n_1820, n_1822, n_1824, n_1825, n_1827, n_1828, n_1830;
  wire n_1832, n_1834, n_1835, n_1837, n_1838, n_1840, n_1842, n_1844;
  wire n_1845, n_1847, n_1848, n_1850, n_1854, n_1855, n_1856, n_1858;
  wire n_1859, n_1860, n_1862, n_1863, n_1864, n_1865, n_1867, n_1869;
  wire n_1871, n_1872, n_1873, n_1875, n_1876, n_1877, n_1879, n_1880;
  wire n_1882, n_1884, n_1886, n_1887, n_1888, n_1890, n_1891, n_1892;
  wire n_1894, n_1895, n_1897, n_1899, n_1901, n_1902, n_1903, n_1905;
  wire n_1906, n_1907, n_1909, n_1910, n_1912, n_1914, n_1916, n_1917;
  wire n_1918, n_1920, n_1921, n_1922, n_1924, n_1925, n_1927, n_1929;
  wire n_1931, n_1932, n_1933, n_1935, n_1937, n_1938, n_1939, n_1941;
  wire n_1942, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950;
  wire n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958;
  wire n_1960, n_1963, n_1965, n_1966, n_1967, n_1970, n_1973, n_1975;
  wire n_1976, n_1978, n_1980, n_1981, n_1983, n_1985, n_1986, n_1988;
  wire n_1990, n_1991, n_1993, n_1994, n_1996, n_1999, n_2001, n_2002;
  wire n_2003, n_2006, n_2009, n_2011, n_2012, n_2014, n_2016, n_2017;
  wire n_2019, n_2021, n_2022, n_2024, n_2026, n_2027, n_2028, n_2030;
  wire n_2031, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039;
  wire n_2040, n_2041, n_2042, n_2043, n_2044, n_2046, n_2047, n_2048;
  wire n_2050, n_2051, n_2052, n_2054, n_2055, n_2056, n_2058, n_2059;
  wire n_2060, n_2062, n_2063, n_2064, n_2066, n_2067, n_2068, n_2070;
  wire n_2071, n_2072, n_2074, n_2075, n_2076, n_2078, n_2079, n_2080;
  wire n_2082, n_2083, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090;
  wire n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2098, n_2099;
  wire n_2100, n_2102, n_2103, n_2104, n_2106, n_2107, n_2108, n_2110;
  wire n_2111, n_2112, n_2114, n_2115, n_2116, n_2118, n_2119, n_2120;
  wire n_2122, n_2123, n_2125, n_2128, n_2129, n_2131, n_2132, n_2133;
  wire n_2134, n_2136, n_2137, n_2138, n_2140, n_2141, n_2142, n_2143;
  wire n_2145, n_2146, n_2148, n_2149, n_2151, n_2152, n_2153, n_2154;
  wire n_2156, n_2157, n_2158, n_2160, n_2161, n_2162, n_2163, n_2165;
  wire n_2166, n_2168, n_2169, n_2171, n_2172, n_2173, n_2174, n_2176;
  wire n_2177, n_2178, n_2179, n_2181, n_2182, n_2183, n_2184, n_2186;
  wire n_2187, n_2189, n_2190, n_2192, n_2193, n_2194, n_2195, n_2197;
  wire n_2198, n_2199, n_2201, n_2202, n_2203, n_2204, n_2206, n_2207;
  wire n_2209, n_2210, n_2212, n_2213, n_2214, n_2215, n_2217, n_2218;
  wire n_2219, n_2220, n_2222, n_2223, n_2224, n_2225, n_2227, n_2228;
  wire n_2230, n_2231, n_2233, n_2234, n_2235, n_2236, n_2238, n_2239;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_70, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_623, A[1], n_171);
  xor g270 (n_69, n_623, A[2]);
  nand g3 (n_624, A[1], n_171);
  nand g271 (n_625, A[2], n_171);
  nand g272 (n_626, A[1], A[2]);
  nand g273 (n_172, n_624, n_625, n_626);
  xor g274 (n_627, A[2], n_172);
  xor g275 (n_116, n_627, A[3]);
  nand g276 (n_628, A[2], n_172);
  nand g4 (n_629, A[3], n_172);
  nand g277 (n_630, A[2], A[3]);
  nand g278 (n_174, n_628, n_629, n_630);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_71, A[0], A[3]);
  xor g281 (n_631, A[4], n_173);
  xor g282 (n_115, n_631, n_174);
  nand g283 (n_632, A[4], n_173);
  nand g284 (n_633, n_174, n_173);
  nand g5 (n_634, A[4], n_174);
  nand g6 (n_73, n_632, n_633, n_634);
  xor g287 (n_635, n_70, A[4]);
  xor g288 (n_72, n_635, n_71);
  nand g289 (n_636, n_70, A[4]);
  nand g290 (n_637, n_71, A[4]);
  nand g291 (n_638, n_70, n_71);
  nand g292 (n_181, n_636, n_637, n_638);
  xor g293 (n_639, A[5], n_72);
  xor g294 (n_114, n_639, n_73);
  nand g295 (n_640, A[5], n_72);
  nand g296 (n_641, n_73, n_72);
  nand g297 (n_642, A[5], n_73);
  nand g298 (n_65, n_640, n_641, n_642);
  xor g305 (n_647, n_69, A[5]);
  xor g306 (n_182, n_647, A[6]);
  nand g307 (n_648, n_69, A[5]);
  nand g308 (n_649, A[6], A[5]);
  nand g309 (n_650, n_69, A[6]);
  nand g310 (n_185, n_648, n_649, n_650);
  xor g311 (n_651, n_181, n_182);
  xor g312 (n_113, n_651, A[8]);
  nand g313 (n_652, n_181, n_182);
  nand g314 (n_653, A[8], n_182);
  nand g315 (n_654, n_181, A[8]);
  nand g316 (n_64, n_652, n_653, n_654);
  xor g317 (n_655, A[2], A[3]);
  xor g318 (n_184, n_655, n_172);
  xor g323 (n_659, A[6], n_184);
  xor g324 (n_186, n_659, A[7]);
  nand g325 (n_660, A[6], n_184);
  nand g326 (n_661, A[7], n_184);
  nand g327 (n_662, A[6], A[7]);
  nand g328 (n_190, n_660, n_661, n_662);
  xor g329 (n_663, n_185, A[9]);
  xor g330 (n_112, n_663, n_186);
  nand g331 (n_664, n_185, A[9]);
  nand g332 (n_665, n_186, A[9]);
  nand g333 (n_666, n_185, n_186);
  nand g334 (n_63, n_664, n_665, n_666);
  xor g343 (n_671, A[7], n_115);
  xor g344 (n_191, n_671, A[8]);
  nand g345 (n_672, A[7], n_115);
  nand g346 (n_673, A[8], n_115);
  nand g347 (n_674, A[7], A[8]);
  nand g348 (n_197, n_672, n_673, n_674);
  xor g349 (n_675, A[10], n_190);
  xor g350 (n_111, n_675, n_191);
  nand g351 (n_676, A[10], n_190);
  nand g352 (n_677, n_191, n_190);
  nand g353 (n_678, A[10], n_191);
  nand g354 (n_62, n_676, n_677, n_678);
  xor g369 (n_687, A[8], A[9]);
  xor g370 (n_198, n_687, n_114);
  nand g371 (n_688, A[8], A[9]);
  nand g372 (n_689, n_114, A[9]);
  nand g373 (n_690, A[8], n_114);
  nand g374 (n_205, n_688, n_689, n_690);
  xor g375 (n_691, A[11], n_197);
  xor g376 (n_110, n_691, n_198);
  nand g377 (n_692, A[11], n_197);
  nand g378 (n_693, n_198, n_197);
  nand g379 (n_694, A[11], n_198);
  nand g380 (n_61, n_692, n_693, n_694);
  xor g394 (n_204, n_651, A[9]);
  nand g396 (n_705, A[9], n_182);
  nand g397 (n_706, n_181, A[9]);
  nand g398 (n_211, n_652, n_705, n_706);
  xor g399 (n_707, A[10], n_65);
  xor g400 (n_206, n_707, A[12]);
  nand g401 (n_708, A[10], n_65);
  nand g402 (n_709, A[12], n_65);
  nand g403 (n_710, A[10], A[12]);
  nand g404 (n_212, n_708, n_709, n_710);
  xor g405 (n_711, n_204, n_205);
  xor g406 (n_109, n_711, n_206);
  nand g407 (n_712, n_204, n_205);
  nand g408 (n_713, n_206, n_205);
  nand g409 (n_714, n_204, n_206);
  nand g410 (n_60, n_712, n_713, n_714);
  xor g417 (n_719, A[6], n_116);
  xor g418 (n_210, n_719, A[7]);
  nand g419 (n_720, A[6], n_116);
  nand g420 (n_721, A[7], n_116);
  nand g422 (n_218, n_720, n_721, n_662);
  xor g423 (n_723, n_185, A[10]);
  xor g424 (n_213, n_723, n_210);
  nand g425 (n_724, n_185, A[10]);
  nand g426 (n_725, n_210, A[10]);
  nand g427 (n_726, n_185, n_210);
  nand g428 (n_220, n_724, n_725, n_726);
  xor g429 (n_727, A[11], n_211);
  xor g430 (n_214, n_727, n_212);
  nand g431 (n_728, A[11], n_211);
  nand g432 (n_729, n_212, n_211);
  nand g433 (n_730, A[11], n_212);
  nand g434 (n_221, n_728, n_729, n_730);
  xor g435 (n_731, A[13], n_213);
  xor g436 (n_108, n_731, n_214);
  nand g437 (n_732, A[13], n_213);
  nand g438 (n_733, n_214, n_213);
  nand g439 (n_734, A[13], n_214);
  nand g440 (n_59, n_732, n_733, n_734);
  xor g455 (n_743, n_218, n_191);
  xor g456 (n_67, n_743, A[12]);
  nand g457 (n_744, n_218, n_191);
  nand g458 (n_745, A[12], n_191);
  nand g459 (n_746, n_218, A[12]);
  nand g460 (n_226, n_744, n_745, n_746);
  xor g461 (n_747, A[11], n_220);
  xor g462 (n_68, n_747, A[14]);
  nand g463 (n_748, A[11], n_220);
  nand g464 (n_749, A[14], n_220);
  nand g465 (n_750, A[11], A[14]);
  nand g466 (n_228, n_748, n_749, n_750);
  xor g467 (n_751, n_67, n_68);
  xor g468 (n_107, n_751, n_221);
  nand g469 (n_752, n_67, n_68);
  nand g470 (n_753, n_221, n_68);
  nand g471 (n_754, n_67, n_221);
  nand g472 (n_58, n_752, n_753, n_754);
  xor g493 (n_767, A[12], n_197);
  xor g494 (n_227, n_767, n_198);
  nand g495 (n_768, A[12], n_197);
  nand g497 (n_770, A[12], n_198);
  nand g498 (n_238, n_768, n_693, n_770);
  xor g499 (n_771, A[13], n_226);
  xor g500 (n_229, n_771, A[15]);
  nand g501 (n_772, A[13], n_226);
  nand g502 (n_773, A[15], n_226);
  nand g503 (n_774, A[13], A[15]);
  nand g504 (n_240, n_772, n_773, n_774);
  xor g505 (n_775, n_227, n_228);
  xor g506 (n_106, n_775, n_229);
  nand g507 (n_776, n_227, n_228);
  nand g508 (n_777, n_229, n_228);
  nand g509 (n_778, n_227, n_229);
  nand g510 (n_57, n_776, n_777, n_778);
  xor g530 (n_237, n_707, n_204);
  nand g532 (n_793, n_204, n_65);
  nand g533 (n_794, A[10], n_204);
  nand g534 (n_248, n_708, n_793, n_794);
  xor g535 (n_795, n_205, A[13]);
  xor g536 (n_239, n_795, A[14]);
  nand g537 (n_796, n_205, A[13]);
  nand g538 (n_797, A[14], A[13]);
  nand g539 (n_798, n_205, A[14]);
  nand g540 (n_250, n_796, n_797, n_798);
  xor g541 (n_799, n_237, n_238);
  xor g542 (n_241, n_799, A[16]);
  nand g543 (n_800, n_237, n_238);
  nand g544 (n_801, A[16], n_238);
  nand g545 (n_802, n_237, A[16]);
  nand g546 (n_252, n_800, n_801, n_802);
  xor g547 (n_803, n_239, n_240);
  xor g548 (n_105, n_803, n_241);
  nand g549 (n_804, n_239, n_240);
  nand g550 (n_805, n_241, n_240);
  nand g551 (n_806, n_239, n_241);
  nand g552 (n_56, n_804, n_805, n_806);
  xor g566 (n_247, n_723, n_186);
  nand g568 (n_817, n_186, A[10]);
  nand g570 (n_259, n_724, n_817, n_666);
  xor g572 (n_249, n_727, A[14]);
  nand g574 (n_821, A[14], n_211);
  nand g576 (n_261, n_728, n_821, n_750);
  xor g577 (n_823, n_247, A[15]);
  xor g578 (n_251, n_823, n_248);
  nand g579 (n_824, n_247, A[15]);
  nand g580 (n_825, n_248, A[15]);
  nand g581 (n_826, n_247, n_248);
  nand g582 (n_117, n_824, n_825, n_826);
  xor g583 (n_827, n_249, A[17]);
  xor g584 (n_253, n_827, n_250);
  nand g585 (n_828, n_249, A[17]);
  nand g586 (n_829, n_250, A[17]);
  nand g587 (n_830, n_249, n_250);
  nand g588 (n_119, n_828, n_829, n_830);
  xor g589 (n_831, n_251, n_252);
  xor g590 (n_104, n_831, n_253);
  nand g591 (n_832, n_251, n_252);
  nand g592 (n_833, n_253, n_252);
  nand g593 (n_834, n_251, n_253);
  nand g594 (n_55, n_832, n_833, n_834);
  xor g609 (n_843, n_190, A[11]);
  xor g610 (n_260, n_843, A[12]);
  nand g611 (n_844, n_190, A[11]);
  nand g612 (n_845, A[12], A[11]);
  nand g613 (n_846, n_190, A[12]);
  nand g614 (n_271, n_844, n_845, n_846);
  xor g615 (n_847, n_191, n_259);
  xor g616 (n_118, n_847, n_260);
  nand g617 (n_848, n_191, n_259);
  nand g618 (n_849, n_260, n_259);
  nand g619 (n_850, n_191, n_260);
  nand g620 (n_273, n_848, n_849, n_850);
  xor g621 (n_851, A[15], A[16]);
  xor g622 (n_262, n_851, n_261);
  nand g623 (n_852, A[15], A[16]);
  nand g624 (n_853, n_261, A[16]);
  nand g625 (n_854, A[15], n_261);
  nand g626 (n_275, n_852, n_853, n_854);
  xor g627 (n_855, A[18], n_117);
  xor g628 (n_263, n_855, n_118);
  nand g629 (n_856, A[18], n_117);
  nand g630 (n_857, n_118, n_117);
  nand g631 (n_858, A[18], n_118);
  nand g632 (n_277, n_856, n_857, n_858);
  xor g633 (n_859, n_119, n_262);
  xor g634 (n_103, n_859, n_263);
  nand g635 (n_860, n_119, n_262);
  nand g636 (n_861, n_263, n_262);
  nand g637 (n_862, n_119, n_263);
  nand g638 (n_54, n_860, n_861, n_862);
  xor g665 (n_879, A[13], n_271);
  xor g666 (n_274, n_879, A[16]);
  nand g667 (n_880, A[13], n_271);
  nand g668 (n_881, A[16], n_271);
  nand g669 (n_882, A[13], A[16]);
  nand g670 (n_289, n_880, n_881, n_882);
  xor g671 (n_883, n_227, A[17]);
  xor g672 (n_276, n_883, A[19]);
  nand g673 (n_884, n_227, A[17]);
  nand g674 (n_885, A[19], A[17]);
  nand g675 (n_886, n_227, A[19]);
  nand g676 (n_291, n_884, n_885, n_886);
  xor g677 (n_887, n_273, n_274);
  xor g678 (n_278, n_887, n_275);
  nand g679 (n_888, n_273, n_274);
  nand g680 (n_889, n_275, n_274);
  nand g681 (n_890, n_273, n_275);
  nand g682 (n_293, n_888, n_889, n_890);
  xor g683 (n_891, n_276, n_277);
  xor g684 (n_102, n_891, n_278);
  nand g685 (n_892, n_276, n_277);
  nand g686 (n_893, n_278, n_277);
  nand g687 (n_894, n_276, n_278);
  nand g688 (n_53, n_892, n_893, n_894);
  xor g720 (n_290, n_799, A[17]);
  nand g722 (n_917, A[17], n_238);
  nand g723 (n_918, n_237, A[17]);
  nand g724 (n_305, n_800, n_917, n_918);
  xor g725 (n_919, A[18], n_239);
  xor g726 (n_292, n_919, n_289);
  nand g727 (n_920, A[18], n_239);
  nand g728 (n_921, n_289, n_239);
  nand g729 (n_922, A[18], n_289);
  nand g730 (n_307, n_920, n_921, n_922);
  xor g731 (n_923, A[20], n_290);
  xor g732 (n_294, n_923, n_291);
  nand g733 (n_924, A[20], n_290);
  nand g734 (n_925, n_291, n_290);
  nand g735 (n_926, A[20], n_291);
  nand g736 (n_309, n_924, n_925, n_926);
  xor g737 (n_927, n_292, n_293);
  xor g738 (n_101, n_927, n_294);
  nand g739 (n_928, n_292, n_293);
  nand g740 (n_929, n_294, n_293);
  nand g741 (n_930, n_292, n_294);
  nand g742 (n_52, n_928, n_929, n_930);
  xor g762 (n_303, n_727, n_247);
  nand g764 (n_945, n_247, n_211);
  nand g765 (n_946, A[11], n_247);
  nand g766 (n_318, n_728, n_945, n_946);
  xor g767 (n_947, A[14], n_248);
  xor g768 (n_304, n_947, A[15]);
  nand g769 (n_948, A[14], n_248);
  nand g771 (n_950, A[14], A[15]);
  nand g772 (n_319, n_948, n_825, n_950);
  xor g773 (n_951, n_250, n_303);
  xor g774 (n_306, n_951, A[19]);
  nand g775 (n_952, n_250, n_303);
  nand g776 (n_953, A[19], n_303);
  nand g777 (n_954, n_250, A[19]);
  nand g778 (n_322, n_952, n_953, n_954);
  xor g779 (n_955, A[18], A[21]);
  xor g780 (n_308, n_955, n_304);
  nand g781 (n_956, A[18], A[21]);
  nand g782 (n_957, n_304, A[21]);
  nand g783 (n_958, A[18], n_304);
  nand g784 (n_324, n_956, n_957, n_958);
  xor g785 (n_959, n_305, n_306);
  xor g786 (n_310, n_959, n_307);
  nand g787 (n_960, n_305, n_306);
  nand g788 (n_961, n_307, n_306);
  nand g789 (n_962, n_305, n_307);
  nand g790 (n_326, n_960, n_961, n_962);
  xor g791 (n_963, n_308, n_309);
  xor g792 (n_100, n_963, n_310);
  nand g793 (n_964, n_308, n_309);
  nand g794 (n_965, n_310, n_309);
  nand g795 (n_966, n_308, n_310);
  nand g796 (n_51, n_964, n_965, n_966);
  xor g811 (n_975, n_190, A[12]);
  xor g812 (n_317, n_975, n_191);
  nand g816 (n_335, n_846, n_745, n_677);
  xor g817 (n_979, A[11], n_259);
  xor g818 (n_320, n_979, n_317);
  nand g819 (n_980, A[11], n_259);
  nand g820 (n_981, n_317, n_259);
  nand g821 (n_982, A[11], n_317);
  nand g822 (n_337, n_980, n_981, n_982);
  xor g824 (n_321, n_851, n_318);
  nand g826 (n_985, n_318, A[16]);
  nand g827 (n_986, A[15], n_318);
  nand g828 (n_339, n_852, n_985, n_986);
  xor g829 (n_987, n_319, A[19]);
  xor g830 (n_323, n_987, n_320);
  nand g831 (n_988, n_319, A[19]);
  nand g832 (n_989, n_320, A[19]);
  nand g833 (n_990, n_319, n_320);
  nand g834 (n_340, n_988, n_989, n_990);
  xor g835 (n_991, A[20], A[22]);
  xor g836 (n_325, n_991, n_321);
  nand g837 (n_992, A[20], A[22]);
  nand g838 (n_993, n_321, A[22]);
  nand g839 (n_994, A[20], n_321);
  nand g840 (n_343, n_992, n_993, n_994);
  xor g841 (n_995, n_322, n_323);
  xor g842 (n_327, n_995, n_324);
  nand g843 (n_996, n_322, n_323);
  nand g844 (n_997, n_324, n_323);
  nand g845 (n_998, n_322, n_324);
  nand g846 (n_345, n_996, n_997, n_998);
  xor g847 (n_999, n_325, n_326);
  xor g848 (n_99, n_999, n_327);
  nand g849 (n_1000, n_325, n_326);
  nand g850 (n_1001, n_327, n_326);
  nand g851 (n_1002, n_325, n_327);
  nand g852 (n_50, n_1000, n_1001, n_1002);
  xor g879 (n_1019, n_335, A[13]);
  xor g880 (n_338, n_1019, n_227);
  nand g881 (n_1020, n_335, A[13]);
  nand g882 (n_1021, n_227, A[13]);
  nand g883 (n_1022, n_335, n_227);
  nand g884 (n_359, n_1020, n_1021, n_1022);
  xor g885 (n_1023, A[16], A[17]);
  xor g886 (n_341, n_1023, n_337);
  nand g887 (n_1024, A[16], A[17]);
  nand g888 (n_1025, n_337, A[17]);
  nand g889 (n_1026, A[16], n_337);
  nand g890 (n_361, n_1024, n_1025, n_1026);
  xor g891 (n_1027, A[21], A[20]);
  xor g892 (n_342, n_1027, n_338);
  nand g893 (n_1028, A[21], A[20]);
  nand g894 (n_1029, n_338, A[20]);
  nand g895 (n_1030, A[21], n_338);
  nand g896 (n_362, n_1028, n_1029, n_1030);
  xor g897 (n_1031, A[23], n_339);
  xor g898 (n_344, n_1031, n_340);
  nand g899 (n_1032, A[23], n_339);
  nand g900 (n_1033, n_340, n_339);
  nand g901 (n_1034, A[23], n_340);
  nand g902 (n_365, n_1032, n_1033, n_1034);
  xor g903 (n_1035, n_341, n_342);
  xor g904 (n_346, n_1035, n_343);
  nand g905 (n_1036, n_341, n_342);
  nand g906 (n_1037, n_343, n_342);
  nand g907 (n_1038, n_341, n_343);
  nand g908 (n_367, n_1036, n_1037, n_1038);
  xor g909 (n_1039, n_344, n_345);
  xor g910 (n_98, n_1039, n_346);
  nand g911 (n_1040, n_344, n_345);
  nand g912 (n_1041, n_346, n_345);
  nand g913 (n_1042, n_344, n_346);
  nand g914 (n_49, n_1040, n_1041, n_1042);
  nand g922 (n_372, n_1044, n_1045, n_625);
  nand g928 (n_374, n_1048, n_649, n_1050);
  nand g934 (n_376, n_1052, n_1053, n_706);
  nand g940 (n_378, n_708, n_1057, n_1058);
  xor g941 (n_1059, n_205, A[14]);
  xor g942 (n_358, n_1059, A[13]);
  nand g952 (n_383, n_1064, n_917, n_1066);
  xor g953 (n_1067, A[18], n_358);
  nand g955 (n_1068, A[18], n_358);
  nand g958 (n_385, n_1068, n_1069, n_1070);
  xor g959 (n_1071, n_359, A[21]);
  xor g960 (n_364, n_1071, A[22]);
  nand g961 (n_1072, n_359, A[21]);
  nand g962 (n_1073, A[22], A[21]);
  nand g963 (n_1074, n_359, A[22]);
  nand g964 (n_386, n_1072, n_1073, n_1074);
  xor g966 (n_366, n_1075, n_362);
  nand g968 (n_1077, n_362, n_361);
  nand g970 (n_388, n_1076, n_1077, n_1078);
  xor g971 (n_1079, n_363, n_364);
  xor g972 (n_368, n_1079, n_365);
  nand g973 (n_1080, n_363, n_364);
  nand g974 (n_1081, n_365, n_364);
  nand g975 (n_1082, n_363, n_365);
  nand g976 (n_390, n_1080, n_1081, n_1082);
  xor g977 (n_1083, n_366, n_367);
  xor g978 (n_97, n_1083, n_368);
  nand g979 (n_1084, n_366, n_367);
  nand g980 (n_1085, n_368, n_367);
  nand g981 (n_1086, n_366, n_368);
  nand g982 (n_48, n_1084, n_1085, n_1086);
  xor g986 (n_373, n_1087, A[3]);
  nand g990 (n_393, n_1045, n_1089, n_630);
  xor g991 (n_1091, n_372, n_373);
  xor g992 (n_375, n_1091, A[6]);
  nand g993 (n_1092, n_372, n_373);
  nand g994 (n_1093, A[6], n_373);
  nand g995 (n_1094, n_372, A[6]);
  nand g996 (n_395, n_1092, n_1093, n_1094);
  xor g997 (n_1095, A[7], n_374);
  xor g998 (n_377, n_1095, n_375);
  nand g999 (n_1096, A[7], n_374);
  nand g1000 (n_1097, n_375, n_374);
  nand g1001 (n_1098, A[7], n_375);
  nand g1002 (n_397, n_1096, n_1097, n_1098);
  xor g1003 (n_1099, A[10], A[11]);
  xor g1004 (n_379, n_1099, n_376);
  nand g1005 (n_1100, A[10], A[11]);
  nand g1006 (n_1101, n_376, A[11]);
  nand g1007 (n_1102, A[10], n_376);
  nand g1008 (n_399, n_1100, n_1101, n_1102);
  xor g1009 (n_1103, n_377, A[14]);
  xor g1010 (n_381, n_1103, n_378);
  nand g1011 (n_1104, n_377, A[14]);
  nand g1012 (n_1105, n_378, A[14]);
  nand g1013 (n_1106, n_377, n_378);
  nand g1014 (n_401, n_1104, n_1105, n_1106);
  xor g1015 (n_1107, n_379, A[15]);
  xor g1016 (n_382, n_1107, n_250);
  nand g1017 (n_1108, n_379, A[15]);
  nand g1018 (n_1109, n_250, A[15]);
  nand g1019 (n_1110, n_379, n_250);
  nand g1020 (n_403, n_1108, n_1109, n_1110);
  xor g1021 (n_1111, A[19], A[18]);
  xor g1022 (n_384, n_1111, n_381);
  nand g1023 (n_1112, A[19], A[18]);
  nand g1024 (n_1113, n_381, A[18]);
  nand g1025 (n_1114, A[19], n_381);
  nand g1026 (n_404, n_1112, n_1113, n_1114);
  xor g1027 (n_1115, n_382, n_383);
  xor g1028 (n_387, n_1115, A[23]);
  nand g1029 (n_1116, n_382, n_383);
  nand g1030 (n_1117, A[23], n_383);
  nand g1031 (n_1118, n_382, A[23]);
  nand g1032 (n_407, n_1116, n_1117, n_1118);
  xor g1033 (n_1119, A[22], n_384);
  xor g1034 (n_389, n_1119, n_385);
  nand g1035 (n_1120, A[22], n_384);
  nand g1036 (n_1121, n_385, n_384);
  nand g1037 (n_1122, A[22], n_385);
  nand g1038 (n_409, n_1120, n_1121, n_1122);
  xor g1039 (n_1123, n_386, n_387);
  xor g1040 (n_391, n_1123, n_388);
  nand g1041 (n_1124, n_386, n_387);
  nand g1042 (n_1125, n_388, n_387);
  nand g1043 (n_1126, n_386, n_388);
  nand g1044 (n_412, n_1124, n_1125, n_1126);
  xor g1045 (n_1127, n_389, n_390);
  xor g1046 (n_96, n_1127, n_391);
  nand g1047 (n_1128, n_389, n_390);
  nand g1048 (n_1129, n_391, n_390);
  nand g1049 (n_1130, n_389, n_391);
  nand g1050 (n_47, n_1128, n_1129, n_1130);
  xor g1051 (n_1131, A[1], A[3]);
  xor g1052 (n_394, n_1131, A[4]);
  nand g1053 (n_1132, A[1], A[3]);
  nand g1054 (n_1133, A[4], A[3]);
  nand g1055 (n_1134, A[1], A[4]);
  nand g1056 (n_413, n_1132, n_1133, n_1134);
  xor g1057 (n_1135, n_393, n_394);
  xor g1058 (n_396, n_1135, A[7]);
  nand g1059 (n_1136, n_393, n_394);
  nand g1060 (n_1137, A[7], n_394);
  nand g1061 (n_1138, n_393, A[7]);
  nand g1062 (n_415, n_1136, n_1137, n_1138);
  xor g1063 (n_1139, A[8], n_395);
  xor g1064 (n_398, n_1139, n_396);
  nand g1065 (n_1140, A[8], n_395);
  nand g1066 (n_1141, n_396, n_395);
  nand g1067 (n_1142, A[8], n_396);
  nand g1068 (n_417, n_1140, n_1141, n_1142);
  xor g1069 (n_1143, n_397, A[11]);
  xor g1070 (n_400, n_1143, A[12]);
  nand g1071 (n_1144, n_397, A[11]);
  nand g1073 (n_1146, n_397, A[12]);
  nand g1074 (n_418, n_1144, n_845, n_1146);
  xor g1075 (n_1147, n_398, n_399);
  xor g1076 (n_402, n_1147, n_400);
  nand g1077 (n_1148, n_398, n_399);
  nand g1078 (n_1149, n_400, n_399);
  nand g1079 (n_1150, n_398, n_400);
  nand g1080 (n_420, n_1148, n_1149, n_1150);
  xor g1082 (n_405, n_851, A[19]);
  nand g1084 (n_1153, A[19], A[16]);
  nand g1085 (n_1154, A[15], A[19]);
  nand g1086 (n_423, n_852, n_1153, n_1154);
  xor g1088 (n_406, n_1155, A[20]);
  nand g1091 (n_1158, n_401, A[20]);
  nand g1092 (n_424, n_1156, n_1157, n_1158);
  xor g1093 (n_1159, n_402, n_403);
  xor g1094 (n_408, n_1159, A[23]);
  nand g1095 (n_1160, n_402, n_403);
  nand g1096 (n_1161, A[23], n_403);
  nand g1097 (n_1162, n_402, A[23]);
  nand g1098 (n_426, n_1160, n_1161, n_1162);
  xor g1099 (n_1163, n_404, n_405);
  xor g1100 (n_410, n_1163, n_406);
  nand g1101 (n_1164, n_404, n_405);
  nand g1102 (n_1165, n_406, n_405);
  nand g1103 (n_1166, n_404, n_406);
  nand g1104 (n_429, n_1164, n_1165, n_1166);
  xor g1105 (n_1167, n_407, n_408);
  xor g1106 (n_411, n_1167, n_409);
  nand g1107 (n_1168, n_407, n_408);
  nand g1108 (n_1169, n_409, n_408);
  nand g1109 (n_1170, n_407, n_409);
  nand g1110 (n_430, n_1168, n_1169, n_1170);
  xor g1111 (n_1171, n_410, n_411);
  xor g1112 (n_95, n_1171, n_412);
  nand g1113 (n_1172, n_410, n_411);
  nand g1114 (n_1173, n_412, n_411);
  nand g1115 (n_1174, n_410, n_412);
  nand g1116 (n_46, n_1172, n_1173, n_1174);
  xor g1117 (n_1175, A[4], A[5]);
  xor g1118 (n_414, n_1175, n_413);
  nand g1119 (n_1176, A[4], A[5]);
  nand g1120 (n_1177, n_413, A[5]);
  nand g1121 (n_1178, A[4], n_413);
  nand g1122 (n_434, n_1176, n_1177, n_1178);
  xor g1123 (n_1179, A[8], n_414);
  xor g1124 (n_416, n_1179, A[9]);
  nand g1125 (n_1180, A[8], n_414);
  nand g1126 (n_1181, A[9], n_414);
  nand g1128 (n_436, n_1180, n_1181, n_688);
  xor g1129 (n_1183, n_415, A[12]);
  xor g1130 (n_419, n_1183, n_416);
  nand g1131 (n_1184, n_415, A[12]);
  nand g1132 (n_1185, n_416, A[12]);
  nand g1133 (n_1186, n_415, n_416);
  nand g1134 (n_438, n_1184, n_1185, n_1186);
  xor g1135 (n_1187, n_417, A[13]);
  xor g1136 (n_421, n_1187, n_418);
  nand g1137 (n_1188, n_417, A[13]);
  nand g1138 (n_1189, n_418, A[13]);
  nand g1139 (n_1190, n_417, n_418);
  nand g1140 (n_439, n_1188, n_1189, n_1190);
  xor g1141 (n_1191, n_419, A[16]);
  xor g1142 (n_422, n_1191, A[17]);
  nand g1143 (n_1192, n_419, A[16]);
  nand g1145 (n_1194, n_419, A[17]);
  nand g1146 (n_442, n_1192, n_1024, n_1194);
  xor g1147 (n_1195, n_420, n_421);
  nand g1149 (n_1196, n_420, n_421);
  nand g1152 (n_444, n_1196, n_1197, n_1198);
  xor g1154 (n_427, n_1027, n_422);
  nand g1156 (n_1201, n_422, A[21]);
  nand g1157 (n_1202, A[20], n_422);
  nand g1158 (n_445, n_1028, n_1201, n_1202);
  xor g1159 (n_1203, n_423, n_424);
  xor g1160 (n_428, n_1203, n_425);
  nand g1161 (n_1204, n_423, n_424);
  nand g1162 (n_1205, n_425, n_424);
  nand g1163 (n_1206, n_423, n_425);
  nand g1164 (n_447, n_1204, n_1205, n_1206);
  xor g1165 (n_1207, n_426, n_427);
  xor g1166 (n_431, n_1207, n_428);
  nand g1167 (n_1208, n_426, n_427);
  nand g1168 (n_1209, n_428, n_427);
  nand g1169 (n_1210, n_426, n_428);
  nand g1170 (n_450, n_1208, n_1209, n_1210);
  xor g1171 (n_1211, n_429, n_430);
  xor g1172 (n_94, n_1211, n_431);
  nand g1173 (n_1212, n_429, n_430);
  nand g1174 (n_1213, n_431, n_430);
  nand g1175 (n_1214, n_429, n_431);
  nand g1176 (n_45, n_1212, n_1213, n_1214);
  xor g1180 (n_435, n_1215, n_434);
  nand g1183 (n_1218, A[6], n_434);
  nand g1184 (n_455, n_1216, n_1217, n_1218);
  xor g1185 (n_1219, A[9], A[10]);
  xor g1186 (n_437, n_1219, n_435);
  nand g1187 (n_1220, A[9], A[10]);
  nand g1188 (n_1221, n_435, A[10]);
  nand g1189 (n_1222, A[9], n_435);
  nand g1190 (n_456, n_1220, n_1221, n_1222);
  xor g1191 (n_1223, n_436, n_437);
  xor g1192 (n_440, n_1223, A[14]);
  nand g1193 (n_1224, n_436, n_437);
  nand g1194 (n_1225, A[14], n_437);
  nand g1195 (n_1226, n_436, A[14]);
  nand g1196 (n_458, n_1224, n_1225, n_1226);
  xor g1197 (n_1227, A[13], n_438);
  xor g1198 (n_441, n_1227, A[17]);
  nand g1199 (n_1228, A[13], n_438);
  nand g1200 (n_1229, A[17], n_438);
  nand g1201 (n_1230, A[13], A[17]);
  nand g1202 (n_461, n_1228, n_1229, n_1230);
  xor g1203 (n_1231, n_439, A[18]);
  xor g1204 (n_443, n_1231, n_440);
  nand g1205 (n_1232, n_439, A[18]);
  nand g1206 (n_1233, n_440, A[18]);
  nand g1207 (n_1234, n_439, n_440);
  nand g1208 (n_462, n_1232, n_1233, n_1234);
  xor g1209 (n_1235, A[21], n_441);
  xor g1210 (n_446, n_1235, n_442);
  nand g1211 (n_1236, A[21], n_441);
  nand g1212 (n_1237, n_442, n_441);
  nand g1213 (n_1238, A[21], n_442);
  nand g1214 (n_464, n_1236, n_1237, n_1238);
  xor g1215 (n_1239, A[22], n_443);
  xor g1216 (n_448, n_1239, n_444);
  nand g1217 (n_1240, A[22], n_443);
  nand g1218 (n_1241, n_444, n_443);
  nand g1219 (n_1242, A[22], n_444);
  nand g1220 (n_467, n_1240, n_1241, n_1242);
  xor g1221 (n_1243, n_445, n_446);
  xor g1222 (n_449, n_1243, n_447);
  nand g1223 (n_1244, n_445, n_446);
  nand g1224 (n_1245, n_447, n_446);
  nand g1225 (n_1246, n_445, n_447);
  nand g1226 (n_469, n_1244, n_1245, n_1246);
  xor g1227 (n_1247, n_448, n_449);
  xor g1228 (n_93, n_1247, n_450);
  nand g1229 (n_1248, n_448, n_449);
  nand g1230 (n_1249, n_450, n_449);
  nand g1231 (n_1250, n_448, n_450);
  nand g1232 (n_44, n_1248, n_1249, n_1250);
  xor g1235 (n_1251, A[5], A[7]);
  nand g1237 (n_1252, A[5], A[7]);
  nand g1240 (n_471, n_1252, n_1253, n_1254);
  xor g1242 (n_457, n_1099, n_454);
  nand g1244 (n_1257, n_454, A[11]);
  nand g1245 (n_1258, A[10], n_454);
  nand g1246 (n_473, n_1100, n_1257, n_1258);
  xor g1247 (n_1259, n_455, A[14]);
  xor g1248 (n_459, n_1259, n_456);
  nand g1249 (n_1260, n_455, A[14]);
  nand g1250 (n_1261, n_456, A[14]);
  nand g1251 (n_1262, n_455, n_456);
  nand g1252 (n_475, n_1260, n_1261, n_1262);
  xor g1253 (n_1263, n_457, A[15]);
  xor g1254 (n_460, n_1263, n_458);
  nand g1255 (n_1264, n_457, A[15]);
  nand g1256 (n_1265, n_458, A[15]);
  nand g1257 (n_1266, n_457, n_458);
  nand g1258 (n_477, n_1264, n_1265, n_1266);
  xor g1260 (n_463, n_1111, n_459);
  nand g1262 (n_1269, n_459, A[18]);
  nand g1263 (n_1270, A[19], n_459);
  nand g1264 (n_479, n_1112, n_1269, n_1270);
  xor g1265 (n_1271, n_460, n_461);
  xor g1266 (n_465, n_1271, A[22]);
  nand g1267 (n_1272, n_460, n_461);
  nand g1268 (n_1273, A[22], n_461);
  nand g1269 (n_1274, n_460, A[22]);
  nand g1270 (n_481, n_1272, n_1273, n_1274);
  xor g1271 (n_1275, A[23], n_462);
  xor g1272 (n_466, n_1275, n_463);
  nand g1273 (n_1276, A[23], n_462);
  nand g1274 (n_1277, n_463, n_462);
  nand g1275 (n_1278, A[23], n_463);
  nand g1276 (n_483, n_1276, n_1277, n_1278);
  xor g1277 (n_1279, n_464, n_465);
  xor g1278 (n_468, n_1279, n_466);
  nand g1279 (n_1280, n_464, n_465);
  nand g1280 (n_1281, n_466, n_465);
  nand g1281 (n_1282, n_464, n_466);
  nand g1282 (n_486, n_1280, n_1281, n_1282);
  xor g1283 (n_1283, n_467, n_468);
  xor g1284 (n_92, n_1283, n_469);
  nand g1285 (n_1284, n_467, n_468);
  nand g1286 (n_1285, n_469, n_468);
  nand g1287 (n_1286, n_467, n_469);
  nand g1288 (n_43, n_1284, n_1285, n_1286);
  xor g1289 (n_1287, A[7], A[6]);
  xor g1290 (n_472, n_1287, A[8]);
  nand g1292 (n_1289, A[8], A[6]);
  nand g1294 (n_487, n_662, n_1289, n_674);
  xor g1295 (n_1291, n_471, A[11]);
  xor g1296 (n_474, n_1291, n_472);
  nand g1297 (n_1292, n_471, A[11]);
  nand g1298 (n_1293, n_472, A[11]);
  nand g1299 (n_1294, n_471, n_472);
  nand g1300 (n_488, n_1292, n_1293, n_1294);
  xor g1301 (n_1295, A[12], n_473);
  xor g1302 (n_476, n_1295, n_474);
  nand g1303 (n_1296, A[12], n_473);
  nand g1304 (n_1297, n_474, n_473);
  nand g1305 (n_1298, A[12], n_474);
  nand g1306 (n_490, n_1296, n_1297, n_1298);
  xor g1308 (n_478, n_851, n_475);
  nand g1310 (n_1301, n_475, A[16]);
  nand g1311 (n_1302, A[15], n_475);
  nand g1312 (n_492, n_852, n_1301, n_1302);
  xor g1313 (n_1303, A[19], n_476);
  nand g1315 (n_1304, A[19], n_476);
  nand g1318 (n_495, n_1304, n_1305, n_1306);
  xor g1319 (n_1307, A[20], n_477);
  xor g1320 (n_482, n_1307, A[23]);
  nand g1321 (n_1308, A[20], n_477);
  nand g1322 (n_1309, A[23], n_477);
  nand g1323 (n_1310, A[20], A[23]);
  nand g1324 (n_497, n_1308, n_1309, n_1310);
  xor g1325 (n_1311, n_478, n_479);
  xor g1326 (n_484, n_1311, n_480);
  nand g1327 (n_1312, n_478, n_479);
  nand g1328 (n_1313, n_480, n_479);
  nand g1329 (n_1314, n_478, n_480);
  nand g1330 (n_498, n_1312, n_1313, n_1314);
  xor g1331 (n_1315, n_481, n_482);
  xor g1332 (n_485, n_1315, n_483);
  nand g1333 (n_1316, n_481, n_482);
  nand g1334 (n_1317, n_483, n_482);
  nand g1335 (n_1318, n_481, n_483);
  nand g1336 (n_501, n_1316, n_1317, n_1318);
  xor g1337 (n_1319, n_484, n_485);
  xor g1338 (n_91, n_1319, n_486);
  nand g1339 (n_1320, n_484, n_485);
  nand g1340 (n_1321, n_486, n_485);
  nand g1341 (n_1322, n_484, n_486);
  nand g1342 (n_42, n_1320, n_1321, n_1322);
  xor g1344 (n_489, n_687, A[12]);
  nand g1346 (n_1325, A[12], A[9]);
  nand g1347 (n_1326, A[8], A[12]);
  nand g1348 (n_504, n_688, n_1325, n_1326);
  xor g1349 (n_1327, n_487, n_488);
  xor g1350 (n_491, n_1327, n_489);
  nand g1351 (n_1328, n_487, n_488);
  nand g1352 (n_1329, n_489, n_488);
  nand g1353 (n_1330, n_487, n_489);
  nand g1354 (n_505, n_1328, n_1329, n_1330);
  xor g1355 (n_1331, A[13], A[16]);
  xor g1356 (n_493, n_1331, A[17]);
  nand g1360 (n_507, n_882, n_1024, n_1230);
  xor g1361 (n_1335, n_490, n_491);
  xor g1362 (n_494, n_1335, A[21]);
  nand g1363 (n_1336, n_490, n_491);
  nand g1364 (n_1337, A[21], n_491);
  nand g1365 (n_1338, n_490, A[21]);
  nand g1366 (n_510, n_1336, n_1337, n_1338);
  xor g1368 (n_496, n_1339, n_492);
  nand g1370 (n_1341, n_492, A[20]);
  nand g1372 (n_511, n_1157, n_1341, n_1342);
  xor g1373 (n_1343, n_493, n_494);
  xor g1374 (n_499, n_1343, n_495);
  nand g1375 (n_1344, n_493, n_494);
  nand g1376 (n_1345, n_495, n_494);
  nand g1377 (n_1346, n_493, n_495);
  nand g1378 (n_513, n_1344, n_1345, n_1346);
  xor g1379 (n_1347, n_496, n_497);
  xor g1380 (n_500, n_1347, n_498);
  nand g1381 (n_1348, n_496, n_497);
  nand g1382 (n_1349, n_498, n_497);
  nand g1383 (n_1350, n_496, n_498);
  nand g1384 (n_516, n_1348, n_1349, n_1350);
  xor g1385 (n_1351, n_499, n_500);
  xor g1386 (n_90, n_1351, n_501);
  nand g1387 (n_1352, n_499, n_500);
  nand g1388 (n_1353, n_501, n_500);
  nand g1389 (n_1354, n_499, n_501);
  nand g1390 (n_41, n_1352, n_1353, n_1354);
  nand g1397 (n_1358, A[10], n_504);
  nand g1398 (n_521, n_1356, n_1357, n_1358);
  xor g1399 (n_1359, A[14], A[13]);
  xor g1400 (n_508, n_1359, A[17]);
  nand g1403 (n_1362, A[14], A[17]);
  nand g1404 (n_523, n_797, n_1230, n_1362);
  xor g1405 (n_1363, n_505, n_506);
  xor g1406 (n_509, n_1363, A[18]);
  nand g1407 (n_1364, n_505, n_506);
  nand g1408 (n_1365, A[18], n_506);
  nand g1409 (n_1366, n_505, A[18]);
  nand g1410 (n_524, n_1364, n_1365, n_1366);
  xor g1411 (n_1367, A[21], A[22]);
  xor g1412 (n_512, n_1367, n_507);
  nand g1414 (n_1369, n_507, A[22]);
  nand g1415 (n_1370, A[21], n_507);
  nand g1416 (n_526, n_1073, n_1369, n_1370);
  xor g1417 (n_1371, n_508, n_509);
  xor g1418 (n_514, n_1371, n_510);
  nand g1419 (n_1372, n_508, n_509);
  nand g1420 (n_1373, n_510, n_509);
  nand g1421 (n_1374, n_508, n_510);
  nand g1422 (n_529, n_1372, n_1373, n_1374);
  xor g1423 (n_1375, n_511, n_512);
  xor g1424 (n_515, n_1375, n_513);
  nand g1425 (n_1376, n_511, n_512);
  nand g1426 (n_1377, n_513, n_512);
  nand g1427 (n_1378, n_511, n_513);
  nand g1428 (n_531, n_1376, n_1377, n_1378);
  xor g1429 (n_1379, n_514, n_515);
  xor g1430 (n_89, n_1379, n_516);
  nand g1431 (n_1380, n_514, n_515);
  nand g1432 (n_1381, n_516, n_515);
  nand g1433 (n_1382, n_514, n_516);
  nand g1434 (n_40, n_1380, n_1381, n_1382);
  xor g1437 (n_1383, A[11], A[9]);
  nand g1439 (n_1384, A[11], A[9]);
  nand g1442 (n_533, n_1384, n_1385, n_1386);
  xor g1443 (n_1387, A[14], A[15]);
  xor g1444 (n_522, n_1387, n_520);
  nand g1446 (n_1389, n_520, A[15]);
  nand g1447 (n_1390, A[14], n_520);
  nand g1448 (n_535, n_950, n_1389, n_1390);
  xor g1449 (n_1391, n_521, A[19]);
  xor g1450 (n_525, n_1391, A[18]);
  nand g1451 (n_1392, n_521, A[19]);
  nand g1453 (n_1394, n_521, A[18]);
  nand g1454 (n_537, n_1392, n_1112, n_1394);
  xor g1455 (n_1395, n_522, A[22]);
  xor g1456 (n_527, n_1395, n_523);
  nand g1457 (n_1396, n_522, A[22]);
  nand g1458 (n_1397, n_523, A[22]);
  nand g1459 (n_1398, n_522, n_523);
  nand g1460 (n_540, n_1396, n_1397, n_1398);
  xor g1461 (n_1399, A[23], n_524);
  xor g1462 (n_528, n_1399, n_525);
  nand g1463 (n_1400, A[23], n_524);
  nand g1464 (n_1401, n_525, n_524);
  nand g1465 (n_1402, A[23], n_525);
  nand g1466 (n_541, n_1400, n_1401, n_1402);
  xor g1467 (n_1403, n_526, n_527);
  xor g1468 (n_530, n_1403, n_528);
  nand g1469 (n_1404, n_526, n_527);
  nand g1470 (n_1405, n_528, n_527);
  nand g1471 (n_1406, n_526, n_528);
  nand g1472 (n_544, n_1404, n_1405, n_1406);
  xor g1473 (n_1407, n_529, n_530);
  xor g1474 (n_88, n_1407, n_531);
  nand g1475 (n_1408, n_529, n_530);
  nand g1476 (n_1409, n_531, n_530);
  nand g1477 (n_1410, n_529, n_531);
  nand g1478 (n_39, n_1408, n_1409, n_1410);
  xor g1479 (n_1411, A[12], A[11]);
  xor g1480 (n_534, n_1411, A[10]);
  nand g1484 (n_545, n_845, n_1100, n_710);
  xor g1485 (n_1415, n_533, A[15]);
  xor g1486 (n_536, n_1415, n_534);
  nand g1487 (n_1416, n_533, A[15]);
  nand g1488 (n_1417, n_534, A[15]);
  nand g1489 (n_1418, n_533, n_534);
  nand g1490 (n_546, n_1416, n_1417, n_1418);
  xor g1491 (n_1419, A[16], A[19]);
  xor g1492 (n_538, n_1419, n_535);
  nand g1494 (n_1421, n_535, A[19]);
  nand g1495 (n_1422, A[16], n_535);
  nand g1496 (n_549, n_1153, n_1421, n_1422);
  xor g1498 (n_539, n_1339, n_536);
  nand g1500 (n_1425, n_536, A[20]);
  nand g1502 (n_550, n_1157, n_1425, n_1426);
  xor g1503 (n_1427, A[23], n_537);
  xor g1504 (n_542, n_1427, n_538);
  nand g1505 (n_1428, A[23], n_537);
  nand g1506 (n_1429, n_538, n_537);
  nand g1507 (n_1430, A[23], n_538);
  nand g1508 (n_553, n_1428, n_1429, n_1430);
  xor g1509 (n_1431, n_539, n_540);
  xor g1510 (n_543, n_1431, n_541);
  nand g1511 (n_1432, n_539, n_540);
  nand g1512 (n_1433, n_541, n_540);
  nand g1513 (n_1434, n_539, n_541);
  nand g1514 (n_555, n_1432, n_1433, n_1434);
  xor g1515 (n_1435, n_542, n_543);
  xor g1516 (n_87, n_1435, n_544);
  nand g1517 (n_1436, n_542, n_543);
  nand g1518 (n_1437, n_544, n_543);
  nand g1519 (n_1438, n_542, n_544);
  nand g1520 (n_38, n_1436, n_1437, n_1438);
  xor g1521 (n_1439, A[12], A[13]);
  xor g1522 (n_547, n_1439, n_545);
  nand g1523 (n_1440, A[12], A[13]);
  nand g1524 (n_1441, n_545, A[13]);
  nand g1525 (n_1442, A[12], n_545);
  nand g1526 (n_558, n_1440, n_1441, n_1442);
  xor g1528 (n_548, n_1023, n_546);
  nand g1530 (n_1445, n_546, A[17]);
  nand g1531 (n_1446, A[16], n_546);
  nand g1532 (n_560, n_1024, n_1445, n_1446);
  xor g1533 (n_1447, n_547, A[21]);
  nand g1535 (n_1448, n_547, A[21]);
  nand g1538 (n_562, n_1448, n_1449, n_1450);
  xor g1539 (n_1451, A[20], n_548);
  xor g1540 (n_552, n_1451, n_549);
  nand g1541 (n_1452, A[20], n_548);
  nand g1542 (n_1453, n_549, n_548);
  nand g1543 (n_1454, A[20], n_549);
  nand g1544 (n_563, n_1452, n_1453, n_1454);
  xor g1545 (n_1455, n_550, n_551);
  xor g1546 (n_554, n_1455, n_552);
  nand g1547 (n_1456, n_550, n_551);
  nand g1548 (n_1457, n_552, n_551);
  nand g1549 (n_1458, n_550, n_552);
  nand g1550 (n_566, n_1456, n_1457, n_1458);
  xor g1551 (n_1459, n_553, n_554);
  xor g1552 (n_86, n_1459, n_555);
  nand g1553 (n_1460, n_553, n_554);
  nand g1554 (n_1461, n_555, n_554);
  nand g1555 (n_1462, n_553, n_555);
  nand g1556 (n_37, n_1460, n_1461, n_1462);
  nand g1564 (n_570, n_1464, n_1465, n_1230);
  xor g1565 (n_1467, n_558, A[18]);
  xor g1566 (n_561, n_1467, A[21]);
  nand g1567 (n_1468, n_558, A[18]);
  nand g1569 (n_1470, n_558, A[21]);
  nand g1570 (n_572, n_1468, n_956, n_1470);
  xor g1572 (n_564, n_1471, n_560);
  nand g1575 (n_1474, A[22], n_560);
  nand g1576 (n_575, n_1472, n_1473, n_1474);
  xor g1577 (n_1475, n_561, n_562);
  xor g1578 (n_565, n_1475, n_563);
  nand g1579 (n_1476, n_561, n_562);
  nand g1580 (n_1477, n_563, n_562);
  nand g1581 (n_1478, n_561, n_563);
  nand g1582 (n_577, n_1476, n_1477, n_1478);
  xor g1583 (n_1479, n_564, n_565);
  xor g1584 (n_85, n_1479, n_566);
  nand g1585 (n_1480, n_564, n_565);
  nand g1586 (n_1481, n_566, n_565);
  nand g1587 (n_1482, n_564, n_566);
  nand g1588 (n_36, n_1480, n_1481, n_1482);
  xor g1598 (n_573, n_1111, A[22]);
  nand g1600 (n_1489, A[22], A[18]);
  nand g1601 (n_1490, A[19], A[22]);
  nand g1602 (n_581, n_1112, n_1489, n_1490);
  xor g1603 (n_1491, n_570, n_571);
  xor g1604 (n_574, n_1491, A[23]);
  nand g1605 (n_1492, n_570, n_571);
  nand g1606 (n_1493, A[23], n_571);
  nand g1607 (n_1494, n_570, A[23]);
  nand g1608 (n_583, n_1492, n_1493, n_1494);
  xor g1609 (n_1495, n_572, n_573);
  xor g1610 (n_576, n_1495, n_574);
  nand g1611 (n_1496, n_572, n_573);
  nand g1612 (n_1497, n_574, n_573);
  nand g1613 (n_1498, n_572, n_574);
  nand g1614 (n_586, n_1496, n_1497, n_1498);
  xor g1615 (n_1499, n_575, n_576);
  xor g1616 (n_84, n_1499, n_577);
  nand g1617 (n_1500, n_575, n_576);
  nand g1618 (n_1501, n_577, n_576);
  nand g1619 (n_1502, n_575, n_577);
  nand g1620 (n_35, n_1500, n_1501, n_1502);
  xor g1622 (n_580, n_851, A[14]);
  nand g1624 (n_1505, A[14], A[16]);
  nand g1626 (n_587, n_852, n_1505, n_950);
  xor g1627 (n_1507, A[19], n_579);
  nand g1629 (n_1508, A[19], n_579);
  nand g1632 (n_589, n_1508, n_1509, n_1306);
  xor g1633 (n_1511, A[20], A[23]);
  xor g1634 (n_584, n_1511, n_580);
  nand g1636 (n_1513, n_580, A[23]);
  nand g1637 (n_1514, A[20], n_580);
  nand g1638 (n_590, n_1310, n_1513, n_1514);
  xor g1639 (n_1515, n_581, n_582);
  xor g1640 (n_585, n_1515, n_583);
  nand g1641 (n_1516, n_581, n_582);
  nand g1642 (n_1517, n_583, n_582);
  nand g1643 (n_1518, n_581, n_583);
  nand g1644 (n_593, n_1516, n_1517, n_1518);
  xor g1645 (n_1519, n_584, n_585);
  xor g1646 (n_83, n_1519, n_586);
  nand g1647 (n_1520, n_584, n_585);
  nand g1648 (n_1521, n_586, n_585);
  nand g1649 (n_1522, n_584, n_586);
  nand g1650 (n_34, n_1520, n_1521, n_1522);
  xor g1652 (n_588, n_1023, A[21]);
  nand g1654 (n_1525, A[21], A[17]);
  nand g1655 (n_1526, A[16], A[21]);
  nand g1656 (n_596, n_1024, n_1525, n_1526);
  xor g1658 (n_591, n_1339, n_587);
  nand g1660 (n_1529, n_587, A[20]);
  nand g1662 (n_597, n_1157, n_1529, n_1530);
  xor g1663 (n_1531, n_588, n_589);
  xor g1664 (n_592, n_1531, n_590);
  nand g1665 (n_1532, n_588, n_589);
  nand g1666 (n_1533, n_590, n_589);
  nand g1667 (n_1534, n_588, n_590);
  nand g1668 (n_600, n_1532, n_1533, n_1534);
  xor g1669 (n_1535, n_591, n_592);
  xor g1670 (n_82, n_1535, n_593);
  nand g1671 (n_1536, n_591, n_592);
  nand g1672 (n_1537, n_593, n_592);
  nand g1673 (n_1538, n_591, n_593);
  nand g1674 (n_33, n_1536, n_1537, n_1538);
  xor g1678 (n_598, n_1539, A[21]);
  nand g1682 (n_604, n_1540, n_1541, n_956);
  xor g1683 (n_1543, A[22], n_596);
  xor g1684 (n_599, n_1543, n_597);
  nand g1685 (n_1544, A[22], n_596);
  nand g1686 (n_1545, n_597, n_596);
  nand g1687 (n_1546, A[22], n_597);
  nand g1688 (n_607, n_1544, n_1545, n_1546);
  xor g1689 (n_1547, n_598, n_599);
  xor g1690 (n_81, n_1547, n_600);
  nand g1691 (n_1548, n_598, n_599);
  nand g1692 (n_1549, n_600, n_599);
  nand g1693 (n_1550, n_598, n_600);
  nand g1694 (n_32, n_1548, n_1549, n_1550);
  nand g1699 (n_1552, A[18], A[17]);
  nand g1700 (n_1553, A[22], A[17]);
  nand g1702 (n_610, n_1552, n_1553, n_1489);
  xor g1704 (n_606, n_1555, n_604);
  nand g1706 (n_1557, n_604, A[23]);
  nand g1708 (n_611, n_1556, n_1557, n_1558);
  xor g1709 (n_1559, n_605, n_606);
  xor g1710 (n_80, n_1559, n_607);
  nand g1711 (n_1560, n_605, n_606);
  nand g1712 (n_1561, n_607, n_606);
  nand g1713 (n_1562, n_605, n_607);
  nand g1714 (n_31, n_1560, n_1561, n_1562);
  xor g1716 (n_609, n_1563, A[20]);
  nand g1719 (n_1566, A[19], A[20]);
  nand g1720 (n_613, n_1306, n_1157, n_1566);
  nand g1723 (n_1568, A[23], A[19]);
  nand g1724 (n_1569, n_609, A[19]);
  nand g1725 (n_1570, A[23], n_609);
  nand g1726 (n_615, n_1568, n_1569, n_1570);
  xor g1727 (n_1571, n_610, n_611);
  xor g1728 (n_79, n_1571, n_612);
  nand g1729 (n_1572, n_610, n_611);
  nand g1730 (n_1573, n_612, n_611);
  nand g1731 (n_1574, n_610, n_612);
  nand g1732 (n_30, n_1572, n_1573, n_1574);
  xor g1734 (n_614, n_1575, A[20]);
  nand g1738 (n_618, n_1449, n_1028, n_1157);
  xor g1739 (n_1579, n_613, n_614);
  xor g1740 (n_78, n_1579, n_615);
  nand g1741 (n_1580, n_613, n_614);
  nand g1742 (n_1581, n_615, n_614);
  nand g1743 (n_1582, n_613, n_615);
  nand g1744 (n_77, n_1580, n_1581, n_1582);
  nand g1751 (n_1586, A[22], n_618);
  nand g1752 (n_28, n_1584, n_1585, n_1586);
  xor g1755 (n_1587, A[23], A[21]);
  nand g1757 (n_1588, A[23], A[21]);
  nand g1760 (n_27, n_1588, n_1589, n_1590);
  xor g1762 (n_75, n_1591, A[22]);
  nand g1764 (n_1593, A[22], A[23]);
  nand g1766 (n_74, n_1592, n_1593, n_1594);
  nor g11 (n_1610, A[0], A[2]);
  nand g12 (n_1605, A[0], A[2]);
  nor g13 (n_1606, n_70, A[3]);
  nand g14 (n_1607, n_70, A[3]);
  nor g15 (n_1616, n_69, A[4]);
  nand g16 (n_1611, n_69, A[4]);
  nor g17 (n_1612, A[5], n_116);
  nand g18 (n_1613, A[5], n_116);
  nor g19 (n_1622, A[6], n_115);
  nand g20 (n_1617, A[6], n_115);
  nor g21 (n_1618, A[7], n_114);
  nand g22 (n_1619, A[7], n_114);
  nor g23 (n_1628, n_65, n_113);
  nand g24 (n_1623, n_65, n_113);
  nor g25 (n_1624, n_64, n_112);
  nand g26 (n_1625, n_64, n_112);
  nor g27 (n_1634, n_63, n_111);
  nand g28 (n_1629, n_63, n_111);
  nor g29 (n_1630, n_62, n_110);
  nand g30 (n_1631, n_62, n_110);
  nor g31 (n_1640, n_61, n_109);
  nand g32 (n_1635, n_61, n_109);
  nor g33 (n_1636, n_60, n_108);
  nand g34 (n_1637, n_60, n_108);
  nor g35 (n_1646, n_59, n_107);
  nand g36 (n_1641, n_59, n_107);
  nor g37 (n_1642, n_58, n_106);
  nand g38 (n_1643, n_58, n_106);
  nor g39 (n_1652, n_57, n_105);
  nand g40 (n_1647, n_57, n_105);
  nor g41 (n_1648, n_56, n_104);
  nand g42 (n_1649, n_56, n_104);
  nor g43 (n_1658, n_55, n_103);
  nand g44 (n_1653, n_55, n_103);
  nor g45 (n_1654, n_54, n_102);
  nand g46 (n_1655, n_54, n_102);
  nor g47 (n_1664, n_53, n_101);
  nand g48 (n_1659, n_53, n_101);
  nor g49 (n_1660, n_52, n_100);
  nand g50 (n_1661, n_52, n_100);
  nor g51 (n_1670, n_51, n_99);
  nand g52 (n_1665, n_51, n_99);
  nor g53 (n_1666, n_50, n_98);
  nand g54 (n_1667, n_50, n_98);
  nor g55 (n_1676, n_49, n_97);
  nand g56 (n_1671, n_49, n_97);
  nor g57 (n_1672, n_48, n_96);
  nand g58 (n_1673, n_48, n_96);
  nor g59 (n_1682, n_47, n_95);
  nand g60 (n_1677, n_47, n_95);
  nor g61 (n_1678, n_46, n_94);
  nand g62 (n_1679, n_46, n_94);
  nor g63 (n_1688, n_45, n_93);
  nand g64 (n_1683, n_45, n_93);
  nor g65 (n_1684, n_44, n_92);
  nand g66 (n_1685, n_44, n_92);
  nor g67 (n_1694, n_43, n_91);
  nand g68 (n_1689, n_43, n_91);
  nor g69 (n_1690, n_42, n_90);
  nand g70 (n_1691, n_42, n_90);
  nor g71 (n_1700, n_41, n_89);
  nand g72 (n_1695, n_41, n_89);
  nor g73 (n_1696, n_40, n_88);
  nand g74 (n_1697, n_40, n_88);
  nor g75 (n_1706, n_39, n_87);
  nand g76 (n_1701, n_39, n_87);
  nor g77 (n_1702, n_38, n_86);
  nand g78 (n_1703, n_38, n_86);
  nor g79 (n_1712, n_37, n_85);
  nand g80 (n_1707, n_37, n_85);
  nor g81 (n_1708, n_36, n_84);
  nand g82 (n_1709, n_36, n_84);
  nor g83 (n_1718, n_35, n_83);
  nand g84 (n_1713, n_35, n_83);
  nor g85 (n_1714, n_34, n_82);
  nand g86 (n_1715, n_34, n_82);
  nor g87 (n_1724, n_33, n_81);
  nand g88 (n_1719, n_33, n_81);
  nor g89 (n_1720, n_32, n_80);
  nand g90 (n_1721, n_32, n_80);
  nor g91 (n_1730, n_31, n_79);
  nand g92 (n_1725, n_31, n_79);
  nor g93 (n_1726, n_30, n_78);
  nand g94 (n_1727, n_30, n_78);
  nor g95 (n_1736, n_29, n_77);
  nand g96 (n_1731, n_29, n_77);
  nor g97 (n_1732, n_28, n_76);
  nand g98 (n_1733, n_28, n_76);
  nor g99 (n_1740, n_27, n_75);
  nand g100 (n_1737, n_27, n_75);
  nor g106 (n_1608, n_1605, n_1606);
  nor g110 (n_1614, n_1611, n_1612);
  nor g113 (n_1750, n_1616, n_1612);
  nor g114 (n_1620, n_1617, n_1618);
  nor g117 (n_1752, n_1622, n_1618);
  nor g118 (n_1626, n_1623, n_1624);
  nor g121 (n_1760, n_1628, n_1624);
  nor g122 (n_1632, n_1629, n_1630);
  nor g125 (n_1762, n_1634, n_1630);
  nor g126 (n_1638, n_1635, n_1636);
  nor g129 (n_1770, n_1640, n_1636);
  nor g130 (n_1644, n_1641, n_1642);
  nor g133 (n_1772, n_1646, n_1642);
  nor g134 (n_1650, n_1647, n_1648);
  nor g137 (n_1780, n_1652, n_1648);
  nor g138 (n_1656, n_1653, n_1654);
  nor g141 (n_1782, n_1658, n_1654);
  nor g142 (n_1662, n_1659, n_1660);
  nor g145 (n_1790, n_1664, n_1660);
  nor g146 (n_1668, n_1665, n_1666);
  nor g149 (n_1792, n_1670, n_1666);
  nor g150 (n_1674, n_1671, n_1672);
  nor g153 (n_1800, n_1676, n_1672);
  nor g154 (n_1680, n_1677, n_1678);
  nor g157 (n_1802, n_1682, n_1678);
  nor g158 (n_1686, n_1683, n_1684);
  nor g161 (n_1810, n_1688, n_1684);
  nor g162 (n_1692, n_1689, n_1690);
  nor g165 (n_1812, n_1694, n_1690);
  nor g166 (n_1698, n_1695, n_1696);
  nor g169 (n_1820, n_1700, n_1696);
  nor g170 (n_1704, n_1701, n_1702);
  nor g173 (n_1822, n_1706, n_1702);
  nor g174 (n_1710, n_1707, n_1708);
  nor g177 (n_1830, n_1712, n_1708);
  nor g178 (n_1716, n_1713, n_1714);
  nor g181 (n_1832, n_1718, n_1714);
  nor g182 (n_1722, n_1719, n_1720);
  nor g185 (n_1840, n_1724, n_1720);
  nor g186 (n_1728, n_1725, n_1726);
  nor g189 (n_1842, n_1730, n_1726);
  nor g190 (n_1734, n_1731, n_1732);
  nor g193 (n_1850, n_1736, n_1732);
  nor g203 (n_1748, n_1622, n_1747);
  nand g212 (n_1860, n_1750, n_1752);
  nor g213 (n_1758, n_1634, n_1757);
  nand g222 (n_1867, n_1760, n_1762);
  nor g223 (n_1768, n_1646, n_1767);
  nand g232 (n_1875, n_1770, n_1772);
  nor g233 (n_1778, n_1658, n_1777);
  nand g242 (n_1882, n_1780, n_1782);
  nor g243 (n_1788, n_1670, n_1787);
  nand g252 (n_1890, n_1790, n_1792);
  nor g253 (n_1798, n_1682, n_1797);
  nand g262 (n_1897, n_1800, n_1802);
  nor g263 (n_1808, n_1694, n_1807);
  nand g1776 (n_1905, n_1810, n_1812);
  nor g1777 (n_1818, n_1706, n_1817);
  nand g1786 (n_1912, n_1820, n_1822);
  nor g1787 (n_1828, n_1718, n_1827);
  nand g1796 (n_1920, n_1830, n_1832);
  nor g1797 (n_1838, n_1730, n_1837);
  nand g1806 (n_1927, n_1840, n_1842);
  nor g1807 (n_1848, n_1740, n_1847);
  nand g1814 (n_2131, n_1611, n_1854);
  nand g1816 (n_2133, n_1747, n_1855);
  nand g1819 (n_2136, n_1858, n_1859);
  nand g1822 (n_1935, n_1862, n_1863);
  nor g1823 (n_1865, n_1640, n_1864);
  nor g1826 (n_1945, n_1640, n_1867);
  nor g1832 (n_1873, n_1871, n_1864);
  nor g1835 (n_1951, n_1867, n_1871);
  nor g1836 (n_1877, n_1875, n_1864);
  nor g1839 (n_1954, n_1867, n_1875);
  nor g1840 (n_1880, n_1664, n_1879);
  nor g1843 (n_2034, n_1664, n_1882);
  nor g1849 (n_1888, n_1886, n_1879);
  nor g1852 (n_2040, n_1882, n_1886);
  nor g1853 (n_1892, n_1890, n_1879);
  nor g1856 (n_1960, n_1882, n_1890);
  nor g1857 (n_1895, n_1688, n_1894);
  nor g1860 (n_1973, n_1688, n_1897);
  nor g1866 (n_1903, n_1901, n_1894);
  nor g1869 (n_1983, n_1897, n_1901);
  nor g1870 (n_1907, n_1905, n_1894);
  nor g1873 (n_1988, n_1897, n_1905);
  nor g1874 (n_1910, n_1712, n_1909);
  nor g1877 (n_2086, n_1712, n_1912);
  nor g1883 (n_1918, n_1916, n_1909);
  nor g1886 (n_2092, n_1912, n_1916);
  nor g1887 (n_1922, n_1920, n_1909);
  nor g1890 (n_1996, n_1912, n_1920);
  nor g1891 (n_1925, n_1736, n_1924);
  nor g1894 (n_2009, n_1736, n_1927);
  nor g1900 (n_1933, n_1931, n_1924);
  nor g1903 (n_2019, n_1927, n_1931);
  nand g1906 (n_2140, n_1623, n_1937);
  nand g1907 (n_1938, n_1760, n_1935);
  nand g1908 (n_2142, n_1757, n_1938);
  nand g1911 (n_2145, n_1941, n_1942);
  nand g1914 (n_2148, n_1864, n_1944);
  nand g1915 (n_1947, n_1945, n_1935);
  nand g1916 (n_2151, n_1946, n_1947);
  nand g1917 (n_1950, n_1948, n_1935);
  nand g1918 (n_2153, n_1949, n_1950);
  nand g1919 (n_1953, n_1951, n_1935);
  nand g1920 (n_2156, n_1952, n_1953);
  nand g1921 (n_1956, n_1954, n_1935);
  nand g1922 (n_2024, n_1955, n_1956);
  nor g1923 (n_1958, n_1676, n_1957);
  nand g1932 (n_2048, n_1800, n_1960);
  nor g1933 (n_1967, n_1965, n_1957);
  nor g1938 (n_1970, n_1897, n_1957);
  nand g1947 (n_2060, n_1960, n_1973);
  nand g1952 (n_2064, n_1960, n_1978);
  nand g1957 (n_2068, n_1960, n_1983);
  nand g1962 (n_2072, n_1960, n_1988);
  nor g1963 (n_1994, n_1724, n_1993);
  nand g1972 (n_2100, n_1840, n_1996);
  nor g1973 (n_2003, n_2001, n_1993);
  nor g1978 (n_2006, n_1927, n_1993);
  nand g1987 (n_2112, n_1996, n_2009);
  nand g1992 (n_2116, n_1996, n_2014);
  nand g1997 (n_2120, n_1996, n_2019);
  nand g2000 (n_2160, n_1647, n_2026);
  nand g2001 (n_2027, n_1780, n_2024);
  nand g2002 (n_2162, n_1777, n_2027);
  nand g2005 (n_2165, n_2030, n_2031);
  nand g2008 (n_2168, n_1879, n_2033);
  nand g2009 (n_2036, n_2034, n_2024);
  nand g2010 (n_2171, n_2035, n_2036);
  nand g2011 (n_2039, n_2037, n_2024);
  nand g2012 (n_2173, n_2038, n_2039);
  nand g2013 (n_2042, n_2040, n_2024);
  nand g2014 (n_2176, n_2041, n_2042);
  nand g2015 (n_2043, n_1960, n_2024);
  nand g2016 (n_2178, n_1957, n_2043);
  nand g2019 (n_2181, n_2046, n_2047);
  nand g2022 (n_2183, n_2050, n_2051);
  nand g2025 (n_2186, n_2054, n_2055);
  nand g2028 (n_2189, n_2058, n_2059);
  nand g2031 (n_2192, n_2062, n_2063);
  nand g2034 (n_2194, n_2066, n_2067);
  nand g2037 (n_2197, n_2070, n_2071);
  nand g2040 (n_2076, n_2074, n_2075);
  nand g2043 (n_2201, n_1695, n_2078);
  nand g2044 (n_2079, n_1820, n_2076);
  nand g2045 (n_2203, n_1817, n_2079);
  nand g2048 (n_2206, n_2082, n_2083);
  nand g2051 (n_2209, n_1909, n_2085);
  nand g2052 (n_2088, n_2086, n_2076);
  nand g2053 (n_2212, n_2087, n_2088);
  nand g2054 (n_2091, n_2089, n_2076);
  nand g2055 (n_2214, n_2090, n_2091);
  nand g2056 (n_2094, n_2092, n_2076);
  nand g2057 (n_2217, n_2093, n_2094);
  nand g2058 (n_2095, n_1996, n_2076);
  nand g2059 (n_2219, n_1993, n_2095);
  nand g2062 (n_2222, n_2098, n_2099);
  nand g2065 (n_2224, n_2102, n_2103);
  nand g2068 (n_2227, n_2106, n_2107);
  nand g2071 (n_2230, n_2110, n_2111);
  nand g2074 (n_2233, n_2114, n_2115);
  nand g2077 (n_2235, n_2118, n_2119);
  nand g2080 (n_2238, n_2122, n_2123);
  xnor g2092 (Z[5], n_2131, n_2132);
  xnor g2094 (Z[6], n_2133, n_2134);
  xnor g2097 (Z[7], n_2136, n_2137);
  xnor g2099 (Z[8], n_1935, n_2138);
  xnor g2102 (Z[9], n_2140, n_2141);
  xnor g2104 (Z[10], n_2142, n_2143);
  xnor g2107 (Z[11], n_2145, n_2146);
  xnor g2110 (Z[12], n_2148, n_2149);
  xnor g2113 (Z[13], n_2151, n_2152);
  xnor g2115 (Z[14], n_2153, n_2154);
  xnor g2118 (Z[15], n_2156, n_2157);
  xnor g2120 (Z[16], n_2024, n_2158);
  xnor g2123 (Z[17], n_2160, n_2161);
  xnor g2125 (Z[18], n_2162, n_2163);
  xnor g2128 (Z[19], n_2165, n_2166);
  xnor g2131 (Z[20], n_2168, n_2169);
  xnor g2134 (Z[21], n_2171, n_2172);
  xnor g2136 (Z[22], n_2173, n_2174);
  xnor g2139 (Z[23], n_2176, n_2177);
  xnor g2141 (Z[24], n_2178, n_2179);
  xnor g2144 (Z[25], n_2181, n_2182);
  xnor g2146 (Z[26], n_2183, n_2184);
  xnor g2149 (Z[27], n_2186, n_2187);
  xnor g2152 (Z[28], n_2189, n_2190);
  xnor g2155 (Z[29], n_2192, n_2193);
  xnor g2157 (Z[30], n_2194, n_2195);
  xnor g2160 (Z[31], n_2197, n_2198);
  xnor g2162 (Z[32], n_2076, n_2199);
  xnor g2165 (Z[33], n_2201, n_2202);
  xnor g2167 (Z[34], n_2203, n_2204);
  xnor g2170 (Z[35], n_2206, n_2207);
  xnor g2173 (Z[36], n_2209, n_2210);
  xnor g2176 (Z[37], n_2212, n_2213);
  xnor g2178 (Z[38], n_2214, n_2215);
  xnor g2181 (Z[39], n_2217, n_2218);
  xnor g2183 (Z[40], n_2219, n_2220);
  xnor g2186 (Z[41], n_2222, n_2223);
  xnor g2188 (Z[42], n_2224, n_2225);
  xnor g2191 (Z[43], n_2227, n_2228);
  xnor g2194 (Z[44], n_2230, n_2231);
  xnor g2197 (Z[45], n_2233, n_2234);
  xnor g2199 (Z[46], n_2235, n_2236);
  xnor g2202 (Z[47], n_2238, n_2239);
  or g2215 (n_1044, A[1], wc);
  not gc (wc, n_171);
  or g2216 (n_1045, A[1], wc0);
  not gc0 (wc0, A[2]);
  or g2217 (n_1070, wc1, A[24]);
  not gc1 (wc1, A[18]);
  or g2219 (n_1157, wc2, A[24]);
  not gc2 (wc2, A[20]);
  xnor g2220 (n_1215, A[6], A[5]);
  or g2221 (n_1216, A[5], wc3);
  not gc3 (wc3, A[6]);
  or g2222 (n_1253, A[6], wc4);
  not gc4 (wc4, A[7]);
  or g2223 (n_1254, wc5, A[6]);
  not gc5 (wc5, A[5]);
  or g2224 (n_1306, wc6, A[24]);
  not gc6 (wc6, A[19]);
  xnor g2225 (n_1339, A[24], A[20]);
  or g2227 (n_1356, A[9], wc7);
  not gc7 (wc7, A[10]);
  or g2228 (n_1385, wc8, A[10]);
  not gc8 (wc8, A[9]);
  or g2229 (n_1386, A[10], wc9);
  not gc9 (wc9, A[11]);
  or g2230 (n_1449, wc10, A[24]);
  not gc10 (wc10, A[21]);
  or g2232 (n_1464, wc11, A[14]);
  not gc11 (wc11, A[13]);
  or g2233 (n_1465, A[14], wc12);
  not gc12 (wc12, A[17]);
  or g2234 (n_1486, A[14], wc13);
  not gc13 (wc13, A[15]);
  xnor g2235 (n_1539, A[18], A[17]);
  or g2236 (n_1540, A[17], wc14);
  not gc14 (wc14, A[18]);
  or g2237 (n_1541, A[17], wc15);
  not gc15 (wc15, A[21]);
  xnor g2239 (n_1555, A[23], A[19]);
  or g2240 (n_1556, A[19], wc16);
  not gc16 (wc16, A[23]);
  xnor g2241 (n_1563, A[24], A[19]);
  xnor g2243 (n_1575, A[24], A[21]);
  or g2245 (n_1584, A[21], wc17);
  not gc17 (wc17, A[22]);
  or g2246 (n_1589, wc18, A[22]);
  not gc18 (wc18, A[21]);
  or g2247 (n_1590, A[22], wc19);
  not gc19 (wc19, A[23]);
  xnor g2248 (n_1591, A[24], A[23]);
  or g2249 (n_1592, wc20, A[24]);
  not gc20 (wc20, A[23]);
  or g2250 (n_1594, wc21, A[24]);
  not gc21 (wc21, A[22]);
  xnor g2252 (n_1087, A[2], A[1]);
  or g2253 (n_1089, A[1], wc22);
  not gc22 (wc22, A[3]);
  xnor g2254 (n_454, n_1251, A[6]);
  xnor g2255 (n_506, n_1219, n_504);
  or g2256 (n_1357, A[9], wc23);
  not gc23 (wc23, n_504);
  xnor g2257 (n_520, n_1383, A[10]);
  xnor g2259 (n_571, n_1387, A[14]);
  nand g2260 (n_579, n_950, n_1486);
  xnor g2261 (n_605, n_1539, A[22]);
  xnor g2262 (n_76, n_1587, A[22]);
  or g2264 (n_2125, wc24, n_1610);
  not gc24 (wc24, n_1605);
  or g2266 (n_1048, wc25, n_69);
  not gc25 (wc25, A[5]);
  or g2267 (n_1050, wc26, n_69);
  not gc26 (wc26, A[6]);
  xnor g2268 (n_1471, n_508, A[22]);
  or g2269 (n_1472, wc27, n_508);
  not gc27 (wc27, A[22]);
  or g2270 (n_1509, A[24], wc28);
  not gc28 (wc28, n_579);
  or g2271 (n_1530, A[24], wc29);
  not gc29 (wc29, n_587);
  or g2272 (n_1558, A[19], wc30);
  not gc30 (wc30, n_604);
  xnor g2273 (n_612, n_609, n_1555);
  xnor g2274 (n_29, n_1367, n_618);
  or g2275 (n_1585, A[21], wc31);
  not gc31 (wc31, n_618);
  and g2276 (n_1745, wc32, n_1607);
  not gc32 (wc32, n_1608);
  or g2277 (n_2128, wc33, n_1606);
  not gc33 (wc33, n_1607);
  or g2279 (n_1450, A[24], wc34);
  not gc34 (wc34, n_547);
  xnor g2280 (n_582, n_1507, A[24]);
  and g2281 (n_1738, wc35, n_74);
  not gc35 (wc35, A[24]);
  or g2282 (n_1739, wc36, n_74);
  not gc36 (wc36, A[24]);
  not g2283 (Z[2], n_2125);
  or g2285 (n_1052, n_182, wc37);
  not gc37 (wc37, n_181);
  or g2286 (n_1053, wc38, n_182);
  not gc38 (wc38, A[9]);
  or g2287 (n_1426, A[24], wc39);
  not gc39 (wc39, n_536);
  xnor g2288 (n_551, n_1447, A[24]);
  or g2291 (n_2129, wc40, n_1616);
  not gc40 (wc40, n_1611);
  or g2292 (n_2236, wc41, n_1740);
  not gc41 (wc41, n_1737);
  or g2294 (n_1217, A[5], wc42);
  not gc42 (wc42, n_434);
  or g2295 (n_1854, n_1616, n_1745);
  xor g2296 (Z[3], n_1605, n_2128);
  xor g2297 (Z[4], n_1745, n_2129);
  or g2298 (n_2239, wc43, n_1738);
  not gc43 (wc43, n_1739);
  or g2299 (n_1057, wc44, n_204);
  not gc44 (wc44, A[10]);
  or g2300 (n_1305, A[24], wc45);
  not gc45 (wc45, n_476);
  or g2301 (n_1473, wc46, n_508);
  not gc46 (wc46, n_560);
  and g2302 (n_1747, wc47, n_1613);
  not gc47 (wc47, n_1614);
  or g2303 (n_1855, n_1745, wc48);
  not gc48 (wc48, n_1750);
  or g2304 (n_2132, wc49, n_1612);
  not gc49 (wc49, n_1613);
  or g2305 (n_2234, wc50, n_1732);
  not gc50 (wc50, n_1733);
  xnor g2306 (n_480, n_1303, A[24]);
  or g2307 (n_1856, wc51, n_1622);
  not gc51 (wc51, n_1750);
  or g2308 (n_2134, wc52, n_1622);
  not gc52 (wc52, n_1617);
  or g2309 (n_1058, n_204, wc53);
  not gc53 (wc53, n_65);
  and g2310 (n_1847, wc54, n_1733);
  not gc54 (wc54, n_1734);
  and g2311 (n_1858, wc55, n_1617);
  not gc55 (wc55, n_1748);
  or g2312 (n_1931, wc56, n_1740);
  not gc56 (wc56, n_1850);
  or g2313 (n_2141, wc57, n_1624);
  not gc57 (wc57, n_1625);
  or g2314 (n_2228, wc58, n_1726);
  not gc58 (wc58, n_1727);
  or g2315 (n_2231, wc59, n_1736);
  not gc59 (wc59, n_1731);
  and g2317 (n_1754, wc60, n_1619);
  not gc60 (wc60, n_1620);
  or g2318 (n_1859, n_1745, n_1856);
  or g2319 (n_2137, wc61, n_1618);
  not gc61 (wc61, n_1619);
  or g2321 (n_1064, n_237, wc62);
  not gc62 (wc62, n_238);
  or g2322 (n_1066, wc63, n_237);
  not gc63 (wc63, A[17]);
  or g2323 (n_1197, A[24], wc64);
  not gc64 (wc64, n_421);
  and g2324 (n_1757, wc65, n_1625);
  not gc65 (wc65, n_1626);
  and g2325 (n_1837, wc66, n_1721);
  not gc66 (wc66, n_1722);
  and g2326 (n_1844, wc67, n_1727);
  not gc67 (wc67, n_1728);
  and g2327 (n_1755, wc68, n_1752);
  not gc68 (wc68, n_1747);
  or g2328 (n_1939, wc69, n_1634);
  not gc69 (wc69, n_1760);
  or g2329 (n_2001, wc70, n_1730);
  not gc70 (wc70, n_1840);
  and g2330 (n_1932, wc71, n_1737);
  not gc71 (wc71, n_1848);
  or g2331 (n_2138, wc72, n_1628);
  not gc72 (wc72, n_1623);
  or g2332 (n_2143, wc73, n_1634);
  not gc73 (wc73, n_1629);
  or g2333 (n_2220, wc74, n_1724);
  not gc74 (wc74, n_1719);
  or g2334 (n_2223, wc75, n_1720);
  not gc75 (wc75, n_1721);
  or g2335 (n_2225, wc76, n_1730);
  not gc76 (wc76, n_1725);
  or g2337 (n_1069, A[24], wc77);
  not gc77 (wc77, n_358);
  or g2338 (n_1198, A[24], wc78);
  not gc78 (wc78, n_420);
  and g2339 (n_1764, wc79, n_1631);
  not gc79 (wc79, n_1632);
  and g2340 (n_1862, wc80, n_1754);
  not gc80 (wc80, n_1755);
  and g2341 (n_1845, wc81, n_1842);
  not gc81 (wc81, n_1837);
  or g2342 (n_1863, n_1860, n_1745);
  and g2343 (n_2014, wc82, n_1850);
  not gc82 (wc82, n_1927);
  or g2344 (n_2146, wc83, n_1630);
  not gc83 (wc83, n_1631);
  xnor g2345 (n_363, n_1067, A[24]);
  xnor g2346 (n_1075, n_290, n_361);
  or g2347 (n_1076, wc84, n_290);
  not gc84 (wc84, n_361);
  xnor g2348 (n_1155, n_401, A[24]);
  or g2349 (n_1156, A[24], wc85);
  not gc85 (wc85, n_401);
  xnor g2350 (n_425, n_1195, A[24]);
  or g2351 (n_1342, A[24], wc86);
  not gc86 (wc86, n_492);
  and g2352 (n_1941, wc87, n_1629);
  not gc87 (wc87, n_1758);
  and g2353 (n_1765, wc88, n_1762);
  not gc88 (wc88, n_1757);
  and g2354 (n_2002, wc89, n_1725);
  not gc89 (wc89, n_1838);
  and g2355 (n_1924, wc90, n_1844);
  not gc90 (wc90, n_1845);
  or g2356 (n_2218, wc91, n_1714);
  not gc91 (wc91, n_1715);
  or g2357 (n_1078, wc92, n_290);
  not gc92 (wc92, n_362);
  and g2358 (n_1864, wc93, n_1764);
  not gc93 (wc93, n_1765);
  and g2359 (n_1929, wc94, n_1850);
  not gc94 (wc94, n_1924);
  or g2360 (n_1937, wc95, n_1628);
  not gc95 (wc95, n_1935);
  or g2361 (n_1942, n_1939, wc96);
  not gc96 (wc96, n_1935);
  or g2362 (n_1944, wc97, n_1867);
  not gc97 (wc97, n_1935);
  or g2363 (n_2149, wc98, n_1640);
  not gc98 (wc98, n_1635);
  or g2364 (n_2213, wc99, n_1708);
  not gc99 (wc99, n_1709);
  and g2365 (n_1767, wc100, n_1637);
  not gc100 (wc100, n_1638);
  and g2366 (n_1834, wc101, n_1715);
  not gc101 (wc101, n_1716);
  and g2367 (n_2011, wc102, n_1731);
  not gc102 (wc102, n_1925);
  and g2368 (n_2016, wc103, n_1847);
  not gc103 (wc103, n_1929);
  and g2369 (n_2021, n_1932, wc104);
  not gc104 (wc104, n_1933);
  or g2370 (n_2152, wc105, n_1636);
  not gc105 (wc105, n_1637);
  or g2371 (n_2215, wc106, n_1718);
  not gc106 (wc106, n_1713);
  or g2372 (n_1871, wc107, n_1646);
  not gc107 (wc107, n_1770);
  and g2373 (n_1946, wc108, n_1635);
  not gc108 (wc108, n_1865);
  and g2374 (n_1869, wc109, n_1770);
  not gc109 (wc109, n_1864);
  and g2375 (n_1948, wc110, n_1770);
  not gc110 (wc110, n_1867);
  or g2376 (n_2154, wc111, n_1646);
  not gc111 (wc111, n_1641);
  or g2377 (n_2158, wc112, n_1652);
  not gc112 (wc112, n_1647);
  and g2378 (n_1774, wc113, n_1643);
  not gc113 (wc113, n_1644);
  and g2379 (n_1777, wc114, n_1649);
  not gc114 (wc114, n_1650);
  and g2380 (n_1827, wc115, n_1709);
  not gc115 (wc115, n_1710);
  and g2381 (n_1872, wc116, n_1641);
  not gc116 (wc116, n_1768);
  or g2382 (n_1916, wc117, n_1718);
  not gc117 (wc117, n_1830);
  and g2383 (n_1949, wc118, n_1767);
  not gc118 (wc118, n_1869);
  or g2384 (n_2157, wc119, n_1642);
  not gc119 (wc119, n_1643);
  or g2385 (n_2161, wc120, n_1648);
  not gc120 (wc120, n_1649);
  or g2386 (n_2207, wc121, n_1702);
  not gc121 (wc121, n_1703);
  or g2387 (n_2210, wc122, n_1712);
  not gc122 (wc122, n_1707);
  and g2388 (n_1775, wc123, n_1772);
  not gc123 (wc123, n_1767);
  or g2389 (n_2028, wc124, n_1658);
  not gc124 (wc124, n_1780);
  and g2390 (n_1835, wc125, n_1832);
  not gc125 (wc125, n_1827);
  or g2391 (n_2163, wc126, n_1658);
  not gc126 (wc126, n_1653);
  and g2392 (n_1784, wc127, n_1655);
  not gc127 (wc127, n_1656);
  and g2393 (n_1787, wc128, n_1661);
  not gc128 (wc128, n_1662);
  and g2394 (n_1876, wc129, n_1774);
  not gc129 (wc129, n_1775);
  and g2395 (n_2030, wc130, n_1653);
  not gc130 (wc130, n_1778);
  and g2396 (n_1917, wc131, n_1713);
  not gc131 (wc131, n_1828);
  and g2397 (n_1921, wc132, n_1834);
  not gc132 (wc132, n_1835);
  and g2398 (n_1952, n_1872, wc133);
  not gc133 (wc133, n_1873);
  or g2399 (n_2166, wc134, n_1654);
  not gc134 (wc134, n_1655);
  or g2400 (n_2169, wc135, n_1664);
  not gc135 (wc135, n_1659);
  or g2401 (n_2172, wc136, n_1660);
  not gc136 (wc136, n_1661);
  and g2402 (n_1785, wc137, n_1782);
  not gc137 (wc137, n_1777);
  or g2403 (n_1886, wc138, n_1670);
  not gc138 (wc138, n_1790);
  and g2404 (n_2037, wc139, n_1790);
  not gc139 (wc139, n_1882);
  or g2405 (n_2174, wc140, n_1670);
  not gc140 (wc140, n_1665);
  and g2406 (n_1794, wc141, n_1667);
  not gc141 (wc141, n_1668);
  and g2407 (n_1824, wc142, n_1703);
  not gc142 (wc142, n_1704);
  and g2408 (n_1879, wc143, n_1784);
  not gc143 (wc143, n_1785);
  and g2409 (n_1887, wc144, n_1665);
  not gc144 (wc144, n_1788);
  and g2410 (n_1955, n_1876, wc145);
  not gc145 (wc145, n_1877);
  or g2411 (n_2177, wc146, n_1666);
  not gc146 (wc146, n_1667);
  or g2412 (n_2179, wc147, n_1676);
  not gc147 (wc147, n_1671);
  or g2413 (n_2202, wc148, n_1696);
  not gc148 (wc148, n_1697);
  or g2414 (n_2204, wc149, n_1706);
  not gc149 (wc149, n_1701);
  and g2415 (n_1817, wc150, n_1697);
  not gc150 (wc150, n_1698);
  and g2416 (n_1795, wc151, n_1792);
  not gc151 (wc151, n_1787);
  or g2417 (n_2080, wc152, n_1706);
  not gc152 (wc152, n_1820);
  and g2418 (n_1884, wc153, n_1790);
  not gc153 (wc153, n_1879);
  or g2419 (n_2187, wc154, n_1678);
  not gc154 (wc154, n_1679);
  or g2420 (n_2190, wc155, n_1688);
  not gc155 (wc155, n_1683);
  or g2421 (n_2198, wc156, n_1690);
  not gc156 (wc156, n_1691);
  or g2422 (n_2199, wc157, n_1700);
  not gc157 (wc157, n_1695);
  and g2423 (n_1797, wc158, n_1673);
  not gc158 (wc158, n_1674);
  and g2424 (n_1804, wc159, n_1679);
  not gc159 (wc159, n_1680);
  and g2425 (n_1807, wc160, n_1685);
  not gc160 (wc160, n_1686);
  and g2426 (n_1814, wc161, n_1691);
  not gc161 (wc161, n_1692);
  and g2427 (n_1891, wc162, n_1794);
  not gc162 (wc162, n_1795);
  or g2428 (n_1965, wc163, n_1682);
  not gc163 (wc163, n_1800);
  or g2429 (n_1901, wc164, n_1694);
  not gc164 (wc164, n_1810);
  and g2430 (n_1825, wc165, n_1822);
  not gc165 (wc165, n_1817);
  and g2431 (n_2035, wc166, n_1659);
  not gc166 (wc166, n_1880);
  and g2432 (n_2038, wc167, n_1787);
  not gc167 (wc167, n_1884);
  and g2433 (n_2041, n_1887, wc168);
  not gc168 (wc168, n_1888);
  and g2434 (n_2089, wc169, n_1830);
  not gc169 (wc169, n_1912);
  or g2435 (n_2044, wc170, n_1676);
  not gc170 (wc170, n_1960);
  or g2436 (n_2026, wc171, n_1652);
  not gc171 (wc171, n_2024);
  or g2437 (n_2031, n_2028, wc172);
  not gc172 (wc172, n_2024);
  or g2438 (n_2033, wc173, n_1882);
  not gc173 (wc173, n_2024);
  or g2439 (n_2182, wc174, n_1672);
  not gc174 (wc174, n_1673);
  or g2440 (n_2184, wc175, n_1682);
  not gc175 (wc175, n_1677);
  or g2441 (n_2193, wc176, n_1684);
  not gc176 (wc176, n_1685);
  or g2442 (n_2195, wc177, n_1694);
  not gc177 (wc177, n_1689);
  and g2443 (n_1805, wc178, n_1802);
  not gc178 (wc178, n_1797);
  and g2444 (n_1815, wc179, n_1812);
  not gc179 (wc179, n_1807);
  and g2445 (n_2082, wc180, n_1701);
  not gc180 (wc180, n_1818);
  and g2446 (n_1909, wc181, n_1824);
  not gc181 (wc181, n_1825);
  and g2447 (n_1978, wc182, n_1810);
  not gc182 (wc182, n_1897);
  or g2448 (n_2096, wc183, n_1724);
  not gc183 (wc183, n_1996);
  or g2449 (n_2104, n_2001, wc184);
  not gc184 (wc184, n_1996);
  or g2450 (n_2108, wc185, n_1927);
  not gc185 (wc185, n_1996);
  and g2451 (n_1966, wc186, n_1677);
  not gc186 (wc186, n_1798);
  and g2452 (n_1894, wc187, n_1804);
  not gc187 (wc187, n_1805);
  and g2453 (n_1902, wc188, n_1689);
  not gc188 (wc188, n_1808);
  and g2454 (n_1906, wc189, n_1814);
  not gc189 (wc189, n_1815);
  and g2455 (n_1957, n_1891, wc190);
  not gc190 (wc190, n_1892);
  and g2456 (n_1914, wc191, n_1830);
  not gc191 (wc191, n_1909);
  or g2457 (n_2052, n_1965, wc192);
  not gc192 (wc192, n_1960);
  or g2458 (n_2056, wc193, n_1897);
  not gc193 (wc193, n_1960);
  or g2459 (n_2047, n_2044, wc194);
  not gc194 (wc194, n_2024);
  or g2460 (n_2051, n_2048, wc195);
  not gc195 (wc195, n_2024);
  and g2461 (n_1899, wc196, n_1810);
  not gc196 (wc196, n_1894);
  and g2462 (n_2087, wc197, n_1707);
  not gc197 (wc197, n_1910);
  and g2463 (n_2090, wc198, n_1827);
  not gc198 (wc198, n_1914);
  and g2464 (n_2093, n_1917, wc199);
  not gc199 (wc199, n_1918);
  and g2465 (n_1993, n_1921, wc200);
  not gc200 (wc200, n_1922);
  and g2466 (n_1963, wc201, n_1800);
  not gc201 (wc201, n_1957);
  and g2467 (n_1976, wc202, n_1973);
  not gc202 (wc202, n_1957);
  and g2468 (n_1981, wc203, n_1978);
  not gc203 (wc203, n_1957);
  and g2469 (n_1986, wc204, n_1983);
  not gc204 (wc204, n_1957);
  and g2470 (n_1991, wc205, n_1988);
  not gc205 (wc205, n_1957);
  and g2471 (n_1975, wc206, n_1683);
  not gc206 (wc206, n_1895);
  and g2472 (n_1980, wc207, n_1807);
  not gc207 (wc207, n_1899);
  and g2473 (n_1985, n_1902, wc208);
  not gc208 (wc208, n_1903);
  and g2474 (n_1990, n_1906, wc209);
  not gc209 (wc209, n_1907);
  and g2475 (n_2046, wc210, n_1671);
  not gc210 (wc210, n_1958);
  and g2476 (n_2050, wc211, n_1797);
  not gc211 (wc211, n_1963);
  and g2477 (n_2054, n_1966, wc212);
  not gc212 (wc212, n_1967);
  and g2478 (n_2058, n_1894, wc213);
  not gc213 (wc213, n_1970);
  and g2479 (n_1999, wc214, n_1840);
  not gc214 (wc214, n_1993);
  and g2480 (n_2012, wc215, n_2009);
  not gc215 (wc215, n_1993);
  and g2481 (n_2017, wc216, n_2014);
  not gc216 (wc216, n_1993);
  and g2482 (n_2022, wc217, n_2019);
  not gc217 (wc217, n_1993);
  or g2483 (n_2055, n_2052, wc218);
  not gc218 (wc218, n_2024);
  or g2484 (n_2059, n_2056, wc219);
  not gc219 (wc219, n_2024);
  or g2485 (n_2063, n_2060, wc220);
  not gc220 (wc220, n_2024);
  or g2486 (n_2067, n_2064, wc221);
  not gc221 (wc221, n_2024);
  or g2487 (n_2071, n_2068, wc222);
  not gc222 (wc222, n_2024);
  or g2488 (n_2075, n_2072, wc223);
  not gc223 (wc223, n_2024);
  and g2489 (n_2098, wc224, n_1719);
  not gc224 (wc224, n_1994);
  and g2490 (n_2102, wc225, n_1837);
  not gc225 (wc225, n_1999);
  and g2491 (n_2106, n_2002, wc226);
  not gc226 (wc226, n_2003);
  and g2492 (n_2110, n_1924, wc227);
  not gc227 (wc227, n_2006);
  and g2493 (n_2114, wc228, n_2011);
  not gc228 (wc228, n_2012);
  and g2494 (n_2118, wc229, n_2016);
  not gc229 (wc229, n_2017);
  and g2495 (n_2122, wc230, n_2021);
  not gc230 (wc230, n_2022);
  and g2496 (n_2062, n_1975, wc231);
  not gc231 (wc231, n_1976);
  and g2497 (n_2066, n_1980, wc232);
  not gc232 (wc232, n_1981);
  and g2498 (n_2070, n_1985, wc233);
  not gc233 (wc233, n_1986);
  and g2499 (n_2074, n_1990, wc234);
  not gc234 (wc234, n_1991);
  or g2500 (n_2078, wc235, n_1700);
  not gc235 (wc235, n_2076);
  or g2501 (n_2083, n_2080, wc236);
  not gc236 (wc236, n_2076);
  or g2502 (n_2085, wc237, n_1912);
  not gc237 (wc237, n_2076);
  or g2503 (n_2099, n_2096, wc238);
  not gc238 (wc238, n_2076);
  or g2504 (n_2103, wc239, n_2100);
  not gc239 (wc239, n_2076);
  or g2505 (n_2107, n_2104, wc240);
  not gc240 (wc240, n_2076);
  or g2506 (n_2111, n_2108, wc241);
  not gc241 (wc241, n_2076);
  or g2507 (n_2115, wc242, n_2112);
  not gc242 (wc242, n_2076);
  or g2508 (n_2119, wc243, n_2116);
  not gc243 (wc243, n_2076);
  or g2509 (n_2123, wc244, n_2120);
  not gc244 (wc244, n_2076);
endmodule

module mult_signed_const_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_3884_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_171, n_172, n_174, n_178, n_179;
  wire n_181, n_182, n_183, n_185, n_186, n_187, n_188, n_193;
  wire n_194, n_195, n_199, n_200, n_201, n_202, n_203, n_205;
  wire n_207, n_208, n_209, n_210, n_211, n_213, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_223, n_224, n_225, n_226;
  wire n_227, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_245, n_246, n_247, n_248, n_249, n_250, n_251;
  wire n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263;
  wire n_264, n_266, n_268, n_269, n_270, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_278, n_281, n_283, n_284;
  wire n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_298, n_299, n_300, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_314, n_315;
  wire n_316, n_317, n_318, n_319, n_320, n_321, n_322, n_323;
  wire n_324, n_325, n_326, n_327, n_332, n_333, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_350, n_352, n_353, n_354, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_372, n_373, n_374, n_375, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444;
  wire n_445, n_446, n_447, n_448, n_449, n_450, n_454, n_455;
  wire n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463;
  wire n_464, n_465, n_466, n_467, n_468, n_469, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_501, n_505, n_506, n_507, n_508;
  wire n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516;
  wire n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_530, n_531, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_558, n_559, n_560, n_561, n_562, n_563;
  wire n_564, n_565, n_566, n_570, n_571, n_572, n_573, n_574;
  wire n_575, n_576, n_577, n_579, n_580, n_581, n_582, n_583;
  wire n_584, n_585, n_586, n_588, n_589, n_590, n_591, n_592;
  wire n_593, n_598, n_599, n_600, n_606, n_607, n_609, n_611;
  wire n_612, n_613, n_614, n_615, n_618, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_642, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
  wire n_654, n_657, n_658, n_659, n_660, n_661, n_662, n_663;
  wire n_664, n_665, n_666, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_678, n_685, n_686, n_687;
  wire n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_699;
  wire n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710;
  wire n_711, n_712, n_713, n_714, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_739, n_740;
  wire n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748;
  wire n_749, n_750, n_751, n_752, n_753, n_754, n_761, n_762;
  wire n_763, n_764, n_765, n_766, n_767, n_768, n_769, n_770;
  wire n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778;
  wire n_787, n_791, n_792, n_793, n_794, n_795, n_796, n_797;
  wire n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805;
  wire n_806, n_815, n_816, n_817, n_818, n_819, n_820, n_821;
  wire n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829;
  wire n_830, n_831, n_832, n_833, n_834, n_842, n_843, n_844;
  wire n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860;
  wire n_861, n_862, n_865, n_866, n_867, n_868, n_869, n_870;
  wire n_871, n_874, n_875, n_876, n_877, n_878, n_879, n_880;
  wire n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888;
  wire n_889, n_890, n_891, n_892, n_893, n_894, n_903, n_904;
  wire n_906, n_907, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_937, n_938;
  wire n_939, n_940, n_941, n_945, n_946, n_947, n_948, n_949;
  wire n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957;
  wire n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965;
  wire n_966, n_973, n_975, n_979, n_980, n_981, n_982, n_983;
  wire n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991;
  wire n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999;
  wire n_1000, n_1001, n_1002, n_1009, n_1010, n_1015, n_1016, n_1017;
  wire n_1019, n_1020, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027;
  wire n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035;
  wire n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043;
  wire n_1045, n_1046, n_1049, n_1050, n_1051, n_1055, n_1056, n_1057;
  wire n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066;
  wire n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074;
  wire n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082;
  wire n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090;
  wire n_1091, n_1092, n_1093, n_1094, n_1095, n_1098, n_1099, n_1100;
  wire n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108;
  wire n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116;
  wire n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124;
  wire n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132;
  wire n_1133, n_1135, n_1136, n_1137, n_1138, n_1141, n_1143, n_1144;
  wire n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1153, n_1154;
  wire n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162;
  wire n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170;
  wire n_1171, n_1172, n_1173, n_1174, n_1175, n_1177, n_1178, n_1179;
  wire n_1180, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1190;
  wire n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200;
  wire n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208;
  wire n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1216, n_1217;
  wire n_1218, n_1219, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226;
  wire n_1227, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237;
  wire n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
  wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1253, n_1254;
  wire n_1259, n_1261, n_1262, n_1265, n_1266, n_1267, n_1268, n_1269;
  wire n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
  wire n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285;
  wire n_1286, n_1289, n_1290, n_1291, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1298, n_1301, n_1303, n_1304, n_1305, n_1306, n_1307;
  wire n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315;
  wire n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1327;
  wire n_1330, n_1333, n_1334, n_1335, n_1337, n_1338, n_1339, n_1340;
  wire n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348;
  wire n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356;
  wire n_1359, n_1360, n_1362, n_1363, n_1365, n_1366, n_1367, n_1368;
  wire n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376;
  wire n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1387, n_1388;
  wire n_1390, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399;
  wire n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407;
  wire n_1408, n_1409, n_1410, n_1414, n_1415, n_1418, n_1419, n_1422;
  wire n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430;
  wire n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438;
  wire n_1439, n_1442, n_1445, n_1447, n_1448, n_1449, n_1450, n_1451;
  wire n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1460, n_1461, n_1462, n_1466, n_1467, n_1468, n_1469, n_1471;
  wire n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479;
  wire n_1480, n_1481, n_1482, n_1485, n_1486, n_1489, n_1491, n_1492;
  wire n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500;
  wire n_1501, n_1502, n_1506, n_1507, n_1511, n_1512, n_1513, n_1514;
  wire n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522;
  wire n_1523, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535;
  wire n_1536, n_1537, n_1538, n_1543, n_1544, n_1546, n_1547, n_1548;
  wire n_1549, n_1550, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560;
  wire n_1561, n_1562, n_1563, n_1567, n_1569, n_1570, n_1571, n_1572;
  wire n_1573, n_1574, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583;
  wire n_1584, n_1585, n_1586, n_1587, n_1588, n_1605, n_1606, n_1607;
  wire n_1608, n_1610, n_1611, n_1612, n_1613, n_1614, n_1616, n_1617;
  wire n_1618, n_1619, n_1620, n_1622, n_1623, n_1624, n_1625, n_1626;
  wire n_1628, n_1629, n_1630, n_1631, n_1632, n_1634, n_1635, n_1636;
  wire n_1637, n_1638, n_1640, n_1641, n_1642, n_1643, n_1644, n_1646;
  wire n_1647, n_1648, n_1649, n_1650, n_1652, n_1653, n_1654, n_1655;
  wire n_1656, n_1658, n_1659, n_1660, n_1661, n_1662, n_1664, n_1665;
  wire n_1666, n_1667, n_1668, n_1670, n_1671, n_1672, n_1673, n_1674;
  wire n_1676, n_1677, n_1678, n_1679, n_1680, n_1682, n_1683, n_1684;
  wire n_1685, n_1686, n_1688, n_1689, n_1690, n_1691, n_1692, n_1694;
  wire n_1695, n_1696, n_1697, n_1698, n_1700, n_1701, n_1702, n_1703;
  wire n_1704, n_1706, n_1707, n_1708, n_1709, n_1710, n_1712, n_1713;
  wire n_1714, n_1715, n_1716, n_1718, n_1719, n_1720, n_1721, n_1722;
  wire n_1724, n_1725, n_1726, n_1727, n_1728, n_1730, n_1731, n_1732;
  wire n_1733, n_1734, n_1736, n_1737, n_1738, n_1739, n_1740, n_1745;
  wire n_1747, n_1748, n_1750, n_1752, n_1754, n_1755, n_1757, n_1758;
  wire n_1760, n_1762, n_1764, n_1765, n_1767, n_1768, n_1770, n_1772;
  wire n_1774, n_1775, n_1777, n_1778, n_1780, n_1782, n_1784, n_1785;
  wire n_1787, n_1788, n_1790, n_1792, n_1794, n_1795, n_1797, n_1798;
  wire n_1800, n_1802, n_1804, n_1805, n_1807, n_1808, n_1810, n_1812;
  wire n_1814, n_1815, n_1817, n_1818, n_1820, n_1822, n_1824, n_1825;
  wire n_1827, n_1828, n_1830, n_1832, n_1834, n_1835, n_1837, n_1838;
  wire n_1840, n_1842, n_1844, n_1845, n_1847, n_1848, n_1850, n_1854;
  wire n_1855, n_1856, n_1858, n_1859, n_1860, n_1862, n_1863, n_1864;
  wire n_1865, n_1867, n_1869, n_1871, n_1872, n_1873, n_1875, n_1876;
  wire n_1877, n_1879, n_1880, n_1882, n_1884, n_1886, n_1887, n_1888;
  wire n_1890, n_1891, n_1892, n_1894, n_1895, n_1897, n_1899, n_1901;
  wire n_1902, n_1903, n_1905, n_1906, n_1907, n_1909, n_1910, n_1912;
  wire n_1914, n_1916, n_1917, n_1918, n_1920, n_1921, n_1922, n_1924;
  wire n_1925, n_1927, n_1929, n_1931, n_1932, n_1933, n_1935, n_1937;
  wire n_1938, n_1939, n_1941, n_1942, n_1944, n_1945, n_1946, n_1947;
  wire n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955;
  wire n_1956, n_1957, n_1958, n_1960, n_1963, n_1965, n_1966, n_1967;
  wire n_1970, n_1973, n_1975, n_1976, n_1978, n_1980, n_1981, n_1983;
  wire n_1985, n_1986, n_1988, n_1990, n_1991, n_1993, n_1994, n_1996;
  wire n_1999, n_2001, n_2002, n_2003, n_2006, n_2009, n_2011, n_2012;
  wire n_2014, n_2016, n_2017, n_2019, n_2021, n_2022, n_2024, n_2026;
  wire n_2027, n_2028, n_2030, n_2031, n_2033, n_2034, n_2035, n_2036;
  wire n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044;
  wire n_2046, n_2047, n_2048, n_2050, n_2051, n_2052, n_2054, n_2055;
  wire n_2056, n_2058, n_2059, n_2060, n_2062, n_2063, n_2064, n_2066;
  wire n_2067, n_2068, n_2070, n_2071, n_2072, n_2074, n_2075, n_2076;
  wire n_2078, n_2079, n_2080, n_2082, n_2083, n_2085, n_2086, n_2087;
  wire n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095;
  wire n_2096, n_2098, n_2099, n_2100, n_2102, n_2103, n_2104, n_2106;
  wire n_2107, n_2108, n_2110, n_2111, n_2112, n_2114, n_2115, n_2116;
  wire n_2118, n_2119, n_2120, n_2122, n_2123, n_2125, n_2128, n_2129;
  wire n_2131, n_2132, n_2133, n_2134, n_2136, n_2137, n_2138, n_2140;
  wire n_2141, n_2142, n_2143, n_2145, n_2146, n_2148, n_2149, n_2151;
  wire n_2152, n_2153, n_2154, n_2156, n_2157, n_2158, n_2160, n_2161;
  wire n_2162, n_2163, n_2165, n_2166, n_2168, n_2169, n_2171, n_2172;
  wire n_2173, n_2174, n_2176, n_2177, n_2178, n_2179, n_2181, n_2182;
  wire n_2183, n_2184, n_2186, n_2187, n_2189, n_2190, n_2192, n_2193;
  wire n_2194, n_2195, n_2197, n_2198, n_2199, n_2201, n_2202, n_2203;
  wire n_2204, n_2206, n_2207, n_2209, n_2210, n_2212, n_2213, n_2214;
  wire n_2215, n_2217, n_2218, n_2219, n_2220, n_2222, n_2223, n_2224;
  wire n_2225, n_2227, n_2228, n_2230, n_2231, n_2233, n_2234, n_2235;
  wire n_2236, n_2238, n_2239;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_118, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_623, A[1], A[2]);
  xor g270 (n_117, n_623, n_171);
  nand g3 (n_624, A[1], A[2]);
  nand g271 (n_625, n_171, A[2]);
  nand g272 (n_626, A[1], n_171);
  nand g273 (n_68, n_624, n_625, n_626);
  xor g274 (n_627, A[2], A[3]);
  xor g275 (n_116, n_627, A[5]);
  nand g276 (n_628, A[2], A[3]);
  nand g4 (n_629, A[5], A[3]);
  nand g277 (n_630, A[2], A[5]);
  nand g278 (n_67, n_628, n_629, n_630);
  xor g279 (n_172, A[0], A[3]);
  and g280 (n_174, A[0], A[3]);
  xor g281 (n_631, A[4], n_172);
  xor g282 (n_115, n_631, A[6]);
  nand g283 (n_632, A[4], n_172);
  nand g284 (n_633, A[6], n_172);
  nand g5 (n_634, A[4], A[6]);
  nand g6 (n_66, n_632, n_633, n_634);
  xor g287 (n_635, n_118, A[4]);
  xor g288 (n_69, n_635, n_174);
  nand g289 (n_636, n_118, A[4]);
  nand g290 (n_637, n_174, A[4]);
  nand g291 (n_638, n_118, n_174);
  nand g292 (n_178, n_636, n_637, n_638);
  xor g293 (n_639, A[5], n_69);
  xor g294 (n_114, n_639, A[7]);
  nand g295 (n_640, A[5], n_69);
  nand g296 (n_641, A[7], n_69);
  nand g297 (n_642, A[5], A[7]);
  nand g298 (n_65, n_640, n_641, n_642);
  xor g305 (n_647, A[5], n_117);
  xor g306 (n_179, n_647, A[6]);
  nand g307 (n_648, A[5], n_117);
  nand g308 (n_649, A[6], n_117);
  nand g309 (n_650, A[5], A[6]);
  nand g310 (n_181, n_648, n_649, n_650);
  xor g311 (n_651, n_178, A[8]);
  xor g312 (n_113, n_651, n_179);
  nand g313 (n_652, n_178, A[8]);
  nand g314 (n_653, n_179, A[8]);
  nand g315 (n_654, n_178, n_179);
  nand g316 (n_64, n_652, n_653, n_654);
  xor g318 (n_182, n_627, A[6]);
  nand g320 (n_657, A[6], A[3]);
  nand g321 (n_658, A[2], A[6]);
  nand g322 (n_185, n_628, n_657, n_658);
  xor g323 (n_659, n_68, A[7]);
  xor g324 (n_183, n_659, n_181);
  nand g325 (n_660, n_68, A[7]);
  nand g326 (n_661, n_181, A[7]);
  nand g327 (n_662, n_68, n_181);
  nand g328 (n_187, n_660, n_661, n_662);
  xor g329 (n_663, A[9], n_182);
  xor g330 (n_112, n_663, n_183);
  nand g331 (n_664, A[9], n_182);
  nand g332 (n_665, n_183, n_182);
  nand g333 (n_666, A[9], n_183);
  nand g334 (n_63, n_664, n_665, n_666);
  xor g338 (n_186, n_631, A[7]);
  nand g340 (n_669, A[7], n_172);
  nand g341 (n_670, A[4], A[7]);
  nand g342 (n_71, n_632, n_669, n_670);
  xor g343 (n_671, n_185, A[8]);
  xor g344 (n_188, n_671, A[10]);
  nand g345 (n_672, n_185, A[8]);
  nand g346 (n_673, A[10], A[8]);
  nand g347 (n_674, n_185, A[10]);
  nand g348 (n_194, n_672, n_673, n_674);
  xor g349 (n_675, n_186, n_187);
  xor g350 (n_111, n_675, n_188);
  nand g351 (n_676, n_186, n_187);
  nand g352 (n_677, n_188, n_187);
  nand g353 (n_678, n_186, n_188);
  nand g354 (n_62, n_676, n_677, n_678);
  xor g364 (n_193, n_639, A[9]);
  nand g366 (n_685, A[9], n_69);
  nand g367 (n_686, A[5], A[9]);
  nand g368 (n_200, n_640, n_685, n_686);
  xor g369 (n_687, A[8], A[11]);
  xor g370 (n_195, n_687, n_71);
  nand g371 (n_688, A[8], A[11]);
  nand g372 (n_689, n_71, A[11]);
  nand g373 (n_690, A[8], n_71);
  nand g374 (n_202, n_688, n_689, n_690);
  xor g375 (n_691, n_193, n_194);
  xor g376 (n_110, n_691, n_195);
  nand g377 (n_692, n_193, n_194);
  nand g378 (n_693, n_195, n_194);
  nand g379 (n_694, n_193, n_195);
  nand g380 (n_61, n_692, n_693, n_694);
  xor g387 (n_699, A[5], A[6]);
  xor g388 (n_199, n_699, n_117);
  xor g393 (n_703, n_178, A[10]);
  xor g394 (n_201, n_703, A[9]);
  nand g395 (n_704, n_178, A[10]);
  nand g396 (n_705, A[9], A[10]);
  nand g397 (n_706, n_178, A[9]);
  nand g398 (n_208, n_704, n_705, n_706);
  xor g399 (n_707, n_199, A[12]);
  xor g400 (n_203, n_707, n_200);
  nand g401 (n_708, n_199, A[12]);
  nand g402 (n_709, n_200, A[12]);
  nand g403 (n_710, n_199, n_200);
  nand g404 (n_210, n_708, n_709, n_710);
  xor g405 (n_711, n_201, n_202);
  xor g406 (n_109, n_711, n_203);
  nand g407 (n_712, n_201, n_202);
  nand g408 (n_713, n_203, n_202);
  nand g409 (n_714, n_201, n_203);
  nand g410 (n_60, n_712, n_713, n_714);
  xor g412 (n_205, n_627, n_68);
  nand g414 (n_717, n_68, A[3]);
  nand g415 (n_718, A[2], n_68);
  nand g416 (n_213, n_628, n_717, n_718);
  xor g417 (n_719, A[6], A[7]);
  xor g418 (n_207, n_719, n_205);
  nand g419 (n_720, A[6], A[7]);
  nand g420 (n_721, n_205, A[7]);
  nand g421 (n_722, A[6], n_205);
  nand g422 (n_215, n_720, n_721, n_722);
  xor g423 (n_723, n_181, A[10]);
  xor g424 (n_209, n_723, A[11]);
  nand g425 (n_724, n_181, A[10]);
  nand g426 (n_725, A[11], A[10]);
  nand g427 (n_726, n_181, A[11]);
  nand g428 (n_216, n_724, n_725, n_726);
  xor g429 (n_727, A[13], n_207);
  xor g430 (n_211, n_727, n_208);
  nand g431 (n_728, A[13], n_207);
  nand g432 (n_729, n_208, n_207);
  nand g433 (n_730, A[13], n_208);
  nand g434 (n_219, n_728, n_729, n_730);
  xor g435 (n_731, n_209, n_210);
  xor g436 (n_108, n_731, n_211);
  nand g437 (n_732, n_209, n_210);
  nand g438 (n_733, n_211, n_210);
  nand g439 (n_734, n_209, n_211);
  nand g440 (n_59, n_732, n_733, n_734);
  xor g449 (n_739, A[8], n_213);
  xor g450 (n_217, n_739, A[12]);
  nand g451 (n_740, A[8], n_213);
  nand g452 (n_741, A[12], n_213);
  nand g453 (n_742, A[8], A[12]);
  nand g454 (n_73, n_740, n_741, n_742);
  xor g455 (n_743, A[14], A[11]);
  xor g456 (n_218, n_743, n_186);
  nand g457 (n_744, A[14], A[11]);
  nand g458 (n_745, n_186, A[11]);
  nand g459 (n_746, A[14], n_186);
  nand g460 (n_224, n_744, n_745, n_746);
  xor g461 (n_747, n_215, n_216);
  xor g462 (n_220, n_747, n_217);
  nand g463 (n_748, n_215, n_216);
  nand g464 (n_749, n_217, n_216);
  nand g465 (n_750, n_215, n_217);
  nand g466 (n_226, n_748, n_749, n_750);
  xor g467 (n_751, n_218, n_219);
  xor g468 (n_107, n_751, n_220);
  nand g469 (n_752, n_218, n_219);
  nand g470 (n_753, n_220, n_219);
  nand g471 (n_754, n_218, n_220);
  nand g472 (n_58, n_752, n_753, n_754);
  xor g482 (n_72, n_639, A[8]);
  nand g484 (n_761, A[8], n_69);
  nand g485 (n_762, A[5], A[8]);
  nand g486 (n_232, n_640, n_761, n_762);
  xor g487 (n_763, A[9], A[13]);
  xor g488 (n_223, n_763, A[12]);
  nand g489 (n_764, A[9], A[13]);
  nand g490 (n_765, A[12], A[13]);
  nand g491 (n_766, A[9], A[12]);
  nand g492 (n_234, n_764, n_765, n_766);
  xor g493 (n_767, A[15], n_71);
  xor g494 (n_225, n_767, n_72);
  nand g495 (n_768, A[15], n_71);
  nand g496 (n_769, n_72, n_71);
  nand g497 (n_770, A[15], n_72);
  nand g498 (n_236, n_768, n_769, n_770);
  xor g499 (n_771, n_73, n_223);
  xor g500 (n_227, n_771, n_224);
  nand g501 (n_772, n_73, n_223);
  nand g502 (n_773, n_224, n_223);
  nand g503 (n_774, n_73, n_224);
  nand g504 (n_238, n_772, n_773, n_774);
  xor g505 (n_775, n_225, n_226);
  xor g506 (n_106, n_775, n_227);
  nand g507 (n_776, n_225, n_226);
  nand g508 (n_777, n_227, n_226);
  nand g509 (n_778, n_225, n_227);
  nand g510 (n_57, n_776, n_777, n_778);
  xor g523 (n_787, n_178, A[9]);
  xor g524 (n_233, n_787, A[10]);
  xor g529 (n_791, n_199, A[14]);
  xor g530 (n_235, n_791, A[13]);
  nand g531 (n_792, n_199, A[14]);
  nand g532 (n_793, A[13], A[14]);
  nand g533 (n_794, n_199, A[13]);
  nand g534 (n_245, n_792, n_793, n_794);
  xor g535 (n_795, n_232, A[16]);
  xor g536 (n_237, n_795, n_233);
  nand g537 (n_796, n_232, A[16]);
  nand g538 (n_797, n_233, A[16]);
  nand g539 (n_798, n_232, n_233);
  nand g540 (n_249, n_796, n_797, n_798);
  xor g541 (n_799, n_234, n_235);
  xor g542 (n_239, n_799, n_236);
  nand g543 (n_800, n_234, n_235);
  nand g544 (n_801, n_236, n_235);
  nand g545 (n_802, n_234, n_236);
  nand g546 (n_250, n_800, n_801, n_802);
  xor g547 (n_803, n_237, n_238);
  xor g548 (n_105, n_803, n_239);
  nand g549 (n_804, n_237, n_238);
  nand g550 (n_805, n_239, n_238);
  nand g551 (n_806, n_237, n_239);
  nand g552 (n_56, n_804, n_805, n_806);
  xor g565 (n_815, n_182, A[10]);
  xor g566 (n_246, n_815, A[14]);
  nand g567 (n_816, n_182, A[10]);
  nand g568 (n_817, A[14], A[10]);
  nand g569 (n_818, n_182, A[14]);
  nand g570 (n_257, n_816, n_817, n_818);
  xor g571 (n_819, A[11], A[15]);
  xor g572 (n_247, n_819, A[17]);
  nand g573 (n_820, A[11], A[15]);
  nand g574 (n_821, A[17], A[15]);
  nand g575 (n_822, A[11], A[17]);
  nand g576 (n_258, n_820, n_821, n_822);
  xor g577 (n_823, n_183, n_208);
  xor g578 (n_248, n_823, n_245);
  nand g579 (n_824, n_183, n_208);
  nand g580 (n_825, n_245, n_208);
  nand g581 (n_826, n_183, n_245);
  nand g582 (n_261, n_824, n_825, n_826);
  xor g583 (n_827, n_246, n_247);
  xor g584 (n_251, n_827, n_248);
  nand g585 (n_828, n_246, n_247);
  nand g586 (n_829, n_248, n_247);
  nand g587 (n_830, n_246, n_248);
  nand g588 (n_263, n_828, n_829, n_830);
  xor g589 (n_831, n_249, n_250);
  xor g590 (n_104, n_831, n_251);
  nand g591 (n_832, n_249, n_250);
  nand g592 (n_833, n_251, n_250);
  nand g593 (n_834, n_249, n_251);
  nand g594 (n_55, n_832, n_833, n_834);
  xor g604 (n_256, n_671, A[11]);
  nand g607 (n_842, n_185, A[11]);
  nand g608 (n_269, n_672, n_688, n_842);
  xor g609 (n_843, A[12], A[15]);
  xor g610 (n_259, n_843, n_186);
  nand g611 (n_844, A[12], A[15]);
  nand g612 (n_845, n_186, A[15]);
  nand g613 (n_846, A[12], n_186);
  nand g614 (n_270, n_844, n_845, n_846);
  xor g615 (n_847, A[16], A[18]);
  xor g616 (n_260, n_847, n_187);
  nand g617 (n_848, A[16], A[18]);
  nand g618 (n_849, n_187, A[18]);
  nand g619 (n_850, A[16], n_187);
  nand g620 (n_272, n_848, n_849, n_850);
  xor g621 (n_851, n_256, n_257);
  xor g622 (n_262, n_851, n_258);
  nand g623 (n_852, n_256, n_257);
  nand g624 (n_853, n_258, n_257);
  nand g625 (n_854, n_256, n_258);
  nand g626 (n_275, n_852, n_853, n_854);
  xor g627 (n_855, n_259, n_260);
  xor g628 (n_264, n_855, n_261);
  nand g629 (n_856, n_259, n_260);
  nand g630 (n_857, n_261, n_260);
  nand g631 (n_858, n_259, n_261);
  nand g632 (n_277, n_856, n_857, n_858);
  xor g633 (n_859, n_262, n_263);
  xor g634 (n_103, n_859, n_264);
  nand g635 (n_860, n_262, n_263);
  nand g636 (n_861, n_264, n_263);
  nand g637 (n_862, n_262, n_264);
  nand g638 (n_54, n_860, n_861, n_862);
  xor g642 (n_266, n_635, A[5]);
  nand g644 (n_865, A[5], A[4]);
  nand g645 (n_866, n_118, A[5]);
  nand g646 (n_281, n_636, n_865, n_866);
  xor g647 (n_867, n_174, n_266);
  xor g648 (n_268, n_867, A[9]);
  nand g649 (n_868, n_174, n_266);
  nand g650 (n_869, A[9], n_266);
  nand g651 (n_870, n_174, A[9]);
  nand g652 (n_283, n_868, n_869, n_870);
  xor g653 (n_871, A[8], A[12]);
  xor g654 (n_271, n_871, A[13]);
  nand g657 (n_874, A[8], A[13]);
  nand g658 (n_285, n_742, n_765, n_874);
  xor g659 (n_875, n_71, A[17]);
  xor g660 (n_274, n_875, A[19]);
  nand g661 (n_876, n_71, A[17]);
  nand g662 (n_877, A[19], A[17]);
  nand g663 (n_878, n_71, A[19]);
  nand g664 (n_287, n_876, n_877, n_878);
  xor g665 (n_879, A[16], n_268);
  xor g666 (n_273, n_879, n_269);
  nand g667 (n_880, A[16], n_268);
  nand g668 (n_881, n_269, n_268);
  nand g669 (n_882, A[16], n_269);
  nand g670 (n_288, n_880, n_881, n_882);
  xor g671 (n_883, n_270, n_271);
  xor g672 (n_276, n_883, n_272);
  nand g673 (n_884, n_270, n_271);
  nand g674 (n_885, n_272, n_271);
  nand g675 (n_886, n_270, n_272);
  nand g676 (n_291, n_884, n_885, n_886);
  xor g677 (n_887, n_273, n_274);
  xor g678 (n_278, n_887, n_275);
  nand g679 (n_888, n_273, n_274);
  nand g680 (n_889, n_275, n_274);
  nand g681 (n_890, n_273, n_275);
  nand g682 (n_294, n_888, n_889, n_890);
  xor g683 (n_891, n_276, n_277);
  xor g684 (n_102, n_891, n_278);
  nand g685 (n_892, n_276, n_277);
  nand g686 (n_893, n_278, n_277);
  nand g687 (n_894, n_276, n_278);
  nand g688 (n_53, n_892, n_893, n_894);
  xor g701 (n_903, n_281, A[10]);
  xor g702 (n_284, n_903, A[9]);
  nand g703 (n_904, n_281, A[10]);
  nand g705 (n_906, n_281, A[9]);
  nand g706 (n_299, n_904, n_705, n_906);
  xor g707 (n_907, A[13], n_199);
  xor g708 (n_286, n_907, A[14]);
  xor g713 (n_911, A[18], A[20]);
  xor g714 (n_289, n_911, A[17]);
  nand g715 (n_912, A[18], A[20]);
  nand g716 (n_913, A[17], A[20]);
  nand g717 (n_914, A[18], A[17]);
  nand g718 (n_303, n_912, n_913, n_914);
  xor g719 (n_915, n_283, n_284);
  xor g720 (n_290, n_915, n_285);
  nand g721 (n_916, n_283, n_284);
  nand g722 (n_917, n_285, n_284);
  nand g723 (n_918, n_283, n_285);
  nand g724 (n_305, n_916, n_917, n_918);
  xor g725 (n_919, n_286, n_287);
  xor g726 (n_292, n_919, n_288);
  nand g727 (n_920, n_286, n_287);
  nand g728 (n_921, n_288, n_287);
  nand g729 (n_922, n_286, n_288);
  nand g730 (n_307, n_920, n_921, n_922);
  xor g731 (n_923, n_289, n_290);
  xor g732 (n_293, n_923, n_291);
  nand g733 (n_924, n_289, n_290);
  nand g734 (n_925, n_291, n_290);
  nand g735 (n_926, n_289, n_291);
  nand g736 (n_309, n_924, n_925, n_926);
  xor g737 (n_927, n_292, n_293);
  xor g738 (n_101, n_927, n_294);
  nand g739 (n_928, n_292, n_293);
  nand g740 (n_929, n_294, n_293);
  nand g741 (n_930, n_292, n_294);
  nand g742 (n_52, n_928, n_929, n_930);
  xor g750 (n_298, n_659, A[10]);
  nand g752 (n_937, A[10], A[7]);
  nand g753 (n_938, n_68, A[10]);
  nand g754 (n_314, n_660, n_937, n_938);
  xor g755 (n_939, n_182, n_181);
  xor g756 (n_300, n_939, A[14]);
  nand g757 (n_940, n_182, n_181);
  nand g758 (n_941, A[14], n_181);
  nand g760 (n_316, n_940, n_941, n_818);
  xor g762 (n_302, n_819, A[19]);
  nand g764 (n_945, A[19], A[15]);
  nand g765 (n_946, A[11], A[19]);
  nand g766 (n_319, n_820, n_945, n_946);
  xor g767 (n_947, n_298, A[21]);
  xor g768 (n_304, n_947, A[18]);
  nand g769 (n_948, n_298, A[21]);
  nand g770 (n_949, A[18], A[21]);
  nand g771 (n_950, n_298, A[18]);
  nand g772 (n_318, n_948, n_949, n_950);
  xor g773 (n_951, n_299, n_300);
  xor g774 (n_306, n_951, n_245);
  nand g775 (n_952, n_299, n_300);
  nand g776 (n_953, n_245, n_300);
  nand g777 (n_954, n_299, n_245);
  nand g778 (n_321, n_952, n_953, n_954);
  xor g779 (n_955, n_302, n_303);
  xor g780 (n_308, n_955, n_304);
  nand g781 (n_956, n_302, n_303);
  nand g782 (n_957, n_304, n_303);
  nand g783 (n_958, n_302, n_304);
  nand g784 (n_324, n_956, n_957, n_958);
  xor g785 (n_959, n_305, n_306);
  xor g786 (n_310, n_959, n_307);
  nand g787 (n_960, n_305, n_306);
  nand g788 (n_961, n_307, n_306);
  nand g789 (n_962, n_305, n_307);
  nand g790 (n_326, n_960, n_961, n_962);
  xor g791 (n_963, n_308, n_309);
  xor g792 (n_100, n_963, n_310);
  nand g793 (n_964, n_308, n_309);
  nand g794 (n_965, n_310, n_309);
  nand g795 (n_966, n_308, n_310);
  nand g796 (n_51, n_964, n_965, n_966);
  xor g806 (n_315, n_671, A[12]);
  nand g808 (n_973, A[12], n_185);
  nand g810 (n_333, n_672, n_973, n_742);
  xor g811 (n_975, A[11], n_186);
  xor g812 (n_317, n_975, A[15]);
  nand g816 (n_335, n_745, n_845, n_820);
  xor g817 (n_979, A[20], A[16]);
  xor g818 (n_320, n_979, A[19]);
  nand g819 (n_980, A[20], A[16]);
  nand g820 (n_981, A[19], A[16]);
  nand g821 (n_982, A[20], A[19]);
  nand g822 (n_336, n_980, n_981, n_982);
  xor g823 (n_983, n_314, n_315);
  xor g824 (n_322, n_983, A[22]);
  nand g825 (n_984, n_314, n_315);
  nand g826 (n_985, A[22], n_315);
  nand g827 (n_986, n_314, A[22]);
  nand g828 (n_338, n_984, n_985, n_986);
  xor g829 (n_987, n_316, n_317);
  xor g830 (n_323, n_987, n_318);
  nand g831 (n_988, n_316, n_317);
  nand g832 (n_989, n_318, n_317);
  nand g833 (n_990, n_316, n_318);
  nand g834 (n_341, n_988, n_989, n_990);
  xor g835 (n_991, n_319, n_320);
  xor g836 (n_325, n_991, n_321);
  nand g837 (n_992, n_319, n_320);
  nand g838 (n_993, n_321, n_320);
  nand g839 (n_994, n_319, n_321);
  nand g840 (n_343, n_992, n_993, n_994);
  xor g841 (n_995, n_322, n_323);
  xor g842 (n_327, n_995, n_324);
  nand g843 (n_996, n_322, n_323);
  nand g844 (n_997, n_324, n_323);
  nand g845 (n_998, n_322, n_324);
  nand g846 (n_345, n_996, n_997, n_998);
  xor g847 (n_999, n_325, n_326);
  xor g848 (n_99, n_999, n_327);
  nand g849 (n_1000, n_325, n_326);
  nand g850 (n_1001, n_327, n_326);
  nand g851 (n_1002, n_325, n_327);
  nand g852 (n_50, n_1000, n_1001, n_1002);
  xor g862 (n_332, n_867, A[8]);
  nand g864 (n_1009, A[8], n_266);
  nand g865 (n_1010, n_174, A[8]);
  nand g866 (n_353, n_868, n_1009, n_1010);
  xor g873 (n_1015, n_71, n_332);
  xor g874 (n_337, n_1015, A[17]);
  nand g875 (n_1016, n_71, n_332);
  nand g876 (n_1017, A[17], n_332);
  nand g878 (n_358, n_1016, n_1017, n_876);
  xor g879 (n_1019, A[21], A[16]);
  xor g880 (n_339, n_1019, A[20]);
  nand g881 (n_1020, A[21], A[16]);
  nand g883 (n_1022, A[21], A[20]);
  nand g884 (n_357, n_1020, n_980, n_1022);
  xor g885 (n_1023, A[23], n_333);
  xor g886 (n_340, n_1023, n_223);
  nand g887 (n_1024, A[23], n_333);
  nand g888 (n_1025, n_223, n_333);
  nand g889 (n_1026, A[23], n_223);
  nand g890 (n_361, n_1024, n_1025, n_1026);
  xor g891 (n_1027, n_335, n_336);
  xor g892 (n_342, n_1027, n_337);
  nand g893 (n_1028, n_335, n_336);
  nand g894 (n_1029, n_337, n_336);
  nand g895 (n_1030, n_335, n_337);
  nand g896 (n_364, n_1028, n_1029, n_1030);
  xor g897 (n_1031, n_338, n_339);
  xor g898 (n_344, n_1031, n_340);
  nand g899 (n_1032, n_338, n_339);
  nand g900 (n_1033, n_340, n_339);
  nand g901 (n_1034, n_338, n_340);
  nand g902 (n_365, n_1032, n_1033, n_1034);
  xor g903 (n_1035, n_341, n_342);
  xor g904 (n_346, n_1035, n_343);
  nand g905 (n_1036, n_341, n_342);
  nand g906 (n_1037, n_343, n_342);
  nand g907 (n_1038, n_341, n_343);
  nand g908 (n_367, n_1036, n_1037, n_1038);
  xor g909 (n_1039, n_344, n_345);
  xor g910 (n_98, n_1039, n_346);
  nand g911 (n_1040, n_344, n_345);
  nand g912 (n_1041, n_346, n_345);
  nand g913 (n_1042, n_344, n_346);
  nand g914 (n_49, n_1040, n_1041, n_1042);
  xor g917 (n_1043, A[2], n_171);
  nand g922 (n_372, n_625, n_1045, n_1046);
  xor g924 (n_352, n_699, n_350);
  nand g926 (n_1049, n_350, A[6]);
  nand g927 (n_1050, A[5], n_350);
  nand g928 (n_374, n_650, n_1049, n_1050);
  xor g929 (n_1051, n_281, A[9]);
  xor g930 (n_354, n_1051, A[10]);
  xor g935 (n_1055, A[14], n_352);
  xor g936 (n_356, n_1055, A[13]);
  nand g937 (n_1056, A[14], n_352);
  nand g938 (n_1057, A[13], n_352);
  nand g940 (n_378, n_1056, n_1057, n_793);
  xor g942 (n_360, n_1059, A[18]);
  nand g944 (n_1061, A[18], n_353);
  nand g946 (n_380, n_1060, n_1061, n_1062);
  xor g947 (n_1063, A[17], A[21]);
  xor g948 (n_359, n_1063, A[22]);
  nand g949 (n_1064, A[17], A[21]);
  nand g950 (n_1065, A[22], A[21]);
  nand g951 (n_1066, A[17], A[22]);
  nand g952 (n_383, n_1064, n_1065, n_1066);
  xor g953 (n_1067, n_354, n_234);
  xor g954 (n_362, n_1067, n_356);
  nand g955 (n_1068, n_354, n_234);
  nand g956 (n_1069, n_356, n_234);
  nand g957 (n_1070, n_354, n_356);
  nand g958 (n_385, n_1068, n_1069, n_1070);
  xor g959 (n_1071, n_357, n_358);
  xor g960 (n_363, n_1071, n_359);
  nand g961 (n_1072, n_357, n_358);
  nand g962 (n_1073, n_359, n_358);
  nand g963 (n_1074, n_357, n_359);
  nand g964 (n_386, n_1072, n_1073, n_1074);
  xor g965 (n_1075, n_360, n_361);
  xor g966 (n_366, n_1075, n_362);
  nand g967 (n_1076, n_360, n_361);
  nand g968 (n_1077, n_362, n_361);
  nand g969 (n_1078, n_360, n_362);
  nand g970 (n_388, n_1076, n_1077, n_1078);
  xor g971 (n_1079, n_363, n_364);
  xor g972 (n_368, n_1079, n_365);
  nand g973 (n_1080, n_363, n_364);
  nand g974 (n_1081, n_365, n_364);
  nand g975 (n_1082, n_363, n_365);
  nand g976 (n_390, n_1080, n_1081, n_1082);
  xor g977 (n_1083, n_366, n_367);
  xor g978 (n_97, n_1083, n_368);
  nand g979 (n_1084, n_366, n_367);
  nand g980 (n_1085, n_368, n_367);
  nand g981 (n_1086, n_366, n_368);
  nand g982 (n_48, n_1084, n_1085, n_1086);
  xor g985 (n_1087, A[3], A[1]);
  nand g987 (n_1088, A[3], A[1]);
  nand g990 (n_393, n_1088, n_1089, n_1090);
  xor g991 (n_1091, A[6], n_372);
  xor g992 (n_375, n_1091, n_373);
  nand g993 (n_1092, A[6], n_372);
  nand g994 (n_1093, n_373, n_372);
  nand g995 (n_1094, A[6], n_373);
  nand g996 (n_395, n_1092, n_1093, n_1094);
  xor g997 (n_1095, A[7], A[10]);
  xor g998 (n_377, n_1095, A[14]);
  nand g1001 (n_1098, A[7], A[14]);
  nand g1002 (n_397, n_937, n_817, n_1098);
  xor g1003 (n_1099, n_374, n_375);
  xor g1004 (n_379, n_1099, A[11]);
  nand g1005 (n_1100, n_374, n_375);
  nand g1006 (n_1101, A[11], n_375);
  nand g1007 (n_1102, n_374, A[11]);
  nand g1008 (n_398, n_1100, n_1101, n_1102);
  xor g1009 (n_1103, A[15], n_299);
  xor g1010 (n_382, n_1103, A[23]);
  nand g1011 (n_1104, A[15], n_299);
  nand g1012 (n_1105, A[23], n_299);
  nand g1013 (n_1106, A[15], A[23]);
  nand g1014 (n_401, n_1104, n_1105, n_1106);
  xor g1015 (n_1107, A[18], A[19]);
  xor g1016 (n_381, n_1107, A[22]);
  nand g1017 (n_1108, A[18], A[19]);
  nand g1018 (n_1109, A[22], A[19]);
  nand g1019 (n_1110, A[18], A[22]);
  nand g1020 (n_404, n_1108, n_1109, n_1110);
  xor g1021 (n_1111, n_377, n_378);
  xor g1022 (n_384, n_1111, n_379);
  nand g1023 (n_1112, n_377, n_378);
  nand g1024 (n_1113, n_379, n_378);
  nand g1025 (n_1114, n_377, n_379);
  nand g1026 (n_405, n_1112, n_1113, n_1114);
  xor g1027 (n_1115, n_380, n_381);
  xor g1028 (n_387, n_1115, n_382);
  nand g1029 (n_1116, n_380, n_381);
  nand g1030 (n_1117, n_382, n_381);
  nand g1031 (n_1118, n_380, n_382);
  nand g1032 (n_407, n_1116, n_1117, n_1118);
  xor g1033 (n_1119, n_383, n_384);
  xor g1034 (n_389, n_1119, n_385);
  nand g1035 (n_1120, n_383, n_384);
  nand g1036 (n_1121, n_385, n_384);
  nand g1037 (n_1122, n_383, n_385);
  nand g1038 (n_409, n_1120, n_1121, n_1122);
  xor g1039 (n_1123, n_386, n_387);
  xor g1040 (n_391, n_1123, n_388);
  nand g1041 (n_1124, n_386, n_387);
  nand g1042 (n_1125, n_388, n_387);
  nand g1043 (n_1126, n_386, n_388);
  nand g1044 (n_411, n_1124, n_1125, n_1126);
  xor g1045 (n_1127, n_389, n_390);
  xor g1046 (n_96, n_1127, n_391);
  nand g1047 (n_1128, n_389, n_390);
  nand g1048 (n_1129, n_391, n_390);
  nand g1049 (n_1130, n_389, n_391);
  nand g1050 (n_47, n_1128, n_1129, n_1130);
  xor g1051 (n_1131, A[3], A[4]);
  xor g1052 (n_394, n_1131, A[2]);
  nand g1053 (n_1132, A[3], A[4]);
  nand g1054 (n_1133, A[2], A[4]);
  nand g1056 (n_413, n_1132, n_1133, n_628);
  xor g1057 (n_1135, n_393, A[7]);
  xor g1058 (n_396, n_1135, n_394);
  nand g1059 (n_1136, n_393, A[7]);
  nand g1060 (n_1137, n_394, A[7]);
  nand g1061 (n_1138, n_393, n_394);
  nand g1062 (n_415, n_1136, n_1137, n_1138);
  xor g1064 (n_399, n_687, A[12]);
  nand g1066 (n_1141, A[12], A[11]);
  nand g1068 (n_417, n_688, n_1141, n_742);
  xor g1070 (n_400, n_1143, A[15]);
  nand g1073 (n_1146, n_395, A[15]);
  nand g1074 (n_419, n_1144, n_1145, n_1146);
  xor g1075 (n_1147, A[19], A[23]);
  xor g1076 (n_403, n_1147, n_396);
  nand g1077 (n_1148, A[19], A[23]);
  nand g1078 (n_1149, n_396, A[23]);
  nand g1079 (n_1150, A[19], n_396);
  nand g1080 (n_420, n_1148, n_1149, n_1150);
  xor g1082 (n_402, n_979, n_397);
  nand g1084 (n_1153, n_397, A[20]);
  nand g1085 (n_1154, A[16], n_397);
  nand g1086 (n_421, n_980, n_1153, n_1154);
  xor g1087 (n_1155, n_398, n_399);
  xor g1088 (n_406, n_1155, n_400);
  nand g1089 (n_1156, n_398, n_399);
  nand g1090 (n_1157, n_400, n_399);
  nand g1091 (n_1158, n_398, n_400);
  nand g1092 (n_425, n_1156, n_1157, n_1158);
  xor g1093 (n_1159, n_401, n_402);
  xor g1094 (n_408, n_1159, n_403);
  nand g1095 (n_1160, n_401, n_402);
  nand g1096 (n_1161, n_403, n_402);
  nand g1097 (n_1162, n_401, n_403);
  nand g1098 (n_426, n_1160, n_1161, n_1162);
  xor g1099 (n_1163, n_404, n_405);
  xor g1100 (n_410, n_1163, n_406);
  nand g1101 (n_1164, n_404, n_405);
  nand g1102 (n_1165, n_406, n_405);
  nand g1103 (n_1166, n_404, n_406);
  nand g1104 (n_428, n_1164, n_1165, n_1166);
  xor g1105 (n_1167, n_407, n_408);
  xor g1106 (n_412, n_1167, n_409);
  nand g1107 (n_1168, n_407, n_408);
  nand g1108 (n_1169, n_409, n_408);
  nand g1109 (n_1170, n_407, n_409);
  nand g1110 (n_430, n_1168, n_1169, n_1170);
  xor g1111 (n_1171, n_410, n_411);
  xor g1112 (n_95, n_1171, n_412);
  nand g1113 (n_1172, n_410, n_411);
  nand g1114 (n_1173, n_412, n_411);
  nand g1115 (n_1174, n_410, n_412);
  nand g1116 (n_46, n_1172, n_1173, n_1174);
  xor g1117 (n_1175, A[4], A[5]);
  xor g1118 (n_414, n_1175, n_413);
  nand g1120 (n_1177, n_413, A[5]);
  nand g1121 (n_1178, A[4], n_413);
  nand g1122 (n_434, n_865, n_1177, n_1178);
  xor g1123 (n_1179, A[9], A[8]);
  xor g1124 (n_416, n_1179, A[13]);
  nand g1125 (n_1180, A[9], A[8]);
  nand g1128 (n_436, n_1180, n_874, n_764);
  xor g1129 (n_1183, n_414, A[12]);
  xor g1130 (n_418, n_1183, n_415);
  nand g1131 (n_1184, n_414, A[12]);
  nand g1132 (n_1185, n_415, A[12]);
  nand g1133 (n_1186, n_414, n_415);
  nand g1134 (n_438, n_1184, n_1185, n_1186);
  xor g1136 (n_422, n_1187, A[21]);
  nand g1140 (n_439, n_1188, n_1064, n_1190);
  xor g1142 (n_423, n_979, n_416);
  nand g1144 (n_1193, n_416, A[20]);
  nand g1145 (n_1194, A[16], n_416);
  nand g1146 (n_440, n_980, n_1193, n_1194);
  xor g1147 (n_1195, n_417, n_418);
  xor g1148 (n_424, n_1195, n_419);
  nand g1149 (n_1196, n_417, n_418);
  nand g1150 (n_1197, n_419, n_418);
  nand g1151 (n_1198, n_417, n_419);
  nand g1152 (n_443, n_1196, n_1197, n_1198);
  xor g1153 (n_1199, n_420, n_421);
  xor g1154 (n_427, n_1199, n_422);
  nand g1155 (n_1200, n_420, n_421);
  nand g1156 (n_1201, n_422, n_421);
  nand g1157 (n_1202, n_420, n_422);
  nand g1158 (n_445, n_1200, n_1201, n_1202);
  xor g1159 (n_1203, n_423, n_424);
  xor g1160 (n_429, n_1203, n_425);
  nand g1161 (n_1204, n_423, n_424);
  nand g1162 (n_1205, n_425, n_424);
  nand g1163 (n_1206, n_423, n_425);
  nand g1164 (n_447, n_1204, n_1205, n_1206);
  xor g1165 (n_1207, n_426, n_427);
  xor g1166 (n_431, n_1207, n_428);
  nand g1167 (n_1208, n_426, n_427);
  nand g1168 (n_1209, n_428, n_427);
  nand g1169 (n_1210, n_426, n_428);
  nand g1170 (n_450, n_1208, n_1209, n_1210);
  xor g1171 (n_1211, n_429, n_430);
  xor g1172 (n_94, n_1211, n_431);
  nand g1173 (n_1212, n_429, n_430);
  nand g1174 (n_1213, n_431, n_430);
  nand g1175 (n_1214, n_429, n_431);
  nand g1176 (n_45, n_1212, n_1213, n_1214);
  nand g1183 (n_1218, A[6], A[9]);
  nand g1184 (n_455, n_1216, n_1217, n_1218);
  xor g1185 (n_1219, A[10], A[14]);
  xor g1186 (n_437, n_1219, n_434);
  nand g1188 (n_1221, n_434, A[14]);
  nand g1189 (n_1222, A[10], n_434);
  nand g1190 (n_456, n_817, n_1221, n_1222);
  xor g1191 (n_1223, A[13], A[21]);
  xor g1192 (n_442, n_1223, n_435);
  nand g1193 (n_1224, A[13], A[21]);
  nand g1194 (n_1225, n_435, A[21]);
  nand g1195 (n_1226, A[13], n_435);
  nand g1196 (n_458, n_1224, n_1225, n_1226);
  xor g1197 (n_1227, A[17], A[18]);
  xor g1198 (n_441, n_1227, A[22]);
  nand g1202 (n_461, n_914, n_1110, n_1066);
  xor g1203 (n_1231, n_436, n_437);
  xor g1204 (n_444, n_1231, n_438);
  nand g1205 (n_1232, n_436, n_437);
  nand g1206 (n_1233, n_438, n_437);
  nand g1207 (n_1234, n_436, n_438);
  nand g1208 (n_462, n_1232, n_1233, n_1234);
  xor g1209 (n_1235, n_439, n_440);
  xor g1210 (n_446, n_1235, n_441);
  nand g1211 (n_1236, n_439, n_440);
  nand g1212 (n_1237, n_441, n_440);
  nand g1213 (n_1238, n_439, n_441);
  nand g1214 (n_464, n_1236, n_1237, n_1238);
  xor g1215 (n_1239, n_442, n_443);
  xor g1216 (n_448, n_1239, n_444);
  nand g1217 (n_1240, n_442, n_443);
  nand g1218 (n_1241, n_444, n_443);
  nand g1219 (n_1242, n_442, n_444);
  nand g1220 (n_467, n_1240, n_1241, n_1242);
  xor g1221 (n_1243, n_445, n_446);
  xor g1222 (n_449, n_1243, n_447);
  nand g1223 (n_1244, n_445, n_446);
  nand g1224 (n_1245, n_447, n_446);
  nand g1225 (n_1246, n_445, n_447);
  nand g1226 (n_469, n_1244, n_1245, n_1246);
  xor g1227 (n_1247, n_448, n_449);
  xor g1228 (n_93, n_1247, n_450);
  nand g1229 (n_1248, n_448, n_449);
  nand g1230 (n_1249, n_450, n_449);
  nand g1231 (n_1250, n_448, n_450);
  nand g1232 (n_44, n_1248, n_1249, n_1250);
  xor g1235 (n_1251, A[5], A[7]);
  nand g1240 (n_471, n_642, n_1253, n_1254);
  xor g1242 (n_457, n_1219, A[11]);
  nand g1246 (n_473, n_817, n_744, n_725);
  xor g1247 (n_1259, A[15], A[23]);
  xor g1248 (n_460, n_1259, n_454);
  nand g1250 (n_1261, n_454, A[23]);
  nand g1251 (n_1262, A[15], n_454);
  nand g1252 (n_477, n_1106, n_1261, n_1262);
  xor g1254 (n_459, n_1107, n_455);
  nand g1256 (n_1265, n_455, A[19]);
  nand g1257 (n_1266, A[18], n_455);
  nand g1258 (n_475, n_1108, n_1265, n_1266);
  xor g1259 (n_1267, A[22], n_456);
  xor g1260 (n_463, n_1267, n_457);
  nand g1261 (n_1268, A[22], n_456);
  nand g1262 (n_1269, n_457, n_456);
  nand g1263 (n_1270, A[22], n_457);
  nand g1264 (n_479, n_1268, n_1269, n_1270);
  xor g1265 (n_1271, n_458, n_459);
  xor g1266 (n_465, n_1271, n_460);
  nand g1267 (n_1272, n_458, n_459);
  nand g1268 (n_1273, n_460, n_459);
  nand g1269 (n_1274, n_458, n_460);
  nand g1270 (n_482, n_1272, n_1273, n_1274);
  xor g1271 (n_1275, n_461, n_462);
  xor g1272 (n_466, n_1275, n_463);
  nand g1273 (n_1276, n_461, n_462);
  nand g1274 (n_1277, n_463, n_462);
  nand g1275 (n_1278, n_461, n_463);
  nand g1276 (n_483, n_1276, n_1277, n_1278);
  xor g1277 (n_1279, n_464, n_465);
  xor g1278 (n_468, n_1279, n_466);
  nand g1279 (n_1280, n_464, n_465);
  nand g1280 (n_1281, n_466, n_465);
  nand g1281 (n_1282, n_464, n_466);
  nand g1282 (n_486, n_1280, n_1281, n_1282);
  xor g1283 (n_1283, n_467, n_468);
  xor g1284 (n_92, n_1283, n_469);
  nand g1285 (n_1284, n_467, n_468);
  nand g1286 (n_1285, n_469, n_468);
  nand g1287 (n_1286, n_467, n_469);
  nand g1288 (n_43, n_1284, n_1285, n_1286);
  xor g1290 (n_472, n_719, A[8]);
  nand g1292 (n_1289, A[8], A[6]);
  nand g1293 (n_1290, A[7], A[8]);
  nand g1294 (n_487, n_720, n_1289, n_1290);
  xor g1295 (n_1291, A[11], A[12]);
  nand g1300 (n_489, n_1141, n_1293, n_1294);
  xor g1301 (n_1295, n_471, A[15]);
  xor g1302 (n_476, n_1295, n_472);
  nand g1303 (n_1296, n_471, A[15]);
  nand g1304 (n_1297, n_472, A[15]);
  nand g1305 (n_1298, n_471, n_472);
  nand g1306 (n_491, n_1296, n_1297, n_1298);
  xor g1308 (n_478, n_1147, A[16]);
  nand g1310 (n_1301, A[16], A[23]);
  nand g1312 (n_490, n_1148, n_1301, n_981);
  xor g1313 (n_1303, A[20], n_473);
  xor g1314 (n_480, n_1303, n_474);
  nand g1315 (n_1304, A[20], n_473);
  nand g1316 (n_1305, n_474, n_473);
  nand g1317 (n_1306, A[20], n_474);
  nand g1318 (n_494, n_1304, n_1305, n_1306);
  xor g1319 (n_1307, n_475, n_476);
  xor g1320 (n_481, n_1307, n_477);
  nand g1321 (n_1308, n_475, n_476);
  nand g1322 (n_1309, n_477, n_476);
  nand g1323 (n_1310, n_475, n_477);
  nand g1324 (n_496, n_1308, n_1309, n_1310);
  xor g1325 (n_1311, n_478, n_479);
  xor g1326 (n_484, n_1311, n_480);
  nand g1327 (n_1312, n_478, n_479);
  nand g1328 (n_1313, n_480, n_479);
  nand g1329 (n_1314, n_478, n_480);
  nand g1330 (n_498, n_1312, n_1313, n_1314);
  xor g1331 (n_1315, n_481, n_482);
  xor g1332 (n_485, n_1315, n_483);
  nand g1333 (n_1316, n_481, n_482);
  nand g1334 (n_1317, n_483, n_482);
  nand g1335 (n_1318, n_481, n_483);
  nand g1336 (n_501, n_1316, n_1317, n_1318);
  xor g1337 (n_1319, n_484, n_485);
  xor g1338 (n_91, n_1319, n_486);
  nand g1339 (n_1320, n_484, n_485);
  nand g1340 (n_1321, n_486, n_485);
  nand g1341 (n_1322, n_484, n_486);
  nand g1342 (n_42, n_1320, n_1321, n_1322);
  xor g1350 (n_492, n_1327, A[17]);
  nand g1353 (n_1330, A[12], A[17]);
  nand g1354 (n_506, n_1293, n_1188, n_1330);
  xor g1356 (n_493, n_1019, n_487);
  nand g1358 (n_1333, n_487, A[16]);
  nand g1359 (n_1334, A[21], n_487);
  nand g1360 (n_507, n_1020, n_1333, n_1334);
  xor g1361 (n_1335, A[20], n_416);
  xor g1362 (n_495, n_1335, n_489);
  nand g1364 (n_1337, n_489, n_416);
  nand g1365 (n_1338, A[20], n_489);
  nand g1366 (n_509, n_1193, n_1337, n_1338);
  xor g1367 (n_1339, n_490, n_491);
  xor g1368 (n_497, n_1339, n_492);
  nand g1369 (n_1340, n_490, n_491);
  nand g1370 (n_1341, n_492, n_491);
  nand g1371 (n_1342, n_490, n_492);
  nand g1372 (n_511, n_1340, n_1341, n_1342);
  xor g1373 (n_1343, n_493, n_494);
  xor g1374 (n_499, n_1343, n_495);
  nand g1375 (n_1344, n_493, n_494);
  nand g1376 (n_1345, n_495, n_494);
  nand g1377 (n_1346, n_493, n_495);
  nand g1378 (n_513, n_1344, n_1345, n_1346);
  xor g1379 (n_1347, n_496, n_497);
  xor g1380 (n_500, n_1347, n_498);
  nand g1381 (n_1348, n_496, n_497);
  nand g1382 (n_1349, n_498, n_497);
  nand g1383 (n_1350, n_496, n_498);
  nand g1384 (n_516, n_1348, n_1349, n_1350);
  xor g1385 (n_1351, n_499, n_500);
  xor g1386 (n_90, n_1351, n_501);
  nand g1387 (n_1352, n_499, n_500);
  nand g1388 (n_1353, n_501, n_500);
  nand g1389 (n_1354, n_499, n_501);
  nand g1390 (n_41, n_1352, n_1353, n_1354);
  xor g1393 (n_1355, A[9], A[14]);
  xor g1394 (n_505, n_1355, A[13]);
  nand g1395 (n_1356, A[9], A[14]);
  nand g1398 (n_520, n_1356, n_793, n_764);
  xor g1400 (n_508, n_1359, A[17]);
  nand g1404 (n_522, n_1360, n_1064, n_1362);
  xor g1405 (n_1363, A[18], A[22]);
  xor g1406 (n_510, n_1363, n_436);
  nand g1408 (n_1365, n_436, A[22]);
  nand g1409 (n_1366, A[18], n_436);
  nand g1410 (n_524, n_1110, n_1365, n_1366);
  xor g1411 (n_1367, n_505, n_506);
  xor g1412 (n_512, n_1367, n_507);
  nand g1413 (n_1368, n_505, n_506);
  nand g1414 (n_1369, n_507, n_506);
  nand g1415 (n_1370, n_505, n_507);
  nand g1416 (n_527, n_1368, n_1369, n_1370);
  xor g1417 (n_1371, n_508, n_509);
  xor g1418 (n_514, n_1371, n_510);
  nand g1419 (n_1372, n_508, n_509);
  nand g1420 (n_1373, n_510, n_509);
  nand g1421 (n_1374, n_508, n_510);
  nand g1422 (n_529, n_1372, n_1373, n_1374);
  xor g1423 (n_1375, n_511, n_512);
  xor g1424 (n_515, n_1375, n_513);
  nand g1425 (n_1376, n_511, n_512);
  nand g1426 (n_1377, n_513, n_512);
  nand g1427 (n_1378, n_511, n_513);
  nand g1428 (n_531, n_1376, n_1377, n_1378);
  xor g1429 (n_1379, n_514, n_515);
  xor g1430 (n_89, n_1379, n_516);
  nand g1431 (n_1380, n_514, n_515);
  nand g1432 (n_1381, n_516, n_515);
  nand g1433 (n_1382, n_514, n_516);
  nand g1434 (n_40, n_1380, n_1381, n_1382);
  xor g1438 (n_521, n_743, A[10]);
  xor g1444 (n_523, n_1387, A[23]);
  nand g1448 (n_535, n_1388, n_1106, n_1390);
  xor g1450 (n_525, n_1107, n_520);
  nand g1452 (n_1393, n_520, A[19]);
  nand g1453 (n_1394, A[18], n_520);
  nand g1454 (n_538, n_1108, n_1393, n_1394);
  xor g1455 (n_1395, A[22], n_521);
  xor g1456 (n_526, n_1395, n_522);
  nand g1457 (n_1396, A[22], n_521);
  nand g1458 (n_1397, n_522, n_521);
  nand g1459 (n_1398, A[22], n_522);
  nand g1460 (n_540, n_1396, n_1397, n_1398);
  xor g1461 (n_1399, n_523, n_524);
  xor g1462 (n_528, n_1399, n_525);
  nand g1463 (n_1400, n_523, n_524);
  nand g1464 (n_1401, n_525, n_524);
  nand g1465 (n_1402, n_523, n_525);
  nand g1466 (n_541, n_1400, n_1401, n_1402);
  xor g1467 (n_1403, n_526, n_527);
  xor g1468 (n_530, n_1403, n_528);
  nand g1469 (n_1404, n_526, n_527);
  nand g1470 (n_1405, n_528, n_527);
  nand g1471 (n_1406, n_526, n_528);
  nand g1472 (n_544, n_1404, n_1405, n_1406);
  xor g1473 (n_1407, n_529, n_530);
  xor g1474 (n_88, n_1407, n_531);
  nand g1475 (n_1408, n_529, n_530);
  nand g1476 (n_1409, n_531, n_530);
  nand g1477 (n_1410, n_529, n_531);
  nand g1478 (n_39, n_1408, n_1409, n_1410);
  xor g1480 (n_534, n_1291, A[10]);
  nand g1483 (n_1414, A[12], A[10]);
  nand g1484 (n_545, n_1141, n_725, n_1414);
  xor g1486 (n_536, n_1415, A[19]);
  nand g1490 (n_547, n_1145, n_945, n_1418);
  xor g1491 (n_1419, A[23], A[16]);
  xor g1492 (n_537, n_1419, A[20]);
  nand g1495 (n_1422, A[23], A[20]);
  nand g1496 (n_548, n_1301, n_980, n_1422);
  xor g1497 (n_1423, n_473, n_534);
  xor g1498 (n_539, n_1423, n_535);
  nand g1499 (n_1424, n_473, n_534);
  nand g1500 (n_1425, n_535, n_534);
  nand g1501 (n_1426, n_473, n_535);
  nand g1502 (n_551, n_1424, n_1425, n_1426);
  xor g1503 (n_1427, n_536, n_537);
  xor g1504 (n_542, n_1427, n_538);
  nand g1505 (n_1428, n_536, n_537);
  nand g1506 (n_1429, n_538, n_537);
  nand g1507 (n_1430, n_536, n_538);
  nand g1508 (n_552, n_1428, n_1429, n_1430);
  xor g1509 (n_1431, n_539, n_540);
  xor g1510 (n_543, n_1431, n_541);
  nand g1511 (n_1432, n_539, n_540);
  nand g1512 (n_1433, n_541, n_540);
  nand g1513 (n_1434, n_539, n_541);
  nand g1514 (n_555, n_1432, n_1433, n_1434);
  xor g1515 (n_1435, n_542, n_543);
  xor g1516 (n_87, n_1435, n_544);
  nand g1517 (n_1436, n_542, n_543);
  nand g1518 (n_1437, n_544, n_543);
  nand g1519 (n_1438, n_542, n_544);
  nand g1520 (n_38, n_1436, n_1437, n_1438);
  xor g1521 (n_1439, A[13], A[12]);
  nand g1526 (n_558, n_765, n_1293, n_1442);
  xor g1528 (n_549, n_1063, A[16]);
  nand g1530 (n_1445, A[16], A[17]);
  nand g1532 (n_559, n_1064, n_1445, n_1020);
  xor g1533 (n_1447, A[20], n_545);
  xor g1534 (n_550, n_1447, n_546);
  nand g1535 (n_1448, A[20], n_545);
  nand g1536 (n_1449, n_546, n_545);
  nand g1537 (n_1450, A[20], n_546);
  nand g1538 (n_562, n_1448, n_1449, n_1450);
  xor g1539 (n_1451, n_547, n_548);
  xor g1540 (n_553, n_1451, n_549);
  nand g1541 (n_1452, n_547, n_548);
  nand g1542 (n_1453, n_549, n_548);
  nand g1543 (n_1454, n_547, n_549);
  nand g1544 (n_563, n_1452, n_1453, n_1454);
  xor g1545 (n_1455, n_550, n_551);
  xor g1546 (n_554, n_1455, n_552);
  nand g1547 (n_1456, n_550, n_551);
  nand g1548 (n_1457, n_552, n_551);
  nand g1549 (n_1458, n_550, n_552);
  nand g1550 (n_566, n_1456, n_1457, n_1458);
  xor g1551 (n_1459, n_553, n_554);
  xor g1552 (n_86, n_1459, n_555);
  nand g1553 (n_1460, n_553, n_554);
  nand g1554 (n_1461, n_555, n_554);
  nand g1555 (n_1462, n_553, n_555);
  nand g1556 (n_37, n_1460, n_1461, n_1462);
  xor g1560 (n_561, n_1223, A[17]);
  nand g1563 (n_1466, A[13], A[17]);
  nand g1564 (n_570, n_1224, n_1064, n_1466);
  xor g1566 (n_560, n_1467, A[22]);
  nand g1570 (n_572, n_1468, n_1469, n_1110);
  xor g1571 (n_1471, n_558, n_559);
  xor g1572 (n_564, n_1471, n_560);
  nand g1573 (n_1472, n_558, n_559);
  nand g1574 (n_1473, n_560, n_559);
  nand g1575 (n_1474, n_558, n_560);
  nand g1576 (n_574, n_1472, n_1473, n_1474);
  xor g1577 (n_1475, n_561, n_562);
  xor g1578 (n_565, n_1475, n_563);
  nand g1579 (n_1476, n_561, n_562);
  nand g1580 (n_1477, n_563, n_562);
  nand g1581 (n_1478, n_561, n_563);
  nand g1582 (n_577, n_1476, n_1477, n_1478);
  xor g1583 (n_1479, n_564, n_565);
  xor g1584 (n_85, n_1479, n_566);
  nand g1585 (n_1480, n_564, n_565);
  nand g1586 (n_1481, n_566, n_565);
  nand g1587 (n_1482, n_564, n_566);
  nand g1588 (n_36, n_1480, n_1481, n_1482);
  xor g1592 (n_573, n_1259, A[14]);
  nand g1594 (n_1485, A[14], A[23]);
  nand g1595 (n_1486, A[15], A[14]);
  nand g1596 (n_579, n_1106, n_1485, n_1486);
  nand g1602 (n_580, n_1108, n_1489, n_1468);
  xor g1603 (n_1491, A[22], n_570);
  xor g1604 (n_575, n_1491, n_571);
  nand g1605 (n_1492, A[22], n_570);
  nand g1606 (n_1493, n_571, n_570);
  nand g1607 (n_1494, A[22], n_571);
  nand g1608 (n_584, n_1492, n_1493, n_1494);
  xor g1609 (n_1495, n_572, n_573);
  xor g1610 (n_576, n_1495, n_574);
  nand g1611 (n_1496, n_572, n_573);
  nand g1612 (n_1497, n_574, n_573);
  nand g1613 (n_1498, n_572, n_574);
  nand g1614 (n_586, n_1496, n_1497, n_1498);
  xor g1615 (n_1499, n_575, n_576);
  xor g1616 (n_84, n_1499, n_577);
  nand g1617 (n_1500, n_575, n_576);
  nand g1618 (n_1501, n_577, n_576);
  nand g1619 (n_1502, n_575, n_577);
  nand g1620 (n_35, n_1500, n_1501, n_1502);
  xor g1622 (n_581, n_1415, A[23]);
  nand g1626 (n_588, n_1145, n_1106, n_1506);
  xor g1627 (n_1507, A[19], A[16]);
  xor g1628 (n_582, n_1507, A[20]);
  xor g1633 (n_1511, A[14], n_579);
  xor g1634 (n_583, n_1511, n_580);
  nand g1635 (n_1512, A[14], n_579);
  nand g1636 (n_1513, n_580, n_579);
  nand g1637 (n_1514, A[14], n_580);
  nand g1638 (n_590, n_1512, n_1513, n_1514);
  xor g1639 (n_1515, n_581, n_582);
  xor g1640 (n_585, n_1515, n_583);
  nand g1641 (n_1516, n_581, n_582);
  nand g1642 (n_1517, n_583, n_582);
  nand g1643 (n_1518, n_581, n_583);
  nand g1644 (n_593, n_1516, n_1517, n_1518);
  xor g1645 (n_1519, n_584, n_585);
  xor g1646 (n_83, n_1519, n_586);
  nand g1647 (n_1520, n_584, n_585);
  nand g1648 (n_1521, n_586, n_585);
  nand g1649 (n_1522, n_584, n_586);
  nand g1650 (n_34, n_1520, n_1521, n_1522);
  xor g1652 (n_589, n_1523, A[17]);
  xor g1658 (n_591, n_979, n_336);
  nand g1660 (n_1529, n_336, A[20]);
  nand g1661 (n_1530, A[16], n_336);
  nand g1662 (n_598, n_980, n_1529, n_1530);
  xor g1663 (n_1531, n_588, n_589);
  xor g1664 (n_592, n_1531, n_590);
  nand g1665 (n_1532, n_588, n_589);
  nand g1666 (n_1533, n_590, n_589);
  nand g1667 (n_1534, n_588, n_590);
  nand g1668 (n_600, n_1532, n_1533, n_1534);
  xor g1669 (n_1535, n_591, n_592);
  xor g1670 (n_82, n_1535, n_593);
  nand g1671 (n_1536, n_591, n_592);
  nand g1672 (n_1537, n_593, n_592);
  nand g1673 (n_1538, n_591, n_593);
  nand g1674 (n_81, n_1536, n_1537, n_1538);
  xor g1684 (n_599, n_1543, n_441);
  nand g1688 (n_607, n_1544, n_1238, n_1546);
  xor g1689 (n_1547, n_598, n_599);
  xor g1690 (n_33, n_1547, n_600);
  nand g1691 (n_1548, n_598, n_599);
  nand g1692 (n_1549, n_600, n_599);
  nand g1693 (n_1550, n_598, n_600);
  nand g1694 (n_80, n_1548, n_1549, n_1550);
  xor g1704 (n_606, n_1555, n_461);
  nand g1706 (n_1557, n_461, A[21]);
  nand g1708 (n_612, n_1556, n_1557, n_1558);
  xor g1709 (n_1559, n_381, n_606);
  xor g1710 (n_32, n_1559, n_607);
  nand g1711 (n_1560, n_381, n_606);
  nand g1712 (n_1561, n_607, n_606);
  nand g1713 (n_1562, n_381, n_607);
  nand g1714 (n_31, n_1560, n_1561, n_1562);
  xor g1716 (n_609, n_1563, A[19]);
  nand g1720 (n_613, n_1506, n_1148, n_1418);
  xor g1721 (n_1567, A[20], A[23]);
  xor g1722 (n_611, n_1567, n_609);
  nand g1724 (n_1569, n_609, A[23]);
  nand g1725 (n_1570, A[20], n_609);
  nand g1726 (n_615, n_1422, n_1569, n_1570);
  xor g1727 (n_1571, n_404, n_611);
  xor g1728 (n_79, n_1571, n_612);
  nand g1729 (n_1572, n_404, n_611);
  nand g1730 (n_1573, n_612, n_611);
  nand g1731 (n_1574, n_404, n_612);
  nand g1732 (n_30, n_1572, n_1573, n_1574);
  xor g1734 (n_614, n_1523, A[20]);
  nand g1738 (n_618, n_1190, n_1022, n_1578);
  xor g1739 (n_1579, n_613, n_614);
  xor g1740 (n_78, n_1579, n_615);
  nand g1741 (n_1580, n_613, n_614);
  nand g1742 (n_1581, n_615, n_614);
  nand g1743 (n_1582, n_613, n_615);
  nand g1744 (n_77, n_1580, n_1581, n_1582);
  xor g1748 (n_29, n_1583, n_618);
  nand g1751 (n_1586, A[22], n_618);
  nand g1752 (n_28, n_1584, n_1585, n_1586);
  xor g1756 (n_76, n_1587, A[21]);
  nand g1760 (n_27, n_1588, n_1556, n_1065);
  xor g1762 (n_75, n_1563, A[23]);
  nor g11 (n_1610, A[0], A[2]);
  nand g12 (n_1605, A[0], A[2]);
  nor g13 (n_1606, A[3], n_118);
  nand g14 (n_1607, A[3], n_118);
  nor g15 (n_1616, A[4], n_117);
  nand g16 (n_1611, A[4], n_117);
  nor g17 (n_1612, n_68, n_116);
  nand g18 (n_1613, n_68, n_116);
  nor g19 (n_1622, n_67, n_115);
  nand g20 (n_1617, n_67, n_115);
  nor g21 (n_1618, n_66, n_114);
  nand g22 (n_1619, n_66, n_114);
  nor g23 (n_1628, n_65, n_113);
  nand g24 (n_1623, n_65, n_113);
  nor g25 (n_1624, n_64, n_112);
  nand g26 (n_1625, n_64, n_112);
  nor g27 (n_1634, n_63, n_111);
  nand g28 (n_1629, n_63, n_111);
  nor g29 (n_1630, n_62, n_110);
  nand g30 (n_1631, n_62, n_110);
  nor g31 (n_1640, n_61, n_109);
  nand g32 (n_1635, n_61, n_109);
  nor g33 (n_1636, n_60, n_108);
  nand g34 (n_1637, n_60, n_108);
  nor g35 (n_1646, n_59, n_107);
  nand g36 (n_1641, n_59, n_107);
  nor g37 (n_1642, n_58, n_106);
  nand g38 (n_1643, n_58, n_106);
  nor g39 (n_1652, n_57, n_105);
  nand g40 (n_1647, n_57, n_105);
  nor g41 (n_1648, n_56, n_104);
  nand g42 (n_1649, n_56, n_104);
  nor g43 (n_1658, n_55, n_103);
  nand g44 (n_1653, n_55, n_103);
  nor g45 (n_1654, n_54, n_102);
  nand g46 (n_1655, n_54, n_102);
  nor g47 (n_1664, n_53, n_101);
  nand g48 (n_1659, n_53, n_101);
  nor g49 (n_1660, n_52, n_100);
  nand g50 (n_1661, n_52, n_100);
  nor g51 (n_1670, n_51, n_99);
  nand g52 (n_1665, n_51, n_99);
  nor g53 (n_1666, n_50, n_98);
  nand g54 (n_1667, n_50, n_98);
  nor g55 (n_1676, n_49, n_97);
  nand g56 (n_1671, n_49, n_97);
  nor g57 (n_1672, n_48, n_96);
  nand g58 (n_1673, n_48, n_96);
  nor g59 (n_1682, n_47, n_95);
  nand g60 (n_1677, n_47, n_95);
  nor g61 (n_1678, n_46, n_94);
  nand g62 (n_1679, n_46, n_94);
  nor g63 (n_1688, n_45, n_93);
  nand g64 (n_1683, n_45, n_93);
  nor g65 (n_1684, n_44, n_92);
  nand g66 (n_1685, n_44, n_92);
  nor g67 (n_1694, n_43, n_91);
  nand g68 (n_1689, n_43, n_91);
  nor g69 (n_1690, n_42, n_90);
  nand g70 (n_1691, n_42, n_90);
  nor g71 (n_1700, n_41, n_89);
  nand g72 (n_1695, n_41, n_89);
  nor g73 (n_1696, n_40, n_88);
  nand g74 (n_1697, n_40, n_88);
  nor g75 (n_1706, n_39, n_87);
  nand g76 (n_1701, n_39, n_87);
  nor g77 (n_1702, n_38, n_86);
  nand g78 (n_1703, n_38, n_86);
  nor g79 (n_1712, n_37, n_85);
  nand g80 (n_1707, n_37, n_85);
  nor g81 (n_1708, n_36, n_84);
  nand g82 (n_1709, n_36, n_84);
  nor g83 (n_1718, n_35, n_83);
  nand g84 (n_1713, n_35, n_83);
  nor g85 (n_1714, n_34, n_82);
  nand g86 (n_1715, n_34, n_82);
  nor g87 (n_1724, n_33, n_81);
  nand g88 (n_1719, n_33, n_81);
  nor g89 (n_1720, n_32, n_80);
  nand g90 (n_1721, n_32, n_80);
  nor g91 (n_1730, n_31, n_79);
  nand g92 (n_1725, n_31, n_79);
  nor g93 (n_1726, n_30, n_78);
  nand g94 (n_1727, n_30, n_78);
  nor g95 (n_1736, n_29, n_77);
  nand g96 (n_1731, n_29, n_77);
  nor g97 (n_1732, n_28, n_76);
  nand g98 (n_1733, n_28, n_76);
  nor g99 (n_1740, n_27, n_75);
  nand g100 (n_1737, n_27, n_75);
  nor g106 (n_1608, n_1605, n_1606);
  nor g110 (n_1614, n_1611, n_1612);
  nor g113 (n_1750, n_1616, n_1612);
  nor g114 (n_1620, n_1617, n_1618);
  nor g117 (n_1752, n_1622, n_1618);
  nor g118 (n_1626, n_1623, n_1624);
  nor g121 (n_1760, n_1628, n_1624);
  nor g122 (n_1632, n_1629, n_1630);
  nor g125 (n_1762, n_1634, n_1630);
  nor g126 (n_1638, n_1635, n_1636);
  nor g129 (n_1770, n_1640, n_1636);
  nor g130 (n_1644, n_1641, n_1642);
  nor g133 (n_1772, n_1646, n_1642);
  nor g134 (n_1650, n_1647, n_1648);
  nor g137 (n_1780, n_1652, n_1648);
  nor g138 (n_1656, n_1653, n_1654);
  nor g141 (n_1782, n_1658, n_1654);
  nor g142 (n_1662, n_1659, n_1660);
  nor g145 (n_1790, n_1664, n_1660);
  nor g146 (n_1668, n_1665, n_1666);
  nor g149 (n_1792, n_1670, n_1666);
  nor g150 (n_1674, n_1671, n_1672);
  nor g153 (n_1800, n_1676, n_1672);
  nor g154 (n_1680, n_1677, n_1678);
  nor g157 (n_1802, n_1682, n_1678);
  nor g158 (n_1686, n_1683, n_1684);
  nor g161 (n_1810, n_1688, n_1684);
  nor g162 (n_1692, n_1689, n_1690);
  nor g165 (n_1812, n_1694, n_1690);
  nor g166 (n_1698, n_1695, n_1696);
  nor g169 (n_1820, n_1700, n_1696);
  nor g170 (n_1704, n_1701, n_1702);
  nor g173 (n_1822, n_1706, n_1702);
  nor g174 (n_1710, n_1707, n_1708);
  nor g177 (n_1830, n_1712, n_1708);
  nor g178 (n_1716, n_1713, n_1714);
  nor g181 (n_1832, n_1718, n_1714);
  nor g182 (n_1722, n_1719, n_1720);
  nor g185 (n_1840, n_1724, n_1720);
  nor g186 (n_1728, n_1725, n_1726);
  nor g189 (n_1842, n_1730, n_1726);
  nor g190 (n_1734, n_1731, n_1732);
  nor g193 (n_1850, n_1736, n_1732);
  nor g203 (n_1748, n_1622, n_1747);
  nand g212 (n_1860, n_1750, n_1752);
  nor g213 (n_1758, n_1634, n_1757);
  nand g222 (n_1867, n_1760, n_1762);
  nor g223 (n_1768, n_1646, n_1767);
  nand g232 (n_1875, n_1770, n_1772);
  nor g233 (n_1778, n_1658, n_1777);
  nand g242 (n_1882, n_1780, n_1782);
  nor g243 (n_1788, n_1670, n_1787);
  nand g252 (n_1890, n_1790, n_1792);
  nor g253 (n_1798, n_1682, n_1797);
  nand g262 (n_1897, n_1800, n_1802);
  nor g263 (n_1808, n_1694, n_1807);
  nand g1776 (n_1905, n_1810, n_1812);
  nor g1777 (n_1818, n_1706, n_1817);
  nand g1786 (n_1912, n_1820, n_1822);
  nor g1787 (n_1828, n_1718, n_1827);
  nand g1796 (n_1920, n_1830, n_1832);
  nor g1797 (n_1838, n_1730, n_1837);
  nand g1806 (n_1927, n_1840, n_1842);
  nor g1807 (n_1848, n_1740, n_1847);
  nand g1814 (n_2131, n_1611, n_1854);
  nand g1816 (n_2133, n_1747, n_1855);
  nand g1819 (n_2136, n_1858, n_1859);
  nand g1822 (n_1935, n_1862, n_1863);
  nor g1823 (n_1865, n_1640, n_1864);
  nor g1826 (n_1945, n_1640, n_1867);
  nor g1832 (n_1873, n_1871, n_1864);
  nor g1835 (n_1951, n_1867, n_1871);
  nor g1836 (n_1877, n_1875, n_1864);
  nor g1839 (n_1954, n_1867, n_1875);
  nor g1840 (n_1880, n_1664, n_1879);
  nor g1843 (n_2034, n_1664, n_1882);
  nor g1849 (n_1888, n_1886, n_1879);
  nor g1852 (n_2040, n_1882, n_1886);
  nor g1853 (n_1892, n_1890, n_1879);
  nor g1856 (n_1960, n_1882, n_1890);
  nor g1857 (n_1895, n_1688, n_1894);
  nor g1860 (n_1973, n_1688, n_1897);
  nor g1866 (n_1903, n_1901, n_1894);
  nor g1869 (n_1983, n_1897, n_1901);
  nor g1870 (n_1907, n_1905, n_1894);
  nor g1873 (n_1988, n_1897, n_1905);
  nor g1874 (n_1910, n_1712, n_1909);
  nor g1877 (n_2086, n_1712, n_1912);
  nor g1883 (n_1918, n_1916, n_1909);
  nor g1886 (n_2092, n_1912, n_1916);
  nor g1887 (n_1922, n_1920, n_1909);
  nor g1890 (n_1996, n_1912, n_1920);
  nor g1891 (n_1925, n_1736, n_1924);
  nor g1894 (n_2009, n_1736, n_1927);
  nor g1900 (n_1933, n_1931, n_1924);
  nor g1903 (n_2019, n_1927, n_1931);
  nand g1906 (n_2140, n_1623, n_1937);
  nand g1907 (n_1938, n_1760, n_1935);
  nand g1908 (n_2142, n_1757, n_1938);
  nand g1911 (n_2145, n_1941, n_1942);
  nand g1914 (n_2148, n_1864, n_1944);
  nand g1915 (n_1947, n_1945, n_1935);
  nand g1916 (n_2151, n_1946, n_1947);
  nand g1917 (n_1950, n_1948, n_1935);
  nand g1918 (n_2153, n_1949, n_1950);
  nand g1919 (n_1953, n_1951, n_1935);
  nand g1920 (n_2156, n_1952, n_1953);
  nand g1921 (n_1956, n_1954, n_1935);
  nand g1922 (n_2024, n_1955, n_1956);
  nor g1923 (n_1958, n_1676, n_1957);
  nand g1932 (n_2048, n_1800, n_1960);
  nor g1933 (n_1967, n_1965, n_1957);
  nor g1938 (n_1970, n_1897, n_1957);
  nand g1947 (n_2060, n_1960, n_1973);
  nand g1952 (n_2064, n_1960, n_1978);
  nand g1957 (n_2068, n_1960, n_1983);
  nand g1962 (n_2072, n_1960, n_1988);
  nor g1963 (n_1994, n_1724, n_1993);
  nand g1972 (n_2100, n_1840, n_1996);
  nor g1973 (n_2003, n_2001, n_1993);
  nor g1978 (n_2006, n_1927, n_1993);
  nand g1987 (n_2112, n_1996, n_2009);
  nand g1992 (n_2116, n_1996, n_2014);
  nand g1997 (n_2120, n_1996, n_2019);
  nand g2000 (n_2160, n_1647, n_2026);
  nand g2001 (n_2027, n_1780, n_2024);
  nand g2002 (n_2162, n_1777, n_2027);
  nand g2005 (n_2165, n_2030, n_2031);
  nand g2008 (n_2168, n_1879, n_2033);
  nand g2009 (n_2036, n_2034, n_2024);
  nand g2010 (n_2171, n_2035, n_2036);
  nand g2011 (n_2039, n_2037, n_2024);
  nand g2012 (n_2173, n_2038, n_2039);
  nand g2013 (n_2042, n_2040, n_2024);
  nand g2014 (n_2176, n_2041, n_2042);
  nand g2015 (n_2043, n_1960, n_2024);
  nand g2016 (n_2178, n_1957, n_2043);
  nand g2019 (n_2181, n_2046, n_2047);
  nand g2022 (n_2183, n_2050, n_2051);
  nand g2025 (n_2186, n_2054, n_2055);
  nand g2028 (n_2189, n_2058, n_2059);
  nand g2031 (n_2192, n_2062, n_2063);
  nand g2034 (n_2194, n_2066, n_2067);
  nand g2037 (n_2197, n_2070, n_2071);
  nand g2040 (n_2076, n_2074, n_2075);
  nand g2043 (n_2201, n_1695, n_2078);
  nand g2044 (n_2079, n_1820, n_2076);
  nand g2045 (n_2203, n_1817, n_2079);
  nand g2048 (n_2206, n_2082, n_2083);
  nand g2051 (n_2209, n_1909, n_2085);
  nand g2052 (n_2088, n_2086, n_2076);
  nand g2053 (n_2212, n_2087, n_2088);
  nand g2054 (n_2091, n_2089, n_2076);
  nand g2055 (n_2214, n_2090, n_2091);
  nand g2056 (n_2094, n_2092, n_2076);
  nand g2057 (n_2217, n_2093, n_2094);
  nand g2058 (n_2095, n_1996, n_2076);
  nand g2059 (n_2219, n_1993, n_2095);
  nand g2062 (n_2222, n_2098, n_2099);
  nand g2065 (n_2224, n_2102, n_2103);
  nand g2068 (n_2227, n_2106, n_2107);
  nand g2071 (n_2230, n_2110, n_2111);
  nand g2074 (n_2233, n_2114, n_2115);
  nand g2077 (n_2235, n_2118, n_2119);
  nand g2080 (n_2238, n_2122, n_2123);
  xnor g2092 (Z[5], n_2131, n_2132);
  xnor g2094 (Z[6], n_2133, n_2134);
  xnor g2097 (Z[7], n_2136, n_2137);
  xnor g2099 (Z[8], n_1935, n_2138);
  xnor g2102 (Z[9], n_2140, n_2141);
  xnor g2104 (Z[10], n_2142, n_2143);
  xnor g2107 (Z[11], n_2145, n_2146);
  xnor g2110 (Z[12], n_2148, n_2149);
  xnor g2113 (Z[13], n_2151, n_2152);
  xnor g2115 (Z[14], n_2153, n_2154);
  xnor g2118 (Z[15], n_2156, n_2157);
  xnor g2120 (Z[16], n_2024, n_2158);
  xnor g2123 (Z[17], n_2160, n_2161);
  xnor g2125 (Z[18], n_2162, n_2163);
  xnor g2128 (Z[19], n_2165, n_2166);
  xnor g2131 (Z[20], n_2168, n_2169);
  xnor g2134 (Z[21], n_2171, n_2172);
  xnor g2136 (Z[22], n_2173, n_2174);
  xnor g2139 (Z[23], n_2176, n_2177);
  xnor g2141 (Z[24], n_2178, n_2179);
  xnor g2144 (Z[25], n_2181, n_2182);
  xnor g2146 (Z[26], n_2183, n_2184);
  xnor g2149 (Z[27], n_2186, n_2187);
  xnor g2152 (Z[28], n_2189, n_2190);
  xnor g2155 (Z[29], n_2192, n_2193);
  xnor g2157 (Z[30], n_2194, n_2195);
  xnor g2160 (Z[31], n_2197, n_2198);
  xnor g2162 (Z[32], n_2076, n_2199);
  xnor g2165 (Z[33], n_2201, n_2202);
  xnor g2167 (Z[34], n_2203, n_2204);
  xnor g2170 (Z[35], n_2206, n_2207);
  xnor g2173 (Z[36], n_2209, n_2210);
  xnor g2176 (Z[37], n_2212, n_2213);
  xnor g2178 (Z[38], n_2214, n_2215);
  xnor g2181 (Z[39], n_2217, n_2218);
  xnor g2183 (Z[40], n_2219, n_2220);
  xnor g2186 (Z[41], n_2222, n_2223);
  xnor g2188 (Z[42], n_2224, n_2225);
  xnor g2191 (Z[43], n_2227, n_2228);
  xnor g2194 (Z[44], n_2230, n_2231);
  xnor g2197 (Z[45], n_2233, n_2234);
  xnor g2199 (Z[46], n_2235, n_2236);
  xnor g2202 (Z[47], n_2238, n_2239);
  or g2212 (n_1045, A[1], wc);
  not gc (wc, n_171);
  or g2213 (n_1046, A[1], wc0);
  not gc0 (wc0, A[2]);
  or g2214 (n_1062, wc1, A[24]);
  not gc1 (wc1, A[18]);
  or g2215 (n_1089, wc2, A[2]);
  not gc2 (wc2, A[1]);
  or g2216 (n_1090, A[2], wc3);
  not gc3 (wc3, A[3]);
  or g2217 (n_1145, wc4, A[24]);
  not gc4 (wc4, A[15]);
  xnor g2218 (n_1187, A[24], A[17]);
  or g2219 (n_1188, wc5, A[24]);
  not gc5 (wc5, A[17]);
  or g2220 (n_1190, wc6, A[24]);
  not gc6 (wc6, A[21]);
  or g2222 (n_1216, A[5], wc7);
  not gc7 (wc7, A[6]);
  or g2223 (n_1217, A[5], wc8);
  not gc8 (wc8, A[9]);
  or g2224 (n_1253, A[6], wc9);
  not gc9 (wc9, A[7]);
  or g2225 (n_1254, wc10, A[6]);
  not gc10 (wc10, A[5]);
  xnor g2226 (n_474, n_1291, A[24]);
  or g2227 (n_1293, wc11, A[24]);
  not gc11 (wc11, A[12]);
  or g2228 (n_1294, wc12, A[24]);
  not gc12 (wc12, A[11]);
  xnor g2229 (n_1327, A[24], A[12]);
  xnor g2230 (n_1359, A[21], A[10]);
  or g2231 (n_1360, A[10], wc13);
  not gc13 (wc13, A[21]);
  or g2232 (n_1362, A[10], wc14);
  not gc14 (wc14, A[17]);
  xnor g2233 (n_1387, A[15], A[10]);
  or g2234 (n_1388, A[10], wc15);
  not gc15 (wc15, A[15]);
  or g2235 (n_1390, A[10], wc16);
  not gc16 (wc16, A[23]);
  xnor g2236 (n_1415, A[24], A[15]);
  or g2237 (n_1418, wc17, A[24]);
  not gc17 (wc17, A[19]);
  xnor g2238 (n_546, n_1439, A[24]);
  or g2239 (n_1442, wc18, A[24]);
  not gc18 (wc18, A[13]);
  xnor g2240 (n_1467, A[18], A[14]);
  or g2241 (n_1468, A[14], wc19);
  not gc19 (wc19, A[18]);
  or g2242 (n_1469, A[14], wc20);
  not gc20 (wc20, A[22]);
  xnor g2243 (n_571, n_1107, A[14]);
  or g2244 (n_1489, A[14], wc21);
  not gc21 (wc21, A[19]);
  or g2245 (n_1506, wc22, A[24]);
  not gc22 (wc22, A[23]);
  xnor g2246 (n_1523, A[24], A[21]);
  xnor g2247 (n_1555, A[23], A[21]);
  or g2248 (n_1556, wc23, A[23]);
  not gc23 (wc23, A[21]);
  xnor g2249 (n_1563, A[24], A[23]);
  or g2250 (n_1578, wc24, A[24]);
  not gc24 (wc24, A[20]);
  xnor g2251 (n_1583, A[22], A[21]);
  or g2252 (n_1584, A[21], wc25);
  not gc25 (wc25, A[22]);
  xnor g2253 (n_1587, A[23], A[22]);
  or g2254 (n_1588, wc26, A[23]);
  not gc26 (wc26, A[22]);
  xnor g2255 (n_350, n_1043, A[1]);
  xnor g2256 (n_373, n_1087, A[2]);
  xnor g2257 (n_435, n_699, A[9]);
  xnor g2258 (n_454, n_1251, A[6]);
  or g2259 (n_1546, A[21], wc27);
  not gc27 (wc27, n_441);
  or g2260 (n_1558, A[23], wc28);
  not gc28 (wc28, n_461);
  or g2261 (n_74, A[23], wc29);
  not gc29 (wc29, n_1506);
  or g2263 (n_2125, wc30, n_1610);
  not gc30 (wc30, n_1605);
  xnor g2264 (n_1543, n_439, A[21]);
  or g2265 (n_1544, A[21], wc31);
  not gc31 (wc31, n_439);
  or g2266 (n_1585, A[21], wc32);
  not gc32 (wc32, n_618);
  and g2267 (n_1745, wc33, n_1607);
  not gc33 (wc33, n_1608);
  or g2268 (n_2128, wc34, n_1606);
  not gc34 (wc34, n_1607);
  and g2269 (n_1738, wc35, n_74);
  not gc35 (wc35, A[24]);
  or g2270 (n_1739, wc36, n_74);
  not gc36 (wc36, A[24]);
  not g2271 (Z[2], n_2125);
  or g2272 (n_2129, wc37, n_1616);
  not gc37 (wc37, n_1611);
  xnor g2273 (n_1059, n_353, A[24]);
  or g2274 (n_1060, A[24], wc38);
  not gc38 (wc38, n_353);
  xnor g2275 (n_1143, n_395, A[24]);
  or g2276 (n_1144, A[24], wc39);
  not gc39 (wc39, n_395);
  and g2277 (n_1747, wc40, n_1613);
  not gc40 (wc40, n_1614);
  or g2280 (n_1856, wc41, n_1622);
  not gc41 (wc41, n_1750);
  or g2281 (n_2132, wc42, n_1612);
  not gc42 (wc42, n_1613);
  or g2282 (n_2134, wc43, n_1622);
  not gc43 (wc43, n_1617);
  or g2283 (n_2236, wc44, n_1740);
  not gc44 (wc44, n_1737);
  or g2284 (n_1854, n_1616, n_1745);
  or g2285 (n_1855, n_1745, wc45);
  not gc45 (wc45, n_1750);
  xor g2286 (Z[3], n_1605, n_2128);
  xor g2287 (Z[4], n_1745, n_2129);
  or g2288 (n_2239, wc46, n_1738);
  not gc46 (wc46, n_1739);
  and g2289 (n_1754, wc47, n_1619);
  not gc47 (wc47, n_1620);
  and g2290 (n_1858, wc48, n_1617);
  not gc48 (wc48, n_1748);
  or g2291 (n_1859, n_1745, n_1856);
  or g2292 (n_2137, wc49, n_1618);
  not gc49 (wc49, n_1619);
  or g2293 (n_2138, wc50, n_1628);
  not gc50 (wc50, n_1623);
  or g2294 (n_2234, wc51, n_1732);
  not gc51 (wc51, n_1733);
  and g2295 (n_1757, wc52, n_1625);
  not gc52 (wc52, n_1626);
  and g2296 (n_1755, wc53, n_1752);
  not gc53 (wc53, n_1747);
  or g2297 (n_2141, wc54, n_1624);
  not gc54 (wc54, n_1625);
  or g2298 (n_2228, wc55, n_1726);
  not gc55 (wc55, n_1727);
  and g2299 (n_1844, wc56, n_1727);
  not gc56 (wc56, n_1728);
  and g2300 (n_1847, wc57, n_1733);
  not gc57 (wc57, n_1734);
  and g2301 (n_1862, wc58, n_1754);
  not gc58 (wc58, n_1755);
  or g2302 (n_1931, wc59, n_1740);
  not gc59 (wc59, n_1850);
  or g2303 (n_1863, n_1860, n_1745);
  or g2304 (n_2149, wc60, n_1640);
  not gc60 (wc60, n_1635);
  or g2305 (n_2225, wc61, n_1730);
  not gc61 (wc61, n_1725);
  or g2306 (n_2231, wc62, n_1736);
  not gc62 (wc62, n_1731);
  and g2307 (n_1764, wc63, n_1631);
  not gc63 (wc63, n_1632);
  and g2308 (n_1941, wc64, n_1629);
  not gc64 (wc64, n_1758);
  or g2309 (n_1939, wc65, n_1634);
  not gc65 (wc65, n_1760);
  or g2310 (n_2143, wc66, n_1634);
  not gc66 (wc66, n_1629);
  or g2311 (n_2146, wc67, n_1630);
  not gc67 (wc67, n_1631);
  and g2312 (n_1767, wc68, n_1637);
  not gc68 (wc68, n_1638);
  and g2313 (n_1834, wc69, n_1715);
  not gc69 (wc69, n_1716);
  and g2314 (n_1837, wc70, n_1721);
  not gc70 (wc70, n_1722);
  and g2315 (n_1765, wc71, n_1762);
  not gc71 (wc71, n_1757);
  or g2316 (n_1871, wc72, n_1646);
  not gc72 (wc72, n_1770);
  or g2317 (n_2001, wc73, n_1730);
  not gc73 (wc73, n_1840);
  and g2318 (n_1932, wc74, n_1737);
  not gc74 (wc74, n_1848);
  or g2319 (n_1937, wc75, n_1628);
  not gc75 (wc75, n_1935);
  or g2320 (n_2152, wc76, n_1636);
  not gc76 (wc76, n_1637);
  or g2321 (n_2154, wc77, n_1646);
  not gc77 (wc77, n_1641);
  or g2322 (n_2215, wc78, n_1718);
  not gc78 (wc78, n_1713);
  or g2323 (n_2218, wc79, n_1714);
  not gc79 (wc79, n_1715);
  or g2324 (n_2220, wc80, n_1724);
  not gc80 (wc80, n_1719);
  or g2325 (n_2223, wc81, n_1720);
  not gc81 (wc81, n_1721);
  and g2326 (n_1827, wc82, n_1709);
  not gc82 (wc82, n_1710);
  and g2327 (n_1864, wc83, n_1764);
  not gc83 (wc83, n_1765);
  or g2328 (n_1916, wc84, n_1718);
  not gc84 (wc84, n_1830);
  and g2329 (n_1845, wc85, n_1842);
  not gc85 (wc85, n_1837);
  and g2330 (n_1948, wc86, n_1770);
  not gc86 (wc86, n_1867);
  and g2331 (n_2014, wc87, n_1850);
  not gc87 (wc87, n_1927);
  or g2332 (n_1942, n_1939, wc88);
  not gc88 (wc88, n_1935);
  or g2333 (n_1944, wc89, n_1867);
  not gc89 (wc89, n_1935);
  or g2334 (n_2210, wc90, n_1712);
  not gc90 (wc90, n_1707);
  or g2335 (n_2213, wc91, n_1708);
  not gc91 (wc91, n_1709);
  and g2336 (n_1774, wc92, n_1643);
  not gc92 (wc92, n_1644);
  and g2337 (n_1777, wc93, n_1649);
  not gc93 (wc93, n_1650);
  and g2338 (n_1784, wc94, n_1655);
  not gc94 (wc94, n_1656);
  and g2339 (n_1824, wc95, n_1703);
  not gc95 (wc95, n_1704);
  and g2340 (n_1872, wc96, n_1641);
  not gc96 (wc96, n_1768);
  or g2341 (n_2028, wc97, n_1658);
  not gc97 (wc97, n_1780);
  and g2342 (n_1835, wc98, n_1832);
  not gc98 (wc98, n_1827);
  and g2343 (n_2002, wc99, n_1725);
  not gc99 (wc99, n_1838);
  and g2344 (n_1924, wc100, n_1844);
  not gc100 (wc100, n_1845);
  and g2345 (n_1869, wc101, n_1770);
  not gc101 (wc101, n_1864);
  or g2346 (n_2157, wc102, n_1642);
  not gc102 (wc102, n_1643);
  or g2347 (n_2158, wc103, n_1652);
  not gc103 (wc103, n_1647);
  or g2348 (n_2161, wc104, n_1648);
  not gc104 (wc104, n_1649);
  or g2349 (n_2163, wc105, n_1658);
  not gc105 (wc105, n_1653);
  or g2350 (n_2166, wc106, n_1654);
  not gc106 (wc106, n_1655);
  or g2351 (n_2204, wc107, n_1706);
  not gc107 (wc107, n_1701);
  or g2352 (n_2207, wc108, n_1702);
  not gc108 (wc108, n_1703);
  and g2353 (n_1775, wc109, n_1772);
  not gc109 (wc109, n_1767);
  and g2354 (n_1785, wc110, n_1782);
  not gc110 (wc110, n_1777);
  and g2355 (n_1917, wc111, n_1713);
  not gc111 (wc111, n_1828);
  and g2356 (n_1921, wc112, n_1834);
  not gc112 (wc112, n_1835);
  and g2357 (n_1946, wc113, n_1635);
  not gc113 (wc113, n_1865);
  and g2358 (n_1949, wc114, n_1767);
  not gc114 (wc114, n_1869);
  and g2359 (n_1929, wc115, n_1850);
  not gc115 (wc115, n_1924);
  and g2360 (n_1876, wc116, n_1774);
  not gc116 (wc116, n_1775);
  and g2361 (n_2030, wc117, n_1653);
  not gc117 (wc117, n_1778);
  and g2362 (n_1879, wc118, n_1784);
  not gc118 (wc118, n_1785);
  and g2363 (n_1952, n_1872, wc119);
  not gc119 (wc119, n_1873);
  and g2364 (n_2011, wc120, n_1731);
  not gc120 (wc120, n_1925);
  and g2365 (n_2016, wc121, n_1847);
  not gc121 (wc121, n_1929);
  and g2366 (n_2021, n_1932, wc122);
  not gc122 (wc122, n_1933);
  or g2367 (n_2169, wc123, n_1664);
  not gc123 (wc123, n_1659);
  or g2368 (n_2177, wc124, n_1666);
  not gc124 (wc124, n_1667);
  or g2369 (n_2184, wc125, n_1682);
  not gc125 (wc125, n_1677);
  and g2370 (n_1787, wc126, n_1661);
  not gc126 (wc126, n_1662);
  and g2371 (n_1794, wc127, n_1667);
  not gc127 (wc127, n_1668);
  and g2372 (n_1797, wc128, n_1673);
  not gc128 (wc128, n_1674);
  and g2373 (n_1804, wc129, n_1679);
  not gc129 (wc129, n_1680);
  or g2374 (n_1886, wc130, n_1670);
  not gc130 (wc130, n_1790);
  or g2375 (n_1965, wc131, n_1682);
  not gc131 (wc131, n_1800);
  or g2376 (n_2172, wc132, n_1660);
  not gc132 (wc132, n_1661);
  or g2377 (n_2174, wc133, n_1670);
  not gc133 (wc133, n_1665);
  or g2378 (n_2179, wc134, n_1676);
  not gc134 (wc134, n_1671);
  or g2379 (n_2182, wc135, n_1672);
  not gc135 (wc135, n_1673);
  or g2380 (n_2187, wc136, n_1678);
  not gc136 (wc136, n_1679);
  or g2381 (n_2190, wc137, n_1688);
  not gc137 (wc137, n_1683);
  and g2382 (n_1807, wc138, n_1685);
  not gc138 (wc138, n_1686);
  and g2383 (n_1814, wc139, n_1691);
  not gc139 (wc139, n_1692);
  and g2384 (n_1817, wc140, n_1697);
  not gc140 (wc140, n_1698);
  and g2385 (n_1795, wc141, n_1792);
  not gc141 (wc141, n_1787);
  and g2386 (n_1805, wc142, n_1802);
  not gc142 (wc142, n_1797);
  or g2387 (n_1901, wc143, n_1694);
  not gc143 (wc143, n_1810);
  or g2388 (n_2080, wc144, n_1706);
  not gc144 (wc144, n_1820);
  and g2389 (n_1955, n_1876, wc145);
  not gc145 (wc145, n_1877);
  and g2390 (n_2035, wc146, n_1659);
  not gc146 (wc146, n_1880);
  and g2391 (n_1884, wc147, n_1790);
  not gc147 (wc147, n_1879);
  and g2392 (n_2037, wc148, n_1790);
  not gc148 (wc148, n_1882);
  or g2393 (n_2193, wc149, n_1684);
  not gc149 (wc149, n_1685);
  or g2394 (n_2195, wc150, n_1694);
  not gc150 (wc150, n_1689);
  or g2395 (n_2198, wc151, n_1690);
  not gc151 (wc151, n_1691);
  or g2396 (n_2199, wc152, n_1700);
  not gc152 (wc152, n_1695);
  or g2397 (n_2202, wc153, n_1696);
  not gc153 (wc153, n_1697);
  and g2398 (n_1887, wc154, n_1665);
  not gc154 (wc154, n_1788);
  and g2399 (n_1891, wc155, n_1794);
  not gc155 (wc155, n_1795);
  and g2400 (n_1966, wc156, n_1677);
  not gc156 (wc156, n_1798);
  and g2401 (n_1894, wc157, n_1804);
  not gc157 (wc157, n_1805);
  and g2402 (n_1815, wc158, n_1812);
  not gc158 (wc158, n_1807);
  and g2403 (n_1825, wc159, n_1822);
  not gc159 (wc159, n_1817);
  and g2404 (n_2038, wc160, n_1787);
  not gc160 (wc160, n_1884);
  and g2405 (n_1978, wc161, n_1810);
  not gc161 (wc161, n_1897);
  and g2406 (n_2089, wc162, n_1830);
  not gc162 (wc162, n_1912);
  or g2407 (n_2044, wc163, n_1676);
  not gc163 (wc163, n_1960);
  or g2408 (n_2052, n_1965, wc164);
  not gc164 (wc164, n_1960);
  or g2409 (n_2056, wc165, n_1897);
  not gc165 (wc165, n_1960);
  and g2410 (n_1902, wc166, n_1689);
  not gc166 (wc166, n_1808);
  and g2411 (n_1906, wc167, n_1814);
  not gc167 (wc167, n_1815);
  and g2412 (n_2082, wc168, n_1701);
  not gc168 (wc168, n_1818);
  and g2413 (n_1909, wc169, n_1824);
  not gc169 (wc169, n_1825);
  and g2414 (n_1899, wc170, n_1810);
  not gc170 (wc170, n_1894);
  or g2415 (n_2096, wc171, n_1724);
  not gc171 (wc171, n_1996);
  or g2416 (n_2104, n_2001, wc172);
  not gc172 (wc172, n_1996);
  or g2417 (n_2108, wc173, n_1927);
  not gc173 (wc173, n_1996);
  or g2418 (n_2026, wc174, n_1652);
  not gc174 (wc174, n_2024);
  or g2419 (n_2031, n_2028, wc175);
  not gc175 (wc175, n_2024);
  or g2420 (n_2033, wc176, n_1882);
  not gc176 (wc176, n_2024);
  and g2421 (n_2041, n_1887, wc177);
  not gc177 (wc177, n_1888);
  and g2422 (n_1957, n_1891, wc178);
  not gc178 (wc178, n_1892);
  and g2423 (n_1975, wc179, n_1683);
  not gc179 (wc179, n_1895);
  and g2424 (n_1980, wc180, n_1807);
  not gc180 (wc180, n_1899);
  and g2425 (n_1914, wc181, n_1830);
  not gc181 (wc181, n_1909);
  or g2426 (n_2047, n_2044, wc182);
  not gc182 (wc182, n_2024);
  or g2427 (n_2051, n_2048, wc183);
  not gc183 (wc183, n_2024);
  or g2428 (n_2055, n_2052, wc184);
  not gc184 (wc184, n_2024);
  or g2429 (n_2059, n_2056, wc185);
  not gc185 (wc185, n_2024);
  or g2430 (n_2063, n_2060, wc186);
  not gc186 (wc186, n_2024);
  and g2431 (n_1985, n_1902, wc187);
  not gc187 (wc187, n_1903);
  and g2432 (n_1990, n_1906, wc188);
  not gc188 (wc188, n_1907);
  and g2433 (n_2087, wc189, n_1707);
  not gc189 (wc189, n_1910);
  and g2434 (n_2090, wc190, n_1827);
  not gc190 (wc190, n_1914);
  and g2435 (n_2093, n_1917, wc191);
  not gc191 (wc191, n_1918);
  and g2436 (n_1993, n_1921, wc192);
  not gc192 (wc192, n_1922);
  and g2437 (n_1963, wc193, n_1800);
  not gc193 (wc193, n_1957);
  and g2438 (n_1976, wc194, n_1973);
  not gc194 (wc194, n_1957);
  and g2439 (n_1981, wc195, n_1978);
  not gc195 (wc195, n_1957);
  and g2440 (n_1986, wc196, n_1983);
  not gc196 (wc196, n_1957);
  and g2441 (n_1991, wc197, n_1988);
  not gc197 (wc197, n_1957);
  or g2442 (n_2067, n_2064, wc198);
  not gc198 (wc198, n_2024);
  or g2443 (n_2071, n_2068, wc199);
  not gc199 (wc199, n_2024);
  or g2444 (n_2075, n_2072, wc200);
  not gc200 (wc200, n_2024);
  and g2445 (n_2046, wc201, n_1671);
  not gc201 (wc201, n_1958);
  and g2446 (n_2050, wc202, n_1797);
  not gc202 (wc202, n_1963);
  and g2447 (n_2054, n_1966, wc203);
  not gc203 (wc203, n_1967);
  and g2448 (n_2058, n_1894, wc204);
  not gc204 (wc204, n_1970);
  and g2449 (n_2062, wc205, n_1975);
  not gc205 (wc205, n_1976);
  and g2450 (n_2066, wc206, n_1980);
  not gc206 (wc206, n_1981);
  and g2451 (n_1999, wc207, n_1840);
  not gc207 (wc207, n_1993);
  and g2452 (n_2012, wc208, n_2009);
  not gc208 (wc208, n_1993);
  and g2453 (n_2017, wc209, n_2014);
  not gc209 (wc209, n_1993);
  and g2454 (n_2022, wc210, n_2019);
  not gc210 (wc210, n_1993);
  and g2455 (n_2070, wc211, n_1985);
  not gc211 (wc211, n_1986);
  and g2456 (n_2074, wc212, n_1990);
  not gc212 (wc212, n_1991);
  and g2457 (n_2098, wc213, n_1719);
  not gc213 (wc213, n_1994);
  and g2458 (n_2102, wc214, n_1837);
  not gc214 (wc214, n_1999);
  and g2459 (n_2106, n_2002, wc215);
  not gc215 (wc215, n_2003);
  and g2460 (n_2110, n_1924, wc216);
  not gc216 (wc216, n_2006);
  and g2461 (n_2114, wc217, n_2011);
  not gc217 (wc217, n_2012);
  and g2462 (n_2118, wc218, n_2016);
  not gc218 (wc218, n_2017);
  and g2463 (n_2122, wc219, n_2021);
  not gc219 (wc219, n_2022);
  or g2464 (n_2078, wc220, n_1700);
  not gc220 (wc220, n_2076);
  or g2465 (n_2083, n_2080, wc221);
  not gc221 (wc221, n_2076);
  or g2466 (n_2085, wc222, n_1912);
  not gc222 (wc222, n_2076);
  or g2467 (n_2099, n_2096, wc223);
  not gc223 (wc223, n_2076);
  or g2468 (n_2103, wc224, n_2100);
  not gc224 (wc224, n_2076);
  or g2469 (n_2107, n_2104, wc225);
  not gc225 (wc225, n_2076);
  or g2470 (n_2111, n_2108, wc226);
  not gc226 (wc226, n_2076);
  or g2471 (n_2115, wc227, n_2112);
  not gc227 (wc227, n_2076);
  or g2472 (n_2119, wc228, n_2116);
  not gc228 (wc228, n_2076);
  or g2473 (n_2123, wc229, n_2120);
  not gc229 (wc229, n_2076);
endmodule

module mult_signed_const_3884_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_3884_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_4151_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_176;
  wire n_178, n_179, n_180, n_183, n_184, n_187, n_188, n_189;
  wire n_195, n_196, n_200, n_201, n_202, n_203, n_204, n_207;
  wire n_209, n_210, n_211, n_212, n_217, n_218, n_219, n_220;
  wire n_221, n_223, n_224, n_225, n_226, n_227, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_242;
  wire n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_265, n_268;
  wire n_271, n_272, n_273, n_274, n_275, n_276, n_277, n_282;
  wire n_283, n_285, n_286, n_287, n_288, n_289, n_290, n_291;
  wire n_292, n_293, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_315, n_317;
  wire n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_349, n_351, n_353, n_356;
  wire n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364;
  wire n_365, n_366, n_367, n_371, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_453;
  wire n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461;
  wire n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_470;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494;
  wire n_495, n_496, n_497, n_498, n_499, n_500, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_519, n_520, n_521, n_522, n_523;
  wire n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_532;
  wire n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540;
  wire n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548;
  wire n_549, n_550, n_551, n_552, n_553, n_554, n_557, n_558;
  wire n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_569;
  wire n_570, n_571, n_572, n_573, n_574, n_575, n_576, n_578;
  wire n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586;
  wire n_588, n_589, n_590, n_591, n_592, n_596, n_597, n_598;
  wire n_599, n_603, n_604, n_605, n_606, n_609, n_610, n_611;
  wire n_613, n_614, n_617, n_622, n_623, n_624, n_625, n_626;
  wire n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634;
  wire n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642;
  wire n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675;
  wire n_676, n_677, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_698, n_699, n_700, n_701;
  wire n_702, n_703, n_704, n_705, n_706, n_707, n_708, n_709;
  wire n_710, n_711, n_712, n_713, n_722, n_723, n_724, n_725;
  wire n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733;
  wire n_738, n_742, n_743, n_744, n_745, n_746, n_747, n_748;
  wire n_749, n_750, n_751, n_752, n_753, n_760, n_761, n_762;
  wire n_763, n_765, n_766, n_767, n_768, n_769, n_770, n_771;
  wire n_772, n_773, n_774, n_775, n_776, n_777, n_785, n_786;
  wire n_787, n_788, n_789, n_790, n_791, n_792, n_793, n_794;
  wire n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802;
  wire n_803, n_804, n_805, n_814, n_815, n_817, n_818, n_819;
  wire n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827;
  wire n_828, n_829, n_830, n_831, n_832, n_833, n_842, n_846;
  wire n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854;
  wire n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862;
  wire n_866, n_867, n_868, n_874, n_876, n_877, n_878, n_880;
  wire n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888;
  wire n_889, n_890, n_891, n_892, n_893, n_904, n_905, n_906;
  wire n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914;
  wire n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922;
  wire n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_938;
  wire n_939, n_944, n_945, n_946, n_947, n_948, n_949, n_950;
  wire n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958;
  wire n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_978;
  wire n_979, n_980, n_982, n_983, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_996, n_997, n_998, n_999, n_1000, n_1001, n_1014, n_1020;
  wire n_1021, n_1022, n_1023, n_1024, n_1026, n_1027, n_1028, n_1029;
  wire n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037;
  wire n_1038, n_1039, n_1040, n_1041, n_1042, n_1044, n_1045, n_1046;
  wire n_1047, n_1049, n_1050, n_1051, n_1052, n_1056, n_1057, n_1058;
  wire n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066;
  wire n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074;
  wire n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082;
  wire n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090;
  wire n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098;
  wire n_1099, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108;
  wire n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116;
  wire n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124;
  wire n_1125, n_1126, n_1127, n_1128, n_1129, n_1132, n_1133, n_1134;
  wire n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142;
  wire n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151;
  wire n_1152, n_1153, n_1154, n_1155, n_1156, n_1158, n_1159, n_1160;
  wire n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168;
  wire n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176;
  wire n_1177, n_1178, n_1179, n_1180, n_1182, n_1183, n_1184, n_1185;
  wire n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1193, n_1194;
  wire n_1195, n_1196, n_1197, n_1200, n_1201, n_1202, n_1203, n_1204;
  wire n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212;
  wire n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220;
  wire n_1221, n_1222, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229;
  wire n_1230, n_1231, n_1232, n_1234, n_1235, n_1236, n_1237, n_1238;
  wire n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246;
  wire n_1247, n_1248, n_1249, n_1250, n_1252, n_1253, n_1256, n_1257;
  wire n_1258, n_1259, n_1260, n_1262, n_1263, n_1264, n_1265, n_1266;
  wire n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1274, n_1275;
  wire n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283;
  wire n_1284, n_1285, n_1286, n_1288, n_1292, n_1293, n_1294, n_1295;
  wire n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303;
  wire n_1304, n_1306, n_1307, n_1308, n_1310, n_1311, n_1312, n_1313;
  wire n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321;
  wire n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1333;
  wire n_1334, n_1335, n_1336, n_1337, n_1340, n_1341, n_1342, n_1343;
  wire n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351;
  wire n_1352, n_1353, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360;
  wire n_1361, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370;
  wire n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378;
  wire n_1379, n_1380, n_1381, n_1385, n_1386, n_1388, n_1389, n_1390;
  wire n_1391, n_1393, n_1394, n_1395, n_1396, n_1398, n_1399, n_1400;
  wire n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408;
  wire n_1409, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419;
  wire n_1421, n_1422, n_1423, n_1425, n_1426, n_1427, n_1428, n_1429;
  wire n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437;
  wire n_1438, n_1440, n_1441, n_1442, n_1445, n_1446, n_1447, n_1449;
  wire n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457;
  wire n_1458, n_1459, n_1460, n_1461, n_1463, n_1464, n_1465, n_1466;
  wire n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475;
  wire n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1485, n_1486;
  wire n_1488, n_1489, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
  wire n_1498, n_1499, n_1500, n_1501, n_1504, n_1505, n_1506, n_1507;
  wire n_1508, n_1510, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517;
  wire n_1518, n_1519, n_1520, n_1521, n_1526, n_1528, n_1529, n_1530;
  wire n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1541;
  wire n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1553, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560;
  wire n_1561, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572;
  wire n_1573, n_1578, n_1579, n_1580, n_1581, n_1583, n_1584, n_1585;
  wire n_1587, n_1588, n_1590, n_1591, n_1593, n_1604, n_1605, n_1606;
  wire n_1607, n_1609, n_1610, n_1611, n_1612, n_1613, n_1615, n_1616;
  wire n_1617, n_1618, n_1619, n_1621, n_1622, n_1623, n_1624, n_1625;
  wire n_1627, n_1628, n_1629, n_1630, n_1631, n_1633, n_1634, n_1635;
  wire n_1636, n_1637, n_1639, n_1640, n_1641, n_1642, n_1643, n_1645;
  wire n_1646, n_1647, n_1648, n_1649, n_1651, n_1652, n_1653, n_1654;
  wire n_1655, n_1657, n_1658, n_1659, n_1660, n_1661, n_1663, n_1664;
  wire n_1665, n_1666, n_1667, n_1669, n_1670, n_1671, n_1672, n_1673;
  wire n_1675, n_1676, n_1677, n_1678, n_1679, n_1681, n_1682, n_1683;
  wire n_1684, n_1685, n_1687, n_1688, n_1689, n_1690, n_1691, n_1693;
  wire n_1694, n_1695, n_1696, n_1697, n_1699, n_1700, n_1701, n_1702;
  wire n_1703, n_1705, n_1706, n_1707, n_1708, n_1709, n_1711, n_1712;
  wire n_1713, n_1714, n_1715, n_1717, n_1718, n_1719, n_1720, n_1721;
  wire n_1723, n_1724, n_1725, n_1726, n_1727, n_1729, n_1730, n_1731;
  wire n_1732, n_1733, n_1735, n_1736, n_1737, n_1738, n_1739, n_1744;
  wire n_1746, n_1747, n_1749, n_1751, n_1753, n_1754, n_1756, n_1757;
  wire n_1759, n_1761, n_1763, n_1764, n_1766, n_1767, n_1769, n_1771;
  wire n_1773, n_1774, n_1776, n_1777, n_1779, n_1781, n_1783, n_1784;
  wire n_1786, n_1787, n_1789, n_1791, n_1793, n_1794, n_1796, n_1797;
  wire n_1799, n_1801, n_1803, n_1804, n_1806, n_1807, n_1809, n_1811;
  wire n_1813, n_1814, n_1816, n_1817, n_1819, n_1821, n_1823, n_1824;
  wire n_1826, n_1827, n_1829, n_1831, n_1833, n_1834, n_1836, n_1837;
  wire n_1839, n_1841, n_1843, n_1844, n_1846, n_1847, n_1849, n_1853;
  wire n_1854, n_1855, n_1857, n_1858, n_1859, n_1861, n_1862, n_1863;
  wire n_1864, n_1866, n_1868, n_1870, n_1871, n_1872, n_1874, n_1875;
  wire n_1876, n_1878, n_1879, n_1881, n_1883, n_1885, n_1886, n_1887;
  wire n_1889, n_1890, n_1891, n_1893, n_1894, n_1896, n_1898, n_1900;
  wire n_1901, n_1902, n_1904, n_1905, n_1906, n_1908, n_1909, n_1911;
  wire n_1913, n_1915, n_1916, n_1917, n_1919, n_1920, n_1921, n_1923;
  wire n_1924, n_1926, n_1928, n_1930, n_1931, n_1932, n_1934, n_1936;
  wire n_1937, n_1938, n_1940, n_1941, n_1943, n_1944, n_1945, n_1946;
  wire n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954;
  wire n_1955, n_1956, n_1957, n_1959, n_1962, n_1964, n_1965, n_1966;
  wire n_1969, n_1972, n_1974, n_1975, n_1977, n_1979, n_1980, n_1982;
  wire n_1984, n_1985, n_1987, n_1989, n_1990, n_1992, n_1993, n_1995;
  wire n_1998, n_2000, n_2001, n_2002, n_2005, n_2008, n_2010, n_2011;
  wire n_2013, n_2015, n_2016, n_2018, n_2020, n_2021, n_2023, n_2025;
  wire n_2026, n_2027, n_2029, n_2030, n_2032, n_2033, n_2034, n_2035;
  wire n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043;
  wire n_2045, n_2046, n_2047, n_2049, n_2050, n_2051, n_2053, n_2054;
  wire n_2055, n_2057, n_2058, n_2059, n_2061, n_2062, n_2063, n_2065;
  wire n_2066, n_2067, n_2069, n_2070, n_2071, n_2073, n_2074, n_2075;
  wire n_2077, n_2078, n_2079, n_2081, n_2082, n_2084, n_2085, n_2086;
  wire n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094;
  wire n_2095, n_2097, n_2098, n_2099, n_2101, n_2102, n_2103, n_2105;
  wire n_2106, n_2107, n_2109, n_2110, n_2111, n_2113, n_2114, n_2115;
  wire n_2117, n_2118, n_2119, n_2121, n_2122, n_2124, n_2127, n_2128;
  wire n_2130, n_2131, n_2132, n_2133, n_2135, n_2136, n_2137, n_2139;
  wire n_2140, n_2141, n_2142, n_2144, n_2145, n_2147, n_2148, n_2150;
  wire n_2151, n_2152, n_2153, n_2155, n_2156, n_2157, n_2159, n_2160;
  wire n_2161, n_2162, n_2164, n_2165, n_2167, n_2168, n_2170, n_2171;
  wire n_2172, n_2173, n_2175, n_2176, n_2177, n_2178, n_2180, n_2181;
  wire n_2182, n_2183, n_2185, n_2186, n_2188, n_2189, n_2191, n_2192;
  wire n_2193, n_2194, n_2196, n_2197, n_2198, n_2200, n_2201, n_2202;
  wire n_2203, n_2205, n_2206, n_2208, n_2209, n_2211, n_2212, n_2213;
  wire n_2214, n_2216, n_2217, n_2218, n_2219, n_2221, n_2222, n_2223;
  wire n_2224, n_2226, n_2227, n_2229, n_2230, n_2232, n_2233, n_2234;
  wire n_2235, n_2237, n_2238;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], n_171);
  xor g270 (n_117, n_622, A[2]);
  nand g3 (n_623, A[1], n_171);
  nand g271 (n_624, A[2], n_171);
  nand g272 (n_625, A[1], A[2]);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, n_69);
  xor g288 (n_176, n_634, A[4]);
  nand g289 (n_635, n_68, n_69);
  nand g290 (n_636, A[4], n_69);
  nand g291 (n_637, n_68, A[4]);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_176);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_176);
  nand g296 (n_640, A[7], n_176);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g299 (n_642, A[1], A[2]);
  xor g300 (n_178, n_642, n_171);
  xor g305 (n_646, n_178, A[5]);
  xor g306 (n_180, n_646, A[6]);
  nand g307 (n_647, n_178, A[5]);
  nand g308 (n_648, A[6], A[5]);
  nand g309 (n_649, n_178, A[6]);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, n_179, n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, n_179, n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, n_179, A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_188, n_659, n_660, n_661);
  xor g329 (n_662, n_183, n_184);
  xor g330 (n_112, n_662, A[9]);
  nand g331 (n_663, n_183, n_184);
  nand g332 (n_664, A[9], n_184);
  nand g333 (n_665, n_183, A[9]);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_187, n_630, n_67);
  nand g340 (n_668, n_67, n_173);
  nand g341 (n_669, A[4], n_67);
  nand g342 (n_71, n_631, n_668, n_669);
  xor g343 (n_670, A[7], n_187);
  xor g344 (n_189, n_670, A[8]);
  nand g345 (n_671, A[7], n_187);
  nand g346 (n_672, A[8], n_187);
  nand g347 (n_673, A[7], A[8]);
  nand g348 (n_73, n_671, n_672, n_673);
  xor g349 (n_674, A[10], n_188);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, A[10], n_188);
  nand g352 (n_676, n_189, n_188);
  nand g353 (n_677, A[10], n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_195, n_638, n_71);
  nand g366 (n_684, n_71, n_176);
  nand g367 (n_685, A[5], n_71);
  nand g368 (n_201, n_639, n_684, n_685);
  xor g369 (n_686, A[8], A[9]);
  xor g370 (n_196, n_686, A[11]);
  nand g371 (n_687, A[8], A[9]);
  nand g372 (n_688, A[11], A[9]);
  nand g373 (n_689, A[8], A[11]);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, n_73, n_195);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, n_73, n_195);
  nand g378 (n_692, n_196, n_195);
  nand g379 (n_693, n_73, n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g387 (n_698, n_117, A[5]);
  xor g388 (n_200, n_698, n_179);
  nand g389 (n_699, n_117, A[5]);
  nand g390 (n_700, n_179, A[5]);
  nand g391 (n_701, n_117, n_179);
  nand g392 (n_207, n_699, n_700, n_701);
  xor g393 (n_702, A[6], n_200);
  xor g394 (n_202, n_702, A[10]);
  nand g395 (n_703, A[6], n_200);
  nand g396 (n_704, A[10], n_200);
  nand g397 (n_705, A[6], A[10]);
  nand g398 (n_209, n_703, n_704, n_705);
  xor g399 (n_706, A[9], A[12]);
  xor g400 (n_204, n_706, n_201);
  nand g401 (n_707, A[9], A[12]);
  nand g402 (n_708, n_201, A[12]);
  nand g403 (n_709, A[9], n_201);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, n_202, n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, n_202, n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, n_202, n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g423 (n_722, n_207, A[10]);
  xor g424 (n_210, n_722, n_184);
  nand g425 (n_723, n_207, A[10]);
  nand g426 (n_724, n_184, A[10]);
  nand g427 (n_725, n_207, n_184);
  nand g428 (n_217, n_723, n_724, n_725);
  xor g429 (n_726, A[11], A[13]);
  xor g430 (n_212, n_726, n_209);
  nand g431 (n_727, A[11], A[13]);
  nand g432 (n_728, n_209, A[13]);
  nand g433 (n_729, A[11], n_209);
  nand g434 (n_220, n_727, n_728, n_729);
  xor g435 (n_730, n_210, n_211);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, n_210, n_211);
  nand g438 (n_732, n_212, n_211);
  nand g439 (n_733, n_210, n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_218, n_738, n_187);
  xor g455 (n_742, n_188, A[12]);
  xor g456 (n_219, n_742, A[11]);
  nand g457 (n_743, n_188, A[12]);
  nand g458 (n_744, A[11], A[12]);
  nand g459 (n_745, n_188, A[11]);
  nand g460 (n_224, n_743, n_744, n_745);
  xor g461 (n_746, A[14], n_217);
  xor g462 (n_221, n_746, n_218);
  nand g463 (n_747, A[14], n_217);
  nand g464 (n_748, n_218, n_217);
  nand g465 (n_749, A[14], n_218);
  nand g466 (n_225, n_747, n_748, n_749);
  xor g467 (n_750, n_219, n_220);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, n_219, n_220);
  nand g470 (n_752, n_221, n_220);
  nand g471 (n_753, n_219, n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g482 (n_72, n_638, A[8]);
  nand g484 (n_760, A[8], n_176);
  nand g485 (n_761, A[5], A[8]);
  nand g486 (n_232, n_639, n_760, n_761);
  xor g487 (n_762, n_71, A[9]);
  xor g488 (n_223, n_762, A[12]);
  nand g489 (n_763, n_71, A[9]);
  nand g491 (n_765, n_71, A[12]);
  nand g492 (n_234, n_763, n_707, n_765);
  xor g493 (n_766, n_72, A[13]);
  xor g494 (n_226, n_766, n_73);
  nand g495 (n_767, n_72, A[13]);
  nand g496 (n_768, n_73, A[13]);
  nand g497 (n_769, n_72, n_73);
  nand g498 (n_235, n_767, n_768, n_769);
  xor g499 (n_770, A[15], n_223);
  xor g500 (n_227, n_770, n_224);
  nand g501 (n_771, A[15], n_223);
  nand g502 (n_772, n_224, n_223);
  nand g503 (n_773, A[15], n_224);
  nand g504 (n_238, n_771, n_772, n_773);
  xor g505 (n_774, n_225, n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, n_225, n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, n_225, n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g518 (n_231, n_646, n_179);
  nand g521 (n_785, n_178, n_179);
  nand g522 (n_242, n_647, n_700, n_785);
  xor g523 (n_786, A[6], n_231);
  xor g524 (n_233, n_786, A[9]);
  nand g525 (n_787, A[6], n_231);
  nand g526 (n_788, A[9], n_231);
  nand g527 (n_789, A[6], A[9]);
  nand g528 (n_244, n_787, n_788, n_789);
  xor g529 (n_790, A[10], A[14]);
  xor g530 (n_236, n_790, A[13]);
  nand g531 (n_791, A[10], A[14]);
  nand g532 (n_792, A[13], A[14]);
  nand g533 (n_793, A[10], A[13]);
  nand g534 (n_246, n_791, n_792, n_793);
  xor g535 (n_794, n_232, n_233);
  xor g536 (n_237, n_794, n_234);
  nand g537 (n_795, n_232, n_233);
  nand g538 (n_796, n_234, n_233);
  nand g539 (n_797, n_232, n_234);
  nand g540 (n_248, n_795, n_796, n_797);
  xor g541 (n_798, n_235, n_236);
  xor g542 (n_239, n_798, A[16]);
  nand g543 (n_799, n_235, n_236);
  nand g544 (n_800, A[16], n_236);
  nand g545 (n_801, n_235, A[16]);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, n_237, n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, n_237, n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, n_237, n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g565 (n_814, n_242, A[10]);
  xor g566 (n_245, n_814, n_184);
  nand g567 (n_815, n_242, A[10]);
  nand g569 (n_817, n_242, n_184);
  nand g570 (n_257, n_815, n_724, n_817);
  xor g571 (n_818, A[11], A[14]);
  xor g572 (n_247, n_818, n_244);
  nand g573 (n_819, A[11], A[14]);
  nand g574 (n_820, n_244, A[14]);
  nand g575 (n_821, A[11], n_244);
  nand g576 (n_259, n_819, n_820, n_821);
  xor g577 (n_822, A[15], n_245);
  xor g578 (n_249, n_822, n_246);
  nand g579 (n_823, A[15], n_245);
  nand g580 (n_824, n_246, n_245);
  nand g581 (n_825, A[15], n_246);
  nand g582 (n_261, n_823, n_824, n_825);
  xor g583 (n_826, n_247, n_248);
  xor g584 (n_251, n_826, A[17]);
  nand g585 (n_827, n_247, n_248);
  nand g586 (n_828, A[17], n_248);
  nand g587 (n_829, n_247, A[17]);
  nand g588 (n_118, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g609 (n_842, n_188, A[11]);
  xor g610 (n_258, n_842, A[12]);
  xor g615 (n_846, n_218, A[15]);
  xor g616 (n_260, n_846, n_257);
  nand g617 (n_847, n_218, A[15]);
  nand g618 (n_848, n_257, A[15]);
  nand g619 (n_849, n_218, n_257);
  nand g620 (n_271, n_847, n_848, n_849);
  xor g621 (n_850, n_258, n_259);
  xor g622 (n_262, n_850, A[16]);
  nand g623 (n_851, n_258, n_259);
  nand g624 (n_852, A[16], n_259);
  nand g625 (n_853, n_258, A[16]);
  nand g626 (n_274, n_851, n_852, n_853);
  xor g627 (n_854, n_260, A[18]);
  xor g628 (n_119, n_854, n_261);
  nand g629 (n_855, n_260, A[18]);
  nand g630 (n_856, n_261, A[18]);
  nand g631 (n_857, n_260, n_261);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_262, n_118);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_262, n_118);
  nand g636 (n_860, n_119, n_118);
  nand g637 (n_861, n_262, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g641 (n_862, n_68, A[4]);
  xor g642 (n_265, n_862, n_69);
  xor g647 (n_866, A[5], n_265);
  xor g648 (n_268, n_866, A[8]);
  nand g649 (n_867, A[5], n_265);
  nand g650 (n_868, A[8], n_265);
  nand g652 (n_282, n_867, n_868, n_761);
  xor g659 (n_874, A[13], n_73);
  xor g660 (n_272, n_874, n_268);
  nand g662 (n_876, n_268, n_73);
  nand g663 (n_877, A[13], n_268);
  nand g664 (n_285, n_768, n_876, n_877);
  xor g665 (n_878, n_224, n_223);
  xor g666 (n_273, n_878, n_271);
  nand g668 (n_880, n_271, n_223);
  nand g669 (n_881, n_224, n_271);
  nand g670 (n_288, n_772, n_880, n_881);
  xor g671 (n_882, A[16], n_272);
  xor g672 (n_275, n_882, A[17]);
  nand g673 (n_883, A[16], n_272);
  nand g674 (n_884, A[17], n_272);
  nand g675 (n_885, A[16], A[17]);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, A[19], n_273);
  xor g678 (n_277, n_886, n_274);
  nand g679 (n_887, A[19], n_273);
  nand g680 (n_888, n_274, n_273);
  nand g681 (n_889, A[19], n_274);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g702 (n_283, n_650, A[10]);
  nand g704 (n_904, A[10], n_180);
  nand g705 (n_905, n_179, A[10]);
  nand g706 (n_298, n_651, n_904, n_905);
  xor g707 (n_906, A[9], A[13]);
  xor g708 (n_286, n_906, n_282);
  nand g709 (n_907, A[9], A[13]);
  nand g710 (n_908, n_282, A[13]);
  nand g711 (n_909, A[9], n_282);
  nand g712 (n_300, n_907, n_908, n_909);
  xor g713 (n_910, A[14], n_283);
  xor g714 (n_287, n_910, n_234);
  nand g715 (n_911, A[14], n_283);
  nand g716 (n_912, n_234, n_283);
  nand g717 (n_913, A[14], n_234);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, n_285, n_286);
  xor g720 (n_289, n_914, A[18]);
  nand g721 (n_915, n_285, n_286);
  nand g722 (n_916, A[18], n_286);
  nand g723 (n_917, n_285, A[18]);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, n_287, A[17]);
  xor g726 (n_291, n_918, A[20]);
  nand g727 (n_919, n_287, A[17]);
  nand g728 (n_920, A[20], A[17]);
  nand g729 (n_921, n_287, A[20]);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, n_288, n_289);
  xor g732 (n_293, n_922, n_290);
  nand g733 (n_923, n_288, n_289);
  nand g734 (n_924, n_290, n_289);
  nand g735 (n_925, n_288, n_290);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g755 (n_938, n_183, A[10]);
  xor g756 (n_299, n_938, n_184);
  nand g757 (n_939, n_183, A[10]);
  nand g760 (n_315, n_939, n_724, n_663);
  xor g762 (n_301, n_818, A[15]);
  nand g764 (n_944, A[15], A[14]);
  nand g765 (n_945, A[11], A[15]);
  nand g766 (n_317, n_819, n_944, n_945);
  xor g767 (n_946, n_298, n_299);
  xor g768 (n_303, n_946, n_300);
  nand g769 (n_947, n_298, n_299);
  nand g770 (n_948, n_300, n_299);
  nand g771 (n_949, n_298, n_300);
  nand g772 (n_319, n_947, n_948, n_949);
  xor g773 (n_950, n_301, n_302);
  xor g774 (n_305, n_950, A[19]);
  nand g775 (n_951, n_301, n_302);
  nand g776 (n_952, A[19], n_302);
  nand g777 (n_953, n_301, A[19]);
  nand g778 (n_320, n_951, n_952, n_953);
  xor g779 (n_954, A[18], n_303);
  xor g780 (n_307, n_954, A[21]);
  nand g781 (n_955, A[18], n_303);
  nand g782 (n_956, A[21], n_303);
  nand g783 (n_957, A[18], A[21]);
  nand g784 (n_322, n_955, n_956, n_957);
  xor g785 (n_958, n_304, n_305);
  xor g786 (n_309, n_958, n_306);
  nand g787 (n_959, n_304, n_305);
  nand g788 (n_960, n_306, n_305);
  nand g789 (n_961, n_304, n_306);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g817 (n_978, n_218, n_315);
  xor g818 (n_318, n_978, A[15]);
  nand g819 (n_979, n_218, n_315);
  nand g820 (n_980, A[15], n_315);
  nand g822 (n_335, n_979, n_980, n_847);
  xor g823 (n_982, n_219, n_317);
  xor g824 (n_321, n_982, A[16]);
  nand g825 (n_983, n_219, n_317);
  nand g826 (n_984, A[16], n_317);
  nand g827 (n_985, n_219, A[16]);
  nand g828 (n_337, n_983, n_984, n_985);
  xor g829 (n_986, A[19], n_318);
  xor g830 (n_323, n_986, A[20]);
  nand g831 (n_987, A[19], n_318);
  nand g832 (n_988, A[20], n_318);
  nand g833 (n_989, A[19], A[20]);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, n_319, A[22]);
  xor g836 (n_324, n_990, n_320);
  nand g837 (n_991, n_319, A[22]);
  nand g838 (n_992, n_320, A[22]);
  nand g839 (n_993, n_319, n_320);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, n_321, n_322);
  xor g842 (n_326, n_994, n_323);
  nand g843 (n_995, n_321, n_322);
  nand g844 (n_996, n_323, n_322);
  nand g845 (n_997, n_321, n_323);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, n_324, n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, n_324, n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, n_324, n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g873 (n_1014, n_73, n_268);
  xor g874 (n_336, n_1014, A[13]);
  xor g880 (n_338, n_878, n_335);
  nand g882 (n_1020, n_335, n_223);
  nand g883 (n_1021, n_224, n_335);
  nand g884 (n_358, n_772, n_1020, n_1021);
  xor g885 (n_1022, A[16], n_336);
  xor g886 (n_339, n_1022, A[17]);
  nand g887 (n_1023, A[16], n_336);
  nand g888 (n_1024, A[17], n_336);
  nand g890 (n_359, n_1023, n_1024, n_885);
  xor g891 (n_1026, A[21], A[20]);
  xor g892 (n_341, n_1026, A[23]);
  nand g893 (n_1027, A[21], A[20]);
  nand g894 (n_1028, A[23], A[20]);
  nand g895 (n_1029, A[21], A[23]);
  nand g896 (n_363, n_1027, n_1028, n_1029);
  xor g897 (n_1030, n_337, n_338);
  xor g898 (n_343, n_1030, n_339);
  nand g899 (n_1031, n_337, n_338);
  nand g900 (n_1032, n_339, n_338);
  nand g901 (n_1033, n_337, n_339);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, n_340, n_341);
  xor g904 (n_345, n_1034, n_342);
  nand g905 (n_1035, n_340, n_341);
  nand g906 (n_1036, n_342, n_341);
  nand g907 (n_1037, n_340, n_342);
  nand g908 (n_367, n_1035, n_1036, n_1037);
  xor g909 (n_1038, n_343, n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, n_343, n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, n_343, n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  xor g917 (n_1042, A[2], n_171);
  nand g922 (n_371, n_624, n_1044, n_1045);
  xor g923 (n_1046, n_349, A[5]);
  xor g924 (n_351, n_1046, n_179);
  nand g925 (n_1047, n_349, A[5]);
  nand g927 (n_1049, n_349, n_179);
  nand g928 (n_373, n_1047, n_700, n_1049);
  xor g929 (n_1050, A[6], n_351);
  xor g930 (n_353, n_1050, A[9]);
  nand g931 (n_1051, A[6], n_351);
  nand g932 (n_1052, A[9], n_351);
  nand g934 (n_375, n_1051, n_1052, n_789);
  xor g936 (n_356, n_790, n_282);
  nand g938 (n_1056, n_282, A[14]);
  nand g939 (n_1057, A[10], n_282);
  nand g940 (n_377, n_791, n_1056, n_1057);
  xor g941 (n_1058, A[13], n_353);
  xor g942 (n_357, n_1058, n_234);
  nand g943 (n_1059, A[13], n_353);
  nand g944 (n_1060, n_234, n_353);
  nand g945 (n_1061, A[13], n_234);
  nand g946 (n_379, n_1059, n_1060, n_1061);
  xor g947 (n_1062, n_285, n_356);
  xor g948 (n_360, n_1062, A[17]);
  nand g949 (n_1063, n_285, n_356);
  nand g950 (n_1064, A[17], n_356);
  nand g951 (n_1065, n_285, A[17]);
  nand g952 (n_381, n_1063, n_1064, n_1065);
  xor g953 (n_1066, A[18], n_357);
  xor g954 (n_361, n_1066, A[22]);
  nand g955 (n_1067, A[18], n_357);
  nand g956 (n_1068, A[22], n_357);
  nand g957 (n_1069, A[18], A[22]);
  nand g958 (n_384, n_1067, n_1068, n_1069);
  xor g960 (n_362, n_1070, n_358);
  nand g962 (n_1072, n_358, A[21]);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, n_359, n_360);
  xor g966 (n_365, n_1074, n_361);
  nand g967 (n_1075, n_359, n_360);
  nand g968 (n_1076, n_361, n_360);
  nand g969 (n_1077, n_359, n_361);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g971 (n_1078, n_362, n_363);
  xor g972 (n_366, n_1078, n_364);
  nand g973 (n_1079, n_362, n_363);
  nand g974 (n_1080, n_364, n_363);
  nand g975 (n_1081, n_362, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  xor g985 (n_1086, A[1], A[3]);
  nand g987 (n_1087, A[1], A[3]);
  nand g990 (n_392, n_1087, n_1088, n_1089);
  xor g991 (n_1090, n_371, n_372);
  xor g992 (n_374, n_1090, A[6]);
  nand g993 (n_1091, n_371, n_372);
  nand g994 (n_1092, A[6], n_372);
  nand g995 (n_1093, n_371, A[6]);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, n_374);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, n_374, n_373);
  nand g1001 (n_1097, A[7], n_374);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, A[10], A[11]);
  xor g1004 (n_378, n_1098, A[14]);
  nand g1005 (n_1099, A[10], A[11]);
  nand g1008 (n_398, n_1099, n_819, n_791);
  xor g1009 (n_1102, n_375, n_376);
  xor g1010 (n_380, n_1102, A[15]);
  nand g1011 (n_1103, n_375, n_376);
  nand g1012 (n_1104, A[15], n_376);
  nand g1013 (n_1105, n_375, A[15]);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, n_377, n_378);
  xor g1016 (n_382, n_1106, A[19]);
  nand g1017 (n_1107, n_377, n_378);
  nand g1018 (n_1108, A[19], n_378);
  nand g1019 (n_1109, n_377, A[19]);
  nand g1020 (n_403, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, n_379, A[18]);
  xor g1022 (n_383, n_1110, n_380);
  nand g1023 (n_1111, n_379, A[18]);
  nand g1024 (n_1112, n_380, A[18]);
  nand g1025 (n_1113, n_379, n_380);
  nand g1026 (n_402, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, A[22], A[23]);
  xor g1028 (n_386, n_1114, n_381);
  nand g1029 (n_1115, A[22], A[23]);
  nand g1030 (n_1116, n_381, A[23]);
  nand g1031 (n_1117, A[22], n_381);
  nand g1032 (n_407, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_382, n_383);
  xor g1034 (n_388, n_1118, n_384);
  nand g1035 (n_1119, n_382, n_383);
  nand g1036 (n_1120, n_384, n_383);
  nand g1037 (n_1121, n_382, n_384);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, n_385, n_386);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, n_385, n_386);
  nand g1042 (n_1124, n_387, n_386);
  nand g1043 (n_1125, n_385, n_387);
  nand g1044 (n_411, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1052 (n_393, n_626, A[4]);
  nand g1054 (n_1132, A[4], A[2]);
  nand g1055 (n_1133, A[3], A[4]);
  nand g1056 (n_412, n_627, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, A[11], A[12]);
  xor g1070 (n_399, n_1142, n_396);
  nand g1072 (n_1144, n_396, A[12]);
  nand g1073 (n_1145, A[11], n_396);
  nand g1074 (n_418, n_744, n_1144, n_1145);
  xor g1075 (n_1146, n_397, A[15]);
  xor g1076 (n_401, n_1146, n_398);
  nand g1077 (n_1147, n_397, A[15]);
  nand g1078 (n_1148, n_398, A[15]);
  nand g1079 (n_1149, n_397, n_398);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, n_399, n_400);
  xor g1082 (n_404, n_1150, A[16]);
  nand g1083 (n_1151, n_399, n_400);
  nand g1084 (n_1152, A[16], n_400);
  nand g1085 (n_1153, n_399, A[16]);
  nand g1086 (n_421, n_1151, n_1152, n_1153);
  xor g1088 (n_405, n_1154, A[20]);
  nand g1092 (n_423, n_1155, n_1156, n_989);
  xor g1093 (n_1158, n_401, A[23]);
  xor g1094 (n_406, n_1158, n_402);
  nand g1095 (n_1159, n_401, A[23]);
  nand g1096 (n_1160, n_402, A[23]);
  nand g1097 (n_1161, n_401, n_402);
  nand g1098 (n_426, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_403, n_404);
  xor g1100 (n_409, n_1162, n_405);
  nand g1101 (n_1163, n_403, n_404);
  nand g1102 (n_1164, n_405, n_404);
  nand g1103 (n_1165, n_403, n_405);
  nand g1104 (n_427, n_1163, n_1164, n_1165);
  xor g1105 (n_1166, n_406, n_407);
  xor g1106 (n_410, n_1166, n_408);
  nand g1107 (n_1167, n_406, n_407);
  nand g1108 (n_1168, n_408, n_407);
  nand g1109 (n_1169, n_406, n_408);
  nand g1110 (n_429, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1123 (n_1178, A[8], n_413);
  xor g1124 (n_415, n_1178, A[9]);
  nand g1125 (n_1179, A[8], n_413);
  nand g1126 (n_1180, A[9], n_413);
  nand g1128 (n_435, n_1179, n_1180, n_687);
  xor g1129 (n_1182, n_414, A[12]);
  xor g1130 (n_417, n_1182, A[13]);
  nand g1131 (n_1183, n_414, A[12]);
  nand g1132 (n_1184, A[13], A[12]);
  nand g1133 (n_1185, n_414, A[13]);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, n_415, n_416);
  xor g1136 (n_420, n_1186, n_417);
  nand g1137 (n_1187, n_415, n_416);
  nand g1138 (n_1188, n_417, n_416);
  nand g1139 (n_1189, n_415, n_417);
  nand g1140 (n_439, n_1187, n_1188, n_1189);
  xor g1141 (n_1190, n_418, A[16]);
  xor g1142 (n_422, n_1190, A[17]);
  nand g1143 (n_1191, n_418, A[16]);
  nand g1145 (n_1193, n_418, A[17]);
  nand g1146 (n_441, n_1191, n_885, n_1193);
  xor g1148 (n_425, n_1194, n_420);
  nand g1151 (n_1197, n_419, n_420);
  nand g1152 (n_442, n_1195, n_1196, n_1197);
  xor g1154 (n_424, n_1026, n_421);
  nand g1156 (n_1200, n_421, A[21]);
  nand g1157 (n_1201, A[20], n_421);
  nand g1158 (n_445, n_1027, n_1200, n_1201);
  xor g1159 (n_1202, n_422, n_423);
  xor g1160 (n_428, n_1202, n_424);
  nand g1161 (n_1203, n_422, n_423);
  nand g1162 (n_1204, n_424, n_423);
  nand g1163 (n_1205, n_422, n_424);
  nand g1164 (n_446, n_1203, n_1204, n_1205);
  xor g1165 (n_1206, n_425, n_426);
  xor g1166 (n_430, n_1206, n_427);
  nand g1167 (n_1207, n_425, n_426);
  nand g1168 (n_1208, n_427, n_426);
  nand g1169 (n_1209, n_425, n_427);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, n_433);
  nand g1183 (n_1217, A[6], n_433);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, A[9], A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, A[9], A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, A[9], n_434);
  nand g1190 (n_456, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, A[14], A[13]);
  xor g1192 (n_438, n_1222, n_435);
  nand g1194 (n_1224, n_435, A[13]);
  nand g1195 (n_1225, A[14], n_435);
  nand g1196 (n_458, n_792, n_1224, n_1225);
  xor g1197 (n_1226, n_436, n_437);
  xor g1198 (n_440, n_1226, n_438);
  nand g1199 (n_1227, n_436, n_437);
  nand g1200 (n_1228, n_438, n_437);
  nand g1201 (n_1229, n_436, n_438);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, A[18], A[17]);
  xor g1204 (n_443, n_1230, A[21]);
  nand g1205 (n_1231, A[18], A[17]);
  nand g1206 (n_1232, A[21], A[17]);
  nand g1208 (n_462, n_1231, n_1232, n_957);
  xor g1209 (n_1234, A[22], n_439);
  xor g1210 (n_444, n_1234, n_440);
  nand g1211 (n_1235, A[22], n_439);
  nand g1212 (n_1236, n_440, n_439);
  nand g1213 (n_1237, A[22], n_440);
  nand g1214 (n_463, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_441, n_442);
  xor g1216 (n_447, n_1238, n_443);
  nand g1217 (n_1239, n_441, n_442);
  nand g1218 (n_1240, n_443, n_442);
  nand g1219 (n_1241, n_441, n_443);
  nand g1220 (n_465, n_1239, n_1240, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[7], A[5]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1242 (n_455, n_1098, n_453);
  nand g1244 (n_1256, n_453, A[11]);
  nand g1245 (n_1257, A[10], n_453);
  nand g1246 (n_472, n_1099, n_1256, n_1257);
  xor g1247 (n_1258, A[14], n_454);
  xor g1248 (n_457, n_1258, A[15]);
  nand g1249 (n_1259, A[14], n_454);
  nand g1250 (n_1260, A[15], n_454);
  nand g1252 (n_474, n_1259, n_1260, n_944);
  xor g1253 (n_1262, n_455, n_456);
  xor g1254 (n_460, n_1262, n_457);
  nand g1255 (n_1263, n_455, n_456);
  nand g1256 (n_1264, n_457, n_456);
  nand g1257 (n_1265, n_455, n_457);
  nand g1258 (n_476, n_1263, n_1264, n_1265);
  xor g1259 (n_1266, n_458, A[19]);
  xor g1260 (n_461, n_1266, A[18]);
  nand g1261 (n_1267, n_458, A[19]);
  nand g1262 (n_1268, A[18], A[19]);
  nand g1263 (n_1269, n_458, A[18]);
  nand g1264 (n_477, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, A[22], n_459);
  xor g1266 (n_464, n_1270, A[23]);
  nand g1267 (n_1271, A[22], n_459);
  nand g1268 (n_1272, A[23], n_459);
  nand g1270 (n_480, n_1271, n_1272, n_1115);
  xor g1271 (n_1274, n_460, n_461);
  xor g1272 (n_466, n_1274, n_462);
  nand g1273 (n_1275, n_460, n_461);
  nand g1274 (n_1276, n_462, n_461);
  nand g1275 (n_1277, n_460, n_462);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1277 (n_1278, n_463, n_464);
  xor g1278 (n_467, n_1278, n_465);
  nand g1279 (n_1279, n_463, n_464);
  nand g1280 (n_1280, n_465, n_464);
  nand g1281 (n_1281, n_463, n_465);
  nand g1282 (n_485, n_1279, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1289 (n_1286, A[7], A[6]);
  xor g1290 (n_471, n_1286, A[8]);
  nand g1292 (n_1288, A[8], A[6]);
  nand g1294 (n_486, n_661, n_1288, n_673);
  xor g1296 (n_473, n_1142, n_470);
  nand g1298 (n_1292, n_470, A[12]);
  nand g1299 (n_1293, A[11], n_470);
  nand g1300 (n_487, n_744, n_1292, n_1293);
  xor g1301 (n_1294, n_471, A[15]);
  xor g1302 (n_475, n_1294, n_472);
  nand g1303 (n_1295, n_471, A[15]);
  nand g1304 (n_1296, n_472, A[15]);
  nand g1305 (n_1297, n_471, n_472);
  nand g1306 (n_489, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, n_473, A[16]);
  xor g1308 (n_478, n_1298, n_474);
  nand g1309 (n_1299, n_473, A[16]);
  nand g1310 (n_1300, n_474, A[16]);
  nand g1311 (n_1301, n_473, n_474);
  nand g1312 (n_491, n_1299, n_1300, n_1301);
  xor g1313 (n_1302, A[19], n_475);
  nand g1315 (n_1303, A[19], n_475);
  nand g1318 (n_493, n_1303, n_1304, n_1155);
  xor g1319 (n_1306, A[20], n_476);
  xor g1320 (n_481, n_1306, A[23]);
  nand g1321 (n_1307, A[20], n_476);
  nand g1322 (n_1308, A[23], n_476);
  nand g1324 (n_495, n_1307, n_1308, n_1028);
  xor g1325 (n_1310, n_477, n_478);
  xor g1326 (n_483, n_1310, n_479);
  nand g1327 (n_1311, n_477, n_478);
  nand g1328 (n_1312, n_479, n_478);
  nand g1329 (n_1313, n_477, n_479);
  nand g1330 (n_497, n_1311, n_1312, n_1313);
  xor g1331 (n_1314, n_480, n_481);
  xor g1332 (n_484, n_1314, n_482);
  nand g1333 (n_1315, n_480, n_481);
  nand g1334 (n_1316, n_482, n_481);
  nand g1335 (n_1317, n_480, n_482);
  nand g1336 (n_500, n_1315, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1344 (n_488, n_686, A[12]);
  nand g1347 (n_1325, A[8], A[12]);
  nand g1348 (n_503, n_687, n_707, n_1325);
  xor g1349 (n_1326, n_486, A[13]);
  xor g1350 (n_490, n_1326, n_487);
  nand g1351 (n_1327, n_486, A[13]);
  nand g1352 (n_1328, n_487, A[13]);
  nand g1353 (n_1329, n_486, n_487);
  nand g1354 (n_505, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, n_488, A[16]);
  xor g1356 (n_492, n_1330, A[17]);
  nand g1357 (n_1331, n_488, A[16]);
  nand g1359 (n_1333, n_488, A[17]);
  nand g1360 (n_507, n_1331, n_885, n_1333);
  xor g1361 (n_1334, n_489, n_490);
  nand g1363 (n_1335, n_489, n_490);
  nand g1366 (n_509, n_1335, n_1336, n_1337);
  xor g1368 (n_496, n_1026, n_491);
  nand g1370 (n_1340, n_491, A[20]);
  nand g1371 (n_1341, A[21], n_491);
  nand g1372 (n_511, n_1027, n_1340, n_1341);
  xor g1373 (n_1342, n_492, n_493);
  xor g1374 (n_498, n_1342, n_494);
  nand g1375 (n_1343, n_492, n_493);
  nand g1376 (n_1344, n_494, n_493);
  nand g1377 (n_1345, n_492, n_494);
  nand g1378 (n_512, n_1343, n_1344, n_1345);
  xor g1379 (n_1346, n_495, n_496);
  xor g1380 (n_499, n_1346, n_497);
  nand g1381 (n_1347, n_495, n_496);
  nand g1382 (n_1348, n_497, n_496);
  nand g1383 (n_1349, n_495, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  nand g1397 (n_1357, A[9], A[14]);
  nand g1398 (n_519, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], n_503);
  xor g1400 (n_506, n_1358, n_504);
  nand g1401 (n_1359, A[13], n_503);
  nand g1402 (n_1360, n_504, n_503);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_522, n_1359, n_1360, n_1361);
  xor g1406 (n_508, n_1230, n_505);
  nand g1408 (n_1364, n_505, A[17]);
  nand g1409 (n_1365, A[18], n_505);
  nand g1410 (n_523, n_1231, n_1364, n_1365);
  xor g1411 (n_1366, A[21], A[22]);
  xor g1412 (n_510, n_1366, n_506);
  nand g1413 (n_1367, A[21], A[22]);
  nand g1414 (n_1368, n_506, A[22]);
  nand g1415 (n_1369, A[21], n_506);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_507, n_508);
  xor g1418 (n_513, n_1370, n_509);
  nand g1419 (n_1371, n_507, n_508);
  nand g1420 (n_1372, n_509, n_508);
  nand g1421 (n_1373, n_507, n_509);
  nand g1422 (n_527, n_1371, n_1372, n_1373);
  xor g1423 (n_1374, n_510, n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, n_510, n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, n_510, n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1443 (n_1386, A[14], A[15]);
  xor g1444 (n_521, n_1386, n_519);
  nand g1446 (n_1388, n_519, A[15]);
  nand g1447 (n_1389, A[14], n_519);
  nand g1448 (n_534, n_944, n_1388, n_1389);
  xor g1449 (n_1390, n_520, A[19]);
  xor g1450 (n_524, n_1390, A[18]);
  nand g1451 (n_1391, n_520, A[19]);
  nand g1453 (n_1393, n_520, A[18]);
  nand g1454 (n_536, n_1391, n_1268, n_1393);
  xor g1455 (n_1394, A[22], n_521);
  xor g1456 (n_525, n_1394, A[23]);
  nand g1457 (n_1395, A[22], n_521);
  nand g1458 (n_1396, A[23], n_521);
  nand g1460 (n_539, n_1395, n_1396, n_1115);
  xor g1461 (n_1398, n_522, n_523);
  xor g1462 (n_528, n_1398, n_524);
  nand g1463 (n_1399, n_522, n_523);
  nand g1464 (n_1400, n_524, n_523);
  nand g1465 (n_1401, n_522, n_524);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1467 (n_1402, n_525, n_526);
  xor g1468 (n_529, n_1402, n_527);
  nand g1469 (n_1403, n_525, n_526);
  nand g1470 (n_1404, n_527, n_526);
  nand g1471 (n_1405, n_525, n_527);
  nand g1472 (n_543, n_1403, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1480 (n_533, n_1142, A[10]);
  nand g1483 (n_1413, A[12], A[10]);
  nand g1484 (n_544, n_744, n_1099, n_1413);
  xor g1485 (n_1414, A[15], n_532);
  xor g1486 (n_535, n_1414, n_533);
  nand g1487 (n_1415, A[15], n_532);
  nand g1488 (n_1416, n_533, n_532);
  nand g1489 (n_1417, A[15], n_533);
  nand g1490 (n_545, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, A[16], A[19]);
  nand g1493 (n_1419, A[16], A[19]);
  nand g1496 (n_548, n_1419, n_1155, n_1421);
  xor g1497 (n_1422, n_534, A[20]);
  xor g1498 (n_538, n_1422, A[23]);
  nand g1499 (n_1423, n_534, A[20]);
  nand g1501 (n_1425, n_534, A[23]);
  nand g1502 (n_549, n_1423, n_1028, n_1425);
  xor g1503 (n_1426, n_535, n_536);
  xor g1504 (n_541, n_1426, n_537);
  nand g1505 (n_1427, n_535, n_536);
  nand g1506 (n_1428, n_537, n_536);
  nand g1507 (n_1429, n_535, n_537);
  nand g1508 (n_551, n_1427, n_1428, n_1429);
  xor g1509 (n_1430, n_538, n_539);
  xor g1510 (n_542, n_1430, n_540);
  nand g1511 (n_1431, n_538, n_539);
  nand g1512 (n_1432, n_540, n_539);
  nand g1513 (n_1433, n_538, n_540);
  nand g1514 (n_554, n_1431, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1521 (n_1438, A[12], A[13]);
  xor g1522 (n_546, n_1438, n_544);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_1184, n_1440, n_1441);
  xor g1527 (n_1442, A[16], A[17]);
  xor g1528 (n_547, n_1442, A[21]);
  nand g1531 (n_1445, A[16], A[21]);
  nand g1532 (n_560, n_885, n_1232, n_1445);
  xor g1534 (n_550, n_1446, A[20]);
  nand g1537 (n_1449, n_545, A[20]);
  nand g1538 (n_559, n_1447, n_1156, n_1449);
  xor g1539 (n_1450, n_546, n_547);
  xor g1540 (n_552, n_1450, n_548);
  nand g1541 (n_1451, n_546, n_547);
  nand g1542 (n_1452, n_548, n_547);
  nand g1543 (n_1453, n_546, n_548);
  nand g1544 (n_563, n_1451, n_1452, n_1453);
  xor g1545 (n_1454, n_549, n_550);
  xor g1546 (n_553, n_1454, n_551);
  nand g1547 (n_1455, n_549, n_550);
  nand g1548 (n_1456, n_551, n_550);
  nand g1549 (n_1457, n_549, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1563 (n_1465, A[13], A[18]);
  nand g1564 (n_570, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, A[17], A[21]);
  xor g1566 (n_561, n_1466, n_557);
  nand g1568 (n_1468, n_557, A[21]);
  nand g1569 (n_1469, A[17], n_557);
  nand g1570 (n_572, n_1232, n_1468, n_1469);
  xor g1571 (n_1470, A[22], n_558);
  xor g1572 (n_562, n_1470, n_559);
  nand g1573 (n_1471, A[22], n_558);
  nand g1574 (n_1472, n_559, n_558);
  nand g1575 (n_1473, A[22], n_559);
  nand g1576 (n_574, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, n_560, n_561);
  xor g1578 (n_564, n_1474, n_562);
  nand g1579 (n_1475, n_560, n_561);
  nand g1580 (n_1476, n_562, n_561);
  nand g1581 (n_1477, n_560, n_562);
  nand g1582 (n_576, n_1475, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  xor g1597 (n_1486, A[19], A[18]);
  xor g1598 (n_571, n_1486, n_569);
  nand g1600 (n_1488, n_569, A[18]);
  nand g1601 (n_1489, A[19], n_569);
  nand g1602 (n_580, n_1268, n_1488, n_1489);
  xor g1604 (n_573, n_1114, n_570);
  nand g1606 (n_1492, n_570, A[23]);
  nand g1607 (n_1493, A[22], n_570);
  nand g1608 (n_583, n_1115, n_1492, n_1493);
  xor g1609 (n_1494, n_571, n_572);
  xor g1610 (n_575, n_1494, n_573);
  nand g1611 (n_1495, n_571, n_572);
  nand g1612 (n_1496, n_573, n_572);
  nand g1613 (n_1497, n_571, n_573);
  nand g1614 (n_585, n_1495, n_1496, n_1497);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1622 (n_579, n_1386, A[16]);
  nand g1624 (n_1504, A[16], A[14]);
  nand g1625 (n_1505, A[15], A[16]);
  nand g1626 (n_586, n_944, n_1504, n_1505);
  xor g1627 (n_1506, A[19], n_578);
  nand g1629 (n_1507, A[19], n_578);
  nand g1632 (n_588, n_1507, n_1508, n_1155);
  xor g1633 (n_1510, A[20], A[23]);
  xor g1634 (n_582, n_1510, n_579);
  nand g1636 (n_1512, n_579, A[23]);
  nand g1637 (n_1513, A[20], n_579);
  nand g1638 (n_589, n_1028, n_1512, n_1513);
  xor g1639 (n_1514, n_580, n_581);
  xor g1640 (n_584, n_1514, n_582);
  nand g1641 (n_1515, n_580, n_581);
  nand g1642 (n_1516, n_582, n_581);
  nand g1643 (n_1517, n_580, n_582);
  nand g1644 (n_592, n_1515, n_1516, n_1517);
  xor g1645 (n_1518, n_583, n_584);
  xor g1646 (n_83, n_1518, n_585);
  nand g1647 (n_1519, n_583, n_584);
  nand g1648 (n_1520, n_585, n_584);
  nand g1649 (n_1521, n_583, n_585);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1658 (n_590, n_1526, n_586);
  nand g1660 (n_1528, n_586, A[20]);
  nand g1662 (n_596, n_1156, n_1528, n_1529);
  xor g1663 (n_1530, n_547, n_588);
  xor g1664 (n_591, n_1530, n_589);
  nand g1665 (n_1531, n_547, n_588);
  nand g1666 (n_1532, n_589, n_588);
  nand g1667 (n_1533, n_547, n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_33, n_1535, n_1536, n_1537);
  xor g1678 (n_597, n_1466, A[22]);
  nand g1681 (n_1541, A[17], A[22]);
  nand g1682 (n_603, n_1232, n_1367, n_1541);
  xor g1684 (n_598, n_1542, n_596);
  nand g1686 (n_1544, n_596, n_560);
  nand g1688 (n_606, n_1543, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_81, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[18], A[22]);
  xor g1698 (n_604, n_1550, A[23]);
  nand g1701 (n_1553, A[18], A[23]);
  nand g1702 (n_609, n_1069, n_1115, n_1553);
  nand g1706 (n_1556, n_603, A[18]);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, n_604, n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, n_604, n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, n_604, n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1721 (n_1566, A[23], A[19]);
  xor g1722 (n_611, n_1566, n_405);
  nand g1723 (n_1567, A[23], A[19]);
  nand g1724 (n_1568, n_405, A[19]);
  nand g1725 (n_1569, A[23], n_405);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1727 (n_1570, n_609, n_610);
  xor g1728 (n_79, n_1570, n_611);
  nand g1729 (n_1571, n_609, n_610);
  nand g1730 (n_1572, n_611, n_610);
  nand g1731 (n_1573, n_609, n_611);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1734 (n_613, n_1070, A[20]);
  nand g1738 (n_617, n_1071, n_1027, n_1156);
  xor g1739 (n_1578, n_423, n_613);
  xor g1740 (n_78, n_1578, n_614);
  nand g1741 (n_1579, n_423, n_613);
  nand g1742 (n_1580, n_614, n_613);
  nand g1743 (n_1581, n_423, n_614);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_617);
  nand g1752 (n_28, n_1583, n_1584, n_1585);
  nand g1760 (n_27, n_1587, n_1588, n_1029);
  xor g1762 (n_75, n_1590, A[22]);
  nand g1766 (n_74, n_1591, n_1115, n_1593);
  nor g11 (n_1609, A[0], A[2]);
  nand g12 (n_1604, A[0], A[2]);
  nor g13 (n_1605, n_68, A[3]);
  nand g14 (n_1606, n_68, A[3]);
  nor g15 (n_1615, A[4], n_117);
  nand g16 (n_1610, A[4], n_117);
  nor g17 (n_1611, A[5], n_116);
  nand g18 (n_1612, A[5], n_116);
  nor g19 (n_1621, n_67, n_115);
  nand g20 (n_1616, n_67, n_115);
  nor g21 (n_1617, n_66, n_114);
  nand g22 (n_1618, n_66, n_114);
  nor g23 (n_1627, n_65, n_113);
  nand g24 (n_1622, n_65, n_113);
  nor g25 (n_1623, n_64, n_112);
  nand g26 (n_1624, n_64, n_112);
  nor g27 (n_1633, n_63, n_111);
  nand g28 (n_1628, n_63, n_111);
  nor g29 (n_1629, n_62, n_110);
  nand g30 (n_1630, n_62, n_110);
  nor g31 (n_1639, n_61, n_109);
  nand g32 (n_1634, n_61, n_109);
  nor g33 (n_1635, n_60, n_108);
  nand g34 (n_1636, n_60, n_108);
  nor g35 (n_1645, n_59, n_107);
  nand g36 (n_1640, n_59, n_107);
  nor g37 (n_1641, n_58, n_106);
  nand g38 (n_1642, n_58, n_106);
  nor g39 (n_1651, n_57, n_105);
  nand g40 (n_1646, n_57, n_105);
  nor g41 (n_1647, n_56, n_104);
  nand g42 (n_1648, n_56, n_104);
  nor g43 (n_1657, n_55, n_103);
  nand g44 (n_1652, n_55, n_103);
  nor g45 (n_1653, n_54, n_102);
  nand g46 (n_1654, n_54, n_102);
  nor g47 (n_1663, n_53, n_101);
  nand g48 (n_1658, n_53, n_101);
  nor g49 (n_1659, n_52, n_100);
  nand g50 (n_1660, n_52, n_100);
  nor g51 (n_1669, n_51, n_99);
  nand g52 (n_1664, n_51, n_99);
  nor g53 (n_1665, n_50, n_98);
  nand g54 (n_1666, n_50, n_98);
  nor g55 (n_1675, n_49, n_97);
  nand g56 (n_1670, n_49, n_97);
  nor g57 (n_1671, n_48, n_96);
  nand g58 (n_1672, n_48, n_96);
  nor g59 (n_1681, n_47, n_95);
  nand g60 (n_1676, n_47, n_95);
  nor g61 (n_1677, n_46, n_94);
  nand g62 (n_1678, n_46, n_94);
  nor g63 (n_1687, n_45, n_93);
  nand g64 (n_1682, n_45, n_93);
  nor g65 (n_1683, n_44, n_92);
  nand g66 (n_1684, n_44, n_92);
  nor g67 (n_1693, n_43, n_91);
  nand g68 (n_1688, n_43, n_91);
  nor g69 (n_1689, n_42, n_90);
  nand g70 (n_1690, n_42, n_90);
  nor g71 (n_1699, n_41, n_89);
  nand g72 (n_1694, n_41, n_89);
  nor g73 (n_1695, n_40, n_88);
  nand g74 (n_1696, n_40, n_88);
  nor g75 (n_1705, n_39, n_87);
  nand g76 (n_1700, n_39, n_87);
  nor g77 (n_1701, n_38, n_86);
  nand g78 (n_1702, n_38, n_86);
  nor g79 (n_1711, n_37, n_85);
  nand g80 (n_1706, n_37, n_85);
  nor g81 (n_1707, n_36, n_84);
  nand g82 (n_1708, n_36, n_84);
  nor g83 (n_1717, n_35, n_83);
  nand g84 (n_1712, n_35, n_83);
  nor g85 (n_1713, n_34, n_82);
  nand g86 (n_1714, n_34, n_82);
  nor g87 (n_1723, n_33, n_81);
  nand g88 (n_1718, n_33, n_81);
  nor g89 (n_1719, n_32, n_80);
  nand g90 (n_1720, n_32, n_80);
  nor g91 (n_1729, n_31, n_79);
  nand g92 (n_1724, n_31, n_79);
  nor g93 (n_1725, n_30, n_78);
  nand g94 (n_1726, n_30, n_78);
  nor g95 (n_1735, n_29, n_77);
  nand g96 (n_1730, n_29, n_77);
  nor g97 (n_1731, n_28, n_76);
  nand g98 (n_1732, n_28, n_76);
  nor g99 (n_1739, n_27, n_75);
  nand g100 (n_1736, n_27, n_75);
  nor g106 (n_1607, n_1604, n_1605);
  nor g110 (n_1613, n_1610, n_1611);
  nor g113 (n_1749, n_1615, n_1611);
  nor g114 (n_1619, n_1616, n_1617);
  nor g117 (n_1751, n_1621, n_1617);
  nor g118 (n_1625, n_1622, n_1623);
  nor g121 (n_1759, n_1627, n_1623);
  nor g122 (n_1631, n_1628, n_1629);
  nor g125 (n_1761, n_1633, n_1629);
  nor g126 (n_1637, n_1634, n_1635);
  nor g129 (n_1769, n_1639, n_1635);
  nor g130 (n_1643, n_1640, n_1641);
  nor g133 (n_1771, n_1645, n_1641);
  nor g134 (n_1649, n_1646, n_1647);
  nor g137 (n_1779, n_1651, n_1647);
  nor g138 (n_1655, n_1652, n_1653);
  nor g141 (n_1781, n_1657, n_1653);
  nor g142 (n_1661, n_1658, n_1659);
  nor g145 (n_1789, n_1663, n_1659);
  nor g146 (n_1667, n_1664, n_1665);
  nor g149 (n_1791, n_1669, n_1665);
  nor g150 (n_1673, n_1670, n_1671);
  nor g153 (n_1799, n_1675, n_1671);
  nor g154 (n_1679, n_1676, n_1677);
  nor g157 (n_1801, n_1681, n_1677);
  nor g158 (n_1685, n_1682, n_1683);
  nor g161 (n_1809, n_1687, n_1683);
  nor g162 (n_1691, n_1688, n_1689);
  nor g165 (n_1811, n_1693, n_1689);
  nor g166 (n_1697, n_1694, n_1695);
  nor g169 (n_1819, n_1699, n_1695);
  nor g170 (n_1703, n_1700, n_1701);
  nor g173 (n_1821, n_1705, n_1701);
  nor g174 (n_1709, n_1706, n_1707);
  nor g177 (n_1829, n_1711, n_1707);
  nor g178 (n_1715, n_1712, n_1713);
  nor g181 (n_1831, n_1717, n_1713);
  nor g182 (n_1721, n_1718, n_1719);
  nor g185 (n_1839, n_1723, n_1719);
  nor g186 (n_1727, n_1724, n_1725);
  nor g189 (n_1841, n_1729, n_1725);
  nor g190 (n_1733, n_1730, n_1731);
  nor g193 (n_1849, n_1735, n_1731);
  nor g203 (n_1747, n_1621, n_1746);
  nand g212 (n_1859, n_1749, n_1751);
  nor g213 (n_1757, n_1633, n_1756);
  nand g222 (n_1866, n_1759, n_1761);
  nor g223 (n_1767, n_1645, n_1766);
  nand g232 (n_1874, n_1769, n_1771);
  nor g233 (n_1777, n_1657, n_1776);
  nand g242 (n_1881, n_1779, n_1781);
  nor g243 (n_1787, n_1669, n_1786);
  nand g252 (n_1889, n_1789, n_1791);
  nor g253 (n_1797, n_1681, n_1796);
  nand g262 (n_1896, n_1799, n_1801);
  nor g263 (n_1807, n_1693, n_1806);
  nand g1776 (n_1904, n_1809, n_1811);
  nor g1777 (n_1817, n_1705, n_1816);
  nand g1786 (n_1911, n_1819, n_1821);
  nor g1787 (n_1827, n_1717, n_1826);
  nand g1796 (n_1919, n_1829, n_1831);
  nor g1797 (n_1837, n_1729, n_1836);
  nand g1806 (n_1926, n_1839, n_1841);
  nor g1807 (n_1847, n_1739, n_1846);
  nand g1814 (n_2130, n_1610, n_1853);
  nand g1816 (n_2132, n_1746, n_1854);
  nand g1819 (n_2135, n_1857, n_1858);
  nand g1822 (n_1934, n_1861, n_1862);
  nor g1823 (n_1864, n_1639, n_1863);
  nor g1826 (n_1944, n_1639, n_1866);
  nor g1832 (n_1872, n_1870, n_1863);
  nor g1835 (n_1950, n_1866, n_1870);
  nor g1836 (n_1876, n_1874, n_1863);
  nor g1839 (n_1953, n_1866, n_1874);
  nor g1840 (n_1879, n_1663, n_1878);
  nor g1843 (n_2033, n_1663, n_1881);
  nor g1849 (n_1887, n_1885, n_1878);
  nor g1852 (n_2039, n_1881, n_1885);
  nor g1853 (n_1891, n_1889, n_1878);
  nor g1856 (n_1959, n_1881, n_1889);
  nor g1857 (n_1894, n_1687, n_1893);
  nor g1860 (n_1972, n_1687, n_1896);
  nor g1866 (n_1902, n_1900, n_1893);
  nor g1869 (n_1982, n_1896, n_1900);
  nor g1870 (n_1906, n_1904, n_1893);
  nor g1873 (n_1987, n_1896, n_1904);
  nor g1874 (n_1909, n_1711, n_1908);
  nor g1877 (n_2085, n_1711, n_1911);
  nor g1883 (n_1917, n_1915, n_1908);
  nor g1886 (n_2091, n_1911, n_1915);
  nor g1887 (n_1921, n_1919, n_1908);
  nor g1890 (n_1995, n_1911, n_1919);
  nor g1891 (n_1924, n_1735, n_1923);
  nor g1894 (n_2008, n_1735, n_1926);
  nor g1900 (n_1932, n_1930, n_1923);
  nor g1903 (n_2018, n_1926, n_1930);
  nand g1906 (n_2139, n_1622, n_1936);
  nand g1907 (n_1937, n_1759, n_1934);
  nand g1908 (n_2141, n_1756, n_1937);
  nand g1911 (n_2144, n_1940, n_1941);
  nand g1914 (n_2147, n_1863, n_1943);
  nand g1915 (n_1946, n_1944, n_1934);
  nand g1916 (n_2150, n_1945, n_1946);
  nand g1917 (n_1949, n_1947, n_1934);
  nand g1918 (n_2152, n_1948, n_1949);
  nand g1919 (n_1952, n_1950, n_1934);
  nand g1920 (n_2155, n_1951, n_1952);
  nand g1921 (n_1955, n_1953, n_1934);
  nand g1922 (n_2023, n_1954, n_1955);
  nor g1923 (n_1957, n_1675, n_1956);
  nand g1932 (n_2047, n_1799, n_1959);
  nor g1933 (n_1966, n_1964, n_1956);
  nor g1938 (n_1969, n_1896, n_1956);
  nand g1947 (n_2059, n_1959, n_1972);
  nand g1952 (n_2063, n_1959, n_1977);
  nand g1957 (n_2067, n_1959, n_1982);
  nand g1962 (n_2071, n_1959, n_1987);
  nor g1963 (n_1993, n_1723, n_1992);
  nand g1972 (n_2099, n_1839, n_1995);
  nor g1973 (n_2002, n_2000, n_1992);
  nor g1978 (n_2005, n_1926, n_1992);
  nand g1987 (n_2111, n_1995, n_2008);
  nand g1992 (n_2115, n_1995, n_2013);
  nand g1997 (n_2119, n_1995, n_2018);
  nand g2000 (n_2159, n_1646, n_2025);
  nand g2001 (n_2026, n_1779, n_2023);
  nand g2002 (n_2161, n_1776, n_2026);
  nand g2005 (n_2164, n_2029, n_2030);
  nand g2008 (n_2167, n_1878, n_2032);
  nand g2009 (n_2035, n_2033, n_2023);
  nand g2010 (n_2170, n_2034, n_2035);
  nand g2011 (n_2038, n_2036, n_2023);
  nand g2012 (n_2172, n_2037, n_2038);
  nand g2013 (n_2041, n_2039, n_2023);
  nand g2014 (n_2175, n_2040, n_2041);
  nand g2015 (n_2042, n_1959, n_2023);
  nand g2016 (n_2177, n_1956, n_2042);
  nand g2019 (n_2180, n_2045, n_2046);
  nand g2022 (n_2182, n_2049, n_2050);
  nand g2025 (n_2185, n_2053, n_2054);
  nand g2028 (n_2188, n_2057, n_2058);
  nand g2031 (n_2191, n_2061, n_2062);
  nand g2034 (n_2193, n_2065, n_2066);
  nand g2037 (n_2196, n_2069, n_2070);
  nand g2040 (n_2075, n_2073, n_2074);
  nand g2043 (n_2200, n_1694, n_2077);
  nand g2044 (n_2078, n_1819, n_2075);
  nand g2045 (n_2202, n_1816, n_2078);
  nand g2048 (n_2205, n_2081, n_2082);
  nand g2051 (n_2208, n_1908, n_2084);
  nand g2052 (n_2087, n_2085, n_2075);
  nand g2053 (n_2211, n_2086, n_2087);
  nand g2054 (n_2090, n_2088, n_2075);
  nand g2055 (n_2213, n_2089, n_2090);
  nand g2056 (n_2093, n_2091, n_2075);
  nand g2057 (n_2216, n_2092, n_2093);
  nand g2058 (n_2094, n_1995, n_2075);
  nand g2059 (n_2218, n_1992, n_2094);
  nand g2062 (n_2221, n_2097, n_2098);
  nand g2065 (n_2223, n_2101, n_2102);
  nand g2068 (n_2226, n_2105, n_2106);
  nand g2071 (n_2229, n_2109, n_2110);
  nand g2074 (n_2232, n_2113, n_2114);
  nand g2077 (n_2234, n_2117, n_2118);
  nand g2080 (n_2237, n_2121, n_2122);
  xnor g2092 (Z[5], n_2130, n_2131);
  xnor g2094 (Z[6], n_2132, n_2133);
  xnor g2097 (Z[7], n_2135, n_2136);
  xnor g2099 (Z[8], n_1934, n_2137);
  xnor g2102 (Z[9], n_2139, n_2140);
  xnor g2104 (Z[10], n_2141, n_2142);
  xnor g2107 (Z[11], n_2144, n_2145);
  xnor g2110 (Z[12], n_2147, n_2148);
  xnor g2113 (Z[13], n_2150, n_2151);
  xnor g2115 (Z[14], n_2152, n_2153);
  xnor g2118 (Z[15], n_2155, n_2156);
  xnor g2120 (Z[16], n_2023, n_2157);
  xnor g2123 (Z[17], n_2159, n_2160);
  xnor g2125 (Z[18], n_2161, n_2162);
  xnor g2128 (Z[19], n_2164, n_2165);
  xnor g2131 (Z[20], n_2167, n_2168);
  xnor g2134 (Z[21], n_2170, n_2171);
  xnor g2136 (Z[22], n_2172, n_2173);
  xnor g2139 (Z[23], n_2175, n_2176);
  xnor g2141 (Z[24], n_2177, n_2178);
  xnor g2144 (Z[25], n_2180, n_2181);
  xnor g2146 (Z[26], n_2182, n_2183);
  xnor g2149 (Z[27], n_2185, n_2186);
  xnor g2152 (Z[28], n_2188, n_2189);
  xnor g2155 (Z[29], n_2191, n_2192);
  xnor g2157 (Z[30], n_2193, n_2194);
  xnor g2160 (Z[31], n_2196, n_2197);
  xnor g2162 (Z[32], n_2075, n_2198);
  xnor g2165 (Z[33], n_2200, n_2201);
  xnor g2167 (Z[34], n_2202, n_2203);
  xnor g2170 (Z[35], n_2205, n_2206);
  xnor g2173 (Z[36], n_2208, n_2209);
  xnor g2176 (Z[37], n_2211, n_2212);
  xnor g2178 (Z[38], n_2213, n_2214);
  xnor g2181 (Z[39], n_2216, n_2217);
  xnor g2183 (Z[40], n_2218, n_2219);
  xnor g2186 (Z[41], n_2221, n_2222);
  xnor g2188 (Z[42], n_2223, n_2224);
  xnor g2191 (Z[43], n_2226, n_2227);
  xnor g2194 (Z[44], n_2229, n_2230);
  xnor g2197 (Z[45], n_2232, n_2233);
  xnor g2199 (Z[46], n_2234, n_2235);
  xnor g2202 (Z[47], n_2237, n_2238);
  or g2214 (n_1044, A[1], wc);
  not gc (wc, n_171);
  or g2215 (n_1045, A[1], wc0);
  not gc0 (wc0, A[2]);
  xnor g2216 (n_1070, A[24], A[21]);
  or g2217 (n_1071, wc1, A[24]);
  not gc1 (wc1, A[21]);
  or g2218 (n_1088, A[2], wc2);
  not gc2 (wc2, A[3]);
  or g2219 (n_1089, wc3, A[2]);
  not gc3 (wc3, A[1]);
  xnor g2220 (n_1154, A[24], A[19]);
  or g2221 (n_1155, wc4, A[24]);
  not gc4 (wc4, A[19]);
  or g2222 (n_1156, wc5, A[24]);
  not gc5 (wc5, A[20]);
  xnor g2223 (n_1214, A[6], A[5]);
  or g2224 (n_1215, A[5], wc6);
  not gc6 (wc6, A[6]);
  or g2225 (n_1252, wc7, A[6]);
  not gc7 (wc7, A[5]);
  or g2226 (n_1253, A[6], wc8);
  not gc8 (wc8, A[7]);
  or g2228 (n_1355, wc9, A[10]);
  not gc9 (wc9, A[9]);
  or g2229 (n_1356, A[10], wc10);
  not gc10 (wc10, A[14]);
  or g2230 (n_1385, A[10], wc11);
  not gc11 (wc11, A[11]);
  xnor g2231 (n_537, n_1418, A[24]);
  or g2232 (n_1421, wc12, A[24]);
  not gc12 (wc12, A[16]);
  or g2234 (n_1463, wc13, A[14]);
  not gc13 (wc13, A[13]);
  or g2235 (n_1464, A[14], wc14);
  not gc14 (wc14, A[18]);
  or g2236 (n_1485, A[14], wc15);
  not gc15 (wc15, A[15]);
  xnor g2237 (n_1526, A[24], A[20]);
  or g2239 (n_1555, wc16, A[19]);
  not gc16 (wc16, A[18]);
  or g2241 (n_1583, A[21], wc17);
  not gc17 (wc17, A[22]);
  or g2243 (n_1587, A[22], wc18);
  not gc18 (wc18, A[23]);
  or g2244 (n_1588, wc19, A[22]);
  not gc19 (wc19, A[21]);
  xnor g2245 (n_1590, A[24], A[23]);
  or g2246 (n_1591, wc20, A[24]);
  not gc20 (wc20, A[23]);
  or g2247 (n_1593, wc21, A[24]);
  not gc21 (wc21, A[22]);
  xnor g2248 (n_349, n_1042, A[1]);
  xnor g2249 (n_372, n_1086, A[2]);
  xnor g2250 (n_453, n_1250, A[6]);
  xnor g2251 (n_504, n_1218, A[14]);
  xnor g2252 (n_520, n_1098, A[10]);
  nand g2253 (n_532, n_1099, n_1385);
  xnor g2254 (n_558, n_1222, A[18]);
  xnor g2255 (n_569, n_1386, A[14]);
  nand g2256 (n_578, n_944, n_1485);
  xnor g2257 (n_1542, n_560, A[18]);
  or g2258 (n_1543, A[18], wc22);
  not gc22 (wc22, n_560);
  xnor g2259 (n_605, n_1486, n_603);
  or g2260 (n_1557, A[19], wc23);
  not gc23 (wc23, n_603);
  xnor g2261 (n_76, n_1114, A[21]);
  or g2263 (n_2124, wc24, n_1609);
  not gc24 (wc24, n_1604);
  or g2264 (n_1508, A[24], wc25);
  not gc25 (wc25, n_578);
  or g2265 (n_1529, A[24], wc26);
  not gc26 (wc26, n_586);
  xnor g2266 (n_29, n_1366, n_617);
  or g2267 (n_1584, A[21], wc27);
  not gc27 (wc27, n_617);
  and g2268 (n_1744, wc28, n_1606);
  not gc28 (wc28, n_1607);
  or g2269 (n_2127, wc29, n_1605);
  not gc29 (wc29, n_1606);
  xnor g2270 (n_581, n_1506, A[24]);
  and g2271 (n_1737, wc30, n_74);
  not gc30 (wc30, A[24]);
  or g2272 (n_1738, wc31, n_74);
  not gc31 (wc31, A[24]);
  not g2273 (Z[2], n_2124);
  or g2274 (n_1216, A[5], wc32);
  not gc32 (wc32, n_433);
  xnor g2275 (n_1446, n_545, A[24]);
  or g2276 (n_1447, A[24], wc33);
  not gc33 (wc33, n_545);
  or g2277 (n_1545, A[18], wc34);
  not gc34 (wc34, n_596);
  or g2280 (n_2128, wc35, n_1615);
  not gc35 (wc35, n_1610);
  or g2281 (n_2235, wc36, n_1739);
  not gc36 (wc36, n_1736);
  or g2282 (n_1304, A[24], wc37);
  not gc37 (wc37, n_475);
  or g2283 (n_1336, A[24], wc38);
  not gc38 (wc38, n_490);
  and g2284 (n_1746, wc39, n_1612);
  not gc39 (wc39, n_1613);
  or g2285 (n_1853, n_1615, n_1744);
  or g2286 (n_1854, n_1744, wc40);
  not gc40 (wc40, n_1749);
  xor g2287 (Z[3], n_1604, n_2127);
  xor g2288 (Z[4], n_1744, n_2128);
  or g2289 (n_2131, wc41, n_1611);
  not gc41 (wc41, n_1612);
  or g2290 (n_2238, wc42, n_1737);
  not gc42 (wc42, n_1738);
  xnor g2291 (n_479, n_1302, A[24]);
  or g2292 (n_1337, A[24], wc43);
  not gc43 (wc43, n_489);
  and g2293 (n_1753, wc44, n_1618);
  not gc44 (wc44, n_1619);
  or g2294 (n_1855, wc45, n_1621);
  not gc45 (wc45, n_1749);
  or g2295 (n_2133, wc46, n_1621);
  not gc46 (wc46, n_1616);
  or g2296 (n_2136, wc47, n_1617);
  not gc47 (wc47, n_1618);
  or g2297 (n_2233, wc48, n_1731);
  not gc48 (wc48, n_1732);
  xnor g2298 (n_494, n_1334, A[24]);
  and g2299 (n_1857, wc49, n_1616);
  not gc49 (wc49, n_1747);
  and g2300 (n_1754, wc50, n_1751);
  not gc50 (wc50, n_1746);
  or g2301 (n_2137, wc51, n_1627);
  not gc51 (wc51, n_1622);
  or g2302 (n_2227, wc52, n_1725);
  not gc52 (wc52, n_1726);
  xnor g2303 (n_1194, n_419, A[24]);
  or g2304 (n_1195, A[24], wc53);
  not gc53 (wc53, n_419);
  or g2305 (n_1196, A[24], wc54);
  not gc54 (wc54, n_420);
  and g2306 (n_1846, wc55, n_1732);
  not gc55 (wc55, n_1733);
  and g2307 (n_1861, wc56, n_1753);
  not gc56 (wc56, n_1754);
  or g2308 (n_1930, wc57, n_1739);
  not gc57 (wc57, n_1849);
  or g2309 (n_1858, n_1744, n_1855);
  or g2310 (n_1862, n_1859, n_1744);
  or g2311 (n_2230, wc58, n_1735);
  not gc58 (wc58, n_1730);
  and g2312 (n_1756, wc59, n_1624);
  not gc59 (wc59, n_1625);
  or g2313 (n_2140, wc60, n_1623);
  not gc60 (wc60, n_1624);
  and g2314 (n_1836, wc61, n_1720);
  not gc61 (wc61, n_1721);
  and g2315 (n_1843, wc62, n_1726);
  not gc62 (wc62, n_1727);
  or g2316 (n_1938, wc63, n_1633);
  not gc63 (wc63, n_1759);
  or g2317 (n_2000, wc64, n_1729);
  not gc64 (wc64, n_1839);
  and g2318 (n_1931, wc65, n_1736);
  not gc65 (wc65, n_1847);
  or g2319 (n_1936, wc66, n_1627);
  not gc66 (wc66, n_1934);
  or g2320 (n_2142, wc67, n_1633);
  not gc67 (wc67, n_1628);
  or g2321 (n_2219, wc68, n_1723);
  not gc68 (wc68, n_1718);
  or g2322 (n_2222, wc69, n_1719);
  not gc69 (wc69, n_1720);
  or g2323 (n_2224, wc70, n_1729);
  not gc70 (wc70, n_1724);
  or g2324 (n_1073, A[24], wc71);
  not gc71 (wc71, n_358);
  and g2325 (n_1763, wc72, n_1630);
  not gc72 (wc72, n_1631);
  and g2326 (n_1940, wc73, n_1628);
  not gc73 (wc73, n_1757);
  and g2327 (n_1844, wc74, n_1841);
  not gc74 (wc74, n_1836);
  and g2328 (n_2013, wc75, n_1849);
  not gc75 (wc75, n_1926);
  or g2329 (n_2145, wc76, n_1629);
  not gc76 (wc76, n_1630);
  and g2330 (n_1764, wc77, n_1761);
  not gc77 (wc77, n_1756);
  and g2331 (n_2001, wc78, n_1724);
  not gc78 (wc78, n_1837);
  and g2332 (n_1923, wc79, n_1843);
  not gc79 (wc79, n_1844);
  or g2333 (n_1941, n_1938, wc80);
  not gc80 (wc80, n_1934);
  or g2334 (n_2148, wc81, n_1639);
  not gc81 (wc81, n_1634);
  or g2335 (n_2212, wc82, n_1707);
  not gc82 (wc82, n_1708);
  or g2336 (n_2217, wc83, n_1713);
  not gc83 (wc83, n_1714);
  and g2337 (n_1833, wc84, n_1714);
  not gc84 (wc84, n_1715);
  and g2338 (n_1863, wc85, n_1763);
  not gc85 (wc85, n_1764);
  and g2339 (n_1928, wc86, n_1849);
  not gc86 (wc86, n_1923);
  or g2340 (n_1943, wc87, n_1866);
  not gc87 (wc87, n_1934);
  or g2341 (n_2156, wc88, n_1641);
  not gc88 (wc88, n_1642);
  or g2342 (n_2214, wc89, n_1717);
  not gc89 (wc89, n_1712);
  and g2343 (n_1766, wc90, n_1636);
  not gc90 (wc90, n_1637);
  and g2344 (n_1773, wc91, n_1642);
  not gc91 (wc91, n_1643);
  or g2345 (n_1870, wc92, n_1645);
  not gc92 (wc92, n_1769);
  and g2346 (n_2010, wc93, n_1730);
  not gc93 (wc93, n_1924);
  and g2347 (n_2015, wc94, n_1846);
  not gc94 (wc94, n_1928);
  and g2348 (n_2020, n_1931, wc95);
  not gc95 (wc95, n_1932);
  or g2349 (n_2151, wc96, n_1635);
  not gc96 (wc96, n_1636);
  or g2350 (n_2153, wc97, n_1645);
  not gc97 (wc97, n_1640);
  or g2351 (n_2157, wc98, n_1651);
  not gc98 (wc98, n_1646);
  and g2352 (n_1776, wc99, n_1648);
  not gc99 (wc99, n_1649);
  and g2353 (n_1774, wc100, n_1771);
  not gc100 (wc100, n_1766);
  and g2354 (n_1945, wc101, n_1634);
  not gc101 (wc101, n_1864);
  and g2355 (n_1868, wc102, n_1769);
  not gc102 (wc102, n_1863);
  and g2356 (n_1947, wc103, n_1769);
  not gc103 (wc103, n_1866);
  or g2357 (n_2160, wc104, n_1647);
  not gc104 (wc104, n_1648);
  and g2358 (n_1783, wc105, n_1654);
  not gc105 (wc105, n_1655);
  and g2359 (n_1826, wc106, n_1708);
  not gc106 (wc106, n_1709);
  and g2360 (n_1871, wc107, n_1640);
  not gc107 (wc107, n_1767);
  and g2361 (n_1875, wc108, n_1773);
  not gc108 (wc108, n_1774);
  or g2362 (n_2027, wc109, n_1657);
  not gc109 (wc109, n_1779);
  or g2363 (n_1915, wc110, n_1717);
  not gc110 (wc110, n_1829);
  and g2364 (n_1948, wc111, n_1766);
  not gc111 (wc111, n_1868);
  or g2365 (n_2162, wc112, n_1657);
  not gc112 (wc112, n_1652);
  or g2366 (n_2165, wc113, n_1653);
  not gc113 (wc113, n_1654);
  or g2367 (n_2168, wc114, n_1663);
  not gc114 (wc114, n_1658);
  or g2368 (n_2206, wc115, n_1701);
  not gc115 (wc115, n_1702);
  or g2369 (n_2209, wc116, n_1711);
  not gc116 (wc116, n_1706);
  and g2370 (n_1786, wc117, n_1660);
  not gc117 (wc117, n_1661);
  and g2371 (n_2029, wc118, n_1652);
  not gc118 (wc118, n_1777);
  and g2372 (n_1784, wc119, n_1781);
  not gc119 (wc119, n_1776);
  and g2373 (n_1834, wc120, n_1831);
  not gc120 (wc120, n_1826);
  or g2374 (n_2171, wc121, n_1659);
  not gc121 (wc121, n_1660);
  and g2375 (n_1793, wc122, n_1666);
  not gc122 (wc122, n_1667);
  and g2376 (n_1816, wc123, n_1696);
  not gc123 (wc123, n_1697);
  and g2377 (n_1823, wc124, n_1702);
  not gc124 (wc124, n_1703);
  and g2378 (n_1878, wc125, n_1783);
  not gc125 (wc125, n_1784);
  or g2379 (n_1885, wc126, n_1669);
  not gc126 (wc126, n_1789);
  or g2380 (n_2079, wc127, n_1705);
  not gc127 (wc127, n_1819);
  and g2381 (n_1916, wc128, n_1712);
  not gc128 (wc128, n_1827);
  and g2382 (n_1920, wc129, n_1833);
  not gc129 (wc129, n_1834);
  and g2383 (n_1951, n_1871, wc130);
  not gc130 (wc130, n_1872);
  and g2384 (n_1954, n_1875, wc131);
  not gc131 (wc131, n_1876);
  and g2385 (n_2036, wc132, n_1789);
  not gc132 (wc132, n_1881);
  or g2386 (n_2173, wc133, n_1669);
  not gc133 (wc133, n_1664);
  or g2387 (n_2176, wc134, n_1665);
  not gc134 (wc134, n_1666);
  or g2388 (n_2197, wc135, n_1689);
  not gc135 (wc135, n_1690);
  or g2389 (n_2198, wc136, n_1699);
  not gc136 (wc136, n_1694);
  or g2390 (n_2201, wc137, n_1695);
  not gc137 (wc137, n_1696);
  or g2391 (n_2203, wc138, n_1705);
  not gc138 (wc138, n_1700);
  and g2392 (n_1813, wc139, n_1690);
  not gc139 (wc139, n_1691);
  and g2393 (n_1886, wc140, n_1664);
  not gc140 (wc140, n_1787);
  and g2394 (n_1794, wc141, n_1791);
  not gc141 (wc141, n_1786);
  and g2395 (n_1824, wc142, n_1821);
  not gc142 (wc142, n_1816);
  and g2396 (n_1883, wc143, n_1789);
  not gc143 (wc143, n_1878);
  and g2397 (n_2088, wc144, n_1829);
  not gc144 (wc144, n_1911);
  or g2398 (n_2178, wc145, n_1675);
  not gc145 (wc145, n_1670);
  or g2399 (n_2183, wc146, n_1681);
  not gc146 (wc146, n_1676);
  or g2400 (n_2194, wc147, n_1693);
  not gc147 (wc147, n_1688);
  and g2401 (n_1796, wc148, n_1672);
  not gc148 (wc148, n_1673);
  and g2402 (n_1803, wc149, n_1678);
  not gc149 (wc149, n_1679);
  and g2403 (n_1806, wc150, n_1684);
  not gc150 (wc150, n_1685);
  and g2404 (n_1890, wc151, n_1793);
  not gc151 (wc151, n_1794);
  or g2405 (n_1964, wc152, n_1681);
  not gc152 (wc152, n_1799);
  or g2406 (n_1900, wc153, n_1693);
  not gc153 (wc153, n_1809);
  and g2407 (n_2081, wc154, n_1700);
  not gc154 (wc154, n_1817);
  and g2408 (n_1908, wc155, n_1823);
  not gc155 (wc155, n_1824);
  and g2409 (n_2034, wc156, n_1658);
  not gc156 (wc156, n_1879);
  and g2410 (n_2037, wc157, n_1786);
  not gc157 (wc157, n_1883);
  or g2411 (n_2043, wc158, n_1675);
  not gc158 (wc158, n_1959);
  or g2412 (n_2095, wc159, n_1723);
  not gc159 (wc159, n_1995);
  or g2413 (n_2103, n_2000, wc160);
  not gc160 (wc160, n_1995);
  or g2414 (n_2107, wc161, n_1926);
  not gc161 (wc161, n_1995);
  or g2415 (n_2025, wc162, n_1651);
  not gc162 (wc162, n_2023);
  or g2416 (n_2030, n_2027, wc163);
  not gc163 (wc163, n_2023);
  or g2417 (n_2032, wc164, n_1881);
  not gc164 (wc164, n_2023);
  or g2418 (n_2181, wc165, n_1671);
  not gc165 (wc165, n_1672);
  or g2419 (n_2186, wc166, n_1677);
  not gc166 (wc166, n_1678);
  or g2420 (n_2189, wc167, n_1687);
  not gc167 (wc167, n_1682);
  or g2421 (n_2192, wc168, n_1683);
  not gc168 (wc168, n_1684);
  and g2422 (n_1804, wc169, n_1801);
  not gc169 (wc169, n_1796);
  and g2423 (n_1814, wc170, n_1811);
  not gc170 (wc170, n_1806);
  and g2424 (n_2040, n_1886, wc171);
  not gc171 (wc171, n_1887);
  and g2425 (n_1977, wc172, n_1809);
  not gc172 (wc172, n_1896);
  and g2426 (n_1913, wc173, n_1829);
  not gc173 (wc173, n_1908);
  and g2427 (n_1965, wc174, n_1676);
  not gc174 (wc174, n_1797);
  and g2428 (n_1893, wc175, n_1803);
  not gc175 (wc175, n_1804);
  and g2429 (n_1901, wc176, n_1688);
  not gc176 (wc176, n_1807);
  and g2430 (n_1905, wc177, n_1813);
  not gc177 (wc177, n_1814);
  and g2431 (n_1956, n_1890, wc178);
  not gc178 (wc178, n_1891);
  and g2432 (n_2086, wc179, n_1706);
  not gc179 (wc179, n_1909);
  and g2433 (n_2089, wc180, n_1826);
  not gc180 (wc180, n_1913);
  and g2434 (n_2092, n_1916, wc181);
  not gc181 (wc181, n_1917);
  and g2435 (n_1992, n_1920, wc182);
  not gc182 (wc182, n_1921);
  or g2436 (n_2051, n_1964, wc183);
  not gc183 (wc183, n_1959);
  or g2437 (n_2055, wc184, n_1896);
  not gc184 (wc184, n_1959);
  or g2438 (n_2046, n_2043, wc185);
  not gc185 (wc185, n_2023);
  or g2439 (n_2050, n_2047, wc186);
  not gc186 (wc186, n_2023);
  and g2440 (n_1898, wc187, n_1809);
  not gc187 (wc187, n_1893);
  and g2441 (n_1962, wc188, n_1799);
  not gc188 (wc188, n_1956);
  and g2442 (n_1975, wc189, n_1972);
  not gc189 (wc189, n_1956);
  and g2443 (n_1980, wc190, n_1977);
  not gc190 (wc190, n_1956);
  and g2444 (n_1985, wc191, n_1982);
  not gc191 (wc191, n_1956);
  and g2445 (n_1990, wc192, n_1987);
  not gc192 (wc192, n_1956);
  and g2446 (n_1998, wc193, n_1839);
  not gc193 (wc193, n_1992);
  and g2447 (n_2011, wc194, n_2008);
  not gc194 (wc194, n_1992);
  and g2448 (n_2016, wc195, n_2013);
  not gc195 (wc195, n_1992);
  and g2449 (n_2021, wc196, n_2018);
  not gc196 (wc196, n_1992);
  and g2450 (n_1974, wc197, n_1682);
  not gc197 (wc197, n_1894);
  and g2451 (n_1979, wc198, n_1806);
  not gc198 (wc198, n_1898);
  and g2452 (n_1984, n_1901, wc199);
  not gc199 (wc199, n_1902);
  and g2453 (n_1989, n_1905, wc200);
  not gc200 (wc200, n_1906);
  and g2454 (n_2045, wc201, n_1670);
  not gc201 (wc201, n_1957);
  and g2455 (n_2049, wc202, n_1796);
  not gc202 (wc202, n_1962);
  and g2456 (n_2053, n_1965, wc203);
  not gc203 (wc203, n_1966);
  and g2457 (n_2057, n_1893, wc204);
  not gc204 (wc204, n_1969);
  and g2458 (n_2097, wc205, n_1718);
  not gc205 (wc205, n_1993);
  and g2459 (n_2101, wc206, n_1836);
  not gc206 (wc206, n_1998);
  and g2460 (n_2105, n_2001, wc207);
  not gc207 (wc207, n_2002);
  and g2461 (n_2109, n_1923, wc208);
  not gc208 (wc208, n_2005);
  and g2462 (n_2113, wc209, n_2010);
  not gc209 (wc209, n_2011);
  and g2463 (n_2117, wc210, n_2015);
  not gc210 (wc210, n_2016);
  and g2464 (n_2121, wc211, n_2020);
  not gc211 (wc211, n_2021);
  or g2465 (n_2054, n_2051, wc212);
  not gc212 (wc212, n_2023);
  or g2466 (n_2058, n_2055, wc213);
  not gc213 (wc213, n_2023);
  or g2467 (n_2062, n_2059, wc214);
  not gc214 (wc214, n_2023);
  or g2468 (n_2066, n_2063, wc215);
  not gc215 (wc215, n_2023);
  or g2469 (n_2070, n_2067, wc216);
  not gc216 (wc216, n_2023);
  or g2470 (n_2074, n_2071, wc217);
  not gc217 (wc217, n_2023);
  and g2471 (n_2061, n_1974, wc218);
  not gc218 (wc218, n_1975);
  and g2472 (n_2065, n_1979, wc219);
  not gc219 (wc219, n_1980);
  and g2473 (n_2069, n_1984, wc220);
  not gc220 (wc220, n_1985);
  and g2474 (n_2073, n_1989, wc221);
  not gc221 (wc221, n_1990);
  or g2475 (n_2077, wc222, n_1699);
  not gc222 (wc222, n_2075);
  or g2476 (n_2082, n_2079, wc223);
  not gc223 (wc223, n_2075);
  or g2477 (n_2084, wc224, n_1911);
  not gc224 (wc224, n_2075);
  or g2478 (n_2098, n_2095, wc225);
  not gc225 (wc225, n_2075);
  or g2479 (n_2102, wc226, n_2099);
  not gc226 (wc226, n_2075);
  or g2480 (n_2106, n_2103, wc227);
  not gc227 (wc227, n_2075);
  or g2481 (n_2110, n_2107, wc228);
  not gc228 (wc228, n_2075);
  or g2482 (n_2114, wc229, n_2111);
  not gc229 (wc229, n_2075);
  or g2483 (n_2118, wc230, n_2115);
  not gc230 (wc230, n_2075);
  or g2484 (n_2122, wc231, n_2119);
  not gc231 (wc231, n_2075);
endmodule

module mult_signed_const_4151_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_4151_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_4418_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_171, n_172, n_174, n_178, n_179;
  wire n_181, n_182, n_183, n_185, n_186, n_187, n_188, n_193;
  wire n_194, n_195, n_199, n_200, n_201, n_202, n_203, n_206;
  wire n_207, n_208, n_209, n_210, n_211, n_213, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_223, n_224, n_225, n_226;
  wire n_227, n_232, n_233, n_234, n_235, n_236, n_237, n_238;
  wire n_239, n_243, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_255, n_256, n_257, n_258, n_259, n_260, n_261;
  wire n_262, n_263, n_264, n_266, n_268, n_269, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_278, n_283;
  wire n_284, n_286, n_287, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_294, n_298, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_314, n_315;
  wire n_317, n_318, n_319, n_320, n_321, n_322, n_323, n_324;
  wire n_325, n_326, n_327, n_333, n_334, n_335, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_351, n_352, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_391, n_393, n_394;
  wire n_395, n_396, n_397, n_399, n_400, n_401, n_402, n_403;
  wire n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411;
  wire n_412, n_413, n_414, n_415, n_416, n_418, n_419, n_420;
  wire n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_489, n_490, n_491;
  wire n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500;
  wire n_501, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_520, n_521, n_522, n_523;
  wire n_524, n_525, n_526, n_527, n_528, n_529, n_530, n_531;
  wire n_533, n_534, n_535, n_536, n_537, n_538, n_539, n_540;
  wire n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548;
  wire n_549, n_550, n_551, n_552, n_553, n_554, n_555, n_558;
  wire n_559, n_560, n_561, n_562, n_563, n_564, n_565, n_566;
  wire n_570, n_572, n_573, n_574, n_575, n_576, n_577, n_580;
  wire n_581, n_583, n_584, n_585, n_586, n_587, n_588, n_590;
  wire n_591, n_592, n_593, n_596, n_597, n_598, n_599, n_600;
  wire n_604, n_605, n_606, n_607, n_609, n_610, n_611, n_612;
  wire n_613, n_614, n_615, n_618, n_623, n_624, n_625, n_626;
  wire n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634;
  wire n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642;
  wire n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_654;
  wire n_657, n_658, n_659, n_660, n_661, n_662, n_663, n_664;
  wire n_665, n_666, n_669, n_670, n_671, n_672, n_673, n_674;
  wire n_675, n_676, n_677, n_678, n_683, n_684, n_685, n_687;
  wire n_688, n_689, n_690, n_691, n_692, n_693, n_694, n_699;
  wire n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710;
  wire n_711, n_712, n_713, n_714, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_752, n_753, n_754, n_761, n_762, n_763, n_764;
  wire n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772;
  wire n_773, n_774, n_775, n_776, n_777, n_778, n_787, n_791;
  wire n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799;
  wire n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_813;
  wire n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821;
  wire n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829;
  wire n_830, n_831, n_832, n_833, n_834, n_841, n_843, n_844;
  wire n_845, n_846, n_847, n_848, n_849, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860;
  wire n_861, n_862, n_863, n_869, n_870, n_871, n_873, n_874;
  wire n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882;
  wire n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890;
  wire n_891, n_892, n_893, n_894, n_909, n_910, n_911, n_912;
  wire n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920;
  wire n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928;
  wire n_929, n_930, n_938, n_939, n_940, n_942, n_943, n_945;
  wire n_946, n_947, n_948, n_949, n_950, n_951, n_952, n_953;
  wire n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961;
  wire n_962, n_963, n_964, n_965, n_966, n_977, n_978, n_979;
  wire n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1007;
  wire n_1011, n_1012, n_1014, n_1015, n_1016, n_1018, n_1019, n_1020;
  wire n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028;
  wire n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036;
  wire n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1045;
  wire n_1046, n_1049, n_1050, n_1051, n_1052, n_1054, n_1057, n_1058;
  wire n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066;
  wire n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074;
  wire n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082;
  wire n_1083, n_1084, n_1085, n_1086, n_1090, n_1091, n_1092, n_1093;
  wire n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102;
  wire n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110;
  wire n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118;
  wire n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126;
  wire n_1127, n_1128, n_1129, n_1130, n_1133, n_1134, n_1135, n_1136;
  wire n_1137, n_1138, n_1143, n_1145, n_1147, n_1148, n_1149, n_1150;
  wire n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158;
  wire n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166;
  wire n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174;
  wire n_1175, n_1176, n_1177, n_1178, n_1179, n_1182, n_1183, n_1184;
  wire n_1187, n_1188, n_1189, n_1190, n_1191, n_1193, n_1194, n_1195;
  wire n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203;
  wire n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211;
  wire n_1212, n_1213, n_1214, n_1216, n_1217, n_1218, n_1219, n_1225;
  wire n_1226, n_1227, n_1228, n_1229, n_1231, n_1232, n_1233, n_1234;
  wire n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242;
  wire n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250;
  wire n_1253, n_1255, n_1256, n_1257, n_1259, n_1260, n_1263, n_1264;
  wire n_1265, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273;
  wire n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281;
  wire n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1290, n_1291;
  wire n_1292, n_1293, n_1294, n_1295, n_1297, n_1298, n_1299, n_1301;
  wire n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309;
  wire n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317;
  wire n_1318, n_1319, n_1320, n_1321, n_1322, n_1331, n_1332, n_1333;
  wire n_1334, n_1335, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342;
  wire n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350;
  wire n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1359, n_1360;
  wire n_1361, n_1363, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370;
  wire n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378;
  wire n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1387, n_1388;
  wire n_1389, n_1391, n_1392, n_1394, n_1395, n_1396, n_1397, n_1398;
  wire n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406;
  wire n_1407, n_1408, n_1409, n_1410, n_1416, n_1417, n_1419, n_1422;
  wire n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430;
  wire n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438;
  wire n_1439, n_1442, n_1443, n_1446, n_1447, n_1448, n_1449, n_1450;
  wire n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458;
  wire n_1459, n_1460, n_1461, n_1462, n_1463, n_1469, n_1470, n_1471;
  wire n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479;
  wire n_1480, n_1481, n_1482, n_1487, n_1488, n_1489, n_1491, n_1492;
  wire n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500;
  wire n_1501, n_1502, n_1503, n_1506, n_1511, n_1512, n_1513, n_1514;
  wire n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522;
  wire n_1523, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535;
  wire n_1536, n_1537, n_1538, n_1539, n_1540, n_1542, n_1543, n_1544;
  wire n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552;
  wire n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561;
  wire n_1562, n_1563, n_1565, n_1567, n_1568, n_1569, n_1570, n_1571;
  wire n_1572, n_1573, n_1574, n_1579, n_1580, n_1581, n_1582, n_1584;
  wire n_1585, n_1586, n_1587, n_1588, n_1589, n_1594, n_1605, n_1606;
  wire n_1607, n_1608, n_1610, n_1611, n_1612, n_1613, n_1614, n_1616;
  wire n_1617, n_1618, n_1619, n_1620, n_1622, n_1623, n_1624, n_1625;
  wire n_1626, n_1628, n_1629, n_1630, n_1631, n_1632, n_1634, n_1635;
  wire n_1636, n_1637, n_1638, n_1640, n_1641, n_1642, n_1643, n_1644;
  wire n_1646, n_1647, n_1648, n_1649, n_1650, n_1652, n_1653, n_1654;
  wire n_1655, n_1656, n_1658, n_1659, n_1660, n_1661, n_1662, n_1664;
  wire n_1665, n_1666, n_1667, n_1668, n_1670, n_1671, n_1672, n_1673;
  wire n_1674, n_1676, n_1677, n_1678, n_1679, n_1680, n_1682, n_1683;
  wire n_1684, n_1685, n_1686, n_1688, n_1689, n_1690, n_1691, n_1692;
  wire n_1694, n_1695, n_1696, n_1697, n_1698, n_1700, n_1701, n_1702;
  wire n_1703, n_1704, n_1706, n_1707, n_1708, n_1709, n_1710, n_1712;
  wire n_1713, n_1714, n_1715, n_1716, n_1718, n_1719, n_1720, n_1721;
  wire n_1722, n_1724, n_1725, n_1726, n_1727, n_1728, n_1730, n_1731;
  wire n_1732, n_1733, n_1734, n_1736, n_1737, n_1738, n_1739, n_1740;
  wire n_1745, n_1747, n_1748, n_1750, n_1752, n_1754, n_1755, n_1757;
  wire n_1758, n_1760, n_1762, n_1764, n_1765, n_1767, n_1768, n_1770;
  wire n_1772, n_1774, n_1775, n_1777, n_1778, n_1780, n_1782, n_1784;
  wire n_1785, n_1787, n_1788, n_1790, n_1792, n_1794, n_1795, n_1797;
  wire n_1798, n_1800, n_1802, n_1804, n_1805, n_1807, n_1808, n_1810;
  wire n_1812, n_1814, n_1815, n_1817, n_1818, n_1820, n_1822, n_1824;
  wire n_1825, n_1827, n_1828, n_1830, n_1832, n_1834, n_1835, n_1837;
  wire n_1838, n_1840, n_1842, n_1844, n_1845, n_1847, n_1848, n_1850;
  wire n_1854, n_1855, n_1856, n_1858, n_1859, n_1860, n_1862, n_1863;
  wire n_1864, n_1865, n_1867, n_1869, n_1871, n_1872, n_1873, n_1875;
  wire n_1876, n_1877, n_1879, n_1880, n_1882, n_1884, n_1886, n_1887;
  wire n_1888, n_1890, n_1891, n_1892, n_1894, n_1895, n_1897, n_1899;
  wire n_1901, n_1902, n_1903, n_1905, n_1906, n_1907, n_1909, n_1910;
  wire n_1912, n_1914, n_1916, n_1917, n_1918, n_1920, n_1921, n_1922;
  wire n_1924, n_1925, n_1927, n_1929, n_1931, n_1932, n_1933, n_1935;
  wire n_1937, n_1938, n_1939, n_1941, n_1942, n_1944, n_1945, n_1946;
  wire n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954;
  wire n_1955, n_1956, n_1957, n_1958, n_1960, n_1963, n_1965, n_1966;
  wire n_1967, n_1970, n_1973, n_1975, n_1976, n_1978, n_1980, n_1981;
  wire n_1983, n_1985, n_1986, n_1988, n_1990, n_1991, n_1993, n_1994;
  wire n_1996, n_1999, n_2001, n_2002, n_2003, n_2006, n_2009, n_2011;
  wire n_2012, n_2014, n_2016, n_2017, n_2019, n_2021, n_2022, n_2024;
  wire n_2026, n_2027, n_2028, n_2030, n_2031, n_2033, n_2034, n_2035;
  wire n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043;
  wire n_2044, n_2046, n_2047, n_2048, n_2050, n_2051, n_2052, n_2054;
  wire n_2055, n_2056, n_2058, n_2059, n_2060, n_2062, n_2063, n_2064;
  wire n_2066, n_2067, n_2068, n_2070, n_2071, n_2072, n_2074, n_2075;
  wire n_2076, n_2078, n_2079, n_2080, n_2082, n_2083, n_2085, n_2086;
  wire n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094;
  wire n_2095, n_2096, n_2098, n_2099, n_2100, n_2102, n_2103, n_2104;
  wire n_2106, n_2107, n_2108, n_2110, n_2111, n_2112, n_2114, n_2115;
  wire n_2116, n_2118, n_2119, n_2120, n_2122, n_2123, n_2125, n_2128;
  wire n_2129, n_2131, n_2132, n_2133, n_2134, n_2136, n_2137, n_2138;
  wire n_2140, n_2141, n_2142, n_2143, n_2145, n_2146, n_2148, n_2149;
  wire n_2151, n_2152, n_2153, n_2154, n_2156, n_2157, n_2158, n_2160;
  wire n_2161, n_2162, n_2163, n_2165, n_2166, n_2168, n_2169, n_2171;
  wire n_2172, n_2173, n_2174, n_2176, n_2177, n_2178, n_2179, n_2181;
  wire n_2182, n_2183, n_2184, n_2186, n_2187, n_2189, n_2190, n_2192;
  wire n_2193, n_2194, n_2195, n_2197, n_2198, n_2199, n_2201, n_2202;
  wire n_2203, n_2204, n_2206, n_2207, n_2209, n_2210, n_2212, n_2213;
  wire n_2214, n_2215, n_2217, n_2218, n_2219, n_2220, n_2222, n_2223;
  wire n_2224, n_2225, n_2227, n_2228, n_2230, n_2231, n_2233, n_2234;
  wire n_2235, n_2236, n_2238, n_2239;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_118, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_623, A[2], A[1]);
  xor g270 (n_117, n_623, n_171);
  nand g3 (n_624, A[2], A[1]);
  nand g271 (n_625, n_171, A[1]);
  nand g272 (n_626, A[2], n_171);
  nand g273 (n_68, n_624, n_625, n_626);
  xor g274 (n_627, A[2], A[3]);
  xor g275 (n_116, n_627, A[5]);
  nand g276 (n_628, A[2], A[3]);
  nand g4 (n_629, A[5], A[3]);
  nand g277 (n_630, A[2], A[5]);
  nand g278 (n_67, n_628, n_629, n_630);
  xor g279 (n_172, A[0], A[3]);
  and g280 (n_174, A[0], A[3]);
  xor g281 (n_631, A[4], n_172);
  xor g282 (n_115, n_631, A[6]);
  nand g283 (n_632, A[4], n_172);
  nand g284 (n_633, A[6], n_172);
  nand g5 (n_634, A[4], A[6]);
  nand g6 (n_66, n_632, n_633, n_634);
  xor g287 (n_635, n_118, n_174);
  xor g288 (n_69, n_635, A[4]);
  nand g289 (n_636, n_118, n_174);
  nand g290 (n_637, A[4], n_174);
  nand g291 (n_638, n_118, A[4]);
  nand g292 (n_178, n_636, n_637, n_638);
  xor g293 (n_639, A[5], A[7]);
  xor g294 (n_114, n_639, n_69);
  nand g295 (n_640, A[5], A[7]);
  nand g296 (n_641, n_69, A[7]);
  nand g297 (n_642, A[5], n_69);
  nand g298 (n_65, n_640, n_641, n_642);
  xor g305 (n_647, A[5], n_117);
  xor g306 (n_179, n_647, A[6]);
  nand g307 (n_648, A[5], n_117);
  nand g308 (n_649, A[6], n_117);
  nand g309 (n_650, A[5], A[6]);
  nand g310 (n_181, n_648, n_649, n_650);
  xor g311 (n_651, n_178, A[8]);
  xor g312 (n_113, n_651, n_179);
  nand g313 (n_652, n_178, A[8]);
  nand g314 (n_653, n_179, A[8]);
  nand g315 (n_654, n_178, n_179);
  nand g316 (n_64, n_652, n_653, n_654);
  xor g318 (n_182, n_627, A[6]);
  nand g320 (n_657, A[6], A[3]);
  nand g321 (n_658, A[2], A[6]);
  nand g322 (n_185, n_628, n_657, n_658);
  xor g323 (n_659, n_68, A[7]);
  xor g324 (n_183, n_659, A[9]);
  nand g325 (n_660, n_68, A[7]);
  nand g326 (n_661, A[9], A[7]);
  nand g327 (n_662, n_68, A[9]);
  nand g328 (n_187, n_660, n_661, n_662);
  xor g329 (n_663, n_181, n_182);
  xor g330 (n_112, n_663, n_183);
  nand g331 (n_664, n_181, n_182);
  nand g332 (n_665, n_183, n_182);
  nand g333 (n_666, n_181, n_183);
  nand g334 (n_63, n_664, n_665, n_666);
  xor g338 (n_186, n_631, A[7]);
  nand g340 (n_669, A[7], n_172);
  nand g341 (n_670, A[4], A[7]);
  nand g342 (n_71, n_632, n_669, n_670);
  xor g343 (n_671, A[8], A[10]);
  xor g344 (n_188, n_671, n_185);
  nand g345 (n_672, A[8], A[10]);
  nand g346 (n_673, n_185, A[10]);
  nand g347 (n_674, A[8], n_185);
  nand g348 (n_193, n_672, n_673, n_674);
  xor g349 (n_675, n_186, n_187);
  xor g350 (n_111, n_675, n_188);
  nand g351 (n_676, n_186, n_187);
  nand g352 (n_677, n_188, n_187);
  nand g353 (n_678, n_186, n_188);
  nand g354 (n_62, n_676, n_677, n_678);
  xor g363 (n_683, A[5], A[9]);
  xor g364 (n_194, n_683, n_69);
  nand g365 (n_684, A[5], A[9]);
  nand g366 (n_685, n_69, A[9]);
  nand g368 (n_200, n_684, n_685, n_642);
  xor g369 (n_687, A[11], A[8]);
  xor g370 (n_195, n_687, n_71);
  nand g371 (n_688, A[11], A[8]);
  nand g372 (n_689, n_71, A[8]);
  nand g373 (n_690, A[11], n_71);
  nand g374 (n_202, n_688, n_689, n_690);
  xor g375 (n_691, n_193, n_194);
  xor g376 (n_110, n_691, n_195);
  nand g377 (n_692, n_193, n_194);
  nand g378 (n_693, n_195, n_194);
  nand g379 (n_694, n_193, n_195);
  nand g380 (n_61, n_692, n_693, n_694);
  xor g387 (n_699, A[5], A[6]);
  xor g388 (n_199, n_699, n_117);
  xor g393 (n_703, n_178, A[10]);
  xor g394 (n_201, n_703, A[9]);
  nand g395 (n_704, n_178, A[10]);
  nand g396 (n_705, A[9], A[10]);
  nand g397 (n_706, n_178, A[9]);
  nand g398 (n_208, n_704, n_705, n_706);
  xor g399 (n_707, A[12], n_199);
  xor g400 (n_203, n_707, n_200);
  nand g401 (n_708, A[12], n_199);
  nand g402 (n_709, n_200, n_199);
  nand g403 (n_710, A[12], n_200);
  nand g404 (n_210, n_708, n_709, n_710);
  xor g405 (n_711, n_201, n_202);
  xor g406 (n_109, n_711, n_203);
  nand g407 (n_712, n_201, n_202);
  nand g408 (n_713, n_203, n_202);
  nand g409 (n_714, n_201, n_203);
  nand g410 (n_60, n_712, n_713, n_714);
  xor g412 (n_206, n_627, n_68);
  nand g414 (n_717, n_68, A[3]);
  nand g415 (n_718, A[2], n_68);
  nand g416 (n_213, n_628, n_717, n_718);
  xor g417 (n_719, A[6], A[7]);
  xor g418 (n_207, n_719, A[11]);
  nand g419 (n_720, A[6], A[7]);
  nand g420 (n_721, A[11], A[7]);
  nand g421 (n_722, A[6], A[11]);
  nand g422 (n_215, n_720, n_721, n_722);
  xor g423 (n_723, A[10], n_181);
  xor g424 (n_209, n_723, A[13]);
  nand g425 (n_724, A[10], n_181);
  nand g426 (n_725, A[13], n_181);
  nand g427 (n_726, A[10], A[13]);
  nand g428 (n_216, n_724, n_725, n_726);
  xor g429 (n_727, n_206, n_207);
  xor g430 (n_211, n_727, n_208);
  nand g431 (n_728, n_206, n_207);
  nand g432 (n_729, n_208, n_207);
  nand g433 (n_730, n_206, n_208);
  nand g434 (n_219, n_728, n_729, n_730);
  xor g435 (n_731, n_209, n_210);
  xor g436 (n_108, n_731, n_211);
  nand g437 (n_732, n_209, n_210);
  nand g438 (n_733, n_211, n_210);
  nand g439 (n_734, n_209, n_211);
  nand g440 (n_59, n_732, n_733, n_734);
  xor g450 (n_217, n_687, A[12]);
  nand g452 (n_741, A[12], A[8]);
  nand g453 (n_742, A[11], A[12]);
  nand g454 (n_72, n_688, n_741, n_742);
  xor g455 (n_743, n_213, A[14]);
  xor g456 (n_218, n_743, n_186);
  nand g457 (n_744, n_213, A[14]);
  nand g458 (n_745, n_186, A[14]);
  nand g459 (n_746, n_213, n_186);
  nand g460 (n_224, n_744, n_745, n_746);
  xor g461 (n_747, n_215, n_216);
  xor g462 (n_220, n_747, n_217);
  nand g463 (n_748, n_215, n_216);
  nand g464 (n_749, n_217, n_216);
  nand g465 (n_750, n_215, n_217);
  nand g466 (n_225, n_748, n_749, n_750);
  xor g467 (n_751, n_218, n_219);
  xor g468 (n_107, n_751, n_220);
  nand g469 (n_752, n_218, n_219);
  nand g470 (n_753, n_220, n_219);
  nand g471 (n_754, n_218, n_220);
  nand g472 (n_58, n_752, n_753, n_754);
  xor g482 (n_73, n_683, A[8]);
  nand g484 (n_761, A[8], A[9]);
  nand g485 (n_762, A[5], A[8]);
  nand g486 (n_232, n_684, n_761, n_762);
  xor g487 (n_763, n_69, A[13]);
  xor g488 (n_223, n_763, A[15]);
  nand g489 (n_764, n_69, A[13]);
  nand g490 (n_765, A[15], A[13]);
  nand g491 (n_766, n_69, A[15]);
  nand g492 (n_233, n_764, n_765, n_766);
  xor g493 (n_767, A[12], n_71);
  xor g494 (n_226, n_767, n_72);
  nand g495 (n_768, A[12], n_71);
  nand g496 (n_769, n_72, n_71);
  nand g497 (n_770, A[12], n_72);
  nand g498 (n_236, n_768, n_769, n_770);
  xor g499 (n_771, n_73, n_223);
  xor g500 (n_227, n_771, n_224);
  nand g501 (n_772, n_73, n_223);
  nand g502 (n_773, n_224, n_223);
  nand g503 (n_774, n_73, n_224);
  nand g504 (n_238, n_772, n_773, n_774);
  xor g505 (n_775, n_225, n_226);
  xor g506 (n_106, n_775, n_227);
  nand g507 (n_776, n_225, n_226);
  nand g508 (n_777, n_227, n_226);
  nand g509 (n_778, n_225, n_227);
  nand g510 (n_57, n_776, n_777, n_778);
  xor g523 (n_787, n_178, A[9]);
  xor g524 (n_234, n_787, A[10]);
  xor g529 (n_791, A[14], A[13]);
  xor g530 (n_235, n_791, A[16]);
  nand g531 (n_792, A[14], A[13]);
  nand g532 (n_793, A[16], A[13]);
  nand g533 (n_794, A[14], A[16]);
  nand g534 (n_245, n_792, n_793, n_794);
  xor g535 (n_795, n_199, n_232);
  xor g536 (n_237, n_795, n_233);
  nand g537 (n_796, n_199, n_232);
  nand g538 (n_797, n_233, n_232);
  nand g539 (n_798, n_199, n_233);
  nand g540 (n_248, n_796, n_797, n_798);
  xor g541 (n_799, n_234, n_235);
  xor g542 (n_239, n_799, n_236);
  nand g543 (n_800, n_234, n_235);
  nand g544 (n_801, n_236, n_235);
  nand g545 (n_802, n_234, n_236);
  nand g546 (n_251, n_800, n_801, n_802);
  xor g547 (n_803, n_237, n_238);
  xor g548 (n_105, n_803, n_239);
  nand g549 (n_804, n_237, n_238);
  nand g550 (n_805, n_239, n_238);
  nand g551 (n_806, n_237, n_239);
  nand g552 (n_56, n_804, n_805, n_806);
  xor g560 (n_243, n_659, A[10]);
  nand g562 (n_813, A[10], A[7]);
  nand g563 (n_814, n_68, A[10]);
  nand g564 (n_255, n_660, n_813, n_814);
  xor g565 (n_815, A[11], A[15]);
  xor g566 (n_247, n_815, n_181);
  nand g567 (n_816, A[11], A[15]);
  nand g568 (n_817, n_181, A[15]);
  nand g569 (n_818, A[11], n_181);
  nand g570 (n_257, n_816, n_817, n_818);
  xor g571 (n_819, A[14], n_182);
  xor g572 (n_246, n_819, A[17]);
  nand g573 (n_820, A[14], n_182);
  nand g574 (n_821, A[17], n_182);
  nand g575 (n_822, A[14], A[17]);
  nand g576 (n_258, n_820, n_821, n_822);
  xor g577 (n_823, n_243, n_208);
  xor g578 (n_249, n_823, n_245);
  nand g579 (n_824, n_243, n_208);
  nand g580 (n_825, n_245, n_208);
  nand g581 (n_826, n_243, n_245);
  nand g582 (n_261, n_824, n_825, n_826);
  xor g583 (n_827, n_246, n_247);
  xor g584 (n_250, n_827, n_248);
  nand g585 (n_828, n_246, n_247);
  nand g586 (n_829, n_248, n_247);
  nand g587 (n_830, n_246, n_248);
  nand g588 (n_263, n_828, n_829, n_830);
  xor g589 (n_831, n_249, n_250);
  xor g590 (n_104, n_831, n_251);
  nand g591 (n_832, n_249, n_250);
  nand g592 (n_833, n_251, n_250);
  nand g593 (n_834, n_249, n_251);
  nand g594 (n_55, n_832, n_833, n_834);
  xor g604 (n_256, n_687, A[15]);
  nand g606 (n_841, A[15], A[8]);
  nand g608 (n_269, n_688, n_841, n_816);
  xor g609 (n_843, A[12], n_185);
  xor g610 (n_259, n_843, A[16]);
  nand g611 (n_844, A[12], n_185);
  nand g612 (n_845, A[16], n_185);
  nand g613 (n_846, A[12], A[16]);
  nand g614 (n_271, n_844, n_845, n_846);
  xor g615 (n_847, A[18], n_186);
  xor g616 (n_260, n_847, n_255);
  nand g617 (n_848, A[18], n_186);
  nand g618 (n_849, n_255, n_186);
  nand g619 (n_850, A[18], n_255);
  nand g620 (n_273, n_848, n_849, n_850);
  xor g621 (n_851, n_256, n_257);
  xor g622 (n_262, n_851, n_258);
  nand g623 (n_852, n_256, n_257);
  nand g624 (n_853, n_258, n_257);
  nand g625 (n_854, n_256, n_258);
  nand g626 (n_274, n_852, n_853, n_854);
  xor g627 (n_855, n_259, n_260);
  xor g628 (n_264, n_855, n_261);
  nand g629 (n_856, n_259, n_260);
  nand g630 (n_857, n_261, n_260);
  nand g631 (n_858, n_259, n_261);
  nand g632 (n_277, n_856, n_857, n_858);
  xor g633 (n_859, n_262, n_263);
  xor g634 (n_103, n_859, n_264);
  nand g635 (n_860, n_262, n_263);
  nand g636 (n_861, n_264, n_263);
  nand g637 (n_862, n_262, n_264);
  nand g638 (n_54, n_860, n_861, n_862);
  xor g641 (n_863, n_118, A[4]);
  xor g642 (n_266, n_863, n_174);
  xor g648 (n_268, n_683, n_266);
  nand g650 (n_869, n_266, A[9]);
  nand g651 (n_870, A[5], n_266);
  nand g652 (n_283, n_684, n_869, n_870);
  xor g653 (n_871, A[8], A[12]);
  xor g654 (n_270, n_871, A[13]);
  nand g656 (n_873, A[13], A[12]);
  nand g657 (n_874, A[8], A[13]);
  nand g658 (n_284, n_741, n_873, n_874);
  xor g659 (n_875, A[17], A[19]);
  xor g660 (n_272, n_875, n_71);
  nand g661 (n_876, A[17], A[19]);
  nand g662 (n_877, n_71, A[19]);
  nand g663 (n_878, A[17], n_71);
  nand g664 (n_286, n_876, n_877, n_878);
  xor g665 (n_879, A[16], n_268);
  xor g666 (n_275, n_879, n_269);
  nand g667 (n_880, A[16], n_268);
  nand g668 (n_881, n_269, n_268);
  nand g669 (n_882, A[16], n_269);
  nand g670 (n_289, n_880, n_881, n_882);
  xor g671 (n_883, n_270, n_271);
  xor g672 (n_276, n_883, n_272);
  nand g673 (n_884, n_270, n_271);
  nand g674 (n_885, n_272, n_271);
  nand g675 (n_886, n_270, n_272);
  nand g676 (n_291, n_884, n_885, n_886);
  xor g677 (n_887, n_273, n_274);
  xor g678 (n_278, n_887, n_275);
  nand g679 (n_888, n_273, n_274);
  nand g680 (n_889, n_275, n_274);
  nand g681 (n_890, n_273, n_275);
  nand g682 (n_293, n_888, n_889, n_890);
  xor g683 (n_891, n_276, n_277);
  xor g684 (n_102, n_891, n_278);
  nand g685 (n_892, n_276, n_277);
  nand g686 (n_893, n_278, n_277);
  nand g687 (n_894, n_276, n_278);
  nand g688 (n_53, n_892, n_893, n_894);
  xor g708 (n_287, n_791, n_199);
  nand g710 (n_909, n_199, A[14]);
  nand g711 (n_910, A[13], n_199);
  nand g712 (n_301, n_792, n_909, n_910);
  xor g713 (n_911, A[18], A[17]);
  xor g714 (n_288, n_911, A[20]);
  nand g715 (n_912, A[18], A[17]);
  nand g716 (n_913, A[20], A[17]);
  nand g717 (n_914, A[18], A[20]);
  nand g718 (n_303, n_912, n_913, n_914);
  xor g719 (n_915, n_283, n_284);
  xor g720 (n_290, n_915, n_201);
  nand g721 (n_916, n_283, n_284);
  nand g722 (n_917, n_201, n_284);
  nand g723 (n_918, n_283, n_201);
  nand g724 (n_304, n_916, n_917, n_918);
  xor g725 (n_919, n_286, n_287);
  xor g726 (n_292, n_919, n_288);
  nand g727 (n_920, n_286, n_287);
  nand g728 (n_921, n_288, n_287);
  nand g729 (n_922, n_286, n_288);
  nand g730 (n_306, n_920, n_921, n_922);
  xor g731 (n_923, n_289, n_290);
  xor g732 (n_294, n_923, n_291);
  nand g733 (n_924, n_289, n_290);
  nand g734 (n_925, n_291, n_290);
  nand g735 (n_926, n_289, n_291);
  nand g736 (n_309, n_924, n_925, n_926);
  xor g737 (n_927, n_292, n_293);
  xor g738 (n_101, n_927, n_294);
  nand g739 (n_928, n_292, n_293);
  nand g740 (n_929, n_294, n_293);
  nand g741 (n_930, n_292, n_294);
  nand g742 (n_52, n_928, n_929, n_930);
  xor g750 (n_298, n_659, A[11]);
  nand g753 (n_938, n_68, A[11]);
  nand g754 (n_314, n_660, n_721, n_938);
  xor g755 (n_939, A[10], n_182);
  xor g756 (n_302, n_939, A[14]);
  nand g757 (n_940, A[10], n_182);
  nand g759 (n_942, A[10], A[14]);
  nand g760 (n_315, n_940, n_820, n_942);
  xor g761 (n_943, n_181, A[15]);
  xor g762 (n_300, n_943, A[19]);
  nand g764 (n_945, A[19], A[15]);
  nand g765 (n_946, n_181, A[19]);
  nand g766 (n_318, n_817, n_945, n_946);
  xor g767 (n_947, A[18], n_298);
  xor g768 (n_305, n_947, A[21]);
  nand g769 (n_948, A[18], n_298);
  nand g770 (n_949, A[21], n_298);
  nand g771 (n_950, A[18], A[21]);
  nand g772 (n_320, n_948, n_949, n_950);
  xor g773 (n_951, n_208, n_300);
  xor g774 (n_307, n_951, n_301);
  nand g775 (n_952, n_208, n_300);
  nand g776 (n_953, n_301, n_300);
  nand g777 (n_954, n_208, n_301);
  nand g778 (n_322, n_952, n_953, n_954);
  xor g779 (n_955, n_302, n_303);
  xor g780 (n_308, n_955, n_304);
  nand g781 (n_956, n_302, n_303);
  nand g782 (n_957, n_304, n_303);
  nand g783 (n_958, n_302, n_304);
  nand g784 (n_324, n_956, n_957, n_958);
  xor g785 (n_959, n_305, n_306);
  xor g786 (n_310, n_959, n_307);
  nand g787 (n_960, n_305, n_306);
  nand g788 (n_961, n_307, n_306);
  nand g789 (n_962, n_305, n_307);
  nand g790 (n_326, n_960, n_961, n_962);
  xor g791 (n_963, n_308, n_309);
  xor g792 (n_100, n_963, n_310);
  nand g793 (n_964, n_308, n_309);
  nand g794 (n_965, n_310, n_309);
  nand g795 (n_966, n_308, n_310);
  nand g796 (n_51, n_964, n_965, n_966);
  xor g812 (n_317, n_843, A[19]);
  nand g814 (n_977, A[19], A[12]);
  nand g815 (n_978, n_185, A[19]);
  nand g816 (n_335, n_844, n_977, n_978);
  xor g817 (n_979, n_186, A[16]);
  xor g818 (n_319, n_979, A[20]);
  nand g819 (n_980, n_186, A[16]);
  nand g820 (n_981, A[20], A[16]);
  nand g821 (n_982, n_186, A[20]);
  nand g822 (n_337, n_980, n_981, n_982);
  xor g823 (n_983, A[22], n_314);
  xor g824 (n_321, n_983, n_315);
  nand g825 (n_984, A[22], n_314);
  nand g826 (n_985, n_315, n_314);
  nand g827 (n_986, A[22], n_315);
  nand g828 (n_339, n_984, n_985, n_986);
  xor g829 (n_987, n_256, n_317);
  xor g830 (n_323, n_987, n_318);
  nand g831 (n_988, n_256, n_317);
  nand g832 (n_989, n_318, n_317);
  nand g833 (n_990, n_256, n_318);
  nand g834 (n_341, n_988, n_989, n_990);
  xor g835 (n_991, n_319, n_320);
  xor g836 (n_325, n_991, n_321);
  nand g837 (n_992, n_319, n_320);
  nand g838 (n_993, n_321, n_320);
  nand g839 (n_994, n_319, n_321);
  nand g840 (n_343, n_992, n_993, n_994);
  xor g841 (n_995, n_322, n_323);
  xor g842 (n_327, n_995, n_324);
  nand g843 (n_996, n_322, n_323);
  nand g844 (n_997, n_324, n_323);
  nand g845 (n_998, n_322, n_324);
  nand g846 (n_345, n_996, n_997, n_998);
  xor g847 (n_999, n_325, n_326);
  xor g848 (n_99, n_999, n_327);
  nand g849 (n_1000, n_325, n_326);
  nand g850 (n_1001, n_327, n_326);
  nand g851 (n_1002, n_325, n_327);
  nand g852 (n_50, n_1000, n_1001, n_1002);
  xor g861 (n_1007, A[5], A[8]);
  xor g862 (n_333, n_1007, A[9]);
  xor g867 (n_1011, n_266, A[13]);
  xor g868 (n_334, n_1011, A[12]);
  nand g869 (n_1012, n_266, A[13]);
  nand g871 (n_1014, n_266, A[12]);
  nand g872 (n_354, n_1012, n_873, n_1014);
  xor g873 (n_1015, A[16], A[17]);
  xor g874 (n_336, n_1015, n_71);
  nand g875 (n_1016, A[16], A[17]);
  nand g877 (n_1018, A[16], n_71);
  nand g878 (n_357, n_1016, n_878, n_1018);
  xor g879 (n_1019, A[21], A[23]);
  xor g880 (n_338, n_1019, A[20]);
  nand g881 (n_1020, A[21], A[23]);
  nand g882 (n_1021, A[20], A[23]);
  nand g883 (n_1022, A[21], A[20]);
  nand g884 (n_359, n_1020, n_1021, n_1022);
  xor g885 (n_1023, n_269, n_333);
  xor g886 (n_340, n_1023, n_334);
  nand g887 (n_1024, n_269, n_333);
  nand g888 (n_1025, n_334, n_333);
  nand g889 (n_1026, n_269, n_334);
  nand g890 (n_361, n_1024, n_1025, n_1026);
  xor g891 (n_1027, n_335, n_336);
  xor g892 (n_342, n_1027, n_337);
  nand g893 (n_1028, n_335, n_336);
  nand g894 (n_1029, n_337, n_336);
  nand g895 (n_1030, n_335, n_337);
  nand g896 (n_363, n_1028, n_1029, n_1030);
  xor g897 (n_1031, n_338, n_339);
  xor g898 (n_344, n_1031, n_340);
  nand g899 (n_1032, n_338, n_339);
  nand g900 (n_1033, n_340, n_339);
  nand g901 (n_1034, n_338, n_340);
  nand g902 (n_365, n_1032, n_1033, n_1034);
  xor g903 (n_1035, n_341, n_342);
  xor g904 (n_346, n_1035, n_343);
  nand g905 (n_1036, n_341, n_342);
  nand g906 (n_1037, n_343, n_342);
  nand g907 (n_1038, n_341, n_343);
  nand g908 (n_367, n_1036, n_1037, n_1038);
  xor g909 (n_1039, n_344, n_345);
  xor g910 (n_98, n_1039, n_346);
  nand g911 (n_1040, n_344, n_345);
  nand g912 (n_1041, n_346, n_345);
  nand g913 (n_1042, n_344, n_346);
  nand g914 (n_49, n_1040, n_1041, n_1042);
  xor g917 (n_1043, A[1], n_171);
  nand g922 (n_372, n_625, n_1045, n_1046);
  xor g924 (n_352, n_699, n_178);
  nand g926 (n_1049, n_178, A[6]);
  nand g927 (n_1050, A[5], n_178);
  nand g928 (n_374, n_650, n_1049, n_1050);
  xor g929 (n_1051, n_351, A[9]);
  xor g930 (n_355, n_1051, A[10]);
  nand g931 (n_1052, n_351, A[9]);
  nand g933 (n_1054, n_351, A[10]);
  nand g934 (n_376, n_1052, n_705, n_1054);
  xor g936 (n_356, n_791, A[18]);
  nand g938 (n_1057, A[18], A[13]);
  nand g939 (n_1058, A[14], A[18]);
  nand g940 (n_380, n_792, n_1057, n_1058);
  xor g941 (n_1059, n_352, A[17]);
  nand g943 (n_1060, n_352, A[17]);
  nand g946 (n_379, n_1060, n_1061, n_1062);
  xor g947 (n_1063, A[22], n_232);
  xor g948 (n_360, n_1063, A[21]);
  nand g949 (n_1064, A[22], n_232);
  nand g950 (n_1065, A[21], n_232);
  nand g951 (n_1066, A[22], A[21]);
  nand g952 (n_382, n_1064, n_1065, n_1066);
  xor g953 (n_1067, n_354, n_355);
  xor g954 (n_362, n_1067, n_356);
  nand g955 (n_1068, n_354, n_355);
  nand g956 (n_1069, n_356, n_355);
  nand g957 (n_1070, n_354, n_356);
  nand g958 (n_384, n_1068, n_1069, n_1070);
  xor g959 (n_1071, n_357, n_358);
  xor g960 (n_364, n_1071, n_359);
  nand g961 (n_1072, n_357, n_358);
  nand g962 (n_1073, n_359, n_358);
  nand g963 (n_1074, n_357, n_359);
  nand g964 (n_385, n_1072, n_1073, n_1074);
  xor g965 (n_1075, n_360, n_361);
  xor g966 (n_366, n_1075, n_362);
  nand g967 (n_1076, n_360, n_361);
  nand g968 (n_1077, n_362, n_361);
  nand g969 (n_1078, n_360, n_362);
  nand g970 (n_388, n_1076, n_1077, n_1078);
  xor g971 (n_1079, n_363, n_364);
  xor g972 (n_368, n_1079, n_365);
  nand g973 (n_1080, n_363, n_364);
  nand g974 (n_1081, n_365, n_364);
  nand g975 (n_1082, n_363, n_365);
  nand g976 (n_391, n_1080, n_1081, n_1082);
  xor g977 (n_1083, n_366, n_367);
  xor g978 (n_97, n_1083, n_368);
  nand g979 (n_1084, n_366, n_367);
  nand g980 (n_1085, n_368, n_367);
  nand g981 (n_1086, n_366, n_368);
  nand g982 (n_48, n_1084, n_1085, n_1086);
  xor g991 (n_1091, A[6], n_372);
  xor g992 (n_375, n_1091, A[7]);
  nand g993 (n_1092, A[6], n_372);
  nand g994 (n_1093, A[7], n_372);
  nand g996 (n_395, n_1092, n_1093, n_720);
  xor g997 (n_1095, n_373, A[10]);
  xor g998 (n_377, n_1095, A[11]);
  nand g999 (n_1096, n_373, A[10]);
  nand g1000 (n_1097, A[11], A[10]);
  nand g1001 (n_1098, n_373, A[11]);
  nand g1002 (n_396, n_1096, n_1097, n_1098);
  xor g1003 (n_1099, A[15], A[14]);
  xor g1004 (n_378, n_1099, n_374);
  nand g1005 (n_1100, A[15], A[14]);
  nand g1006 (n_1101, n_374, A[14]);
  nand g1007 (n_1102, A[15], n_374);
  nand g1008 (n_399, n_1100, n_1101, n_1102);
  xor g1009 (n_1103, A[19], n_375);
  xor g1010 (n_381, n_1103, A[18]);
  nand g1011 (n_1104, A[19], n_375);
  nand g1012 (n_1105, A[18], n_375);
  nand g1013 (n_1106, A[19], A[18]);
  nand g1014 (n_400, n_1104, n_1105, n_1106);
  xor g1015 (n_1107, n_376, A[22]);
  xor g1016 (n_383, n_1107, A[23]);
  nand g1017 (n_1108, n_376, A[22]);
  nand g1018 (n_1109, A[23], A[22]);
  nand g1019 (n_1110, n_376, A[23]);
  nand g1020 (n_403, n_1108, n_1109, n_1110);
  xor g1021 (n_1111, n_377, n_378);
  xor g1022 (n_386, n_1111, n_379);
  nand g1023 (n_1112, n_377, n_378);
  nand g1024 (n_1113, n_379, n_378);
  nand g1025 (n_1114, n_377, n_379);
  nand g1026 (n_405, n_1112, n_1113, n_1114);
  xor g1027 (n_1115, n_380, n_381);
  xor g1028 (n_387, n_1115, n_382);
  nand g1029 (n_1116, n_380, n_381);
  nand g1030 (n_1117, n_382, n_381);
  nand g1031 (n_1118, n_380, n_382);
  nand g1032 (n_406, n_1116, n_1117, n_1118);
  xor g1033 (n_1119, n_383, n_384);
  xor g1034 (n_389, n_1119, n_385);
  nand g1035 (n_1120, n_383, n_384);
  nand g1036 (n_1121, n_385, n_384);
  nand g1037 (n_1122, n_383, n_385);
  nand g1038 (n_409, n_1120, n_1121, n_1122);
  xor g1039 (n_1123, n_386, n_387);
  xor g1040 (n_390, n_1123, n_388);
  nand g1041 (n_1124, n_386, n_387);
  nand g1042 (n_1125, n_388, n_387);
  nand g1043 (n_1126, n_386, n_388);
  nand g1044 (n_411, n_1124, n_1125, n_1126);
  xor g1045 (n_1127, n_389, n_390);
  xor g1046 (n_96, n_1127, n_391);
  nand g1047 (n_1128, n_389, n_390);
  nand g1048 (n_1129, n_391, n_390);
  nand g1049 (n_1130, n_389, n_391);
  nand g1050 (n_47, n_1128, n_1129, n_1130);
  xor g1052 (n_394, n_627, A[4]);
  nand g1054 (n_1133, A[4], A[2]);
  nand g1055 (n_1134, A[3], A[4]);
  nand g1056 (n_413, n_628, n_1133, n_1134);
  xor g1057 (n_1135, n_393, A[7]);
  xor g1058 (n_397, n_1135, n_394);
  nand g1059 (n_1136, n_393, A[7]);
  nand g1060 (n_1137, n_394, A[7]);
  nand g1061 (n_1138, n_393, n_394);
  nand g1062 (n_415, n_1136, n_1137, n_1138);
  xor g1069 (n_1143, A[12], A[19]);
  xor g1070 (n_402, n_1143, A[16]);
  nand g1072 (n_1145, A[16], A[19]);
  nand g1074 (n_418, n_977, n_1145, n_846);
  xor g1076 (n_401, n_1147, A[23]);
  nand g1078 (n_1149, A[23], n_395);
  nand g1080 (n_420, n_1148, n_1149, n_1150);
  xor g1081 (n_1151, n_396, n_397);
  xor g1082 (n_404, n_1151, A[20]);
  nand g1083 (n_1152, n_396, n_397);
  nand g1084 (n_1153, A[20], n_397);
  nand g1085 (n_1154, n_396, A[20]);
  nand g1086 (n_421, n_1152, n_1153, n_1154);
  xor g1087 (n_1155, n_256, n_399);
  xor g1088 (n_407, n_1155, n_400);
  nand g1089 (n_1156, n_256, n_399);
  nand g1090 (n_1157, n_400, n_399);
  nand g1091 (n_1158, n_256, n_400);
  nand g1092 (n_424, n_1156, n_1157, n_1158);
  xor g1093 (n_1159, n_401, n_402);
  xor g1094 (n_408, n_1159, n_403);
  nand g1095 (n_1160, n_401, n_402);
  nand g1096 (n_1161, n_403, n_402);
  nand g1097 (n_1162, n_401, n_403);
  nand g1098 (n_425, n_1160, n_1161, n_1162);
  xor g1099 (n_1163, n_404, n_405);
  xor g1100 (n_410, n_1163, n_406);
  nand g1101 (n_1164, n_404, n_405);
  nand g1102 (n_1165, n_406, n_405);
  nand g1103 (n_1166, n_404, n_406);
  nand g1104 (n_429, n_1164, n_1165, n_1166);
  xor g1105 (n_1167, n_407, n_408);
  xor g1106 (n_412, n_1167, n_409);
  nand g1107 (n_1168, n_407, n_408);
  nand g1108 (n_1169, n_409, n_408);
  nand g1109 (n_1170, n_407, n_409);
  nand g1110 (n_431, n_1168, n_1169, n_1170);
  xor g1111 (n_1171, n_410, n_411);
  xor g1112 (n_95, n_1171, n_412);
  nand g1113 (n_1172, n_410, n_411);
  nand g1114 (n_1173, n_412, n_411);
  nand g1115 (n_1174, n_410, n_412);
  nand g1116 (n_46, n_1172, n_1173, n_1174);
  xor g1117 (n_1175, A[4], A[5]);
  xor g1118 (n_414, n_1175, n_413);
  nand g1119 (n_1176, A[4], A[5]);
  nand g1120 (n_1177, n_413, A[5]);
  nand g1121 (n_1178, A[4], n_413);
  nand g1122 (n_434, n_1176, n_1177, n_1178);
  xor g1123 (n_1179, A[9], A[8]);
  xor g1124 (n_416, n_1179, A[13]);
  nand g1127 (n_1182, A[9], A[13]);
  nand g1128 (n_436, n_761, n_874, n_1182);
  xor g1129 (n_1183, A[12], A[17]);
  xor g1130 (n_419, n_1183, A[16]);
  nand g1131 (n_1184, A[12], A[17]);
  nand g1134 (n_439, n_1184, n_1016, n_846);
  xor g1135 (n_1187, n_414, n_415);
  nand g1137 (n_1188, n_414, n_415);
  nand g1140 (n_438, n_1188, n_1189, n_1190);
  xor g1141 (n_1191, A[21], A[20]);
  xor g1142 (n_423, n_1191, n_416);
  nand g1144 (n_1193, n_416, A[20]);
  nand g1145 (n_1194, A[21], n_416);
  nand g1146 (n_441, n_1022, n_1193, n_1194);
  xor g1147 (n_1195, n_269, n_418);
  xor g1148 (n_426, n_1195, n_419);
  nand g1149 (n_1196, n_269, n_418);
  nand g1150 (n_1197, n_419, n_418);
  nand g1151 (n_1198, n_269, n_419);
  nand g1152 (n_443, n_1196, n_1197, n_1198);
  xor g1153 (n_1199, n_420, n_421);
  xor g1154 (n_427, n_1199, n_422);
  nand g1155 (n_1200, n_420, n_421);
  nand g1156 (n_1201, n_422, n_421);
  nand g1157 (n_1202, n_420, n_422);
  nand g1158 (n_444, n_1200, n_1201, n_1202);
  xor g1159 (n_1203, n_423, n_424);
  xor g1160 (n_428, n_1203, n_425);
  nand g1161 (n_1204, n_423, n_424);
  nand g1162 (n_1205, n_425, n_424);
  nand g1163 (n_1206, n_423, n_425);
  nand g1164 (n_447, n_1204, n_1205, n_1206);
  xor g1165 (n_1207, n_426, n_427);
  xor g1166 (n_430, n_1207, n_428);
  nand g1167 (n_1208, n_426, n_427);
  nand g1168 (n_1209, n_428, n_427);
  nand g1169 (n_1210, n_426, n_428);
  nand g1170 (n_450, n_1208, n_1209, n_1210);
  xor g1171 (n_1211, n_429, n_430);
  xor g1172 (n_94, n_1211, n_431);
  nand g1173 (n_1212, n_429, n_430);
  nand g1174 (n_1213, n_431, n_430);
  nand g1175 (n_1214, n_429, n_431);
  nand g1176 (n_45, n_1212, n_1213, n_1214);
  nand g1183 (n_1218, A[6], A[9]);
  nand g1184 (n_455, n_1216, n_1217, n_1218);
  xor g1185 (n_1219, A[10], A[14]);
  xor g1186 (n_437, n_1219, A[13]);
  nand g1190 (n_457, n_942, n_792, n_726);
  xor g1192 (n_440, n_911, n_434);
  nand g1194 (n_1225, n_434, A[17]);
  nand g1195 (n_1226, A[18], n_434);
  nand g1196 (n_458, n_912, n_1225, n_1226);
  xor g1197 (n_1227, A[21], n_435);
  xor g1198 (n_442, n_1227, A[22]);
  nand g1199 (n_1228, A[21], n_435);
  nand g1200 (n_1229, A[22], n_435);
  nand g1202 (n_460, n_1228, n_1229, n_1066);
  xor g1203 (n_1231, n_436, n_437);
  xor g1204 (n_445, n_1231, n_438);
  nand g1205 (n_1232, n_436, n_437);
  nand g1206 (n_1233, n_438, n_437);
  nand g1207 (n_1234, n_436, n_438);
  nand g1208 (n_462, n_1232, n_1233, n_1234);
  xor g1209 (n_1235, n_439, n_440);
  xor g1210 (n_446, n_1235, n_441);
  nand g1211 (n_1236, n_439, n_440);
  nand g1212 (n_1237, n_441, n_440);
  nand g1213 (n_1238, n_439, n_441);
  nand g1214 (n_465, n_1236, n_1237, n_1238);
  xor g1215 (n_1239, n_442, n_443);
  xor g1216 (n_448, n_1239, n_444);
  nand g1217 (n_1240, n_442, n_443);
  nand g1218 (n_1241, n_444, n_443);
  nand g1219 (n_1242, n_442, n_444);
  nand g1220 (n_466, n_1240, n_1241, n_1242);
  xor g1221 (n_1243, n_445, n_446);
  xor g1222 (n_449, n_1243, n_447);
  nand g1223 (n_1244, n_445, n_446);
  nand g1224 (n_1245, n_447, n_446);
  nand g1225 (n_1246, n_445, n_447);
  nand g1226 (n_469, n_1244, n_1245, n_1246);
  xor g1227 (n_1247, n_448, n_449);
  xor g1228 (n_93, n_1247, n_450);
  nand g1229 (n_1248, n_448, n_449);
  nand g1230 (n_1249, n_450, n_449);
  nand g1231 (n_1250, n_448, n_450);
  nand g1232 (n_44, n_1248, n_1249, n_1250);
  xor g1236 (n_454, n_639, A[10]);
  nand g1238 (n_1253, A[10], A[5]);
  nand g1240 (n_471, n_640, n_1253, n_813);
  xor g1242 (n_456, n_1255, A[15]);
  nand g1246 (n_473, n_1256, n_1257, n_816);
  xor g1247 (n_1259, A[14], A[19]);
  xor g1248 (n_459, n_1259, A[18]);
  nand g1249 (n_1260, A[14], A[19]);
  nand g1252 (n_475, n_1260, n_1106, n_1058);
  xor g1253 (n_1263, A[22], n_454);
  xor g1254 (n_461, n_1263, A[23]);
  nand g1255 (n_1264, A[22], n_454);
  nand g1256 (n_1265, A[23], n_454);
  nand g1258 (n_476, n_1264, n_1265, n_1109);
  xor g1259 (n_1267, n_455, n_456);
  xor g1260 (n_463, n_1267, n_457);
  nand g1261 (n_1268, n_455, n_456);
  nand g1262 (n_1269, n_457, n_456);
  nand g1263 (n_1270, n_455, n_457);
  nand g1264 (n_478, n_1268, n_1269, n_1270);
  xor g1265 (n_1271, n_458, n_459);
  xor g1266 (n_464, n_1271, n_460);
  nand g1267 (n_1272, n_458, n_459);
  nand g1268 (n_1273, n_460, n_459);
  nand g1269 (n_1274, n_458, n_460);
  nand g1270 (n_481, n_1272, n_1273, n_1274);
  xor g1271 (n_1275, n_461, n_462);
  xor g1272 (n_467, n_1275, n_463);
  nand g1273 (n_1276, n_461, n_462);
  nand g1274 (n_1277, n_463, n_462);
  nand g1275 (n_1278, n_461, n_463);
  nand g1276 (n_483, n_1276, n_1277, n_1278);
  xor g1277 (n_1279, n_464, n_465);
  xor g1278 (n_468, n_1279, n_466);
  nand g1279 (n_1280, n_464, n_465);
  nand g1280 (n_1281, n_466, n_465);
  nand g1281 (n_1282, n_464, n_466);
  nand g1282 (n_486, n_1280, n_1281, n_1282);
  xor g1283 (n_1283, n_467, n_468);
  xor g1284 (n_92, n_1283, n_469);
  nand g1285 (n_1284, n_467, n_468);
  nand g1286 (n_1285, n_469, n_468);
  nand g1287 (n_1286, n_467, n_469);
  nand g1288 (n_43, n_1284, n_1285, n_1286);
  xor g1289 (n_1287, A[7], A[11]);
  xor g1290 (n_472, n_1287, A[8]);
  nand g1293 (n_1290, A[7], A[8]);
  nand g1294 (n_487, n_721, n_688, n_1290);
  xor g1295 (n_1291, A[6], A[15]);
  xor g1296 (n_474, n_1291, A[12]);
  nand g1297 (n_1292, A[6], A[15]);
  nand g1298 (n_1293, A[12], A[15]);
  nand g1299 (n_1294, A[6], A[12]);
  nand g1300 (n_489, n_1292, n_1293, n_1294);
  xor g1301 (n_1295, A[19], A[16]);
  nand g1306 (n_490, n_1145, n_1297, n_1298);
  xor g1307 (n_1299, A[23], A[20]);
  xor g1308 (n_479, n_1299, n_471);
  nand g1310 (n_1301, n_471, A[20]);
  nand g1311 (n_1302, A[23], n_471);
  nand g1312 (n_491, n_1021, n_1301, n_1302);
  xor g1313 (n_1303, n_472, n_473);
  xor g1314 (n_480, n_1303, n_474);
  nand g1315 (n_1304, n_472, n_473);
  nand g1316 (n_1305, n_474, n_473);
  nand g1317 (n_1306, n_472, n_474);
  nand g1318 (n_495, n_1304, n_1305, n_1306);
  xor g1319 (n_1307, n_475, n_476);
  xor g1320 (n_482, n_1307, n_477);
  nand g1321 (n_1308, n_475, n_476);
  nand g1322 (n_1309, n_477, n_476);
  nand g1323 (n_1310, n_475, n_477);
  nand g1324 (n_496, n_1308, n_1309, n_1310);
  xor g1325 (n_1311, n_478, n_479);
  xor g1326 (n_484, n_1311, n_480);
  nand g1327 (n_1312, n_478, n_479);
  nand g1328 (n_1313, n_480, n_479);
  nand g1329 (n_1314, n_478, n_480);
  nand g1330 (n_498, n_1312, n_1313, n_1314);
  xor g1331 (n_1315, n_481, n_482);
  xor g1332 (n_485, n_1315, n_483);
  nand g1333 (n_1316, n_481, n_482);
  nand g1334 (n_1317, n_483, n_482);
  nand g1335 (n_1318, n_481, n_483);
  nand g1336 (n_501, n_1316, n_1317, n_1318);
  xor g1337 (n_1319, n_484, n_485);
  xor g1338 (n_91, n_1319, n_486);
  nand g1339 (n_1320, n_484, n_485);
  nand g1340 (n_1321, n_486, n_485);
  nand g1341 (n_1322, n_484, n_486);
  nand g1342 (n_42, n_1320, n_1321, n_1322);
  xor g1356 (n_493, n_1331, n_487);
  nand g1358 (n_1333, n_487, A[21]);
  nand g1360 (n_507, n_1332, n_1333, n_1334);
  xor g1361 (n_1335, A[20], n_416);
  xor g1362 (n_494, n_1335, n_489);
  nand g1364 (n_1337, n_489, n_416);
  nand g1365 (n_1338, A[20], n_489);
  nand g1366 (n_509, n_1193, n_1337, n_1338);
  xor g1367 (n_1339, n_490, n_491);
  xor g1368 (n_497, n_1339, n_419);
  nand g1369 (n_1340, n_490, n_491);
  nand g1370 (n_1341, n_419, n_491);
  nand g1371 (n_1342, n_490, n_419);
  nand g1372 (n_512, n_1340, n_1341, n_1342);
  xor g1373 (n_1343, n_493, n_494);
  xor g1374 (n_499, n_1343, n_495);
  nand g1375 (n_1344, n_493, n_494);
  nand g1376 (n_1345, n_495, n_494);
  nand g1377 (n_1346, n_493, n_495);
  nand g1378 (n_513, n_1344, n_1345, n_1346);
  xor g1379 (n_1347, n_496, n_497);
  xor g1380 (n_500, n_1347, n_498);
  nand g1381 (n_1348, n_496, n_497);
  nand g1382 (n_1349, n_498, n_497);
  nand g1383 (n_1350, n_496, n_498);
  nand g1384 (n_516, n_1348, n_1349, n_1350);
  xor g1385 (n_1351, n_499, n_500);
  xor g1386 (n_90, n_1351, n_501);
  nand g1387 (n_1352, n_499, n_500);
  nand g1388 (n_1353, n_501, n_500);
  nand g1389 (n_1354, n_499, n_501);
  nand g1390 (n_41, n_1352, n_1353, n_1354);
  xor g1393 (n_1355, A[9], A[14]);
  xor g1394 (n_506, n_1355, A[13]);
  nand g1395 (n_1356, A[9], A[14]);
  nand g1398 (n_520, n_1356, n_792, n_1182);
  xor g1400 (n_508, n_1359, A[17]);
  nand g1404 (n_521, n_1360, n_1361, n_912);
  xor g1405 (n_1363, A[21], A[22]);
  xor g1406 (n_510, n_1363, n_436);
  nand g1408 (n_1365, n_436, A[22]);
  nand g1409 (n_1366, A[21], n_436);
  nand g1410 (n_525, n_1066, n_1365, n_1366);
  xor g1411 (n_1367, n_439, n_506);
  xor g1412 (n_511, n_1367, n_507);
  nand g1413 (n_1368, n_439, n_506);
  nand g1414 (n_1369, n_507, n_506);
  nand g1415 (n_1370, n_439, n_507);
  nand g1416 (n_527, n_1368, n_1369, n_1370);
  xor g1417 (n_1371, n_508, n_509);
  xor g1418 (n_514, n_1371, n_510);
  nand g1419 (n_1372, n_508, n_509);
  nand g1420 (n_1373, n_510, n_509);
  nand g1421 (n_1374, n_508, n_510);
  nand g1422 (n_528, n_1372, n_1373, n_1374);
  xor g1423 (n_1375, n_511, n_512);
  xor g1424 (n_515, n_1375, n_513);
  nand g1425 (n_1376, n_511, n_512);
  nand g1426 (n_1377, n_513, n_512);
  nand g1427 (n_1378, n_511, n_513);
  nand g1428 (n_531, n_1376, n_1377, n_1378);
  xor g1429 (n_1379, n_514, n_515);
  xor g1430 (n_89, n_1379, n_516);
  nand g1431 (n_1380, n_514, n_515);
  nand g1432 (n_1381, n_516, n_515);
  nand g1433 (n_1382, n_514, n_516);
  nand g1434 (n_40, n_1380, n_1381, n_1382);
  xor g1437 (n_1383, A[10], A[15]);
  xor g1438 (n_522, n_1383, A[14]);
  nand g1439 (n_1384, A[10], A[15]);
  nand g1442 (n_533, n_1384, n_1100, n_942);
  xor g1444 (n_523, n_1387, A[18]);
  nand g1448 (n_534, n_1388, n_1389, n_1106);
  xor g1449 (n_1391, A[10], A[22]);
  xor g1450 (n_524, n_1391, A[23]);
  nand g1451 (n_1392, A[10], A[22]);
  nand g1453 (n_1394, A[10], A[23]);
  nand g1454 (n_536, n_1392, n_1109, n_1394);
  xor g1455 (n_1395, n_520, n_521);
  xor g1456 (n_526, n_1395, n_522);
  nand g1457 (n_1396, n_520, n_521);
  nand g1458 (n_1397, n_522, n_521);
  nand g1459 (n_1398, n_520, n_522);
  nand g1460 (n_539, n_1396, n_1397, n_1398);
  xor g1461 (n_1399, n_523, n_524);
  xor g1462 (n_529, n_1399, n_525);
  nand g1463 (n_1400, n_523, n_524);
  nand g1464 (n_1401, n_525, n_524);
  nand g1465 (n_1402, n_523, n_525);
  nand g1466 (n_541, n_1400, n_1401, n_1402);
  xor g1467 (n_1403, n_526, n_527);
  xor g1468 (n_530, n_1403, n_528);
  nand g1469 (n_1404, n_526, n_527);
  nand g1470 (n_1405, n_528, n_527);
  nand g1471 (n_1406, n_526, n_528);
  nand g1472 (n_544, n_1404, n_1405, n_1406);
  xor g1473 (n_1407, n_529, n_530);
  xor g1474 (n_88, n_1407, n_531);
  nand g1475 (n_1408, n_529, n_530);
  nand g1476 (n_1409, n_531, n_530);
  nand g1477 (n_1410, n_529, n_531);
  nand g1478 (n_39, n_1408, n_1409, n_1410);
  xor g1480 (n_535, n_815, A[12]);
  nand g1484 (n_545, n_816, n_1293, n_742);
  nand g1487 (n_1416, A[19], A[11]);
  nand g1488 (n_1417, A[16], A[11]);
  nand g1490 (n_546, n_1416, n_1417, n_1145);
  xor g1492 (n_538, n_1419, A[20]);
  nand g1496 (n_549, n_1150, n_1021, n_1422);
  xor g1497 (n_1423, n_533, n_534);
  xor g1498 (n_540, n_1423, n_535);
  nand g1499 (n_1424, n_533, n_534);
  nand g1500 (n_1425, n_535, n_534);
  nand g1501 (n_1426, n_533, n_535);
  nand g1502 (n_550, n_1424, n_1425, n_1426);
  xor g1503 (n_1427, n_536, n_537);
  xor g1504 (n_542, n_1427, n_538);
  nand g1505 (n_1428, n_536, n_537);
  nand g1506 (n_1429, n_538, n_537);
  nand g1507 (n_1430, n_536, n_538);
  nand g1508 (n_553, n_1428, n_1429, n_1430);
  xor g1509 (n_1431, n_539, n_540);
  xor g1510 (n_543, n_1431, n_541);
  nand g1511 (n_1432, n_539, n_540);
  nand g1512 (n_1433, n_541, n_540);
  nand g1513 (n_1434, n_539, n_541);
  nand g1514 (n_555, n_1432, n_1433, n_1434);
  xor g1515 (n_1435, n_542, n_543);
  xor g1516 (n_87, n_1435, n_544);
  nand g1517 (n_1436, n_542, n_543);
  nand g1518 (n_1437, n_544, n_543);
  nand g1519 (n_1438, n_542, n_544);
  nand g1520 (n_38, n_1436, n_1437, n_1438);
  xor g1521 (n_1439, A[13], A[12]);
  xor g1522 (n_547, n_1439, A[17]);
  nand g1525 (n_1442, A[13], A[17]);
  nand g1526 (n_558, n_873, n_1184, n_1442);
  xor g1528 (n_548, n_1443, A[21]);
  nand g1531 (n_1446, A[16], A[21]);
  nand g1532 (n_559, n_1297, n_1332, n_1446);
  xor g1533 (n_1447, A[20], n_545);
  xor g1534 (n_551, n_1447, n_546);
  nand g1535 (n_1448, A[20], n_545);
  nand g1536 (n_1449, n_546, n_545);
  nand g1537 (n_1450, A[20], n_546);
  nand g1538 (n_562, n_1448, n_1449, n_1450);
  xor g1539 (n_1451, n_547, n_548);
  xor g1540 (n_552, n_1451, n_549);
  nand g1541 (n_1452, n_547, n_548);
  nand g1542 (n_1453, n_549, n_548);
  nand g1543 (n_1454, n_547, n_549);
  nand g1544 (n_563, n_1452, n_1453, n_1454);
  xor g1545 (n_1455, n_550, n_551);
  xor g1546 (n_554, n_1455, n_552);
  nand g1547 (n_1456, n_550, n_551);
  nand g1548 (n_1457, n_552, n_551);
  nand g1549 (n_1458, n_550, n_552);
  nand g1550 (n_566, n_1456, n_1457, n_1458);
  xor g1551 (n_1459, n_553, n_554);
  xor g1552 (n_86, n_1459, n_555);
  nand g1553 (n_1460, n_553, n_554);
  nand g1554 (n_1461, n_555, n_554);
  nand g1555 (n_1462, n_553, n_555);
  nand g1556 (n_37, n_1460, n_1461, n_1462);
  xor g1559 (n_1463, A[13], A[18]);
  xor g1560 (n_560, n_1463, A[17]);
  nand g1564 (n_570, n_1057, n_912, n_1442);
  nand g1570 (n_572, n_1066, n_1469, n_1470);
  xor g1571 (n_1471, n_558, n_559);
  xor g1572 (n_564, n_1471, n_560);
  nand g1573 (n_1472, n_558, n_559);
  nand g1574 (n_1473, n_560, n_559);
  nand g1575 (n_1474, n_558, n_560);
  nand g1576 (n_575, n_1472, n_1473, n_1474);
  xor g1577 (n_1475, n_561, n_562);
  xor g1578 (n_565, n_1475, n_563);
  nand g1579 (n_1476, n_561, n_562);
  nand g1580 (n_1477, n_563, n_562);
  nand g1581 (n_1478, n_561, n_563);
  nand g1582 (n_577, n_1476, n_1477, n_1478);
  xor g1583 (n_1479, n_564, n_565);
  xor g1584 (n_85, n_1479, n_566);
  nand g1585 (n_1480, n_564, n_565);
  nand g1586 (n_1481, n_566, n_565);
  nand g1587 (n_1482, n_564, n_566);
  nand g1588 (n_36, n_1480, n_1481, n_1482);
  xor g1597 (n_1487, A[22], A[14]);
  xor g1598 (n_573, n_1487, A[23]);
  nand g1599 (n_1488, A[22], A[14]);
  nand g1600 (n_1489, A[23], A[14]);
  nand g1602 (n_580, n_1488, n_1489, n_1109);
  xor g1604 (n_574, n_1491, n_459);
  nand g1606 (n_1493, n_459, n_570);
  nand g1608 (n_584, n_1492, n_1493, n_1494);
  xor g1609 (n_1495, n_572, n_573);
  xor g1610 (n_576, n_1495, n_574);
  nand g1611 (n_1496, n_572, n_573);
  nand g1612 (n_1497, n_574, n_573);
  nand g1613 (n_1498, n_572, n_574);
  nand g1614 (n_586, n_1496, n_1497, n_1498);
  xor g1615 (n_1499, n_575, n_576);
  xor g1616 (n_84, n_1499, n_577);
  nand g1617 (n_1500, n_575, n_576);
  nand g1618 (n_1501, n_577, n_576);
  nand g1619 (n_1502, n_575, n_577);
  nand g1620 (n_35, n_1500, n_1501, n_1502);
  xor g1621 (n_1503, A[15], A[19]);
  xor g1622 (n_581, n_1503, A[16]);
  nand g1625 (n_1506, A[15], A[16]);
  nand g1626 (n_587, n_945, n_1145, n_1506);
  xor g1633 (n_1511, A[15], n_475);
  xor g1634 (n_583, n_1511, n_580);
  nand g1635 (n_1512, A[15], n_475);
  nand g1636 (n_1513, n_580, n_475);
  nand g1637 (n_1514, A[15], n_580);
  nand g1638 (n_591, n_1512, n_1513, n_1514);
  xor g1639 (n_1515, n_581, n_538);
  xor g1640 (n_585, n_1515, n_583);
  nand g1641 (n_1516, n_581, n_538);
  nand g1642 (n_1517, n_583, n_538);
  nand g1643 (n_1518, n_581, n_583);
  nand g1644 (n_593, n_1516, n_1517, n_1518);
  xor g1645 (n_1519, n_584, n_585);
  xor g1646 (n_83, n_1519, n_586);
  nand g1647 (n_1520, n_584, n_585);
  nand g1648 (n_1521, n_586, n_585);
  nand g1649 (n_1522, n_584, n_586);
  nand g1650 (n_34, n_1520, n_1521, n_1522);
  xor g1652 (n_588, n_1523, A[16]);
  nand g1656 (n_596, n_1061, n_1016, n_1297);
  xor g1658 (n_590, n_1191, n_587);
  nand g1660 (n_1529, n_587, A[20]);
  nand g1661 (n_1530, A[21], n_587);
  nand g1662 (n_598, n_1022, n_1529, n_1530);
  xor g1663 (n_1531, n_588, n_549);
  xor g1664 (n_592, n_1531, n_590);
  nand g1665 (n_1532, n_588, n_549);
  nand g1666 (n_1533, n_590, n_549);
  nand g1667 (n_1534, n_588, n_590);
  nand g1668 (n_600, n_1532, n_1533, n_1534);
  xor g1669 (n_1535, n_591, n_592);
  xor g1670 (n_82, n_1535, n_593);
  nand g1671 (n_1536, n_591, n_592);
  nand g1672 (n_1537, n_593, n_592);
  nand g1673 (n_1538, n_591, n_593);
  nand g1674 (n_81, n_1536, n_1537, n_1538);
  xor g1677 (n_1539, A[17], A[21]);
  xor g1678 (n_597, n_1539, A[22]);
  nand g1679 (n_1540, A[17], A[21]);
  nand g1681 (n_1542, A[17], A[22]);
  nand g1682 (n_604, n_1540, n_1066, n_1542);
  xor g1684 (n_599, n_1543, n_597);
  nand g1686 (n_1545, n_597, n_596);
  nand g1688 (n_607, n_1544, n_1545, n_1546);
  xor g1689 (n_1547, n_598, n_599);
  xor g1690 (n_33, n_1547, n_600);
  nand g1691 (n_1548, n_598, n_599);
  nand g1692 (n_1549, n_600, n_599);
  nand g1693 (n_1550, n_598, n_600);
  nand g1694 (n_80, n_1548, n_1549, n_1550);
  xor g1697 (n_1551, A[18], A[22]);
  xor g1698 (n_605, n_1551, A[23]);
  nand g1699 (n_1552, A[18], A[22]);
  nand g1701 (n_1554, A[18], A[23]);
  nand g1702 (n_610, n_1552, n_1109, n_1554);
  xor g1704 (n_606, n_1555, n_604);
  nand g1706 (n_1557, n_604, A[18]);
  nand g1708 (n_612, n_1556, n_1557, n_1558);
  xor g1709 (n_1559, n_605, n_606);
  xor g1710 (n_32, n_1559, n_607);
  nand g1711 (n_1560, n_605, n_606);
  nand g1712 (n_1561, n_607, n_606);
  nand g1713 (n_1562, n_605, n_607);
  nand g1714 (n_31, n_1560, n_1561, n_1562);
  xor g1716 (n_609, n_1563, A[23]);
  nand g1718 (n_1565, A[23], A[19]);
  nand g1720 (n_613, n_1298, n_1565, n_1150);
  xor g1721 (n_1567, A[20], A[19]);
  xor g1722 (n_611, n_1567, n_609);
  nand g1723 (n_1568, A[20], A[19]);
  nand g1724 (n_1569, n_609, A[19]);
  nand g1725 (n_1570, A[20], n_609);
  nand g1726 (n_615, n_1568, n_1569, n_1570);
  xor g1727 (n_1571, n_610, n_611);
  xor g1728 (n_79, n_1571, n_612);
  nand g1729 (n_1572, n_610, n_611);
  nand g1730 (n_1573, n_612, n_611);
  nand g1731 (n_1574, n_610, n_612);
  nand g1732 (n_30, n_1572, n_1573, n_1574);
  xor g1734 (n_614, n_1331, A[20]);
  nand g1738 (n_618, n_1332, n_1022, n_1422);
  xor g1739 (n_1579, n_613, n_614);
  xor g1740 (n_78, n_1579, n_615);
  nand g1741 (n_1580, n_613, n_614);
  nand g1742 (n_1581, n_615, n_614);
  nand g1743 (n_1582, n_613, n_615);
  nand g1744 (n_77, n_1580, n_1581, n_1582);
  nand g1751 (n_1586, A[22], n_618);
  nand g1752 (n_28, n_1584, n_1585, n_1586);
  xor g1756 (n_76, n_1587, A[21]);
  nand g1760 (n_27, n_1588, n_1589, n_1020);
  xor g1762 (n_75, n_1419, A[22]);
  nand g1766 (n_74, n_1150, n_1109, n_1594);
  nor g11 (n_1610, A[0], A[2]);
  nand g12 (n_1605, A[0], A[2]);
  nor g13 (n_1606, A[3], n_118);
  nand g14 (n_1607, A[3], n_118);
  nor g15 (n_1616, A[4], n_117);
  nand g16 (n_1611, A[4], n_117);
  nor g17 (n_1612, n_68, n_116);
  nand g18 (n_1613, n_68, n_116);
  nor g19 (n_1622, n_67, n_115);
  nand g20 (n_1617, n_67, n_115);
  nor g21 (n_1618, n_66, n_114);
  nand g22 (n_1619, n_66, n_114);
  nor g23 (n_1628, n_65, n_113);
  nand g24 (n_1623, n_65, n_113);
  nor g25 (n_1624, n_64, n_112);
  nand g26 (n_1625, n_64, n_112);
  nor g27 (n_1634, n_63, n_111);
  nand g28 (n_1629, n_63, n_111);
  nor g29 (n_1630, n_62, n_110);
  nand g30 (n_1631, n_62, n_110);
  nor g31 (n_1640, n_61, n_109);
  nand g32 (n_1635, n_61, n_109);
  nor g33 (n_1636, n_60, n_108);
  nand g34 (n_1637, n_60, n_108);
  nor g35 (n_1646, n_59, n_107);
  nand g36 (n_1641, n_59, n_107);
  nor g37 (n_1642, n_58, n_106);
  nand g38 (n_1643, n_58, n_106);
  nor g39 (n_1652, n_57, n_105);
  nand g40 (n_1647, n_57, n_105);
  nor g41 (n_1648, n_56, n_104);
  nand g42 (n_1649, n_56, n_104);
  nor g43 (n_1658, n_55, n_103);
  nand g44 (n_1653, n_55, n_103);
  nor g45 (n_1654, n_54, n_102);
  nand g46 (n_1655, n_54, n_102);
  nor g47 (n_1664, n_53, n_101);
  nand g48 (n_1659, n_53, n_101);
  nor g49 (n_1660, n_52, n_100);
  nand g50 (n_1661, n_52, n_100);
  nor g51 (n_1670, n_51, n_99);
  nand g52 (n_1665, n_51, n_99);
  nor g53 (n_1666, n_50, n_98);
  nand g54 (n_1667, n_50, n_98);
  nor g55 (n_1676, n_49, n_97);
  nand g56 (n_1671, n_49, n_97);
  nor g57 (n_1672, n_48, n_96);
  nand g58 (n_1673, n_48, n_96);
  nor g59 (n_1682, n_47, n_95);
  nand g60 (n_1677, n_47, n_95);
  nor g61 (n_1678, n_46, n_94);
  nand g62 (n_1679, n_46, n_94);
  nor g63 (n_1688, n_45, n_93);
  nand g64 (n_1683, n_45, n_93);
  nor g65 (n_1684, n_44, n_92);
  nand g66 (n_1685, n_44, n_92);
  nor g67 (n_1694, n_43, n_91);
  nand g68 (n_1689, n_43, n_91);
  nor g69 (n_1690, n_42, n_90);
  nand g70 (n_1691, n_42, n_90);
  nor g71 (n_1700, n_41, n_89);
  nand g72 (n_1695, n_41, n_89);
  nor g73 (n_1696, n_40, n_88);
  nand g74 (n_1697, n_40, n_88);
  nor g75 (n_1706, n_39, n_87);
  nand g76 (n_1701, n_39, n_87);
  nor g77 (n_1702, n_38, n_86);
  nand g78 (n_1703, n_38, n_86);
  nor g79 (n_1712, n_37, n_85);
  nand g80 (n_1707, n_37, n_85);
  nor g81 (n_1708, n_36, n_84);
  nand g82 (n_1709, n_36, n_84);
  nor g83 (n_1718, n_35, n_83);
  nand g84 (n_1713, n_35, n_83);
  nor g85 (n_1714, n_34, n_82);
  nand g86 (n_1715, n_34, n_82);
  nor g87 (n_1724, n_33, n_81);
  nand g88 (n_1719, n_33, n_81);
  nor g89 (n_1720, n_32, n_80);
  nand g90 (n_1721, n_32, n_80);
  nor g91 (n_1730, n_31, n_79);
  nand g92 (n_1725, n_31, n_79);
  nor g93 (n_1726, n_30, n_78);
  nand g94 (n_1727, n_30, n_78);
  nor g95 (n_1736, n_29, n_77);
  nand g96 (n_1731, n_29, n_77);
  nor g97 (n_1732, n_28, n_76);
  nand g98 (n_1733, n_28, n_76);
  nor g99 (n_1740, n_27, n_75);
  nand g100 (n_1737, n_27, n_75);
  nor g106 (n_1608, n_1605, n_1606);
  nor g110 (n_1614, n_1611, n_1612);
  nor g113 (n_1750, n_1616, n_1612);
  nor g114 (n_1620, n_1617, n_1618);
  nor g117 (n_1752, n_1622, n_1618);
  nor g118 (n_1626, n_1623, n_1624);
  nor g121 (n_1760, n_1628, n_1624);
  nor g122 (n_1632, n_1629, n_1630);
  nor g125 (n_1762, n_1634, n_1630);
  nor g126 (n_1638, n_1635, n_1636);
  nor g129 (n_1770, n_1640, n_1636);
  nor g130 (n_1644, n_1641, n_1642);
  nor g133 (n_1772, n_1646, n_1642);
  nor g134 (n_1650, n_1647, n_1648);
  nor g137 (n_1780, n_1652, n_1648);
  nor g138 (n_1656, n_1653, n_1654);
  nor g141 (n_1782, n_1658, n_1654);
  nor g142 (n_1662, n_1659, n_1660);
  nor g145 (n_1790, n_1664, n_1660);
  nor g146 (n_1668, n_1665, n_1666);
  nor g149 (n_1792, n_1670, n_1666);
  nor g150 (n_1674, n_1671, n_1672);
  nor g153 (n_1800, n_1676, n_1672);
  nor g154 (n_1680, n_1677, n_1678);
  nor g157 (n_1802, n_1682, n_1678);
  nor g158 (n_1686, n_1683, n_1684);
  nor g161 (n_1810, n_1688, n_1684);
  nor g162 (n_1692, n_1689, n_1690);
  nor g165 (n_1812, n_1694, n_1690);
  nor g166 (n_1698, n_1695, n_1696);
  nor g169 (n_1820, n_1700, n_1696);
  nor g170 (n_1704, n_1701, n_1702);
  nor g173 (n_1822, n_1706, n_1702);
  nor g174 (n_1710, n_1707, n_1708);
  nor g177 (n_1830, n_1712, n_1708);
  nor g178 (n_1716, n_1713, n_1714);
  nor g181 (n_1832, n_1718, n_1714);
  nor g182 (n_1722, n_1719, n_1720);
  nor g185 (n_1840, n_1724, n_1720);
  nor g186 (n_1728, n_1725, n_1726);
  nor g189 (n_1842, n_1730, n_1726);
  nor g190 (n_1734, n_1731, n_1732);
  nor g193 (n_1850, n_1736, n_1732);
  nor g203 (n_1748, n_1622, n_1747);
  nand g212 (n_1860, n_1750, n_1752);
  nor g213 (n_1758, n_1634, n_1757);
  nand g222 (n_1867, n_1760, n_1762);
  nor g223 (n_1768, n_1646, n_1767);
  nand g232 (n_1875, n_1770, n_1772);
  nor g233 (n_1778, n_1658, n_1777);
  nand g242 (n_1882, n_1780, n_1782);
  nor g243 (n_1788, n_1670, n_1787);
  nand g252 (n_1890, n_1790, n_1792);
  nor g253 (n_1798, n_1682, n_1797);
  nand g262 (n_1897, n_1800, n_1802);
  nor g263 (n_1808, n_1694, n_1807);
  nand g1776 (n_1905, n_1810, n_1812);
  nor g1777 (n_1818, n_1706, n_1817);
  nand g1786 (n_1912, n_1820, n_1822);
  nor g1787 (n_1828, n_1718, n_1827);
  nand g1796 (n_1920, n_1830, n_1832);
  nor g1797 (n_1838, n_1730, n_1837);
  nand g1806 (n_1927, n_1840, n_1842);
  nor g1807 (n_1848, n_1740, n_1847);
  nand g1814 (n_2131, n_1611, n_1854);
  nand g1816 (n_2133, n_1747, n_1855);
  nand g1819 (n_2136, n_1858, n_1859);
  nand g1822 (n_1935, n_1862, n_1863);
  nor g1823 (n_1865, n_1640, n_1864);
  nor g1826 (n_1945, n_1640, n_1867);
  nor g1832 (n_1873, n_1871, n_1864);
  nor g1835 (n_1951, n_1867, n_1871);
  nor g1836 (n_1877, n_1875, n_1864);
  nor g1839 (n_1954, n_1867, n_1875);
  nor g1840 (n_1880, n_1664, n_1879);
  nor g1843 (n_2034, n_1664, n_1882);
  nor g1849 (n_1888, n_1886, n_1879);
  nor g1852 (n_2040, n_1882, n_1886);
  nor g1853 (n_1892, n_1890, n_1879);
  nor g1856 (n_1960, n_1882, n_1890);
  nor g1857 (n_1895, n_1688, n_1894);
  nor g1860 (n_1973, n_1688, n_1897);
  nor g1866 (n_1903, n_1901, n_1894);
  nor g1869 (n_1983, n_1897, n_1901);
  nor g1870 (n_1907, n_1905, n_1894);
  nor g1873 (n_1988, n_1897, n_1905);
  nor g1874 (n_1910, n_1712, n_1909);
  nor g1877 (n_2086, n_1712, n_1912);
  nor g1883 (n_1918, n_1916, n_1909);
  nor g1886 (n_2092, n_1912, n_1916);
  nor g1887 (n_1922, n_1920, n_1909);
  nor g1890 (n_1996, n_1912, n_1920);
  nor g1891 (n_1925, n_1736, n_1924);
  nor g1894 (n_2009, n_1736, n_1927);
  nor g1900 (n_1933, n_1931, n_1924);
  nor g1903 (n_2019, n_1927, n_1931);
  nand g1906 (n_2140, n_1623, n_1937);
  nand g1907 (n_1938, n_1760, n_1935);
  nand g1908 (n_2142, n_1757, n_1938);
  nand g1911 (n_2145, n_1941, n_1942);
  nand g1914 (n_2148, n_1864, n_1944);
  nand g1915 (n_1947, n_1945, n_1935);
  nand g1916 (n_2151, n_1946, n_1947);
  nand g1917 (n_1950, n_1948, n_1935);
  nand g1918 (n_2153, n_1949, n_1950);
  nand g1919 (n_1953, n_1951, n_1935);
  nand g1920 (n_2156, n_1952, n_1953);
  nand g1921 (n_1956, n_1954, n_1935);
  nand g1922 (n_2024, n_1955, n_1956);
  nor g1923 (n_1958, n_1676, n_1957);
  nand g1932 (n_2048, n_1800, n_1960);
  nor g1933 (n_1967, n_1965, n_1957);
  nor g1938 (n_1970, n_1897, n_1957);
  nand g1947 (n_2060, n_1960, n_1973);
  nand g1952 (n_2064, n_1960, n_1978);
  nand g1957 (n_2068, n_1960, n_1983);
  nand g1962 (n_2072, n_1960, n_1988);
  nor g1963 (n_1994, n_1724, n_1993);
  nand g1972 (n_2100, n_1840, n_1996);
  nor g1973 (n_2003, n_2001, n_1993);
  nor g1978 (n_2006, n_1927, n_1993);
  nand g1987 (n_2112, n_1996, n_2009);
  nand g1992 (n_2116, n_1996, n_2014);
  nand g1997 (n_2120, n_1996, n_2019);
  nand g2000 (n_2160, n_1647, n_2026);
  nand g2001 (n_2027, n_1780, n_2024);
  nand g2002 (n_2162, n_1777, n_2027);
  nand g2005 (n_2165, n_2030, n_2031);
  nand g2008 (n_2168, n_1879, n_2033);
  nand g2009 (n_2036, n_2034, n_2024);
  nand g2010 (n_2171, n_2035, n_2036);
  nand g2011 (n_2039, n_2037, n_2024);
  nand g2012 (n_2173, n_2038, n_2039);
  nand g2013 (n_2042, n_2040, n_2024);
  nand g2014 (n_2176, n_2041, n_2042);
  nand g2015 (n_2043, n_1960, n_2024);
  nand g2016 (n_2178, n_1957, n_2043);
  nand g2019 (n_2181, n_2046, n_2047);
  nand g2022 (n_2183, n_2050, n_2051);
  nand g2025 (n_2186, n_2054, n_2055);
  nand g2028 (n_2189, n_2058, n_2059);
  nand g2031 (n_2192, n_2062, n_2063);
  nand g2034 (n_2194, n_2066, n_2067);
  nand g2037 (n_2197, n_2070, n_2071);
  nand g2040 (n_2076, n_2074, n_2075);
  nand g2043 (n_2201, n_1695, n_2078);
  nand g2044 (n_2079, n_1820, n_2076);
  nand g2045 (n_2203, n_1817, n_2079);
  nand g2048 (n_2206, n_2082, n_2083);
  nand g2051 (n_2209, n_1909, n_2085);
  nand g2052 (n_2088, n_2086, n_2076);
  nand g2053 (n_2212, n_2087, n_2088);
  nand g2054 (n_2091, n_2089, n_2076);
  nand g2055 (n_2214, n_2090, n_2091);
  nand g2056 (n_2094, n_2092, n_2076);
  nand g2057 (n_2217, n_2093, n_2094);
  nand g2058 (n_2095, n_1996, n_2076);
  nand g2059 (n_2219, n_1993, n_2095);
  nand g2062 (n_2222, n_2098, n_2099);
  nand g2065 (n_2224, n_2102, n_2103);
  nand g2068 (n_2227, n_2106, n_2107);
  nand g2071 (n_2230, n_2110, n_2111);
  nand g2074 (n_2233, n_2114, n_2115);
  nand g2077 (n_2235, n_2118, n_2119);
  nand g2080 (n_2238, n_2122, n_2123);
  xnor g2092 (Z[5], n_2131, n_2132);
  xnor g2094 (Z[6], n_2133, n_2134);
  xnor g2097 (Z[7], n_2136, n_2137);
  xnor g2099 (Z[8], n_1935, n_2138);
  xnor g2102 (Z[9], n_2140, n_2141);
  xnor g2104 (Z[10], n_2142, n_2143);
  xnor g2107 (Z[11], n_2145, n_2146);
  xnor g2110 (Z[12], n_2148, n_2149);
  xnor g2113 (Z[13], n_2151, n_2152);
  xnor g2115 (Z[14], n_2153, n_2154);
  xnor g2118 (Z[15], n_2156, n_2157);
  xnor g2120 (Z[16], n_2024, n_2158);
  xnor g2123 (Z[17], n_2160, n_2161);
  xnor g2125 (Z[18], n_2162, n_2163);
  xnor g2128 (Z[19], n_2165, n_2166);
  xnor g2131 (Z[20], n_2168, n_2169);
  xnor g2134 (Z[21], n_2171, n_2172);
  xnor g2136 (Z[22], n_2173, n_2174);
  xnor g2139 (Z[23], n_2176, n_2177);
  xnor g2141 (Z[24], n_2178, n_2179);
  xnor g2144 (Z[25], n_2181, n_2182);
  xnor g2146 (Z[26], n_2183, n_2184);
  xnor g2149 (Z[27], n_2186, n_2187);
  xnor g2152 (Z[28], n_2189, n_2190);
  xnor g2155 (Z[29], n_2192, n_2193);
  xnor g2157 (Z[30], n_2194, n_2195);
  xnor g2160 (Z[31], n_2197, n_2198);
  xnor g2162 (Z[32], n_2076, n_2199);
  xnor g2165 (Z[33], n_2201, n_2202);
  xnor g2167 (Z[34], n_2203, n_2204);
  xnor g2170 (Z[35], n_2206, n_2207);
  xnor g2173 (Z[36], n_2209, n_2210);
  xnor g2176 (Z[37], n_2212, n_2213);
  xnor g2178 (Z[38], n_2214, n_2215);
  xnor g2181 (Z[39], n_2217, n_2218);
  xnor g2183 (Z[40], n_2219, n_2220);
  xnor g2186 (Z[41], n_2222, n_2223);
  xnor g2188 (Z[42], n_2224, n_2225);
  xnor g2191 (Z[43], n_2227, n_2228);
  xnor g2194 (Z[44], n_2230, n_2231);
  xnor g2197 (Z[45], n_2233, n_2234);
  xnor g2199 (Z[46], n_2235, n_2236);
  xnor g2202 (Z[47], n_2238, n_2239);
  or g2216 (n_1045, A[2], wc);
  not gc (wc, n_171);
  or g2217 (n_1046, wc0, A[2]);
  not gc0 (wc0, A[1]);
  or g2218 (n_1061, wc1, A[24]);
  not gc1 (wc1, A[17]);
  or g2219 (n_1090, A[2], wc2);
  not gc2 (wc2, A[3]);
  or g2220 (n_1150, wc3, A[24]);
  not gc3 (wc3, A[23]);
  or g2222 (n_1216, A[5], wc4);
  not gc4 (wc4, A[6]);
  or g2223 (n_1217, A[5], wc5);
  not gc5 (wc5, A[9]);
  xnor g2224 (n_1255, A[11], A[6]);
  or g2225 (n_1256, A[6], wc6);
  not gc6 (wc6, A[11]);
  or g2226 (n_1257, A[6], wc7);
  not gc7 (wc7, A[15]);
  xnor g2227 (n_477, n_1295, A[24]);
  or g2228 (n_1297, wc8, A[24]);
  not gc8 (wc8, A[16]);
  or g2229 (n_1298, wc9, A[24]);
  not gc9 (wc9, A[19]);
  xnor g2230 (n_1331, A[24], A[21]);
  or g2231 (n_1332, wc10, A[24]);
  not gc10 (wc10, A[21]);
  xnor g2232 (n_1359, A[18], A[10]);
  or g2233 (n_1360, A[10], wc11);
  not gc11 (wc11, A[18]);
  or g2234 (n_1361, A[10], wc12);
  not gc12 (wc12, A[17]);
  xnor g2235 (n_1387, A[19], A[11]);
  or g2236 (n_1388, A[11], wc13);
  not gc13 (wc13, A[19]);
  or g2237 (n_1389, A[11], wc14);
  not gc14 (wc14, A[18]);
  xnor g2239 (n_1419, A[24], A[23]);
  or g2240 (n_1422, wc15, A[24]);
  not gc15 (wc15, A[20]);
  xnor g2241 (n_1443, A[24], A[16]);
  xnor g2242 (n_561, n_1363, A[14]);
  or g2243 (n_1469, A[14], wc16);
  not gc16 (wc16, A[22]);
  or g2244 (n_1470, A[14], wc17);
  not gc17 (wc17, A[21]);
  xnor g2245 (n_1523, A[24], A[17]);
  xnor g2246 (n_1555, A[19], A[18]);
  or g2247 (n_1556, wc18, A[19]);
  not gc18 (wc18, A[18]);
  xnor g2248 (n_1563, A[24], A[19]);
  or g2250 (n_1584, A[21], wc19);
  not gc19 (wc19, A[22]);
  xnor g2251 (n_1587, A[23], A[22]);
  or g2252 (n_1588, A[22], wc20);
  not gc20 (wc20, A[23]);
  or g2253 (n_1589, wc21, A[22]);
  not gc21 (wc21, A[21]);
  or g2254 (n_1594, wc22, A[24]);
  not gc22 (wc22, A[22]);
  xnor g2255 (n_351, n_1043, A[2]);
  xnor g2256 (n_373, n_627, A[2]);
  nand g2257 (n_393, n_628, n_1090);
  xnor g2258 (n_435, n_699, A[9]);
  or g2259 (n_1334, A[24], wc23);
  not gc23 (wc23, n_487);
  xnor g2260 (n_537, n_1387, A[16]);
  xnor g2261 (n_1491, n_570, A[15]);
  or g2262 (n_1492, A[15], wc24);
  not gc24 (wc24, n_570);
  or g2263 (n_1494, A[15], wc25);
  not gc25 (wc25, n_459);
  or g2264 (n_1546, A[18], wc26);
  not gc26 (wc26, n_597);
  or g2265 (n_1558, A[19], wc27);
  not gc27 (wc27, n_604);
  or g2267 (n_2125, wc28, n_1610);
  not gc28 (wc28, n_1605);
  xnor g2268 (n_1543, n_596, A[18]);
  or g2269 (n_1544, A[18], wc29);
  not gc29 (wc29, n_596);
  xnor g2270 (n_29, n_1363, n_618);
  or g2271 (n_1585, A[21], wc30);
  not gc30 (wc30, n_618);
  and g2272 (n_1745, wc31, n_1607);
  not gc31 (wc31, n_1608);
  or g2273 (n_2128, wc32, n_1606);
  not gc32 (wc32, n_1607);
  or g2274 (n_1062, A[24], wc33);
  not gc33 (wc33, n_352);
  or g2275 (n_1190, A[24], wc34);
  not gc34 (wc34, n_414);
  and g2276 (n_1738, wc35, n_74);
  not gc35 (wc35, A[24]);
  or g2277 (n_1739, wc36, n_74);
  not gc36 (wc36, A[24]);
  not g2278 (Z[2], n_2125);
  or g2279 (n_2129, wc37, n_1616);
  not gc37 (wc37, n_1611);
  xnor g2280 (n_358, n_1059, A[24]);
  xnor g2281 (n_1147, n_395, A[24]);
  or g2282 (n_1148, A[24], wc38);
  not gc38 (wc38, n_395);
  or g2283 (n_1189, A[24], wc39);
  not gc39 (wc39, n_415);
  and g2284 (n_1747, wc40, n_1613);
  not gc40 (wc40, n_1614);
  or g2287 (n_1856, wc41, n_1622);
  not gc41 (wc41, n_1750);
  or g2288 (n_2132, wc42, n_1612);
  not gc42 (wc42, n_1613);
  or g2289 (n_2134, wc43, n_1622);
  not gc43 (wc43, n_1617);
  or g2290 (n_2236, wc44, n_1740);
  not gc44 (wc44, n_1737);
  xnor g2291 (n_422, n_1187, A[24]);
  and g2292 (n_1754, wc45, n_1619);
  not gc45 (wc45, n_1620);
  or g2293 (n_1854, n_1616, n_1745);
  or g2294 (n_1855, n_1745, wc46);
  not gc46 (wc46, n_1750);
  xor g2295 (Z[3], n_1605, n_2128);
  xor g2296 (Z[4], n_1745, n_2129);
  or g2297 (n_2137, wc47, n_1618);
  not gc47 (wc47, n_1619);
  or g2298 (n_2239, wc48, n_1738);
  not gc48 (wc48, n_1739);
  and g2299 (n_1858, wc49, n_1617);
  not gc49 (wc49, n_1748);
  and g2300 (n_1755, wc50, n_1752);
  not gc50 (wc50, n_1747);
  or g2301 (n_1859, n_1745, n_1856);
  or g2302 (n_2138, wc51, n_1628);
  not gc51 (wc51, n_1623);
  or g2303 (n_2234, wc52, n_1732);
  not gc52 (wc52, n_1733);
  and g2304 (n_1757, wc53, n_1625);
  not gc53 (wc53, n_1626);
  and g2305 (n_1862, wc54, n_1754);
  not gc54 (wc54, n_1755);
  or g2306 (n_1863, n_1860, n_1745);
  or g2307 (n_2141, wc55, n_1624);
  not gc55 (wc55, n_1625);
  or g2308 (n_2228, wc56, n_1726);
  not gc56 (wc56, n_1727);
  and g2309 (n_1764, wc57, n_1631);
  not gc57 (wc57, n_1632);
  and g2310 (n_1844, wc58, n_1727);
  not gc58 (wc58, n_1728);
  and g2311 (n_1847, wc59, n_1733);
  not gc59 (wc59, n_1734);
  or g2312 (n_1939, wc60, n_1634);
  not gc60 (wc60, n_1760);
  or g2313 (n_1931, wc61, n_1740);
  not gc61 (wc61, n_1850);
  or g2314 (n_2143, wc62, n_1634);
  not gc62 (wc62, n_1629);
  or g2315 (n_2146, wc63, n_1630);
  not gc63 (wc63, n_1631);
  or g2316 (n_2149, wc64, n_1640);
  not gc64 (wc64, n_1635);
  or g2317 (n_2223, wc65, n_1720);
  not gc65 (wc65, n_1721);
  or g2318 (n_2225, wc66, n_1730);
  not gc66 (wc66, n_1725);
  or g2319 (n_2231, wc67, n_1736);
  not gc67 (wc67, n_1731);
  and g2320 (n_1837, wc68, n_1721);
  not gc68 (wc68, n_1722);
  and g2321 (n_1941, wc69, n_1629);
  not gc69 (wc69, n_1758);
  and g2322 (n_1765, wc70, n_1762);
  not gc70 (wc70, n_1757);
  or g2323 (n_2001, wc71, n_1730);
  not gc71 (wc71, n_1840);
  or g2324 (n_1937, wc72, n_1628);
  not gc72 (wc72, n_1935);
  or g2325 (n_2218, wc73, n_1714);
  not gc73 (wc73, n_1715);
  or g2326 (n_2220, wc74, n_1724);
  not gc74 (wc74, n_1719);
  and g2327 (n_1767, wc75, n_1637);
  not gc75 (wc75, n_1638);
  and g2328 (n_1834, wc76, n_1715);
  not gc76 (wc76, n_1716);
  and g2329 (n_1864, wc77, n_1764);
  not gc77 (wc77, n_1765);
  or g2330 (n_1871, wc78, n_1646);
  not gc78 (wc78, n_1770);
  and g2331 (n_1845, wc79, n_1842);
  not gc79 (wc79, n_1837);
  and g2332 (n_1932, wc80, n_1737);
  not gc80 (wc80, n_1848);
  and g2333 (n_2014, wc81, n_1850);
  not gc81 (wc81, n_1927);
  or g2334 (n_1942, n_1939, wc82);
  not gc82 (wc82, n_1935);
  or g2335 (n_1944, wc83, n_1867);
  not gc83 (wc83, n_1935);
  or g2336 (n_2152, wc84, n_1636);
  not gc84 (wc84, n_1637);
  or g2337 (n_2154, wc85, n_1646);
  not gc85 (wc85, n_1641);
  or g2338 (n_2213, wc86, n_1708);
  not gc86 (wc86, n_1709);
  or g2339 (n_2215, wc87, n_1718);
  not gc87 (wc87, n_1713);
  and g2340 (n_1774, wc88, n_1643);
  not gc88 (wc88, n_1644);
  and g2341 (n_1827, wc89, n_1709);
  not gc89 (wc89, n_1710);
  or g2342 (n_1916, wc90, n_1718);
  not gc90 (wc90, n_1830);
  and g2343 (n_2002, wc91, n_1725);
  not gc91 (wc91, n_1838);
  and g2344 (n_1924, wc92, n_1844);
  not gc92 (wc92, n_1845);
  and g2345 (n_1869, wc93, n_1770);
  not gc93 (wc93, n_1864);
  and g2346 (n_1948, wc94, n_1770);
  not gc94 (wc94, n_1867);
  or g2347 (n_2157, wc95, n_1642);
  not gc95 (wc95, n_1643);
  or g2348 (n_2210, wc96, n_1712);
  not gc96 (wc96, n_1707);
  and g2349 (n_1777, wc97, n_1649);
  not gc97 (wc97, n_1650);
  and g2350 (n_1784, wc98, n_1655);
  not gc98 (wc98, n_1656);
  and g2351 (n_1824, wc99, n_1703);
  not gc99 (wc99, n_1704);
  and g2352 (n_1872, wc100, n_1641);
  not gc100 (wc100, n_1768);
  and g2353 (n_1775, wc101, n_1772);
  not gc101 (wc101, n_1767);
  or g2354 (n_2028, wc102, n_1658);
  not gc102 (wc102, n_1780);
  and g2355 (n_1835, wc103, n_1832);
  not gc103 (wc103, n_1827);
  and g2356 (n_1946, wc104, n_1635);
  not gc104 (wc104, n_1865);
  and g2357 (n_1949, wc105, n_1767);
  not gc105 (wc105, n_1869);
  and g2358 (n_1929, wc106, n_1850);
  not gc106 (wc106, n_1924);
  or g2359 (n_2158, wc107, n_1652);
  not gc107 (wc107, n_1647);
  or g2360 (n_2161, wc108, n_1648);
  not gc108 (wc108, n_1649);
  or g2361 (n_2163, wc109, n_1658);
  not gc109 (wc109, n_1653);
  or g2362 (n_2166, wc110, n_1654);
  not gc110 (wc110, n_1655);
  or g2363 (n_2202, wc111, n_1696);
  not gc111 (wc111, n_1697);
  or g2364 (n_2204, wc112, n_1706);
  not gc112 (wc112, n_1701);
  or g2365 (n_2207, wc113, n_1702);
  not gc113 (wc113, n_1703);
  and g2366 (n_1787, wc114, n_1661);
  not gc114 (wc114, n_1662);
  and g2367 (n_1876, wc115, n_1774);
  not gc115 (wc115, n_1775);
  and g2368 (n_1785, wc116, n_1782);
  not gc116 (wc116, n_1777);
  or g2369 (n_1886, wc117, n_1670);
  not gc117 (wc117, n_1790);
  and g2370 (n_1917, wc118, n_1713);
  not gc118 (wc118, n_1828);
  and g2371 (n_1921, wc119, n_1834);
  not gc119 (wc119, n_1835);
  and g2372 (n_2011, wc120, n_1731);
  not gc120 (wc120, n_1925);
  and g2373 (n_2016, wc121, n_1847);
  not gc121 (wc121, n_1929);
  and g2374 (n_2021, n_1932, wc122);
  not gc122 (wc122, n_1933);
  or g2375 (n_2169, wc123, n_1664);
  not gc123 (wc123, n_1659);
  or g2376 (n_2172, wc124, n_1660);
  not gc124 (wc124, n_1661);
  or g2377 (n_2174, wc125, n_1670);
  not gc125 (wc125, n_1665);
  and g2378 (n_1794, wc126, n_1667);
  not gc126 (wc126, n_1668);
  and g2379 (n_1797, wc127, n_1673);
  not gc127 (wc127, n_1674);
  and g2380 (n_2030, wc128, n_1653);
  not gc128 (wc128, n_1778);
  and g2381 (n_1879, wc129, n_1784);
  not gc129 (wc129, n_1785);
  or g2382 (n_1965, wc130, n_1682);
  not gc130 (wc130, n_1800);
  and g2383 (n_1952, n_1872, wc131);
  not gc131 (wc131, n_1873);
  and g2384 (n_2037, wc132, n_1790);
  not gc132 (wc132, n_1882);
  or g2385 (n_2177, wc133, n_1666);
  not gc133 (wc133, n_1667);
  or g2386 (n_2179, wc134, n_1676);
  not gc134 (wc134, n_1671);
  or g2387 (n_2182, wc135, n_1672);
  not gc135 (wc135, n_1673);
  or g2388 (n_2184, wc136, n_1682);
  not gc136 (wc136, n_1677);
  and g2389 (n_1804, wc137, n_1679);
  not gc137 (wc137, n_1680);
  and g2390 (n_1887, wc138, n_1665);
  not gc138 (wc138, n_1788);
  and g2391 (n_1795, wc139, n_1792);
  not gc139 (wc139, n_1787);
  and g2392 (n_1955, n_1876, wc140);
  not gc140 (wc140, n_1877);
  and g2393 (n_1884, wc141, n_1790);
  not gc141 (wc141, n_1879);
  or g2394 (n_2187, wc142, n_1678);
  not gc142 (wc142, n_1679);
  or g2395 (n_2190, wc143, n_1688);
  not gc143 (wc143, n_1683);
  and g2396 (n_1807, wc144, n_1685);
  not gc144 (wc144, n_1686);
  and g2397 (n_1814, wc145, n_1691);
  not gc145 (wc145, n_1692);
  and g2398 (n_1817, wc146, n_1697);
  not gc146 (wc146, n_1698);
  and g2399 (n_1891, wc147, n_1794);
  not gc147 (wc147, n_1795);
  and g2400 (n_1966, wc148, n_1677);
  not gc148 (wc148, n_1798);
  and g2401 (n_1805, wc149, n_1802);
  not gc149 (wc149, n_1797);
  or g2402 (n_1901, wc150, n_1694);
  not gc150 (wc150, n_1810);
  or g2403 (n_2080, wc151, n_1706);
  not gc151 (wc151, n_1820);
  and g2404 (n_2035, wc152, n_1659);
  not gc152 (wc152, n_1880);
  and g2405 (n_2038, wc153, n_1787);
  not gc153 (wc153, n_1884);
  or g2406 (n_2044, wc154, n_1676);
  not gc154 (wc154, n_1960);
  or g2407 (n_2052, n_1965, wc155);
  not gc155 (wc155, n_1960);
  or g2408 (n_2193, wc156, n_1684);
  not gc156 (wc156, n_1685);
  or g2409 (n_2195, wc157, n_1694);
  not gc157 (wc157, n_1689);
  or g2410 (n_2198, wc158, n_1690);
  not gc158 (wc158, n_1691);
  or g2411 (n_2199, wc159, n_1700);
  not gc159 (wc159, n_1695);
  and g2412 (n_1894, wc160, n_1804);
  not gc160 (wc160, n_1805);
  and g2413 (n_1815, wc161, n_1812);
  not gc161 (wc161, n_1807);
  and g2414 (n_1825, wc162, n_1822);
  not gc162 (wc162, n_1817);
  and g2415 (n_2041, n_1887, wc163);
  not gc163 (wc163, n_1888);
  and g2416 (n_1978, wc164, n_1810);
  not gc164 (wc164, n_1897);
  and g2417 (n_2089, wc165, n_1830);
  not gc165 (wc165, n_1912);
  or g2418 (n_2056, wc166, n_1897);
  not gc166 (wc166, n_1960);
  or g2419 (n_2026, wc167, n_1652);
  not gc167 (wc167, n_2024);
  or g2420 (n_2031, n_2028, wc168);
  not gc168 (wc168, n_2024);
  or g2421 (n_2033, wc169, n_1882);
  not gc169 (wc169, n_2024);
  and g2422 (n_1902, wc170, n_1689);
  not gc170 (wc170, n_1808);
  and g2423 (n_1906, wc171, n_1814);
  not gc171 (wc171, n_1815);
  and g2424 (n_2082, wc172, n_1701);
  not gc172 (wc172, n_1818);
  and g2425 (n_1909, wc173, n_1824);
  not gc173 (wc173, n_1825);
  and g2426 (n_1957, n_1891, wc174);
  not gc174 (wc174, n_1892);
  and g2427 (n_1899, wc175, n_1810);
  not gc175 (wc175, n_1894);
  or g2428 (n_2096, wc176, n_1724);
  not gc176 (wc176, n_1996);
  or g2429 (n_2104, n_2001, wc177);
  not gc177 (wc177, n_1996);
  or g2430 (n_2108, wc178, n_1927);
  not gc178 (wc178, n_1996);
  or g2431 (n_2047, n_2044, wc179);
  not gc179 (wc179, n_2024);
  or g2432 (n_2051, n_2048, wc180);
  not gc180 (wc180, n_2024);
  or g2433 (n_2055, n_2052, wc181);
  not gc181 (wc181, n_2024);
  and g2434 (n_1975, wc182, n_1683);
  not gc182 (wc182, n_1895);
  and g2435 (n_1980, wc183, n_1807);
  not gc183 (wc183, n_1899);
  and g2436 (n_1914, wc184, n_1830);
  not gc184 (wc184, n_1909);
  and g2437 (n_1963, wc185, n_1800);
  not gc185 (wc185, n_1957);
  and g2438 (n_1976, wc186, n_1973);
  not gc186 (wc186, n_1957);
  and g2439 (n_1981, wc187, n_1978);
  not gc187 (wc187, n_1957);
  and g2440 (n_1986, wc188, n_1983);
  not gc188 (wc188, n_1957);
  and g2441 (n_1991, wc189, n_1988);
  not gc189 (wc189, n_1957);
  or g2442 (n_2059, n_2056, wc190);
  not gc190 (wc190, n_2024);
  or g2443 (n_2063, n_2060, wc191);
  not gc191 (wc191, n_2024);
  and g2444 (n_1985, n_1902, wc192);
  not gc192 (wc192, n_1903);
  and g2445 (n_1990, n_1906, wc193);
  not gc193 (wc193, n_1907);
  and g2446 (n_2087, wc194, n_1707);
  not gc194 (wc194, n_1910);
  and g2447 (n_2090, wc195, n_1827);
  not gc195 (wc195, n_1914);
  and g2448 (n_2093, n_1917, wc196);
  not gc196 (wc196, n_1918);
  and g2449 (n_1993, n_1921, wc197);
  not gc197 (wc197, n_1922);
  and g2450 (n_2046, wc198, n_1671);
  not gc198 (wc198, n_1958);
  and g2451 (n_2050, wc199, n_1797);
  not gc199 (wc199, n_1963);
  and g2452 (n_2054, n_1966, wc200);
  not gc200 (wc200, n_1967);
  and g2453 (n_2058, n_1894, wc201);
  not gc201 (wc201, n_1970);
  or g2454 (n_2067, n_2064, wc202);
  not gc202 (wc202, n_2024);
  or g2455 (n_2071, n_2068, wc203);
  not gc203 (wc203, n_2024);
  or g2456 (n_2075, n_2072, wc204);
  not gc204 (wc204, n_2024);
  and g2457 (n_2062, wc205, n_1975);
  not gc205 (wc205, n_1976);
  and g2458 (n_2066, wc206, n_1980);
  not gc206 (wc206, n_1981);
  and g2459 (n_1999, wc207, n_1840);
  not gc207 (wc207, n_1993);
  and g2460 (n_2012, wc208, n_2009);
  not gc208 (wc208, n_1993);
  and g2461 (n_2017, wc209, n_2014);
  not gc209 (wc209, n_1993);
  and g2462 (n_2022, wc210, n_2019);
  not gc210 (wc210, n_1993);
  and g2463 (n_2070, n_1985, wc211);
  not gc211 (wc211, n_1986);
  and g2464 (n_2074, n_1990, wc212);
  not gc212 (wc212, n_1991);
  and g2465 (n_2098, wc213, n_1719);
  not gc213 (wc213, n_1994);
  and g2466 (n_2102, wc214, n_1837);
  not gc214 (wc214, n_1999);
  and g2467 (n_2106, n_2002, wc215);
  not gc215 (wc215, n_2003);
  and g2468 (n_2110, n_1924, wc216);
  not gc216 (wc216, n_2006);
  and g2469 (n_2114, wc217, n_2011);
  not gc217 (wc217, n_2012);
  and g2470 (n_2118, wc218, n_2016);
  not gc218 (wc218, n_2017);
  and g2471 (n_2122, wc219, n_2021);
  not gc219 (wc219, n_2022);
  or g2472 (n_2078, wc220, n_1700);
  not gc220 (wc220, n_2076);
  or g2473 (n_2083, n_2080, wc221);
  not gc221 (wc221, n_2076);
  or g2474 (n_2085, wc222, n_1912);
  not gc222 (wc222, n_2076);
  or g2475 (n_2099, n_2096, wc223);
  not gc223 (wc223, n_2076);
  or g2476 (n_2103, wc224, n_2100);
  not gc224 (wc224, n_2076);
  or g2477 (n_2107, n_2104, wc225);
  not gc225 (wc225, n_2076);
  or g2478 (n_2111, n_2108, wc226);
  not gc226 (wc226, n_2076);
  or g2479 (n_2115, wc227, n_2112);
  not gc227 (wc227, n_2076);
  or g2480 (n_2119, wc228, n_2116);
  not gc228 (wc228, n_2076);
  or g2481 (n_2123, wc229, n_2120);
  not gc229 (wc229, n_2076);
endmodule

module mult_signed_const_4418_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_4418_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_4685_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_176;
  wire n_178, n_179, n_180, n_183, n_184, n_187, n_188, n_189;
  wire n_195, n_196, n_200, n_201, n_202, n_203, n_204, n_207;
  wire n_209, n_210, n_211, n_212, n_217, n_218, n_219, n_220;
  wire n_221, n_223, n_224, n_225, n_226, n_227, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_251, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_265, n_268, n_270, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_280, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_298, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_306, n_307, n_308, n_309, n_317, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_336, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_349, n_351, n_353, n_356, n_357, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_371;
  wire n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_390, n_392, n_393, n_394, n_395, n_396;
  wire n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404;
  wire n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412;
  wire n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420;
  wire n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_489, n_490, n_491;
  wire n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499;
  wire n_500, n_504, n_505, n_506, n_507, n_508, n_509, n_510;
  wire n_511, n_512, n_513, n_514, n_515, n_519, n_520, n_521;
  wire n_522, n_523, n_524, n_525, n_526, n_527, n_528, n_529;
  wire n_530, n_532, n_533, n_534, n_535, n_536, n_537, n_538;
  wire n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_557, n_558, n_559, n_560, n_561, n_562, n_563, n_564;
  wire n_565, n_569, n_570, n_571, n_572, n_573, n_574, n_575;
  wire n_576, n_578, n_579, n_580, n_581, n_582, n_583, n_584;
  wire n_585, n_586, n_588, n_589, n_590, n_591, n_592, n_596;
  wire n_598, n_599, n_604, n_605, n_606, n_608, n_609, n_610;
  wire n_611, n_612, n_614, n_622, n_623, n_624, n_625, n_626;
  wire n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634;
  wire n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642;
  wire n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675;
  wire n_676, n_677, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_698, n_699, n_700, n_702;
  wire n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710;
  wire n_711, n_712, n_713, n_722, n_723, n_724, n_725, n_726;
  wire n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_738;
  wire n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749;
  wire n_750, n_751, n_752, n_753, n_760, n_761, n_762, n_763;
  wire n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772;
  wire n_773, n_774, n_775, n_776, n_777, n_788, n_789, n_790;
  wire n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798;
  wire n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_814;
  wire n_815, n_818, n_819, n_820, n_821, n_822, n_823, n_824;
  wire n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832;
  wire n_833, n_842, n_846, n_847, n_848, n_849, n_850, n_851;
  wire n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859;
  wire n_860, n_861, n_864, n_865, n_866, n_867, n_868, n_869;
  wire n_873, n_874, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_902, n_903, n_904, n_905;
  wire n_906, n_907, n_908, n_909, n_910, n_911, n_912, n_913;
  wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
  wire n_922, n_923, n_924, n_925, n_926, n_927, n_928, n_929;
  wire n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951;
  wire n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959;
  wire n_960, n_961, n_962, n_963, n_964, n_965, n_978, n_982;
  wire n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990;
  wire n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998;
  wire n_999, n_1000, n_1001, n_1014, n_1022, n_1023, n_1024, n_1025;
  wire n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033;
  wire n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041;
  wire n_1042, n_1044, n_1045, n_1046, n_1047, n_1048, n_1050, n_1051;
  wire n_1052, n_1053, n_1054, n_1056, n_1057, n_1058, n_1059, n_1060;
  wire n_1061, n_1062, n_1063, n_1064, n_1066, n_1067, n_1068, n_1069;
  wire n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077;
  wire n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085;
  wire n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093;
  wire n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1101, n_1102;
  wire n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110;
  wire n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118;
  wire n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126;
  wire n_1127, n_1128, n_1129, n_1132, n_1133, n_1134, n_1135, n_1136;
  wire n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1144, n_1145;
  wire n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153;
  wire n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161;
  wire n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169;
  wire n_1170, n_1171, n_1172, n_1173, n_1174, n_1176, n_1177, n_1178;
  wire n_1179, n_1180, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187;
  wire n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195;
  wire n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205;
  wire n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213;
  wire n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221;
  wire n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229;
  wire n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237;
  wire n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
  wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1252, n_1253, n_1254;
  wire n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1262, n_1263;
  wire n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271;
  wire n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279;
  wire n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1288;
  wire n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299;
  wire n_1301, n_1302, n_1303, n_1305, n_1306, n_1307, n_1308, n_1309;
  wire n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317;
  wire n_1318, n_1319, n_1320, n_1321, n_1326, n_1327, n_1328, n_1329;
  wire n_1330, n_1331, n_1333, n_1334, n_1335, n_1336, n_1337, n_1340;
  wire n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348;
  wire n_1349, n_1350, n_1351, n_1352, n_1353, n_1355, n_1356, n_1357;
  wire n_1358, n_1360, n_1361, n_1362, n_1363, n_1364, n_1366, n_1367;
  wire n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375;
  wire n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1385, n_1386;
  wire n_1388, n_1389, n_1390, n_1392, n_1393, n_1394, n_1395, n_1396;
  wire n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405;
  wire n_1406, n_1407, n_1408, n_1409, n_1413, n_1414, n_1415, n_1416;
  wire n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1424, n_1425;
  wire n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433;
  wire n_1434, n_1435, n_1436, n_1437, n_1438, n_1440, n_1441, n_1445;
  wire n_1446, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454;
  wire n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1463;
  wire n_1464, n_1466, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474;
  wire n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1485;
  wire n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
  wire n_1498, n_1499, n_1500, n_1501, n_1504, n_1506, n_1507, n_1508;
  wire n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519;
  wire n_1520, n_1521, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533;
  wire n_1534, n_1535, n_1536, n_1537, n_1542, n_1543, n_1544, n_1545;
  wire n_1546, n_1547, n_1548, n_1549, n_1550, n_1553, n_1555, n_1556;
  wire n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1565, n_1566;
  wire n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1578;
  wire n_1579, n_1580, n_1581, n_1583, n_1584, n_1585, n_1587, n_1588;
  wire n_1590, n_1591, n_1593, n_1604, n_1605, n_1606, n_1607, n_1609;
  wire n_1610, n_1611, n_1612, n_1613, n_1615, n_1616, n_1617, n_1618;
  wire n_1619, n_1621, n_1622, n_1623, n_1624, n_1625, n_1627, n_1628;
  wire n_1629, n_1630, n_1631, n_1633, n_1634, n_1635, n_1636, n_1637;
  wire n_1639, n_1640, n_1641, n_1642, n_1643, n_1645, n_1646, n_1647;
  wire n_1648, n_1649, n_1651, n_1652, n_1653, n_1654, n_1655, n_1657;
  wire n_1658, n_1659, n_1660, n_1661, n_1663, n_1664, n_1665, n_1666;
  wire n_1667, n_1669, n_1670, n_1671, n_1672, n_1673, n_1675, n_1676;
  wire n_1677, n_1678, n_1679, n_1681, n_1682, n_1683, n_1684, n_1685;
  wire n_1687, n_1688, n_1689, n_1690, n_1691, n_1693, n_1694, n_1695;
  wire n_1696, n_1697, n_1699, n_1700, n_1701, n_1702, n_1703, n_1705;
  wire n_1706, n_1707, n_1708, n_1709, n_1711, n_1712, n_1713, n_1714;
  wire n_1715, n_1717, n_1718, n_1719, n_1720, n_1721, n_1723, n_1724;
  wire n_1725, n_1726, n_1727, n_1729, n_1730, n_1731, n_1732, n_1733;
  wire n_1735, n_1736, n_1737, n_1738, n_1739, n_1744, n_1746, n_1747;
  wire n_1749, n_1751, n_1753, n_1754, n_1756, n_1757, n_1759, n_1761;
  wire n_1763, n_1764, n_1766, n_1767, n_1769, n_1771, n_1773, n_1774;
  wire n_1776, n_1777, n_1779, n_1781, n_1783, n_1784, n_1786, n_1787;
  wire n_1789, n_1791, n_1793, n_1794, n_1796, n_1797, n_1799, n_1801;
  wire n_1803, n_1804, n_1806, n_1807, n_1809, n_1811, n_1813, n_1814;
  wire n_1816, n_1817, n_1819, n_1821, n_1823, n_1824, n_1826, n_1827;
  wire n_1829, n_1831, n_1833, n_1834, n_1836, n_1837, n_1839, n_1841;
  wire n_1843, n_1844, n_1846, n_1847, n_1849, n_1853, n_1854, n_1855;
  wire n_1857, n_1858, n_1859, n_1861, n_1862, n_1863, n_1864, n_1866;
  wire n_1868, n_1870, n_1871, n_1872, n_1874, n_1875, n_1876, n_1878;
  wire n_1879, n_1881, n_1883, n_1885, n_1886, n_1887, n_1889, n_1890;
  wire n_1891, n_1893, n_1894, n_1896, n_1898, n_1900, n_1901, n_1902;
  wire n_1904, n_1905, n_1906, n_1908, n_1909, n_1911, n_1913, n_1915;
  wire n_1916, n_1917, n_1919, n_1920, n_1921, n_1923, n_1924, n_1926;
  wire n_1928, n_1930, n_1931, n_1932, n_1934, n_1936, n_1937, n_1938;
  wire n_1940, n_1941, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948;
  wire n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956;
  wire n_1957, n_1959, n_1962, n_1964, n_1965, n_1966, n_1969, n_1972;
  wire n_1974, n_1975, n_1977, n_1979, n_1980, n_1982, n_1984, n_1985;
  wire n_1987, n_1989, n_1990, n_1992, n_1993, n_1995, n_1998, n_2000;
  wire n_2001, n_2002, n_2005, n_2008, n_2010, n_2011, n_2013, n_2015;
  wire n_2016, n_2018, n_2020, n_2021, n_2023, n_2025, n_2026, n_2027;
  wire n_2029, n_2030, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037;
  wire n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2045, n_2046;
  wire n_2047, n_2049, n_2050, n_2051, n_2053, n_2054, n_2055, n_2057;
  wire n_2058, n_2059, n_2061, n_2062, n_2063, n_2065, n_2066, n_2067;
  wire n_2069, n_2070, n_2071, n_2073, n_2074, n_2075, n_2077, n_2078;
  wire n_2079, n_2081, n_2082, n_2084, n_2085, n_2086, n_2087, n_2088;
  wire n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2097;
  wire n_2098, n_2099, n_2101, n_2102, n_2103, n_2105, n_2106, n_2107;
  wire n_2109, n_2110, n_2111, n_2113, n_2114, n_2115, n_2117, n_2118;
  wire n_2119, n_2121, n_2122, n_2124, n_2127, n_2128, n_2130, n_2131;
  wire n_2132, n_2133, n_2135, n_2136, n_2137, n_2139, n_2140, n_2141;
  wire n_2142, n_2144, n_2145, n_2147, n_2148, n_2150, n_2151, n_2152;
  wire n_2153, n_2155, n_2156, n_2157, n_2159, n_2160, n_2161, n_2162;
  wire n_2164, n_2165, n_2167, n_2168, n_2170, n_2171, n_2172, n_2173;
  wire n_2175, n_2176, n_2177, n_2178, n_2180, n_2181, n_2182, n_2183;
  wire n_2185, n_2186, n_2188, n_2189, n_2191, n_2192, n_2193, n_2194;
  wire n_2196, n_2197, n_2198, n_2200, n_2201, n_2202, n_2203, n_2205;
  wire n_2206, n_2208, n_2209, n_2211, n_2212, n_2213, n_2214, n_2216;
  wire n_2217, n_2218, n_2219, n_2221, n_2222, n_2223, n_2224, n_2226;
  wire n_2227, n_2229, n_2230, n_2232, n_2233, n_2234, n_2235, n_2237;
  wire n_2238;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], n_171);
  xor g270 (n_117, n_622, A[2]);
  nand g3 (n_623, A[1], n_171);
  nand g271 (n_624, A[2], n_171);
  nand g272 (n_625, A[1], A[2]);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, A[4]);
  xor g288 (n_176, n_634, n_69);
  nand g289 (n_635, n_68, A[4]);
  nand g290 (n_636, n_69, A[4]);
  nand g291 (n_637, n_68, n_69);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_176);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_176);
  nand g296 (n_640, A[7], n_176);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g299 (n_642, A[1], A[2]);
  xor g300 (n_178, n_642, n_171);
  xor g305 (n_646, A[5], n_178);
  xor g306 (n_180, n_646, A[6]);
  nand g307 (n_647, A[5], n_178);
  nand g308 (n_648, A[6], n_178);
  nand g309 (n_649, A[5], A[6]);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, n_179, n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, n_179, n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, n_179, A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_188, n_659, n_660, n_661);
  xor g329 (n_662, n_183, n_184);
  xor g330 (n_112, n_662, A[9]);
  nand g331 (n_663, n_183, n_184);
  nand g332 (n_664, A[9], n_184);
  nand g333 (n_665, n_183, A[9]);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_187, n_630, n_67);
  nand g340 (n_668, n_67, n_173);
  nand g341 (n_669, A[4], n_67);
  nand g342 (n_71, n_631, n_668, n_669);
  xor g343 (n_670, A[7], n_187);
  xor g344 (n_189, n_670, A[8]);
  nand g345 (n_671, A[7], n_187);
  nand g346 (n_672, A[8], n_187);
  nand g347 (n_673, A[7], A[8]);
  nand g348 (n_73, n_671, n_672, n_673);
  xor g349 (n_674, A[10], n_188);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, A[10], n_188);
  nand g352 (n_676, n_189, n_188);
  nand g353 (n_677, A[10], n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_195, n_638, A[8]);
  nand g366 (n_684, A[8], n_176);
  nand g367 (n_685, A[5], A[8]);
  nand g368 (n_201, n_639, n_684, n_685);
  xor g369 (n_686, n_71, A[9]);
  xor g370 (n_196, n_686, A[11]);
  nand g371 (n_687, n_71, A[9]);
  nand g372 (n_688, A[11], A[9]);
  nand g373 (n_689, n_71, A[11]);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, n_73, n_195);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, n_73, n_195);
  nand g378 (n_692, n_196, n_195);
  nand g379 (n_693, n_73, n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g387 (n_698, A[5], n_117);
  xor g388 (n_200, n_698, A[6]);
  nand g389 (n_699, A[5], n_117);
  nand g390 (n_700, A[6], n_117);
  nand g392 (n_207, n_699, n_700, n_649);
  xor g393 (n_702, n_179, n_200);
  xor g394 (n_202, n_702, A[10]);
  nand g395 (n_703, n_179, n_200);
  nand g396 (n_704, A[10], n_200);
  nand g397 (n_705, n_179, A[10]);
  nand g398 (n_209, n_703, n_704, n_705);
  xor g399 (n_706, A[9], A[12]);
  xor g400 (n_204, n_706, n_201);
  nand g401 (n_707, A[9], A[12]);
  nand g402 (n_708, n_201, A[12]);
  nand g403 (n_709, A[9], n_201);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, n_202, n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, n_202, n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, n_202, n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g423 (n_722, n_207, A[10]);
  xor g424 (n_210, n_722, n_184);
  nand g425 (n_723, n_207, A[10]);
  nand g426 (n_724, n_184, A[10]);
  nand g427 (n_725, n_207, n_184);
  nand g428 (n_217, n_723, n_724, n_725);
  xor g429 (n_726, A[11], A[13]);
  xor g430 (n_212, n_726, n_209);
  nand g431 (n_727, A[11], A[13]);
  nand g432 (n_728, n_209, A[13]);
  nand g433 (n_729, A[11], n_209);
  nand g434 (n_220, n_727, n_728, n_729);
  xor g435 (n_730, n_210, n_211);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, n_210, n_211);
  nand g438 (n_732, n_212, n_211);
  nand g439 (n_733, n_210, n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_218, n_738, n_187);
  xor g455 (n_742, n_188, A[12]);
  xor g456 (n_219, n_742, A[11]);
  nand g457 (n_743, n_188, A[12]);
  nand g458 (n_744, A[11], A[12]);
  nand g459 (n_745, n_188, A[11]);
  nand g460 (n_224, n_743, n_744, n_745);
  xor g461 (n_746, A[14], n_217);
  xor g462 (n_221, n_746, n_218);
  nand g463 (n_747, A[14], n_217);
  nand g464 (n_748, n_218, n_217);
  nand g465 (n_749, A[14], n_218);
  nand g466 (n_225, n_747, n_748, n_749);
  xor g467 (n_750, n_219, n_220);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, n_219, n_220);
  nand g470 (n_752, n_221, n_220);
  nand g471 (n_753, n_219, n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g482 (n_72, n_638, n_71);
  nand g484 (n_760, n_71, n_176);
  nand g485 (n_761, A[5], n_71);
  nand g486 (n_232, n_639, n_760, n_761);
  xor g487 (n_762, A[8], A[9]);
  xor g488 (n_223, n_762, A[12]);
  nand g489 (n_763, A[8], A[9]);
  nand g491 (n_765, A[8], A[12]);
  nand g492 (n_234, n_763, n_707, n_765);
  xor g493 (n_766, n_72, A[13]);
  xor g494 (n_226, n_766, n_73);
  nand g495 (n_767, n_72, A[13]);
  nand g496 (n_768, n_73, A[13]);
  nand g497 (n_769, n_72, n_73);
  nand g498 (n_235, n_767, n_768, n_769);
  xor g499 (n_770, A[15], n_223);
  xor g500 (n_227, n_770, n_224);
  nand g501 (n_771, A[15], n_223);
  nand g502 (n_772, n_224, n_223);
  nand g503 (n_773, A[15], n_224);
  nand g504 (n_237, n_771, n_772, n_773);
  xor g505 (n_774, n_225, n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, n_225, n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, n_225, n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g524 (n_233, n_650, A[9]);
  nand g526 (n_788, A[9], n_180);
  nand g527 (n_789, n_179, A[9]);
  nand g528 (n_244, n_651, n_788, n_789);
  xor g529 (n_790, A[10], n_232);
  xor g530 (n_236, n_790, A[14]);
  nand g531 (n_791, A[10], n_232);
  nand g532 (n_792, A[14], n_232);
  nand g533 (n_793, A[10], A[14]);
  nand g534 (n_246, n_791, n_792, n_793);
  xor g535 (n_794, A[13], n_233);
  xor g536 (n_238, n_794, n_234);
  nand g537 (n_795, A[13], n_233);
  nand g538 (n_796, n_234, n_233);
  nand g539 (n_797, A[13], n_234);
  nand g540 (n_248, n_795, n_796, n_797);
  xor g541 (n_798, A[16], n_235);
  xor g542 (n_239, n_798, n_236);
  nand g543 (n_799, A[16], n_235);
  nand g544 (n_800, n_236, n_235);
  nand g545 (n_801, A[16], n_236);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, n_237, n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, n_237, n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, n_237, n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g565 (n_814, n_183, A[10]);
  xor g566 (n_245, n_814, n_184);
  nand g567 (n_815, n_183, A[10]);
  nand g570 (n_257, n_815, n_724, n_663);
  xor g571 (n_818, A[11], A[14]);
  xor g572 (n_247, n_818, n_244);
  nand g573 (n_819, A[11], A[14]);
  nand g574 (n_820, n_244, A[14]);
  nand g575 (n_821, A[11], n_244);
  nand g576 (n_259, n_819, n_820, n_821);
  xor g577 (n_822, A[15], n_245);
  xor g578 (n_249, n_822, n_246);
  nand g579 (n_823, A[15], n_245);
  nand g580 (n_824, n_246, n_245);
  nand g581 (n_825, A[15], n_246);
  nand g582 (n_261, n_823, n_824, n_825);
  xor g583 (n_826, n_247, A[17]);
  xor g584 (n_251, n_826, n_248);
  nand g585 (n_827, n_247, A[17]);
  nand g586 (n_828, n_248, A[17]);
  nand g587 (n_829, n_247, n_248);
  nand g588 (n_118, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g609 (n_842, n_188, A[11]);
  xor g610 (n_258, n_842, A[12]);
  xor g615 (n_846, n_218, A[15]);
  xor g616 (n_260, n_846, n_257);
  nand g617 (n_847, n_218, A[15]);
  nand g618 (n_848, n_257, A[15]);
  nand g619 (n_849, n_218, n_257);
  nand g620 (n_272, n_847, n_848, n_849);
  xor g621 (n_850, n_258, A[16]);
  xor g622 (n_262, n_850, A[18]);
  nand g623 (n_851, n_258, A[16]);
  nand g624 (n_852, A[18], A[16]);
  nand g625 (n_853, n_258, A[18]);
  nand g626 (n_274, n_851, n_852, n_853);
  xor g627 (n_854, n_259, n_260);
  xor g628 (n_119, n_854, n_261);
  nand g629 (n_855, n_259, n_260);
  nand g630 (n_856, n_261, n_260);
  nand g631 (n_857, n_259, n_261);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_262, n_118);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_262, n_118);
  nand g636 (n_860, n_119, n_118);
  nand g637 (n_861, n_262, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g642 (n_265, n_634, A[5]);
  nand g644 (n_864, A[5], A[4]);
  nand g645 (n_865, n_68, A[5]);
  nand g646 (n_280, n_635, n_864, n_865);
  xor g647 (n_866, n_69, n_265);
  xor g648 (n_268, n_866, A[8]);
  nand g649 (n_867, n_69, n_265);
  nand g650 (n_868, A[8], n_265);
  nand g651 (n_869, n_69, A[8]);
  nand g652 (n_282, n_867, n_868, n_869);
  xor g654 (n_270, n_686, A[12]);
  nand g657 (n_873, n_71, A[12]);
  nand g658 (n_284, n_687, n_707, n_873);
  xor g659 (n_874, A[13], n_73);
  xor g660 (n_271, n_874, n_268);
  nand g662 (n_876, n_268, n_73);
  nand g663 (n_877, A[13], n_268);
  nand g664 (n_285, n_768, n_876, n_877);
  xor g665 (n_878, n_224, n_270);
  xor g666 (n_273, n_878, A[16]);
  nand g667 (n_879, n_224, n_270);
  nand g668 (n_880, A[16], n_270);
  nand g669 (n_881, n_224, A[16]);
  nand g670 (n_288, n_879, n_880, n_881);
  xor g671 (n_882, A[19], A[17]);
  xor g672 (n_275, n_882, n_271);
  nand g673 (n_883, A[19], A[17]);
  nand g674 (n_884, n_271, A[17]);
  nand g675 (n_885, A[19], n_271);
  nand g676 (n_289, n_883, n_884, n_885);
  xor g677 (n_886, n_272, n_273);
  xor g678 (n_277, n_886, n_274);
  nand g679 (n_887, n_272, n_273);
  nand g680 (n_888, n_274, n_273);
  nand g681 (n_889, n_272, n_274);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g701 (n_902, n_280, n_180);
  xor g702 (n_283, n_902, A[10]);
  nand g703 (n_903, n_280, n_180);
  nand g704 (n_904, A[10], n_180);
  nand g705 (n_905, n_280, A[10]);
  nand g706 (n_298, n_903, n_904, n_905);
  xor g707 (n_906, A[9], A[13]);
  xor g708 (n_286, n_906, n_282);
  nand g709 (n_907, A[9], A[13]);
  nand g710 (n_908, n_282, A[13]);
  nand g711 (n_909, A[9], n_282);
  nand g712 (n_300, n_907, n_908, n_909);
  xor g713 (n_910, A[14], n_283);
  xor g714 (n_287, n_910, n_284);
  nand g715 (n_911, A[14], n_283);
  nand g716 (n_912, n_284, n_283);
  nand g717 (n_913, A[14], n_284);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, n_285, A[18]);
  xor g720 (n_290, n_914, A[17]);
  nand g721 (n_915, n_285, A[18]);
  nand g722 (n_916, A[17], A[18]);
  nand g723 (n_917, n_285, A[17]);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, n_286, A[20]);
  xor g726 (n_291, n_918, n_287);
  nand g727 (n_919, n_286, A[20]);
  nand g728 (n_920, n_287, A[20]);
  nand g729 (n_921, n_286, n_287);
  nand g730 (n_305, n_919, n_920, n_921);
  xor g731 (n_922, n_288, n_289);
  xor g732 (n_293, n_922, n_290);
  nand g733 (n_923, n_288, n_289);
  nand g734 (n_924, n_290, n_289);
  nand g735 (n_925, n_288, n_290);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g762 (n_301, n_818, A[15]);
  nand g764 (n_944, A[15], A[14]);
  nand g765 (n_945, A[11], A[15]);
  nand g766 (n_317, n_819, n_944, n_945);
  xor g767 (n_946, n_298, n_245);
  xor g768 (n_303, n_946, n_300);
  nand g769 (n_947, n_298, n_245);
  nand g770 (n_948, n_300, n_245);
  nand g771 (n_949, n_298, n_300);
  nand g772 (n_319, n_947, n_948, n_949);
  xor g773 (n_950, A[19], n_301);
  xor g774 (n_306, n_950, A[18]);
  nand g775 (n_951, A[19], n_301);
  nand g776 (n_952, A[18], n_301);
  nand g777 (n_953, A[19], A[18]);
  nand g778 (n_321, n_951, n_952, n_953);
  xor g779 (n_954, A[21], n_302);
  xor g780 (n_307, n_954, n_303);
  nand g781 (n_955, A[21], n_302);
  nand g782 (n_956, n_303, n_302);
  nand g783 (n_957, A[21], n_303);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, n_304, n_305);
  xor g786 (n_309, n_958, n_306);
  nand g787 (n_959, n_304, n_305);
  nand g788 (n_960, n_306, n_305);
  nand g789 (n_961, n_304, n_306);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g817 (n_978, n_218, n_257);
  xor g818 (n_318, n_978, A[15]);
  xor g823 (n_982, A[16], n_219);
  xor g824 (n_320, n_982, n_317);
  nand g825 (n_983, A[16], n_219);
  nand g826 (n_984, n_317, n_219);
  nand g827 (n_985, A[16], n_317);
  nand g828 (n_338, n_983, n_984, n_985);
  xor g829 (n_986, A[19], A[22]);
  xor g830 (n_322, n_986, n_318);
  nand g831 (n_987, A[19], A[22]);
  nand g832 (n_988, n_318, A[22]);
  nand g833 (n_989, A[19], n_318);
  nand g834 (n_339, n_987, n_988, n_989);
  xor g835 (n_990, A[20], n_319);
  xor g836 (n_324, n_990, n_320);
  nand g837 (n_991, A[20], n_319);
  nand g838 (n_992, n_320, n_319);
  nand g839 (n_993, A[20], n_320);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, n_321, n_322);
  xor g842 (n_326, n_994, n_323);
  nand g843 (n_995, n_321, n_322);
  nand g844 (n_996, n_323, n_322);
  nand g845 (n_997, n_321, n_323);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, n_324, n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, n_324, n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, n_324, n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g873 (n_1014, n_73, n_268);
  xor g874 (n_336, n_1014, A[13]);
  xor g885 (n_1022, A[17], n_272);
  xor g886 (n_340, n_1022, n_336);
  nand g887 (n_1023, A[17], n_272);
  nand g888 (n_1024, n_336, n_272);
  nand g889 (n_1025, A[17], n_336);
  nand g890 (n_359, n_1023, n_1024, n_1025);
  xor g891 (n_1026, A[21], A[20]);
  xor g892 (n_341, n_1026, A[23]);
  nand g893 (n_1027, A[21], A[20]);
  nand g894 (n_1028, A[23], A[20]);
  nand g895 (n_1029, A[21], A[23]);
  nand g896 (n_361, n_1027, n_1028, n_1029);
  xor g897 (n_1030, n_273, n_338);
  xor g898 (n_343, n_1030, n_339);
  nand g899 (n_1031, n_273, n_338);
  nand g900 (n_1032, n_339, n_338);
  nand g901 (n_1033, n_273, n_339);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, n_340, n_341);
  xor g904 (n_345, n_1034, n_342);
  nand g905 (n_1035, n_340, n_341);
  nand g906 (n_1036, n_342, n_341);
  nand g907 (n_1037, n_340, n_342);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, n_343, n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, n_343, n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, n_343, n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  xor g917 (n_1042, A[2], n_171);
  nand g922 (n_371, n_624, n_1044, n_1045);
  xor g923 (n_1046, A[5], n_349);
  xor g924 (n_351, n_1046, A[6]);
  nand g925 (n_1047, A[5], n_349);
  nand g926 (n_1048, A[6], n_349);
  nand g928 (n_373, n_1047, n_1048, n_649);
  xor g929 (n_1050, n_280, n_351);
  xor g930 (n_353, n_1050, A[9]);
  nand g931 (n_1051, n_280, n_351);
  nand g932 (n_1052, A[9], n_351);
  nand g933 (n_1053, n_280, A[9]);
  nand g934 (n_375, n_1051, n_1052, n_1053);
  xor g935 (n_1054, A[10], A[14]);
  xor g936 (n_356, n_1054, n_282);
  nand g938 (n_1056, n_282, A[14]);
  nand g939 (n_1057, A[10], n_282);
  nand g940 (n_377, n_793, n_1056, n_1057);
  xor g941 (n_1058, A[13], n_353);
  xor g942 (n_357, n_1058, n_284);
  nand g943 (n_1059, A[13], n_353);
  nand g944 (n_1060, n_284, n_353);
  nand g945 (n_1061, A[13], n_284);
  nand g946 (n_379, n_1059, n_1060, n_1061);
  xor g947 (n_1062, n_285, n_356);
  xor g948 (n_360, n_1062, A[17]);
  nand g949 (n_1063, n_285, n_356);
  nand g950 (n_1064, A[17], n_356);
  nand g952 (n_381, n_1063, n_1064, n_917);
  xor g953 (n_1066, A[18], n_357);
  nand g955 (n_1067, A[18], n_357);
  nand g958 (n_383, n_1067, n_1068, n_1069);
  xor g959 (n_1070, A[21], A[22]);
  xor g960 (n_362, n_1070, n_288);
  nand g961 (n_1071, A[21], A[22]);
  nand g962 (n_1072, n_288, A[22]);
  nand g963 (n_1073, A[21], n_288);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, n_359, n_360);
  xor g966 (n_365, n_1074, n_361);
  nand g967 (n_1075, n_359, n_360);
  nand g968 (n_1076, n_361, n_360);
  nand g969 (n_1077, n_359, n_361);
  nand g970 (n_388, n_1075, n_1076, n_1077);
  xor g971 (n_1078, n_362, n_363);
  xor g972 (n_367, n_1078, n_364);
  nand g973 (n_1079, n_362, n_363);
  nand g974 (n_1080, n_364, n_363);
  nand g975 (n_1081, n_362, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  xor g985 (n_1086, A[1], A[3]);
  nand g987 (n_1087, A[1], A[3]);
  nand g990 (n_392, n_1087, n_1088, n_1089);
  xor g991 (n_1090, n_371, A[6]);
  xor g992 (n_374, n_1090, n_372);
  nand g993 (n_1091, n_371, A[6]);
  nand g994 (n_1092, n_372, A[6]);
  nand g995 (n_1093, n_371, n_372);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, A[10]);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, A[10], n_373);
  nand g1001 (n_1097, A[7], A[10]);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, n_374, A[11]);
  xor g1004 (n_378, n_1098, A[14]);
  nand g1005 (n_1099, n_374, A[11]);
  nand g1007 (n_1101, n_374, A[14]);
  nand g1008 (n_398, n_1099, n_819, n_1101);
  xor g1009 (n_1102, n_375, n_376);
  xor g1010 (n_380, n_1102, A[15]);
  nand g1011 (n_1103, n_375, n_376);
  nand g1012 (n_1104, A[15], n_376);
  nand g1013 (n_1105, n_375, A[15]);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, n_377, n_378);
  xor g1016 (n_382, n_1106, A[19]);
  nand g1017 (n_1107, n_377, n_378);
  nand g1018 (n_1108, A[19], n_378);
  nand g1019 (n_1109, n_377, A[19]);
  nand g1020 (n_402, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, A[18], n_379);
  xor g1022 (n_384, n_1110, A[22]);
  nand g1023 (n_1111, A[18], n_379);
  nand g1024 (n_1112, A[22], n_379);
  nand g1025 (n_1113, A[18], A[22]);
  nand g1026 (n_403, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, n_380, A[23]);
  xor g1028 (n_386, n_1114, n_381);
  nand g1029 (n_1115, n_380, A[23]);
  nand g1030 (n_1116, n_381, A[23]);
  nand g1031 (n_1117, n_380, n_381);
  nand g1032 (n_407, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_382, n_383);
  xor g1034 (n_387, n_1118, n_384);
  nand g1035 (n_1119, n_382, n_383);
  nand g1036 (n_1120, n_384, n_383);
  nand g1037 (n_1121, n_382, n_384);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, n_385, n_386);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, n_385, n_386);
  nand g1042 (n_1124, n_387, n_386);
  nand g1043 (n_1125, n_385, n_387);
  nand g1044 (n_411, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1052 (n_393, n_626, A[4]);
  nand g1054 (n_1132, A[4], A[2]);
  nand g1055 (n_1133, A[3], A[4]);
  nand g1056 (n_412, n_627, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, A[11], A[12]);
  xor g1070 (n_399, n_1142, n_396);
  nand g1072 (n_1144, n_396, A[12]);
  nand g1073 (n_1145, A[11], n_396);
  nand g1074 (n_418, n_744, n_1144, n_1145);
  xor g1075 (n_1146, n_397, A[15]);
  xor g1076 (n_401, n_1146, n_398);
  nand g1077 (n_1147, n_397, A[15]);
  nand g1078 (n_1148, n_398, A[15]);
  nand g1079 (n_1149, n_397, n_398);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, A[16], A[19]);
  xor g1082 (n_404, n_1150, n_399);
  nand g1083 (n_1151, A[16], A[19]);
  nand g1084 (n_1152, n_399, A[19]);
  nand g1085 (n_1153, A[16], n_399);
  nand g1086 (n_421, n_1151, n_1152, n_1153);
  xor g1088 (n_405, n_1154, A[20]);
  nand g1091 (n_1157, n_400, A[20]);
  nand g1092 (n_422, n_1155, n_1156, n_1157);
  xor g1093 (n_1158, n_401, A[23]);
  xor g1094 (n_406, n_1158, n_402);
  nand g1095 (n_1159, n_401, A[23]);
  nand g1096 (n_1160, n_402, A[23]);
  nand g1097 (n_1161, n_401, n_402);
  nand g1098 (n_425, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_403, n_404);
  xor g1100 (n_409, n_1162, n_405);
  nand g1101 (n_1163, n_403, n_404);
  nand g1102 (n_1164, n_405, n_404);
  nand g1103 (n_1165, n_403, n_405);
  nand g1104 (n_427, n_1163, n_1164, n_1165);
  xor g1105 (n_1166, n_406, n_407);
  xor g1106 (n_410, n_1166, n_408);
  nand g1107 (n_1167, n_406, n_407);
  nand g1108 (n_1168, n_408, n_407);
  nand g1109 (n_1169, n_406, n_408);
  nand g1110 (n_430, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_864, n_1176, n_1177);
  xor g1123 (n_1178, A[8], n_413);
  xor g1124 (n_415, n_1178, A[9]);
  nand g1125 (n_1179, A[8], n_413);
  nand g1126 (n_1180, A[9], n_413);
  nand g1128 (n_435, n_1179, n_1180, n_763);
  xor g1129 (n_1182, n_414, A[12]);
  xor g1130 (n_417, n_1182, A[13]);
  nand g1131 (n_1183, n_414, A[12]);
  nand g1132 (n_1184, A[13], A[12]);
  nand g1133 (n_1185, n_414, A[13]);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, n_415, n_416);
  xor g1136 (n_420, n_1186, n_417);
  nand g1137 (n_1187, n_415, n_416);
  nand g1138 (n_1188, n_417, n_416);
  nand g1139 (n_1189, n_415, n_417);
  nand g1140 (n_439, n_1187, n_1188, n_1189);
  xor g1141 (n_1190, A[16], A[17]);
  xor g1142 (n_423, n_1190, n_418);
  nand g1143 (n_1191, A[16], A[17]);
  nand g1144 (n_1192, n_418, A[17]);
  nand g1145 (n_1193, A[16], n_418);
  nand g1146 (n_440, n_1191, n_1192, n_1193);
  xor g1148 (n_424, n_1194, A[20]);
  nand g1152 (n_442, n_1195, n_1156, n_1027);
  xor g1153 (n_1198, n_419, n_420);
  xor g1154 (n_426, n_1198, n_421);
  nand g1155 (n_1199, n_419, n_420);
  nand g1156 (n_1200, n_421, n_420);
  nand g1157 (n_1201, n_419, n_421);
  nand g1158 (n_444, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_422, n_423);
  xor g1160 (n_428, n_1202, n_424);
  nand g1161 (n_1203, n_422, n_423);
  nand g1162 (n_1204, n_424, n_423);
  nand g1163 (n_1205, n_422, n_424);
  nand g1164 (n_447, n_1203, n_1204, n_1205);
  xor g1165 (n_1206, n_425, n_426);
  xor g1166 (n_429, n_1206, n_427);
  nand g1167 (n_1207, n_425, n_426);
  nand g1168 (n_1208, n_427, n_426);
  nand g1169 (n_1209, n_425, n_427);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, n_433);
  nand g1183 (n_1217, A[6], n_433);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, A[9], A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, A[9], A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, A[9], n_434);
  nand g1190 (n_456, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, A[14], A[13]);
  xor g1192 (n_438, n_1222, n_435);
  nand g1193 (n_1223, A[14], A[13]);
  nand g1194 (n_1224, n_435, A[13]);
  nand g1195 (n_1225, A[14], n_435);
  nand g1196 (n_458, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, n_436, n_437);
  xor g1198 (n_441, n_1226, A[18]);
  nand g1199 (n_1227, n_436, n_437);
  nand g1200 (n_1228, A[18], n_437);
  nand g1201 (n_1229, n_436, A[18]);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, A[17], n_438);
  xor g1204 (n_443, n_1230, A[21]);
  nand g1205 (n_1231, A[17], n_438);
  nand g1206 (n_1232, A[21], n_438);
  nand g1207 (n_1233, A[17], A[21]);
  nand g1208 (n_461, n_1231, n_1232, n_1233);
  xor g1209 (n_1234, A[22], n_439);
  xor g1210 (n_445, n_1234, n_440);
  nand g1211 (n_1235, A[22], n_439);
  nand g1212 (n_1236, n_440, n_439);
  nand g1213 (n_1237, A[22], n_440);
  nand g1214 (n_463, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_441, n_442);
  xor g1216 (n_446, n_1238, n_443);
  nand g1217 (n_1239, n_441, n_442);
  nand g1218 (n_1240, n_443, n_442);
  nand g1219 (n_1241, n_441, n_443);
  nand g1220 (n_465, n_1239, n_1240, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[5], A[7]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], A[11]);
  xor g1242 (n_455, n_1254, n_453);
  nand g1243 (n_1255, A[10], A[11]);
  nand g1244 (n_1256, n_453, A[11]);
  nand g1245 (n_1257, A[10], n_453);
  nand g1246 (n_472, n_1255, n_1256, n_1257);
  xor g1247 (n_1258, A[14], n_454);
  xor g1248 (n_457, n_1258, A[15]);
  nand g1249 (n_1259, A[14], n_454);
  nand g1250 (n_1260, A[15], n_454);
  nand g1252 (n_474, n_1259, n_1260, n_944);
  xor g1253 (n_1262, n_455, n_456);
  xor g1254 (n_460, n_1262, A[19]);
  nand g1255 (n_1263, n_455, n_456);
  nand g1256 (n_1264, A[19], n_456);
  nand g1257 (n_1265, n_455, A[19]);
  nand g1258 (n_477, n_1263, n_1264, n_1265);
  xor g1259 (n_1266, A[18], n_457);
  xor g1260 (n_462, n_1266, n_458);
  nand g1261 (n_1267, A[18], n_457);
  nand g1262 (n_1268, n_458, n_457);
  nand g1263 (n_1269, A[18], n_458);
  nand g1264 (n_478, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, A[22], A[23]);
  xor g1266 (n_464, n_1270, n_459);
  nand g1267 (n_1271, A[22], A[23]);
  nand g1268 (n_1272, n_459, A[23]);
  nand g1269 (n_1273, A[22], n_459);
  nand g1270 (n_480, n_1271, n_1272, n_1273);
  xor g1271 (n_1274, n_460, n_461);
  xor g1272 (n_466, n_1274, n_462);
  nand g1273 (n_1275, n_460, n_461);
  nand g1274 (n_1276, n_462, n_461);
  nand g1275 (n_1277, n_460, n_462);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1277 (n_1278, n_463, n_464);
  xor g1278 (n_467, n_1278, n_465);
  nand g1279 (n_1279, n_463, n_464);
  nand g1280 (n_1280, n_465, n_464);
  nand g1281 (n_1281, n_463, n_465);
  nand g1282 (n_485, n_1279, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1289 (n_1286, A[7], A[6]);
  xor g1290 (n_471, n_1286, A[8]);
  nand g1292 (n_1288, A[8], A[6]);
  nand g1294 (n_486, n_661, n_1288, n_673);
  xor g1296 (n_473, n_1142, n_470);
  nand g1298 (n_1292, n_470, A[12]);
  nand g1299 (n_1293, A[11], n_470);
  nand g1300 (n_487, n_744, n_1292, n_1293);
  xor g1301 (n_1294, n_471, A[15]);
  xor g1302 (n_475, n_1294, n_472);
  nand g1303 (n_1295, n_471, A[15]);
  nand g1304 (n_1296, n_472, A[15]);
  nand g1305 (n_1297, n_471, n_472);
  nand g1306 (n_489, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, n_473, A[16]);
  xor g1308 (n_476, n_1298, A[19]);
  nand g1309 (n_1299, n_473, A[16]);
  nand g1311 (n_1301, n_473, A[19]);
  nand g1312 (n_492, n_1299, n_1151, n_1301);
  xor g1314 (n_479, n_1302, A[20]);
  nand g1317 (n_1305, n_474, A[20]);
  nand g1318 (n_493, n_1303, n_1156, n_1305);
  xor g1319 (n_1306, n_475, A[23]);
  xor g1320 (n_481, n_1306, n_476);
  nand g1321 (n_1307, n_475, A[23]);
  nand g1322 (n_1308, n_476, A[23]);
  nand g1323 (n_1309, n_475, n_476);
  nand g1324 (n_496, n_1307, n_1308, n_1309);
  xor g1325 (n_1310, n_477, n_478);
  xor g1326 (n_483, n_1310, n_479);
  nand g1327 (n_1311, n_477, n_478);
  nand g1328 (n_1312, n_479, n_478);
  nand g1329 (n_1313, n_477, n_479);
  nand g1330 (n_498, n_1311, n_1312, n_1313);
  xor g1331 (n_1314, n_480, n_481);
  xor g1332 (n_484, n_1314, n_482);
  nand g1333 (n_1315, n_480, n_481);
  nand g1334 (n_1316, n_482, n_481);
  nand g1335 (n_1317, n_480, n_482);
  nand g1336 (n_499, n_1315, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1349 (n_1326, n_486, A[13]);
  xor g1350 (n_490, n_1326, n_487);
  nand g1351 (n_1327, n_486, A[13]);
  nand g1352 (n_1328, n_487, A[13]);
  nand g1353 (n_1329, n_486, n_487);
  nand g1354 (n_505, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, n_223, A[16]);
  xor g1356 (n_491, n_1330, A[17]);
  nand g1357 (n_1331, n_223, A[16]);
  nand g1359 (n_1333, n_223, A[17]);
  nand g1360 (n_506, n_1331, n_1191, n_1333);
  xor g1362 (n_494, n_1334, n_490);
  nand g1365 (n_1337, n_489, n_490);
  nand g1366 (n_508, n_1335, n_1336, n_1337);
  xor g1368 (n_495, n_1026, n_491);
  nand g1370 (n_1340, n_491, A[21]);
  nand g1371 (n_1341, A[20], n_491);
  nand g1372 (n_510, n_1027, n_1340, n_1341);
  xor g1373 (n_1342, n_492, n_493);
  xor g1374 (n_497, n_1342, n_494);
  nand g1375 (n_1343, n_492, n_493);
  nand g1376 (n_1344, n_494, n_493);
  nand g1377 (n_1345, n_492, n_494);
  nand g1378 (n_513, n_1343, n_1344, n_1345);
  xor g1379 (n_1346, n_495, n_496);
  xor g1380 (n_500, n_1346, n_497);
  nand g1381 (n_1347, n_495, n_496);
  nand g1382 (n_1348, n_497, n_496);
  nand g1383 (n_1349, n_495, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  nand g1397 (n_1357, A[9], A[14]);
  nand g1398 (n_519, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], n_234);
  xor g1400 (n_507, n_1358, A[18]);
  nand g1402 (n_1360, A[18], n_234);
  nand g1403 (n_1361, A[13], A[18]);
  nand g1404 (n_522, n_797, n_1360, n_1361);
  xor g1405 (n_1362, A[17], n_504);
  xor g1406 (n_509, n_1362, A[21]);
  nand g1407 (n_1363, A[17], n_504);
  nand g1408 (n_1364, A[21], n_504);
  nand g1410 (n_523, n_1363, n_1364, n_1233);
  xor g1411 (n_1366, n_505, A[22]);
  xor g1412 (n_511, n_1366, n_506);
  nand g1413 (n_1367, n_505, A[22]);
  nand g1414 (n_1368, n_506, A[22]);
  nand g1415 (n_1369, n_505, n_506);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_507, n_508);
  xor g1418 (n_512, n_1370, n_509);
  nand g1419 (n_1371, n_507, n_508);
  nand g1420 (n_1372, n_509, n_508);
  nand g1421 (n_1373, n_507, n_509);
  nand g1422 (n_527, n_1371, n_1372, n_1373);
  xor g1423 (n_1374, n_510, n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, n_510, n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, n_510, n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1443 (n_1386, A[14], A[15]);
  xor g1444 (n_521, n_1386, n_519);
  nand g1446 (n_1388, n_519, A[15]);
  nand g1447 (n_1389, A[14], n_519);
  nand g1448 (n_534, n_944, n_1388, n_1389);
  xor g1449 (n_1390, A[19], A[18]);
  xor g1450 (n_524, n_1390, n_520);
  nand g1452 (n_1392, n_520, A[18]);
  nand g1453 (n_1393, A[19], n_520);
  nand g1454 (n_536, n_953, n_1392, n_1393);
  xor g1455 (n_1394, A[22], n_521);
  xor g1456 (n_525, n_1394, A[23]);
  nand g1457 (n_1395, A[22], n_521);
  nand g1458 (n_1396, A[23], n_521);
  nand g1460 (n_538, n_1395, n_1396, n_1271);
  xor g1461 (n_1398, n_522, n_523);
  xor g1462 (n_528, n_1398, n_524);
  nand g1463 (n_1399, n_522, n_523);
  nand g1464 (n_1400, n_524, n_523);
  nand g1465 (n_1401, n_522, n_524);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1467 (n_1402, n_525, n_526);
  xor g1468 (n_529, n_1402, n_527);
  nand g1469 (n_1403, n_525, n_526);
  nand g1470 (n_1404, n_527, n_526);
  nand g1471 (n_1405, n_525, n_527);
  nand g1472 (n_543, n_1403, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1480 (n_533, n_1142, A[10]);
  nand g1483 (n_1413, A[12], A[10]);
  nand g1484 (n_544, n_744, n_1255, n_1413);
  xor g1485 (n_1414, A[15], n_532);
  xor g1486 (n_535, n_1414, A[16]);
  nand g1487 (n_1415, A[15], n_532);
  nand g1488 (n_1416, A[16], n_532);
  nand g1489 (n_1417, A[15], A[16]);
  nand g1490 (n_545, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, n_533, A[19]);
  nand g1493 (n_1419, n_533, A[19]);
  nand g1496 (n_547, n_1419, n_1420, n_1421);
  xor g1497 (n_1422, A[20], A[23]);
  xor g1498 (n_539, n_1422, n_534);
  nand g1500 (n_1424, n_534, A[23]);
  nand g1501 (n_1425, A[20], n_534);
  nand g1502 (n_550, n_1028, n_1424, n_1425);
  xor g1503 (n_1426, n_535, n_536);
  xor g1504 (n_541, n_1426, n_537);
  nand g1505 (n_1427, n_535, n_536);
  nand g1506 (n_1428, n_537, n_536);
  nand g1507 (n_1429, n_535, n_537);
  nand g1508 (n_551, n_1427, n_1428, n_1429);
  xor g1509 (n_1430, n_538, n_539);
  xor g1510 (n_542, n_1430, n_540);
  nand g1511 (n_1431, n_538, n_539);
  nand g1512 (n_1432, n_540, n_539);
  nand g1513 (n_1433, n_538, n_540);
  nand g1514 (n_554, n_1431, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1521 (n_1438, A[12], A[13]);
  xor g1522 (n_546, n_1438, n_544);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_1184, n_1440, n_1441);
  xor g1528 (n_548, n_1190, A[21]);
  nand g1531 (n_1445, A[16], A[21]);
  nand g1532 (n_559, n_1191, n_1233, n_1445);
  xor g1534 (n_549, n_1446, n_545);
  nand g1536 (n_1448, n_545, A[20]);
  nand g1538 (n_561, n_1156, n_1448, n_1449);
  xor g1539 (n_1450, n_546, n_547);
  xor g1540 (n_552, n_1450, n_548);
  nand g1541 (n_1451, n_546, n_547);
  nand g1542 (n_1452, n_548, n_547);
  nand g1543 (n_1453, n_546, n_548);
  nand g1544 (n_562, n_1451, n_1452, n_1453);
  xor g1545 (n_1454, n_549, n_550);
  xor g1546 (n_553, n_1454, n_551);
  nand g1547 (n_1455, n_549, n_550);
  nand g1548 (n_1456, n_551, n_550);
  nand g1549 (n_1457, n_549, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1564 (n_570, n_1463, n_1464, n_1361);
  xor g1565 (n_1466, A[17], A[21]);
  xor g1566 (n_560, n_1466, A[22]);
  nand g1569 (n_1469, A[17], A[22]);
  nand g1570 (n_572, n_1233, n_1071, n_1469);
  xor g1571 (n_1470, n_557, n_558);
  xor g1572 (n_563, n_1470, n_559);
  nand g1573 (n_1471, n_557, n_558);
  nand g1574 (n_1472, n_559, n_558);
  nand g1575 (n_1473, n_557, n_559);
  nand g1576 (n_574, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, n_560, n_561);
  xor g1578 (n_564, n_1474, n_562);
  nand g1579 (n_1475, n_560, n_561);
  nand g1580 (n_1476, n_562, n_561);
  nand g1581 (n_1477, n_560, n_562);
  nand g1582 (n_576, n_1475, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  xor g1598 (n_571, n_1390, A[22]);
  nand g1602 (n_580, n_953, n_1113, n_987);
  xor g1603 (n_1490, A[23], n_569);
  xor g1604 (n_573, n_1490, n_570);
  nand g1605 (n_1491, A[23], n_569);
  nand g1606 (n_1492, n_570, n_569);
  nand g1607 (n_1493, A[23], n_570);
  nand g1608 (n_583, n_1491, n_1492, n_1493);
  xor g1609 (n_1494, n_571, n_572);
  xor g1610 (n_575, n_1494, n_573);
  nand g1611 (n_1495, n_571, n_572);
  nand g1612 (n_1496, n_573, n_572);
  nand g1613 (n_1497, n_571, n_573);
  nand g1614 (n_585, n_1495, n_1496, n_1497);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1622 (n_579, n_1386, A[16]);
  nand g1624 (n_1504, A[16], A[14]);
  nand g1626 (n_586, n_944, n_1504, n_1417);
  xor g1627 (n_1506, A[19], n_578);
  nand g1629 (n_1507, A[19], n_578);
  nand g1632 (n_588, n_1507, n_1508, n_1420);
  xor g1634 (n_582, n_1422, n_579);
  nand g1636 (n_1512, n_579, A[23]);
  nand g1637 (n_1513, A[20], n_579);
  nand g1638 (n_589, n_1028, n_1512, n_1513);
  xor g1639 (n_1514, n_580, n_581);
  xor g1640 (n_584, n_1514, n_582);
  nand g1641 (n_1515, n_580, n_581);
  nand g1642 (n_1516, n_582, n_581);
  nand g1643 (n_1517, n_580, n_582);
  nand g1644 (n_592, n_1515, n_1516, n_1517);
  xor g1645 (n_1518, n_583, n_584);
  xor g1646 (n_83, n_1518, n_585);
  nand g1647 (n_1519, n_583, n_584);
  nand g1648 (n_1520, n_585, n_584);
  nand g1649 (n_1521, n_583, n_585);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1658 (n_590, n_1446, n_586);
  nand g1660 (n_1528, n_586, A[20]);
  nand g1662 (n_596, n_1156, n_1528, n_1529);
  xor g1663 (n_1530, n_548, n_588);
  xor g1664 (n_591, n_1530, n_589);
  nand g1665 (n_1531, n_548, n_588);
  nand g1666 (n_1532, n_589, n_588);
  nand g1667 (n_1533, n_548, n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_33, n_1535, n_1536, n_1537);
  xor g1684 (n_598, n_1542, n_596);
  nand g1686 (n_1544, n_596, n_559);
  nand g1688 (n_606, n_1543, n_1544, n_1545);
  xor g1689 (n_1546, n_560, n_598);
  xor g1690 (n_81, n_1546, n_599);
  nand g1691 (n_1547, n_560, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_560, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[18], A[22]);
  xor g1698 (n_604, n_1550, A[23]);
  nand g1701 (n_1553, A[18], A[23]);
  nand g1702 (n_609, n_1113, n_1271, n_1553);
  nand g1706 (n_1556, n_572, A[18]);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, n_604, n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, n_604, n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, n_604, n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1716 (n_608, n_1562, A[20]);
  nand g1719 (n_1565, A[19], A[20]);
  nand g1720 (n_612, n_1420, n_1156, n_1565);
  xor g1721 (n_1566, A[23], A[19]);
  xor g1722 (n_611, n_1566, n_608);
  nand g1723 (n_1567, A[23], A[19]);
  nand g1724 (n_1568, n_608, A[19]);
  nand g1725 (n_1569, A[23], n_608);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1727 (n_1570, n_609, n_610);
  xor g1728 (n_79, n_1570, n_611);
  nand g1729 (n_1571, n_609, n_610);
  nand g1730 (n_1572, n_611, n_610);
  nand g1731 (n_1573, n_609, n_611);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1739 (n_1578, n_612, n_424);
  xor g1740 (n_78, n_1578, n_614);
  nand g1741 (n_1579, n_612, n_424);
  nand g1742 (n_1580, n_614, n_424);
  nand g1743 (n_1581, n_612, n_614);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_442);
  nand g1752 (n_28, n_1583, n_1584, n_1585);
  nand g1760 (n_27, n_1587, n_1588, n_1029);
  xor g1762 (n_75, n_1590, A[22]);
  nand g1766 (n_74, n_1591, n_1271, n_1593);
  nor g11 (n_1609, A[0], A[2]);
  nand g12 (n_1604, A[0], A[2]);
  nor g13 (n_1605, n_68, A[3]);
  nand g14 (n_1606, n_68, A[3]);
  nor g15 (n_1615, A[4], n_117);
  nand g16 (n_1610, A[4], n_117);
  nor g17 (n_1611, A[5], n_116);
  nand g18 (n_1612, A[5], n_116);
  nor g19 (n_1621, n_67, n_115);
  nand g20 (n_1616, n_67, n_115);
  nor g21 (n_1617, n_66, n_114);
  nand g22 (n_1618, n_66, n_114);
  nor g23 (n_1627, n_65, n_113);
  nand g24 (n_1622, n_65, n_113);
  nor g25 (n_1623, n_64, n_112);
  nand g26 (n_1624, n_64, n_112);
  nor g27 (n_1633, n_63, n_111);
  nand g28 (n_1628, n_63, n_111);
  nor g29 (n_1629, n_62, n_110);
  nand g30 (n_1630, n_62, n_110);
  nor g31 (n_1639, n_61, n_109);
  nand g32 (n_1634, n_61, n_109);
  nor g33 (n_1635, n_60, n_108);
  nand g34 (n_1636, n_60, n_108);
  nor g35 (n_1645, n_59, n_107);
  nand g36 (n_1640, n_59, n_107);
  nor g37 (n_1641, n_58, n_106);
  nand g38 (n_1642, n_58, n_106);
  nor g39 (n_1651, n_57, n_105);
  nand g40 (n_1646, n_57, n_105);
  nor g41 (n_1647, n_56, n_104);
  nand g42 (n_1648, n_56, n_104);
  nor g43 (n_1657, n_55, n_103);
  nand g44 (n_1652, n_55, n_103);
  nor g45 (n_1653, n_54, n_102);
  nand g46 (n_1654, n_54, n_102);
  nor g47 (n_1663, n_53, n_101);
  nand g48 (n_1658, n_53, n_101);
  nor g49 (n_1659, n_52, n_100);
  nand g50 (n_1660, n_52, n_100);
  nor g51 (n_1669, n_51, n_99);
  nand g52 (n_1664, n_51, n_99);
  nor g53 (n_1665, n_50, n_98);
  nand g54 (n_1666, n_50, n_98);
  nor g55 (n_1675, n_49, n_97);
  nand g56 (n_1670, n_49, n_97);
  nor g57 (n_1671, n_48, n_96);
  nand g58 (n_1672, n_48, n_96);
  nor g59 (n_1681, n_47, n_95);
  nand g60 (n_1676, n_47, n_95);
  nor g61 (n_1677, n_46, n_94);
  nand g62 (n_1678, n_46, n_94);
  nor g63 (n_1687, n_45, n_93);
  nand g64 (n_1682, n_45, n_93);
  nor g65 (n_1683, n_44, n_92);
  nand g66 (n_1684, n_44, n_92);
  nor g67 (n_1693, n_43, n_91);
  nand g68 (n_1688, n_43, n_91);
  nor g69 (n_1689, n_42, n_90);
  nand g70 (n_1690, n_42, n_90);
  nor g71 (n_1699, n_41, n_89);
  nand g72 (n_1694, n_41, n_89);
  nor g73 (n_1695, n_40, n_88);
  nand g74 (n_1696, n_40, n_88);
  nor g75 (n_1705, n_39, n_87);
  nand g76 (n_1700, n_39, n_87);
  nor g77 (n_1701, n_38, n_86);
  nand g78 (n_1702, n_38, n_86);
  nor g79 (n_1711, n_37, n_85);
  nand g80 (n_1706, n_37, n_85);
  nor g81 (n_1707, n_36, n_84);
  nand g82 (n_1708, n_36, n_84);
  nor g83 (n_1717, n_35, n_83);
  nand g84 (n_1712, n_35, n_83);
  nor g85 (n_1713, n_34, n_82);
  nand g86 (n_1714, n_34, n_82);
  nor g87 (n_1723, n_33, n_81);
  nand g88 (n_1718, n_33, n_81);
  nor g89 (n_1719, n_32, n_80);
  nand g90 (n_1720, n_32, n_80);
  nor g91 (n_1729, n_31, n_79);
  nand g92 (n_1724, n_31, n_79);
  nor g93 (n_1725, n_30, n_78);
  nand g94 (n_1726, n_30, n_78);
  nor g95 (n_1735, n_29, n_77);
  nand g96 (n_1730, n_29, n_77);
  nor g97 (n_1731, n_28, n_76);
  nand g98 (n_1732, n_28, n_76);
  nor g99 (n_1739, n_27, n_75);
  nand g100 (n_1736, n_27, n_75);
  nor g106 (n_1607, n_1604, n_1605);
  nor g110 (n_1613, n_1610, n_1611);
  nor g113 (n_1749, n_1615, n_1611);
  nor g114 (n_1619, n_1616, n_1617);
  nor g117 (n_1751, n_1621, n_1617);
  nor g118 (n_1625, n_1622, n_1623);
  nor g121 (n_1759, n_1627, n_1623);
  nor g122 (n_1631, n_1628, n_1629);
  nor g125 (n_1761, n_1633, n_1629);
  nor g126 (n_1637, n_1634, n_1635);
  nor g129 (n_1769, n_1639, n_1635);
  nor g130 (n_1643, n_1640, n_1641);
  nor g133 (n_1771, n_1645, n_1641);
  nor g134 (n_1649, n_1646, n_1647);
  nor g137 (n_1779, n_1651, n_1647);
  nor g138 (n_1655, n_1652, n_1653);
  nor g141 (n_1781, n_1657, n_1653);
  nor g142 (n_1661, n_1658, n_1659);
  nor g145 (n_1789, n_1663, n_1659);
  nor g146 (n_1667, n_1664, n_1665);
  nor g149 (n_1791, n_1669, n_1665);
  nor g150 (n_1673, n_1670, n_1671);
  nor g153 (n_1799, n_1675, n_1671);
  nor g154 (n_1679, n_1676, n_1677);
  nor g157 (n_1801, n_1681, n_1677);
  nor g158 (n_1685, n_1682, n_1683);
  nor g161 (n_1809, n_1687, n_1683);
  nor g162 (n_1691, n_1688, n_1689);
  nor g165 (n_1811, n_1693, n_1689);
  nor g166 (n_1697, n_1694, n_1695);
  nor g169 (n_1819, n_1699, n_1695);
  nor g170 (n_1703, n_1700, n_1701);
  nor g173 (n_1821, n_1705, n_1701);
  nor g174 (n_1709, n_1706, n_1707);
  nor g177 (n_1829, n_1711, n_1707);
  nor g178 (n_1715, n_1712, n_1713);
  nor g181 (n_1831, n_1717, n_1713);
  nor g182 (n_1721, n_1718, n_1719);
  nor g185 (n_1839, n_1723, n_1719);
  nor g186 (n_1727, n_1724, n_1725);
  nor g189 (n_1841, n_1729, n_1725);
  nor g190 (n_1733, n_1730, n_1731);
  nor g193 (n_1849, n_1735, n_1731);
  nor g203 (n_1747, n_1621, n_1746);
  nand g212 (n_1859, n_1749, n_1751);
  nor g213 (n_1757, n_1633, n_1756);
  nand g222 (n_1866, n_1759, n_1761);
  nor g223 (n_1767, n_1645, n_1766);
  nand g232 (n_1874, n_1769, n_1771);
  nor g233 (n_1777, n_1657, n_1776);
  nand g242 (n_1881, n_1779, n_1781);
  nor g243 (n_1787, n_1669, n_1786);
  nand g252 (n_1889, n_1789, n_1791);
  nor g253 (n_1797, n_1681, n_1796);
  nand g262 (n_1896, n_1799, n_1801);
  nor g263 (n_1807, n_1693, n_1806);
  nand g1776 (n_1904, n_1809, n_1811);
  nor g1777 (n_1817, n_1705, n_1816);
  nand g1786 (n_1911, n_1819, n_1821);
  nor g1787 (n_1827, n_1717, n_1826);
  nand g1796 (n_1919, n_1829, n_1831);
  nor g1797 (n_1837, n_1729, n_1836);
  nand g1806 (n_1926, n_1839, n_1841);
  nor g1807 (n_1847, n_1739, n_1846);
  nand g1814 (n_2130, n_1610, n_1853);
  nand g1816 (n_2132, n_1746, n_1854);
  nand g1819 (n_2135, n_1857, n_1858);
  nand g1822 (n_1934, n_1861, n_1862);
  nor g1823 (n_1864, n_1639, n_1863);
  nor g1826 (n_1944, n_1639, n_1866);
  nor g1832 (n_1872, n_1870, n_1863);
  nor g1835 (n_1950, n_1866, n_1870);
  nor g1836 (n_1876, n_1874, n_1863);
  nor g1839 (n_1953, n_1866, n_1874);
  nor g1840 (n_1879, n_1663, n_1878);
  nor g1843 (n_2033, n_1663, n_1881);
  nor g1849 (n_1887, n_1885, n_1878);
  nor g1852 (n_2039, n_1881, n_1885);
  nor g1853 (n_1891, n_1889, n_1878);
  nor g1856 (n_1959, n_1881, n_1889);
  nor g1857 (n_1894, n_1687, n_1893);
  nor g1860 (n_1972, n_1687, n_1896);
  nor g1866 (n_1902, n_1900, n_1893);
  nor g1869 (n_1982, n_1896, n_1900);
  nor g1870 (n_1906, n_1904, n_1893);
  nor g1873 (n_1987, n_1896, n_1904);
  nor g1874 (n_1909, n_1711, n_1908);
  nor g1877 (n_2085, n_1711, n_1911);
  nor g1883 (n_1917, n_1915, n_1908);
  nor g1886 (n_2091, n_1911, n_1915);
  nor g1887 (n_1921, n_1919, n_1908);
  nor g1890 (n_1995, n_1911, n_1919);
  nor g1891 (n_1924, n_1735, n_1923);
  nor g1894 (n_2008, n_1735, n_1926);
  nor g1900 (n_1932, n_1930, n_1923);
  nor g1903 (n_2018, n_1926, n_1930);
  nand g1906 (n_2139, n_1622, n_1936);
  nand g1907 (n_1937, n_1759, n_1934);
  nand g1908 (n_2141, n_1756, n_1937);
  nand g1911 (n_2144, n_1940, n_1941);
  nand g1914 (n_2147, n_1863, n_1943);
  nand g1915 (n_1946, n_1944, n_1934);
  nand g1916 (n_2150, n_1945, n_1946);
  nand g1917 (n_1949, n_1947, n_1934);
  nand g1918 (n_2152, n_1948, n_1949);
  nand g1919 (n_1952, n_1950, n_1934);
  nand g1920 (n_2155, n_1951, n_1952);
  nand g1921 (n_1955, n_1953, n_1934);
  nand g1922 (n_2023, n_1954, n_1955);
  nor g1923 (n_1957, n_1675, n_1956);
  nand g1932 (n_2047, n_1799, n_1959);
  nor g1933 (n_1966, n_1964, n_1956);
  nor g1938 (n_1969, n_1896, n_1956);
  nand g1947 (n_2059, n_1959, n_1972);
  nand g1952 (n_2063, n_1959, n_1977);
  nand g1957 (n_2067, n_1959, n_1982);
  nand g1962 (n_2071, n_1959, n_1987);
  nor g1963 (n_1993, n_1723, n_1992);
  nand g1972 (n_2099, n_1839, n_1995);
  nor g1973 (n_2002, n_2000, n_1992);
  nor g1978 (n_2005, n_1926, n_1992);
  nand g1987 (n_2111, n_1995, n_2008);
  nand g1992 (n_2115, n_1995, n_2013);
  nand g1997 (n_2119, n_1995, n_2018);
  nand g2000 (n_2159, n_1646, n_2025);
  nand g2001 (n_2026, n_1779, n_2023);
  nand g2002 (n_2161, n_1776, n_2026);
  nand g2005 (n_2164, n_2029, n_2030);
  nand g2008 (n_2167, n_1878, n_2032);
  nand g2009 (n_2035, n_2033, n_2023);
  nand g2010 (n_2170, n_2034, n_2035);
  nand g2011 (n_2038, n_2036, n_2023);
  nand g2012 (n_2172, n_2037, n_2038);
  nand g2013 (n_2041, n_2039, n_2023);
  nand g2014 (n_2175, n_2040, n_2041);
  nand g2015 (n_2042, n_1959, n_2023);
  nand g2016 (n_2177, n_1956, n_2042);
  nand g2019 (n_2180, n_2045, n_2046);
  nand g2022 (n_2182, n_2049, n_2050);
  nand g2025 (n_2185, n_2053, n_2054);
  nand g2028 (n_2188, n_2057, n_2058);
  nand g2031 (n_2191, n_2061, n_2062);
  nand g2034 (n_2193, n_2065, n_2066);
  nand g2037 (n_2196, n_2069, n_2070);
  nand g2040 (n_2075, n_2073, n_2074);
  nand g2043 (n_2200, n_1694, n_2077);
  nand g2044 (n_2078, n_1819, n_2075);
  nand g2045 (n_2202, n_1816, n_2078);
  nand g2048 (n_2205, n_2081, n_2082);
  nand g2051 (n_2208, n_1908, n_2084);
  nand g2052 (n_2087, n_2085, n_2075);
  nand g2053 (n_2211, n_2086, n_2087);
  nand g2054 (n_2090, n_2088, n_2075);
  nand g2055 (n_2213, n_2089, n_2090);
  nand g2056 (n_2093, n_2091, n_2075);
  nand g2057 (n_2216, n_2092, n_2093);
  nand g2058 (n_2094, n_1995, n_2075);
  nand g2059 (n_2218, n_1992, n_2094);
  nand g2062 (n_2221, n_2097, n_2098);
  nand g2065 (n_2223, n_2101, n_2102);
  nand g2068 (n_2226, n_2105, n_2106);
  nand g2071 (n_2229, n_2109, n_2110);
  nand g2074 (n_2232, n_2113, n_2114);
  nand g2077 (n_2234, n_2117, n_2118);
  nand g2080 (n_2237, n_2121, n_2122);
  xnor g2092 (Z[5], n_2130, n_2131);
  xnor g2094 (Z[6], n_2132, n_2133);
  xnor g2097 (Z[7], n_2135, n_2136);
  xnor g2099 (Z[8], n_1934, n_2137);
  xnor g2102 (Z[9], n_2139, n_2140);
  xnor g2104 (Z[10], n_2141, n_2142);
  xnor g2107 (Z[11], n_2144, n_2145);
  xnor g2110 (Z[12], n_2147, n_2148);
  xnor g2113 (Z[13], n_2150, n_2151);
  xnor g2115 (Z[14], n_2152, n_2153);
  xnor g2118 (Z[15], n_2155, n_2156);
  xnor g2120 (Z[16], n_2023, n_2157);
  xnor g2123 (Z[17], n_2159, n_2160);
  xnor g2125 (Z[18], n_2161, n_2162);
  xnor g2128 (Z[19], n_2164, n_2165);
  xnor g2131 (Z[20], n_2167, n_2168);
  xnor g2134 (Z[21], n_2170, n_2171);
  xnor g2136 (Z[22], n_2172, n_2173);
  xnor g2139 (Z[23], n_2175, n_2176);
  xnor g2141 (Z[24], n_2177, n_2178);
  xnor g2144 (Z[25], n_2180, n_2181);
  xnor g2146 (Z[26], n_2182, n_2183);
  xnor g2149 (Z[27], n_2185, n_2186);
  xnor g2152 (Z[28], n_2188, n_2189);
  xnor g2155 (Z[29], n_2191, n_2192);
  xnor g2157 (Z[30], n_2193, n_2194);
  xnor g2160 (Z[31], n_2196, n_2197);
  xnor g2162 (Z[32], n_2075, n_2198);
  xnor g2165 (Z[33], n_2200, n_2201);
  xnor g2167 (Z[34], n_2202, n_2203);
  xnor g2170 (Z[35], n_2205, n_2206);
  xnor g2173 (Z[36], n_2208, n_2209);
  xnor g2176 (Z[37], n_2211, n_2212);
  xnor g2178 (Z[38], n_2213, n_2214);
  xnor g2181 (Z[39], n_2216, n_2217);
  xnor g2183 (Z[40], n_2218, n_2219);
  xnor g2186 (Z[41], n_2221, n_2222);
  xnor g2188 (Z[42], n_2223, n_2224);
  xnor g2191 (Z[43], n_2226, n_2227);
  xnor g2194 (Z[44], n_2229, n_2230);
  xnor g2197 (Z[45], n_2232, n_2233);
  xnor g2199 (Z[46], n_2234, n_2235);
  xnor g2202 (Z[47], n_2237, n_2238);
  or g2214 (n_1044, A[1], wc);
  not gc (wc, n_171);
  or g2215 (n_1045, A[1], wc0);
  not gc0 (wc0, A[2]);
  or g2216 (n_1069, wc1, A[24]);
  not gc1 (wc1, A[18]);
  or g2217 (n_1088, A[2], wc2);
  not gc2 (wc2, A[3]);
  or g2218 (n_1089, wc3, A[2]);
  not gc3 (wc3, A[1]);
  or g2219 (n_1156, wc4, A[24]);
  not gc4 (wc4, A[20]);
  xnor g2220 (n_1194, A[24], A[21]);
  or g2221 (n_1195, wc5, A[24]);
  not gc5 (wc5, A[21]);
  xnor g2222 (n_1214, A[6], A[5]);
  or g2223 (n_1215, A[5], wc6);
  not gc6 (wc6, A[6]);
  or g2224 (n_1252, A[6], wc7);
  not gc7 (wc7, A[7]);
  or g2225 (n_1253, wc8, A[6]);
  not gc8 (wc8, A[5]);
  or g2227 (n_1355, wc9, A[10]);
  not gc9 (wc9, A[9]);
  or g2228 (n_1356, A[10], wc10);
  not gc10 (wc10, A[14]);
  or g2229 (n_1385, A[10], wc11);
  not gc11 (wc11, A[11]);
  or g2230 (n_1420, wc12, A[24]);
  not gc12 (wc12, A[19]);
  xnor g2231 (n_1446, A[24], A[20]);
  or g2233 (n_1463, wc13, A[14]);
  not gc13 (wc13, A[13]);
  or g2234 (n_1464, A[14], wc14);
  not gc14 (wc14, A[18]);
  or g2235 (n_1485, A[14], wc15);
  not gc15 (wc15, A[15]);
  or g2237 (n_1555, wc16, A[19]);
  not gc16 (wc16, A[18]);
  xnor g2238 (n_1562, A[24], A[19]);
  or g2240 (n_1583, A[21], wc17);
  not gc17 (wc17, A[22]);
  or g2242 (n_1587, A[22], wc18);
  not gc18 (wc18, A[23]);
  or g2243 (n_1588, wc19, A[22]);
  not gc19 (wc19, A[21]);
  xnor g2244 (n_1590, A[24], A[23]);
  or g2245 (n_1591, wc20, A[24]);
  not gc20 (wc20, A[23]);
  or g2246 (n_1593, wc21, A[24]);
  not gc21 (wc21, A[22]);
  xnor g2247 (n_349, n_1042, A[1]);
  xnor g2248 (n_372, n_1086, A[2]);
  xnor g2249 (n_453, n_1250, A[6]);
  xnor g2250 (n_504, n_1218, A[14]);
  xnor g2251 (n_520, n_1254, A[10]);
  nand g2252 (n_532, n_1255, n_1385);
  or g2253 (n_1421, A[24], wc22);
  not gc22 (wc22, n_533);
  xnor g2254 (n_558, n_1222, A[18]);
  xnor g2255 (n_569, n_1386, A[14]);
  nand g2256 (n_578, n_944, n_1485);
  xnor g2257 (n_1542, n_559, A[18]);
  or g2258 (n_1543, A[18], wc23);
  not gc23 (wc23, n_559);
  xnor g2259 (n_605, n_1390, n_572);
  or g2260 (n_1557, A[19], wc24);
  not gc24 (wc24, n_572);
  xnor g2261 (n_76, n_1270, A[21]);
  or g2263 (n_2124, wc25, n_1609);
  not gc25 (wc25, n_1604);
  xnor g2264 (n_537, n_1418, A[24]);
  or g2265 (n_1508, A[24], wc26);
  not gc26 (wc26, n_578);
  or g2266 (n_1529, A[24], wc27);
  not gc27 (wc27, n_586);
  xnor g2267 (n_29, n_1070, n_442);
  or g2268 (n_1584, A[21], wc28);
  not gc28 (wc28, n_442);
  and g2269 (n_1744, wc29, n_1606);
  not gc29 (wc29, n_1607);
  or g2270 (n_2127, wc30, n_1605);
  not gc30 (wc30, n_1606);
  xnor g2271 (n_581, n_1506, A[24]);
  and g2272 (n_1737, wc31, n_74);
  not gc31 (wc31, A[24]);
  or g2273 (n_1738, wc32, n_74);
  not gc32 (wc32, A[24]);
  not g2274 (Z[2], n_2124);
  or g2275 (n_1216, A[5], wc33);
  not gc33 (wc33, n_433);
  or g2276 (n_1449, A[24], wc34);
  not gc34 (wc34, n_545);
  or g2277 (n_1545, A[18], wc35);
  not gc35 (wc35, n_596);
  or g2280 (n_2128, wc36, n_1615);
  not gc36 (wc36, n_1610);
  or g2281 (n_2235, wc37, n_1739);
  not gc37 (wc37, n_1736);
  or g2282 (n_1336, A[24], wc38);
  not gc38 (wc38, n_490);
  and g2283 (n_1746, wc39, n_1612);
  not gc39 (wc39, n_1613);
  or g2284 (n_1853, n_1615, n_1744);
  or g2285 (n_1854, n_1744, wc40);
  not gc40 (wc40, n_1749);
  xor g2286 (Z[3], n_1604, n_2127);
  xor g2287 (Z[4], n_1744, n_2128);
  or g2288 (n_2131, wc41, n_1611);
  not gc41 (wc41, n_1612);
  or g2289 (n_2238, wc42, n_1737);
  not gc42 (wc42, n_1738);
  xnor g2290 (n_1334, n_489, A[24]);
  or g2291 (n_1335, A[24], wc43);
  not gc43 (wc43, n_489);
  and g2292 (n_1753, wc44, n_1618);
  not gc44 (wc44, n_1619);
  or g2293 (n_1855, wc45, n_1621);
  not gc45 (wc45, n_1749);
  or g2294 (n_2133, wc46, n_1621);
  not gc46 (wc46, n_1616);
  or g2295 (n_2136, wc47, n_1617);
  not gc47 (wc47, n_1618);
  or g2296 (n_2233, wc48, n_1731);
  not gc48 (wc48, n_1732);
  and g2297 (n_1857, wc49, n_1616);
  not gc49 (wc49, n_1747);
  and g2298 (n_1754, wc50, n_1751);
  not gc50 (wc50, n_1746);
  or g2299 (n_2137, wc51, n_1627);
  not gc51 (wc51, n_1622);
  or g2300 (n_2227, wc52, n_1725);
  not gc52 (wc52, n_1726);
  xnor g2301 (n_1154, n_400, A[24]);
  or g2302 (n_1155, A[24], wc53);
  not gc53 (wc53, n_400);
  xnor g2303 (n_1302, n_474, A[24]);
  or g2304 (n_1303, A[24], wc54);
  not gc54 (wc54, n_474);
  and g2305 (n_1846, wc55, n_1732);
  not gc55 (wc55, n_1733);
  and g2306 (n_1861, wc56, n_1753);
  not gc56 (wc56, n_1754);
  or g2307 (n_1930, wc57, n_1739);
  not gc57 (wc57, n_1849);
  or g2308 (n_1858, n_1744, n_1855);
  or g2309 (n_1862, n_1859, n_1744);
  or g2310 (n_2230, wc58, n_1735);
  not gc58 (wc58, n_1730);
  or g2311 (n_1068, A[24], wc59);
  not gc59 (wc59, n_357);
  and g2312 (n_1756, wc60, n_1624);
  not gc60 (wc60, n_1625);
  or g2313 (n_2140, wc61, n_1623);
  not gc61 (wc61, n_1624);
  xnor g2314 (n_363, n_1066, A[24]);
  and g2315 (n_1836, wc62, n_1720);
  not gc62 (wc62, n_1721);
  and g2316 (n_1843, wc63, n_1726);
  not gc63 (wc63, n_1727);
  or g2317 (n_1938, wc64, n_1633);
  not gc64 (wc64, n_1759);
  or g2318 (n_2000, wc65, n_1729);
  not gc65 (wc65, n_1839);
  and g2319 (n_1931, wc66, n_1736);
  not gc66 (wc66, n_1847);
  or g2320 (n_1936, wc67, n_1627);
  not gc67 (wc67, n_1934);
  or g2321 (n_2142, wc68, n_1633);
  not gc68 (wc68, n_1628);
  or g2322 (n_2217, wc69, n_1713);
  not gc69 (wc69, n_1714);
  or g2323 (n_2219, wc70, n_1723);
  not gc70 (wc70, n_1718);
  or g2324 (n_2222, wc71, n_1719);
  not gc71 (wc71, n_1720);
  or g2325 (n_2224, wc72, n_1729);
  not gc72 (wc72, n_1724);
  and g2326 (n_1763, wc73, n_1630);
  not gc73 (wc73, n_1631);
  and g2327 (n_1940, wc74, n_1628);
  not gc74 (wc74, n_1757);
  and g2328 (n_1844, wc75, n_1841);
  not gc75 (wc75, n_1836);
  and g2329 (n_2013, wc76, n_1849);
  not gc76 (wc76, n_1926);
  or g2330 (n_2145, wc77, n_1629);
  not gc77 (wc77, n_1630);
  and g2331 (n_1766, wc78, n_1636);
  not gc78 (wc78, n_1637);
  and g2332 (n_1826, wc79, n_1708);
  not gc79 (wc79, n_1709);
  and g2333 (n_1833, wc80, n_1714);
  not gc80 (wc80, n_1715);
  and g2334 (n_1764, wc81, n_1761);
  not gc81 (wc81, n_1756);
  or g2335 (n_1870, wc82, n_1645);
  not gc82 (wc82, n_1769);
  or g2336 (n_1915, wc83, n_1717);
  not gc83 (wc83, n_1829);
  and g2337 (n_2001, wc84, n_1724);
  not gc84 (wc84, n_1837);
  and g2338 (n_1923, wc85, n_1843);
  not gc85 (wc85, n_1844);
  or g2339 (n_1941, n_1938, wc86);
  not gc86 (wc86, n_1934);
  or g2340 (n_2148, wc87, n_1639);
  not gc87 (wc87, n_1634);
  or g2341 (n_2151, wc88, n_1635);
  not gc88 (wc88, n_1636);
  or g2342 (n_2153, wc89, n_1645);
  not gc89 (wc89, n_1640);
  or g2343 (n_2209, wc90, n_1711);
  not gc90 (wc90, n_1706);
  or g2344 (n_2212, wc91, n_1707);
  not gc91 (wc91, n_1708);
  or g2345 (n_2214, wc92, n_1717);
  not gc92 (wc92, n_1712);
  and g2346 (n_1773, wc93, n_1642);
  not gc93 (wc93, n_1643);
  and g2347 (n_1863, wc94, n_1763);
  not gc94 (wc94, n_1764);
  and g2348 (n_1834, wc95, n_1831);
  not gc95 (wc95, n_1826);
  and g2349 (n_1947, wc96, n_1769);
  not gc96 (wc96, n_1866);
  and g2350 (n_1928, wc97, n_1849);
  not gc97 (wc97, n_1923);
  or g2351 (n_1943, wc98, n_1866);
  not gc98 (wc98, n_1934);
  or g2352 (n_2156, wc99, n_1641);
  not gc99 (wc99, n_1642);
  and g2353 (n_1871, wc100, n_1640);
  not gc100 (wc100, n_1767);
  and g2354 (n_1774, wc101, n_1771);
  not gc101 (wc101, n_1766);
  and g2355 (n_1916, wc102, n_1712);
  not gc102 (wc102, n_1827);
  and g2356 (n_1920, wc103, n_1833);
  not gc103 (wc103, n_1834);
  and g2357 (n_1868, wc104, n_1769);
  not gc104 (wc104, n_1863);
  and g2358 (n_2010, wc105, n_1730);
  not gc105 (wc105, n_1924);
  and g2359 (n_2015, wc106, n_1846);
  not gc106 (wc106, n_1928);
  and g2360 (n_2020, n_1931, wc107);
  not gc107 (wc107, n_1932);
  or g2361 (n_2157, wc108, n_1651);
  not gc108 (wc108, n_1646);
  and g2362 (n_1875, wc109, n_1773);
  not gc109 (wc109, n_1774);
  and g2363 (n_1945, wc110, n_1634);
  not gc110 (wc110, n_1864);
  and g2364 (n_1948, wc111, n_1766);
  not gc111 (wc111, n_1868);
  and g2365 (n_1776, wc112, n_1648);
  not gc112 (wc112, n_1649);
  and g2366 (n_1823, wc113, n_1702);
  not gc113 (wc113, n_1703);
  or g2367 (n_2027, wc114, n_1657);
  not gc114 (wc114, n_1779);
  and g2368 (n_1951, n_1871, wc115);
  not gc115 (wc115, n_1872);
  or g2369 (n_2160, wc116, n_1647);
  not gc116 (wc116, n_1648);
  or g2370 (n_2162, wc117, n_1657);
  not gc117 (wc117, n_1652);
  or g2371 (n_2203, wc118, n_1705);
  not gc118 (wc118, n_1700);
  or g2372 (n_2206, wc119, n_1701);
  not gc119 (wc119, n_1702);
  and g2373 (n_1954, n_1875, wc120);
  not gc120 (wc120, n_1876);
  or g2374 (n_2171, wc121, n_1659);
  not gc121 (wc121, n_1660);
  or g2375 (n_2173, wc122, n_1669);
  not gc122 (wc122, n_1664);
  and g2376 (n_1783, wc123, n_1654);
  not gc123 (wc123, n_1655);
  and g2377 (n_1786, wc124, n_1660);
  not gc124 (wc124, n_1661);
  and g2378 (n_1793, wc125, n_1666);
  not gc125 (wc125, n_1667);
  and g2379 (n_1813, wc126, n_1690);
  not gc126 (wc126, n_1691);
  and g2380 (n_1816, wc127, n_1696);
  not gc127 (wc127, n_1697);
  and g2381 (n_2029, wc128, n_1652);
  not gc128 (wc128, n_1777);
  or g2382 (n_1885, wc129, n_1669);
  not gc129 (wc129, n_1789);
  or g2383 (n_2079, wc130, n_1705);
  not gc130 (wc130, n_1819);
  or g2384 (n_2165, wc131, n_1653);
  not gc131 (wc131, n_1654);
  or g2385 (n_2168, wc132, n_1663);
  not gc132 (wc132, n_1658);
  or g2386 (n_2176, wc133, n_1665);
  not gc133 (wc133, n_1666);
  or g2387 (n_2178, wc134, n_1675);
  not gc134 (wc134, n_1670);
  or g2388 (n_2194, wc135, n_1693);
  not gc135 (wc135, n_1688);
  or g2389 (n_2197, wc136, n_1689);
  not gc136 (wc136, n_1690);
  or g2390 (n_2198, wc137, n_1699);
  not gc137 (wc137, n_1694);
  or g2391 (n_2201, wc138, n_1695);
  not gc138 (wc138, n_1696);
  and g2392 (n_1796, wc139, n_1672);
  not gc139 (wc139, n_1673);
  and g2393 (n_1803, wc140, n_1678);
  not gc140 (wc140, n_1679);
  and g2394 (n_1784, wc141, n_1781);
  not gc141 (wc141, n_1776);
  and g2395 (n_1794, wc142, n_1791);
  not gc142 (wc142, n_1786);
  or g2396 (n_1964, wc143, n_1681);
  not gc143 (wc143, n_1799);
  and g2397 (n_1824, wc144, n_1821);
  not gc144 (wc144, n_1816);
  and g2398 (n_2036, wc145, n_1789);
  not gc145 (wc145, n_1881);
  and g2399 (n_2088, wc146, n_1829);
  not gc146 (wc146, n_1911);
  or g2400 (n_2025, wc147, n_1651);
  not gc147 (wc147, n_2023);
  or g2401 (n_2030, n_2027, wc148);
  not gc148 (wc148, n_2023);
  or g2402 (n_2181, wc149, n_1671);
  not gc149 (wc149, n_1672);
  or g2403 (n_2183, wc150, n_1681);
  not gc150 (wc150, n_1676);
  or g2404 (n_2186, wc151, n_1677);
  not gc151 (wc151, n_1678);
  and g2405 (n_1806, wc152, n_1684);
  not gc152 (wc152, n_1685);
  and g2406 (n_1878, wc153, n_1783);
  not gc153 (wc153, n_1784);
  and g2407 (n_1886, wc154, n_1664);
  not gc154 (wc154, n_1787);
  and g2408 (n_1890, wc155, n_1793);
  not gc155 (wc155, n_1794);
  and g2409 (n_1804, wc156, n_1801);
  not gc156 (wc156, n_1796);
  or g2410 (n_1900, wc157, n_1693);
  not gc157 (wc157, n_1809);
  and g2411 (n_2081, wc158, n_1700);
  not gc158 (wc158, n_1817);
  and g2412 (n_1908, wc159, n_1823);
  not gc159 (wc159, n_1824);
  or g2413 (n_2043, wc160, n_1675);
  not gc160 (wc160, n_1959);
  or g2414 (n_2095, wc161, n_1723);
  not gc161 (wc161, n_1995);
  or g2415 (n_2103, n_2000, wc162);
  not gc162 (wc162, n_1995);
  or g2416 (n_2107, wc163, n_1926);
  not gc163 (wc163, n_1995);
  or g2417 (n_2032, wc164, n_1881);
  not gc164 (wc164, n_2023);
  or g2418 (n_2189, wc165, n_1687);
  not gc165 (wc165, n_1682);
  or g2419 (n_2192, wc166, n_1683);
  not gc166 (wc166, n_1684);
  and g2420 (n_1965, wc167, n_1676);
  not gc167 (wc167, n_1797);
  and g2421 (n_1893, wc168, n_1803);
  not gc168 (wc168, n_1804);
  and g2422 (n_1814, wc169, n_1811);
  not gc169 (wc169, n_1806);
  and g2423 (n_1883, wc170, n_1789);
  not gc170 (wc170, n_1878);
  and g2424 (n_1977, wc171, n_1809);
  not gc171 (wc171, n_1896);
  and g2425 (n_1913, wc172, n_1829);
  not gc172 (wc172, n_1908);
  or g2426 (n_2051, n_1964, wc173);
  not gc173 (wc173, n_1959);
  or g2427 (n_2055, wc174, n_1896);
  not gc174 (wc174, n_1959);
  and g2428 (n_1901, wc175, n_1688);
  not gc175 (wc175, n_1807);
  and g2429 (n_1905, wc176, n_1813);
  not gc176 (wc176, n_1814);
  and g2430 (n_2034, wc177, n_1658);
  not gc177 (wc177, n_1879);
  and g2431 (n_2037, wc178, n_1786);
  not gc178 (wc178, n_1883);
  and g2432 (n_2040, n_1886, wc179);
  not gc179 (wc179, n_1887);
  and g2433 (n_1956, n_1890, wc180);
  not gc180 (wc180, n_1891);
  and g2434 (n_1898, wc181, n_1809);
  not gc181 (wc181, n_1893);
  and g2435 (n_2086, wc182, n_1706);
  not gc182 (wc182, n_1909);
  and g2436 (n_2089, wc183, n_1826);
  not gc183 (wc183, n_1913);
  and g2437 (n_2092, n_1916, wc184);
  not gc184 (wc184, n_1917);
  and g2438 (n_1992, n_1920, wc185);
  not gc185 (wc185, n_1921);
  or g2439 (n_2046, n_2043, wc186);
  not gc186 (wc186, n_2023);
  or g2440 (n_2050, n_2047, wc187);
  not gc187 (wc187, n_2023);
  and g2441 (n_1974, wc188, n_1682);
  not gc188 (wc188, n_1894);
  and g2442 (n_1979, wc189, n_1806);
  not gc189 (wc189, n_1898);
  and g2443 (n_1962, wc190, n_1799);
  not gc190 (wc190, n_1956);
  and g2444 (n_1975, wc191, n_1972);
  not gc191 (wc191, n_1956);
  and g2445 (n_1980, wc192, n_1977);
  not gc192 (wc192, n_1956);
  and g2446 (n_1985, wc193, n_1982);
  not gc193 (wc193, n_1956);
  and g2447 (n_1990, wc194, n_1987);
  not gc194 (wc194, n_1956);
  and g2448 (n_1998, wc195, n_1839);
  not gc195 (wc195, n_1992);
  and g2449 (n_2011, wc196, n_2008);
  not gc196 (wc196, n_1992);
  and g2450 (n_2016, wc197, n_2013);
  not gc197 (wc197, n_1992);
  and g2451 (n_2021, wc198, n_2018);
  not gc198 (wc198, n_1992);
  or g2452 (n_2054, n_2051, wc199);
  not gc199 (wc199, n_2023);
  or g2453 (n_2058, n_2055, wc200);
  not gc200 (wc200, n_2023);
  or g2454 (n_2062, n_2059, wc201);
  not gc201 (wc201, n_2023);
  and g2455 (n_1984, n_1901, wc202);
  not gc202 (wc202, n_1902);
  and g2456 (n_1989, n_1905, wc203);
  not gc203 (wc203, n_1906);
  and g2457 (n_2045, wc204, n_1670);
  not gc204 (wc204, n_1957);
  and g2458 (n_2049, wc205, n_1796);
  not gc205 (wc205, n_1962);
  and g2459 (n_2053, n_1965, wc206);
  not gc206 (wc206, n_1966);
  and g2460 (n_2057, n_1893, wc207);
  not gc207 (wc207, n_1969);
  and g2461 (n_2097, wc208, n_1718);
  not gc208 (wc208, n_1993);
  and g2462 (n_2101, wc209, n_1836);
  not gc209 (wc209, n_1998);
  and g2463 (n_2105, n_2001, wc210);
  not gc210 (wc210, n_2002);
  and g2464 (n_2109, n_1923, wc211);
  not gc211 (wc211, n_2005);
  and g2465 (n_2113, wc212, n_2010);
  not gc212 (wc212, n_2011);
  and g2466 (n_2117, wc213, n_2015);
  not gc213 (wc213, n_2016);
  and g2467 (n_2121, wc214, n_2020);
  not gc214 (wc214, n_2021);
  or g2468 (n_2066, n_2063, wc215);
  not gc215 (wc215, n_2023);
  or g2469 (n_2070, n_2067, wc216);
  not gc216 (wc216, n_2023);
  or g2470 (n_2074, n_2071, wc217);
  not gc217 (wc217, n_2023);
  and g2471 (n_2061, wc218, n_1974);
  not gc218 (wc218, n_1975);
  and g2472 (n_2065, wc219, n_1979);
  not gc219 (wc219, n_1980);
  and g2473 (n_2069, n_1984, wc220);
  not gc220 (wc220, n_1985);
  and g2474 (n_2073, n_1989, wc221);
  not gc221 (wc221, n_1990);
  or g2475 (n_2077, wc222, n_1699);
  not gc222 (wc222, n_2075);
  or g2476 (n_2082, n_2079, wc223);
  not gc223 (wc223, n_2075);
  or g2477 (n_2084, wc224, n_1911);
  not gc224 (wc224, n_2075);
  or g2478 (n_2098, n_2095, wc225);
  not gc225 (wc225, n_2075);
  or g2479 (n_2102, wc226, n_2099);
  not gc226 (wc226, n_2075);
  or g2480 (n_2106, n_2103, wc227);
  not gc227 (wc227, n_2075);
  or g2481 (n_2110, n_2107, wc228);
  not gc228 (wc228, n_2075);
  or g2482 (n_2114, wc229, n_2111);
  not gc229 (wc229, n_2075);
  or g2483 (n_2118, wc230, n_2115);
  not gc230 (wc230, n_2075);
  or g2484 (n_2122, wc231, n_2119);
  not gc231 (wc231, n_2075);
endmodule

module mult_signed_const_4685_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_4685_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_4952_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_171, n_172, n_174, n_178, n_179;
  wire n_181, n_182, n_183, n_185, n_186, n_187, n_188, n_193;
  wire n_194, n_195, n_200, n_201, n_202, n_203, n_207, n_208;
  wire n_209, n_210, n_211, n_215, n_216, n_217, n_218, n_219;
  wire n_220, n_223, n_224, n_225, n_226, n_227, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_245, n_246;
  wire n_247, n_249, n_250, n_251, n_256, n_257, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_284, n_285;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_294;
  wire n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308;
  wire n_309, n_310, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_333, n_334;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_351, n_353, n_355, n_356;
  wire n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364;
  wire n_365, n_366, n_367, n_368, n_372, n_373, n_374, n_375;
  wire n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461;
  wire n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469;
  wire n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478;
  wire n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486;
  wire n_487, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_498, n_499, n_500, n_501, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_520, n_521, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_530, n_531, n_533, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550;
  wire n_551, n_552, n_553, n_554, n_555, n_558, n_559, n_560;
  wire n_561, n_562, n_563, n_564, n_565, n_566, n_570, n_571;
  wire n_572, n_573, n_574, n_575, n_576, n_577, n_579, n_581;
  wire n_582, n_583, n_584, n_585, n_586, n_588, n_589, n_590;
  wire n_591, n_592, n_593, n_596, n_597, n_598, n_599, n_600;
  wire n_604, n_605, n_606, n_607, n_609, n_610, n_611, n_612;
  wire n_613, n_615, n_623, n_624, n_625, n_626, n_627, n_628;
  wire n_629, n_630, n_631, n_632, n_633, n_634, n_635, n_636;
  wire n_637, n_638, n_639, n_640, n_641, n_642, n_647, n_648;
  wire n_649, n_650, n_651, n_652, n_653, n_654, n_657, n_658;
  wire n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_666;
  wire n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676;
  wire n_677, n_678, n_683, n_684, n_685, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_694, n_703, n_704, n_705;
  wire n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_714, n_721, n_722, n_723, n_724, n_725, n_726, n_727;
  wire n_728, n_729, n_730, n_731, n_732, n_733, n_734, n_739;
  wire n_740, n_741, n_743, n_744, n_745, n_746, n_747, n_748;
  wire n_749, n_750, n_751, n_752, n_753, n_754, n_759, n_760;
  wire n_761, n_763, n_764, n_765, n_766, n_767, n_768, n_769;
  wire n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777;
  wire n_778, n_787, n_791, n_792, n_793, n_794, n_795, n_796;
  wire n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_804;
  wire n_805, n_806, n_818, n_823, n_824, n_825, n_826, n_827;
  wire n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_841;
  wire n_843, n_844, n_845, n_846, n_847, n_848, n_849, n_850;
  wire n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858;
  wire n_859, n_860, n_861, n_862, n_874, n_875, n_876, n_877;
  wire n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885;
  wire n_886, n_887, n_888, n_889, n_890, n_891, n_892, n_893;
  wire n_894, n_903, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_930, n_939, n_943;
  wire n_944, n_946, n_947, n_948, n_949, n_950, n_951, n_952;
  wire n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960;
  wire n_961, n_962, n_963, n_964, n_965, n_966, n_973, n_975;
  wire n_976, n_977, n_978, n_979, n_980, n_982, n_983, n_984;
  wire n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992;
  wire n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000;
  wire n_1001, n_1002, n_1011, n_1015, n_1017, n_1018, n_1019, n_1020;
  wire n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028;
  wire n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036;
  wire n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1045;
  wire n_1046, n_1049, n_1050, n_1053, n_1054, n_1057, n_1058, n_1059;
  wire n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067;
  wire n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075;
  wire n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083;
  wire n_1084, n_1085, n_1086, n_1090, n_1091, n_1092, n_1093, n_1094;
  wire n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102;
  wire n_1103, n_1104, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111;
  wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119;
  wire n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127;
  wire n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1135, n_1136;
  wire n_1137, n_1138, n_1139, n_1140, n_1142, n_1143, n_1144, n_1145;
  wire n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153;
  wire n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161;
  wire n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169;
  wire n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177;
  wire n_1178, n_1179, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187;
  wire n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1195, n_1196;
  wire n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204;
  wire n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212;
  wire n_1213, n_1214, n_1218, n_1219, n_1220, n_1222, n_1223, n_1224;
  wire n_1225, n_1226, n_1227, n_1229, n_1230, n_1231, n_1232, n_1233;
  wire n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241;
  wire n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249;
  wire n_1250, n_1251, n_1253, n_1254, n_1256, n_1258, n_1259, n_1260;
  wire n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269;
  wire n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
  wire n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285;
  wire n_1286, n_1287, n_1289, n_1291, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1299, n_1300, n_1301, n_1303, n_1304, n_1305, n_1306;
  wire n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314;
  wire n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322;
  wire n_1327, n_1328, n_1329, n_1330, n_1331, n_1333, n_1335, n_1337;
  wire n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345;
  wire n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353;
  wire n_1354, n_1355, n_1356, n_1359, n_1360, n_1361, n_1362, n_1363;
  wire n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372;
  wire n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380;
  wire n_1381, n_1382, n_1385, n_1390, n_1391, n_1392, n_1393, n_1395;
  wire n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403;
  wire n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1414;
  wire n_1415, n_1416, n_1419, n_1421, n_1422, n_1423, n_1424, n_1425;
  wire n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433;
  wire n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1442, n_1446;
  wire n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454;
  wire n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462;
  wire n_1463, n_1465, n_1466, n_1471, n_1472, n_1473, n_1474, n_1475;
  wire n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1485;
  wire n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494;
  wire n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502;
  wire n_1507, n_1508, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515;
  wire n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1526;
  wire n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537;
  wire n_1538, n_1539, n_1540, n_1541, n_1543, n_1544, n_1545, n_1546;
  wire n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1554, n_1555;
  wire n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1565;
  wire n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574;
  wire n_1579, n_1580, n_1581, n_1582, n_1584, n_1585, n_1586, n_1587;
  wire n_1588, n_1589, n_1591, n_1593, n_1594, n_1605, n_1606, n_1607;
  wire n_1608, n_1610, n_1611, n_1612, n_1613, n_1614, n_1616, n_1617;
  wire n_1618, n_1619, n_1620, n_1622, n_1623, n_1624, n_1625, n_1626;
  wire n_1628, n_1629, n_1630, n_1631, n_1632, n_1634, n_1635, n_1636;
  wire n_1637, n_1638, n_1640, n_1641, n_1642, n_1643, n_1644, n_1646;
  wire n_1647, n_1648, n_1649, n_1650, n_1652, n_1653, n_1654, n_1655;
  wire n_1656, n_1658, n_1659, n_1660, n_1661, n_1662, n_1664, n_1665;
  wire n_1666, n_1667, n_1668, n_1670, n_1671, n_1672, n_1673, n_1674;
  wire n_1676, n_1677, n_1678, n_1679, n_1680, n_1682, n_1683, n_1684;
  wire n_1685, n_1686, n_1688, n_1689, n_1690, n_1691, n_1692, n_1694;
  wire n_1695, n_1696, n_1697, n_1698, n_1700, n_1701, n_1702, n_1703;
  wire n_1704, n_1706, n_1707, n_1708, n_1709, n_1710, n_1712, n_1713;
  wire n_1714, n_1715, n_1716, n_1718, n_1719, n_1720, n_1721, n_1722;
  wire n_1724, n_1725, n_1726, n_1727, n_1728, n_1730, n_1731, n_1732;
  wire n_1733, n_1734, n_1736, n_1737, n_1738, n_1739, n_1740, n_1745;
  wire n_1747, n_1748, n_1750, n_1752, n_1754, n_1755, n_1757, n_1758;
  wire n_1760, n_1762, n_1764, n_1765, n_1767, n_1768, n_1770, n_1772;
  wire n_1774, n_1775, n_1777, n_1778, n_1780, n_1782, n_1784, n_1785;
  wire n_1787, n_1788, n_1790, n_1792, n_1794, n_1795, n_1797, n_1798;
  wire n_1800, n_1802, n_1804, n_1805, n_1807, n_1808, n_1810, n_1812;
  wire n_1814, n_1815, n_1817, n_1818, n_1820, n_1822, n_1824, n_1825;
  wire n_1827, n_1828, n_1830, n_1832, n_1834, n_1835, n_1837, n_1838;
  wire n_1840, n_1842, n_1844, n_1845, n_1847, n_1848, n_1850, n_1854;
  wire n_1855, n_1856, n_1858, n_1859, n_1860, n_1862, n_1863, n_1864;
  wire n_1865, n_1867, n_1869, n_1871, n_1872, n_1873, n_1875, n_1876;
  wire n_1877, n_1879, n_1880, n_1882, n_1884, n_1886, n_1887, n_1888;
  wire n_1890, n_1891, n_1892, n_1894, n_1895, n_1897, n_1899, n_1901;
  wire n_1902, n_1903, n_1905, n_1906, n_1907, n_1909, n_1910, n_1912;
  wire n_1914, n_1916, n_1917, n_1918, n_1920, n_1921, n_1922, n_1924;
  wire n_1925, n_1927, n_1929, n_1931, n_1932, n_1933, n_1935, n_1937;
  wire n_1938, n_1939, n_1941, n_1942, n_1944, n_1945, n_1946, n_1947;
  wire n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955;
  wire n_1956, n_1957, n_1958, n_1960, n_1963, n_1965, n_1966, n_1967;
  wire n_1970, n_1973, n_1975, n_1976, n_1978, n_1980, n_1981, n_1983;
  wire n_1985, n_1986, n_1988, n_1990, n_1991, n_1993, n_1994, n_1996;
  wire n_1999, n_2001, n_2002, n_2003, n_2006, n_2009, n_2011, n_2012;
  wire n_2014, n_2016, n_2017, n_2019, n_2021, n_2022, n_2024, n_2026;
  wire n_2027, n_2028, n_2030, n_2031, n_2033, n_2034, n_2035, n_2036;
  wire n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044;
  wire n_2046, n_2047, n_2048, n_2050, n_2051, n_2052, n_2054, n_2055;
  wire n_2056, n_2058, n_2059, n_2060, n_2062, n_2063, n_2064, n_2066;
  wire n_2067, n_2068, n_2070, n_2071, n_2072, n_2074, n_2075, n_2076;
  wire n_2078, n_2079, n_2080, n_2082, n_2083, n_2085, n_2086, n_2087;
  wire n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095;
  wire n_2096, n_2098, n_2099, n_2100, n_2102, n_2103, n_2104, n_2106;
  wire n_2107, n_2108, n_2110, n_2111, n_2112, n_2114, n_2115, n_2116;
  wire n_2118, n_2119, n_2120, n_2122, n_2123, n_2125, n_2128, n_2129;
  wire n_2131, n_2132, n_2133, n_2134, n_2136, n_2137, n_2138, n_2140;
  wire n_2141, n_2142, n_2143, n_2145, n_2146, n_2148, n_2149, n_2151;
  wire n_2152, n_2153, n_2154, n_2156, n_2157, n_2158, n_2160, n_2161;
  wire n_2162, n_2163, n_2165, n_2166, n_2168, n_2169, n_2171, n_2172;
  wire n_2173, n_2174, n_2176, n_2177, n_2178, n_2179, n_2181, n_2182;
  wire n_2183, n_2184, n_2186, n_2187, n_2189, n_2190, n_2192, n_2193;
  wire n_2194, n_2195, n_2197, n_2198, n_2199, n_2201, n_2202, n_2203;
  wire n_2204, n_2206, n_2207, n_2209, n_2210, n_2212, n_2213, n_2214;
  wire n_2215, n_2217, n_2218, n_2219, n_2220, n_2222, n_2223, n_2224;
  wire n_2225, n_2227, n_2228, n_2230, n_2231, n_2233, n_2234, n_2235;
  wire n_2236, n_2238, n_2239;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_118, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_623, A[2], A[1]);
  xor g270 (n_117, n_623, n_171);
  nand g3 (n_624, A[2], A[1]);
  nand g271 (n_625, n_171, A[1]);
  nand g272 (n_626, A[2], n_171);
  nand g273 (n_68, n_624, n_625, n_626);
  xor g274 (n_627, A[2], A[3]);
  xor g275 (n_116, n_627, A[5]);
  nand g276 (n_628, A[2], A[3]);
  nand g4 (n_629, A[5], A[3]);
  nand g277 (n_630, A[2], A[5]);
  nand g278 (n_67, n_628, n_629, n_630);
  xor g279 (n_172, A[0], A[3]);
  and g280 (n_174, A[0], A[3]);
  xor g281 (n_631, A[4], n_172);
  xor g282 (n_115, n_631, A[6]);
  nand g283 (n_632, A[4], n_172);
  nand g284 (n_633, A[6], n_172);
  nand g5 (n_634, A[4], A[6]);
  nand g6 (n_66, n_632, n_633, n_634);
  xor g287 (n_635, A[4], n_118);
  xor g288 (n_69, n_635, n_174);
  nand g289 (n_636, A[4], n_118);
  nand g290 (n_637, n_174, n_118);
  nand g291 (n_638, A[4], n_174);
  nand g292 (n_178, n_636, n_637, n_638);
  xor g293 (n_639, A[5], A[7]);
  xor g294 (n_114, n_639, n_69);
  nand g295 (n_640, A[5], A[7]);
  nand g296 (n_641, n_69, A[7]);
  nand g297 (n_642, A[5], n_69);
  nand g298 (n_65, n_640, n_641, n_642);
  xor g305 (n_647, A[6], A[5]);
  xor g306 (n_179, n_647, n_117);
  nand g307 (n_648, A[6], A[5]);
  nand g308 (n_649, n_117, A[5]);
  nand g309 (n_650, A[6], n_117);
  nand g310 (n_182, n_648, n_649, n_650);
  xor g311 (n_651, A[8], n_178);
  xor g312 (n_113, n_651, n_179);
  nand g313 (n_652, A[8], n_178);
  nand g314 (n_653, n_179, n_178);
  nand g315 (n_654, A[8], n_179);
  nand g316 (n_64, n_652, n_653, n_654);
  xor g318 (n_181, n_627, A[6]);
  nand g320 (n_657, A[6], A[3]);
  nand g321 (n_658, A[2], A[6]);
  nand g322 (n_185, n_628, n_657, n_658);
  xor g323 (n_659, n_68, A[7]);
  xor g324 (n_183, n_659, A[9]);
  nand g325 (n_660, n_68, A[7]);
  nand g326 (n_661, A[9], A[7]);
  nand g327 (n_662, n_68, A[9]);
  nand g328 (n_187, n_660, n_661, n_662);
  xor g329 (n_663, n_181, n_182);
  xor g330 (n_112, n_663, n_183);
  nand g331 (n_664, n_181, n_182);
  nand g332 (n_665, n_183, n_182);
  nand g333 (n_666, n_181, n_183);
  nand g334 (n_63, n_664, n_665, n_666);
  xor g338 (n_186, n_631, A[7]);
  nand g340 (n_669, A[7], n_172);
  nand g341 (n_670, A[4], A[7]);
  nand g342 (n_70, n_632, n_669, n_670);
  xor g343 (n_671, A[8], A[10]);
  xor g344 (n_188, n_671, n_185);
  nand g345 (n_672, A[8], A[10]);
  nand g346 (n_673, n_185, A[10]);
  nand g347 (n_674, A[8], n_185);
  nand g348 (n_194, n_672, n_673, n_674);
  xor g349 (n_675, n_186, n_187);
  xor g350 (n_111, n_675, n_188);
  nand g351 (n_676, n_186, n_187);
  nand g352 (n_677, n_188, n_187);
  nand g353 (n_678, n_186, n_188);
  nand g354 (n_62, n_676, n_677, n_678);
  xor g363 (n_683, A[5], A[9]);
  xor g364 (n_193, n_683, n_69);
  nand g365 (n_684, A[5], A[9]);
  nand g366 (n_685, n_69, A[9]);
  nand g368 (n_200, n_684, n_685, n_642);
  xor g369 (n_687, A[8], A[11]);
  xor g370 (n_195, n_687, n_70);
  nand g371 (n_688, A[8], A[11]);
  nand g372 (n_689, n_70, A[11]);
  nand g373 (n_690, A[8], n_70);
  nand g374 (n_202, n_688, n_689, n_690);
  xor g375 (n_691, n_193, n_194);
  xor g376 (n_110, n_691, n_195);
  nand g377 (n_692, n_193, n_194);
  nand g378 (n_693, n_195, n_194);
  nand g379 (n_694, n_193, n_195);
  nand g380 (n_61, n_692, n_693, n_694);
  xor g393 (n_703, n_178, A[10]);
  xor g394 (n_201, n_703, A[9]);
  nand g395 (n_704, n_178, A[10]);
  nand g396 (n_705, A[9], A[10]);
  nand g397 (n_706, n_178, A[9]);
  nand g398 (n_208, n_704, n_705, n_706);
  xor g399 (n_707, A[12], n_179);
  xor g400 (n_203, n_707, n_200);
  nand g401 (n_708, A[12], n_179);
  nand g402 (n_709, n_200, n_179);
  nand g403 (n_710, A[12], n_200);
  nand g404 (n_210, n_708, n_709, n_710);
  xor g405 (n_711, n_201, n_202);
  xor g406 (n_109, n_711, n_203);
  nand g407 (n_712, n_201, n_202);
  nand g408 (n_713, n_203, n_202);
  nand g409 (n_714, n_201, n_203);
  nand g410 (n_60, n_712, n_713, n_714);
  xor g418 (n_207, n_659, A[10]);
  nand g420 (n_721, A[10], n_68);
  nand g421 (n_722, A[7], A[10]);
  nand g422 (n_215, n_660, n_721, n_722);
  xor g423 (n_723, A[11], n_181);
  xor g424 (n_209, n_723, A[13]);
  nand g425 (n_724, A[11], n_181);
  nand g426 (n_725, A[13], n_181);
  nand g427 (n_726, A[11], A[13]);
  nand g428 (n_216, n_724, n_725, n_726);
  xor g429 (n_727, n_182, n_207);
  xor g430 (n_211, n_727, n_208);
  nand g431 (n_728, n_182, n_207);
  nand g432 (n_729, n_208, n_207);
  nand g433 (n_730, n_182, n_208);
  nand g434 (n_219, n_728, n_729, n_730);
  xor g435 (n_731, n_209, n_210);
  xor g436 (n_108, n_731, n_211);
  nand g437 (n_732, n_209, n_210);
  nand g438 (n_733, n_211, n_210);
  nand g439 (n_734, n_209, n_211);
  nand g440 (n_59, n_732, n_733, n_734);
  xor g449 (n_739, A[8], A[12]);
  xor g450 (n_217, n_739, n_185);
  nand g451 (n_740, A[8], A[12]);
  nand g452 (n_741, n_185, A[12]);
  nand g454 (n_73, n_740, n_741, n_674);
  xor g455 (n_743, A[14], A[11]);
  xor g456 (n_218, n_743, n_186);
  nand g457 (n_744, A[14], A[11]);
  nand g458 (n_745, n_186, A[11]);
  nand g459 (n_746, A[14], n_186);
  nand g460 (n_223, n_744, n_745, n_746);
  xor g461 (n_747, n_215, n_216);
  xor g462 (n_220, n_747, n_217);
  nand g463 (n_748, n_215, n_216);
  nand g464 (n_749, n_217, n_216);
  nand g465 (n_750, n_215, n_217);
  nand g466 (n_226, n_748, n_749, n_750);
  xor g467 (n_751, n_218, n_219);
  xor g468 (n_107, n_751, n_220);
  nand g469 (n_752, n_218, n_219);
  nand g470 (n_753, n_220, n_219);
  nand g471 (n_754, n_218, n_220);
  nand g472 (n_58, n_752, n_753, n_754);
  xor g481 (n_759, A[5], A[8]);
  xor g482 (n_72, n_759, A[9]);
  nand g483 (n_760, A[5], A[8]);
  nand g484 (n_761, A[9], A[8]);
  nand g486 (n_232, n_760, n_761, n_684);
  xor g487 (n_763, n_69, A[12]);
  xor g488 (n_224, n_763, A[13]);
  nand g489 (n_764, n_69, A[12]);
  nand g490 (n_765, A[13], A[12]);
  nand g491 (n_766, n_69, A[13]);
  nand g492 (n_234, n_764, n_765, n_766);
  xor g493 (n_767, n_70, A[15]);
  xor g494 (n_225, n_767, n_72);
  nand g495 (n_768, n_70, A[15]);
  nand g496 (n_769, n_72, A[15]);
  nand g497 (n_770, n_70, n_72);
  nand g498 (n_236, n_768, n_769, n_770);
  xor g499 (n_771, n_73, n_223);
  xor g500 (n_227, n_771, n_224);
  nand g501 (n_772, n_73, n_223);
  nand g502 (n_773, n_224, n_223);
  nand g503 (n_774, n_73, n_224);
  nand g504 (n_238, n_772, n_773, n_774);
  xor g505 (n_775, n_225, n_226);
  xor g506 (n_106, n_775, n_227);
  nand g507 (n_776, n_225, n_226);
  nand g508 (n_777, n_227, n_226);
  nand g509 (n_778, n_225, n_227);
  nand g510 (n_57, n_776, n_777, n_778);
  xor g523 (n_787, A[9], n_178);
  xor g524 (n_233, n_787, A[10]);
  xor g529 (n_791, A[14], A[13]);
  xor g530 (n_235, n_791, n_179);
  nand g531 (n_792, A[14], A[13]);
  nand g532 (n_793, n_179, A[13]);
  nand g533 (n_794, A[14], n_179);
  nand g534 (n_246, n_792, n_793, n_794);
  xor g535 (n_795, n_232, n_233);
  xor g536 (n_237, n_795, n_234);
  nand g537 (n_796, n_232, n_233);
  nand g538 (n_797, n_234, n_233);
  nand g539 (n_798, n_232, n_234);
  nand g540 (n_247, n_796, n_797, n_798);
  xor g541 (n_799, A[16], n_235);
  xor g542 (n_239, n_799, n_236);
  nand g543 (n_800, A[16], n_235);
  nand g544 (n_801, n_236, n_235);
  nand g545 (n_802, A[16], n_236);
  nand g546 (n_250, n_800, n_801, n_802);
  xor g547 (n_803, n_237, n_238);
  xor g548 (n_105, n_803, n_239);
  nand g549 (n_804, n_237, n_238);
  nand g550 (n_805, n_239, n_238);
  nand g551 (n_806, n_237, n_239);
  nand g552 (n_56, n_804, n_805, n_806);
  xor g566 (n_245, n_743, n_181);
  nand g569 (n_818, A[14], n_181);
  nand g570 (n_256, n_744, n_724, n_818);
  xor g577 (n_823, A[15], A[17]);
  xor g578 (n_249, n_823, n_245);
  nand g579 (n_824, A[15], A[17]);
  nand g580 (n_825, n_245, A[17]);
  nand g581 (n_826, A[15], n_245);
  nand g582 (n_261, n_824, n_825, n_826);
  xor g583 (n_827, n_246, n_247);
  xor g584 (n_251, n_827, n_211);
  nand g585 (n_828, n_246, n_247);
  nand g586 (n_829, n_211, n_247);
  nand g587 (n_830, n_246, n_211);
  nand g588 (n_263, n_828, n_829, n_830);
  xor g589 (n_831, n_249, n_250);
  xor g590 (n_104, n_831, n_251);
  nand g591 (n_832, n_249, n_250);
  nand g592 (n_833, n_251, n_250);
  nand g593 (n_834, n_249, n_251);
  nand g594 (n_55, n_832, n_833, n_834);
  xor g604 (n_257, n_687, n_185);
  nand g606 (n_841, n_185, A[11]);
  nand g608 (n_269, n_688, n_841, n_674);
  xor g609 (n_843, A[12], A[18]);
  xor g610 (n_259, n_843, n_186);
  nand g611 (n_844, A[12], A[18]);
  nand g612 (n_845, n_186, A[18]);
  nand g613 (n_846, A[12], n_186);
  nand g614 (n_270, n_844, n_845, n_846);
  xor g615 (n_847, A[15], n_215);
  xor g616 (n_260, n_847, n_256);
  nand g617 (n_848, A[15], n_215);
  nand g618 (n_849, n_256, n_215);
  nand g619 (n_850, A[15], n_256);
  nand g620 (n_273, n_848, n_849, n_850);
  xor g621 (n_851, A[16], n_257);
  xor g622 (n_262, n_851, n_219);
  nand g623 (n_852, A[16], n_257);
  nand g624 (n_853, n_219, n_257);
  nand g625 (n_854, A[16], n_219);
  nand g626 (n_275, n_852, n_853, n_854);
  xor g627 (n_855, n_259, n_260);
  xor g628 (n_264, n_855, n_261);
  nand g629 (n_856, n_259, n_260);
  nand g630 (n_857, n_261, n_260);
  nand g631 (n_858, n_259, n_261);
  nand g632 (n_277, n_856, n_857, n_858);
  xor g633 (n_859, n_262, n_263);
  xor g634 (n_103, n_859, n_264);
  nand g635 (n_860, n_262, n_263);
  nand g636 (n_861, n_264, n_263);
  nand g637 (n_862, n_262, n_264);
  nand g638 (n_54, n_860, n_861, n_862);
  xor g654 (n_271, n_739, A[13]);
  nand g657 (n_874, A[8], A[13]);
  nand g658 (n_284, n_740, n_765, n_874);
  xor g659 (n_875, n_70, A[19]);
  xor g660 (n_272, n_875, n_193);
  nand g661 (n_876, n_70, A[19]);
  nand g662 (n_877, n_193, A[19]);
  nand g663 (n_878, n_70, n_193);
  nand g664 (n_287, n_876, n_877, n_878);
  xor g665 (n_879, n_269, n_270);
  xor g666 (n_274, n_879, A[17]);
  nand g667 (n_880, n_269, n_270);
  nand g668 (n_881, A[17], n_270);
  nand g669 (n_882, n_269, A[17]);
  nand g670 (n_289, n_880, n_881, n_882);
  xor g671 (n_883, n_271, A[16]);
  xor g672 (n_276, n_883, n_272);
  nand g673 (n_884, n_271, A[16]);
  nand g674 (n_885, n_272, A[16]);
  nand g675 (n_886, n_271, n_272);
  nand g676 (n_291, n_884, n_885, n_886);
  xor g677 (n_887, n_273, n_274);
  xor g678 (n_278, n_887, n_275);
  nand g679 (n_888, n_273, n_274);
  nand g680 (n_889, n_275, n_274);
  nand g681 (n_890, n_273, n_275);
  nand g682 (n_293, n_888, n_889, n_890);
  xor g683 (n_891, n_276, n_277);
  xor g684 (n_102, n_891, n_278);
  nand g685 (n_892, n_276, n_277);
  nand g686 (n_893, n_278, n_277);
  nand g687 (n_894, n_276, n_278);
  nand g688 (n_53, n_892, n_893, n_894);
  xor g701 (n_903, A[10], A[9]);
  xor g702 (n_285, n_903, n_178);
  xor g713 (n_911, A[18], n_200);
  xor g714 (n_288, n_911, n_284);
  nand g715 (n_912, A[18], n_200);
  nand g716 (n_913, n_284, n_200);
  nand g717 (n_914, A[18], n_284);
  nand g718 (n_303, n_912, n_913, n_914);
  xor g719 (n_915, A[20], n_285);
  xor g720 (n_290, n_915, A[17]);
  nand g721 (n_916, A[20], n_285);
  nand g722 (n_917, A[17], n_285);
  nand g723 (n_918, A[20], A[17]);
  nand g724 (n_305, n_916, n_917, n_918);
  xor g725 (n_919, n_235, n_287);
  xor g726 (n_292, n_919, n_288);
  nand g727 (n_920, n_235, n_287);
  nand g728 (n_921, n_288, n_287);
  nand g729 (n_922, n_235, n_288);
  nand g730 (n_307, n_920, n_921, n_922);
  xor g731 (n_923, n_289, n_290);
  xor g732 (n_294, n_923, n_291);
  nand g733 (n_924, n_289, n_290);
  nand g734 (n_925, n_291, n_290);
  nand g735 (n_926, n_289, n_291);
  nand g736 (n_310, n_924, n_925, n_926);
  xor g737 (n_927, n_292, n_293);
  xor g738 (n_101, n_927, n_294);
  nand g739 (n_928, n_292, n_293);
  nand g740 (n_929, n_294, n_293);
  nand g741 (n_930, n_292, n_294);
  nand g742 (n_52, n_928, n_929, n_930);
  xor g755 (n_939, n_181, A[14]);
  xor g756 (n_301, n_939, A[11]);
  xor g761 (n_943, A[18], n_182);
  xor g762 (n_302, n_943, n_207);
  nand g763 (n_944, A[18], n_182);
  nand g765 (n_946, A[18], n_207);
  nand g766 (n_319, n_944, n_728, n_946);
  xor g767 (n_947, A[15], A[19]);
  xor g768 (n_304, n_947, n_208);
  nand g769 (n_948, A[15], A[19]);
  nand g770 (n_949, n_208, A[19]);
  nand g771 (n_950, A[15], n_208);
  nand g772 (n_317, n_948, n_949, n_950);
  xor g773 (n_951, A[21], n_246);
  xor g774 (n_306, n_951, n_301);
  nand g775 (n_952, A[21], n_246);
  nand g776 (n_953, n_301, n_246);
  nand g777 (n_954, A[21], n_301);
  nand g778 (n_321, n_952, n_953, n_954);
  xor g779 (n_955, n_302, n_303);
  xor g780 (n_308, n_955, n_304);
  nand g781 (n_956, n_302, n_303);
  nand g782 (n_957, n_304, n_303);
  nand g783 (n_958, n_302, n_304);
  nand g784 (n_323, n_956, n_957, n_958);
  xor g785 (n_959, n_305, n_306);
  xor g786 (n_309, n_959, n_307);
  nand g787 (n_960, n_305, n_306);
  nand g788 (n_961, n_307, n_306);
  nand g789 (n_962, n_305, n_307);
  nand g790 (n_326, n_960, n_961, n_962);
  xor g791 (n_963, n_308, n_309);
  xor g792 (n_100, n_963, n_310);
  nand g793 (n_964, n_308, n_309);
  nand g794 (n_965, n_310, n_309);
  nand g795 (n_966, n_308, n_310);
  nand g796 (n_51, n_964, n_965, n_966);
  xor g806 (n_316, n_739, A[11]);
  nand g808 (n_973, A[11], A[12]);
  nand g810 (n_333, n_740, n_973, n_688);
  xor g811 (n_975, n_185, n_186);
  xor g812 (n_318, n_975, A[15]);
  nand g813 (n_976, n_185, n_186);
  nand g814 (n_977, A[15], n_186);
  nand g815 (n_978, n_185, A[15]);
  nand g816 (n_335, n_976, n_977, n_978);
  xor g817 (n_979, A[19], n_215);
  xor g818 (n_320, n_979, n_256);
  nand g819 (n_980, A[19], n_215);
  nand g821 (n_982, A[19], n_256);
  nand g822 (n_336, n_980, n_849, n_982);
  xor g823 (n_983, A[20], A[22]);
  xor g824 (n_322, n_983, n_316);
  nand g825 (n_984, A[20], A[22]);
  nand g826 (n_985, n_316, A[22]);
  nand g827 (n_986, A[20], n_316);
  nand g828 (n_337, n_984, n_985, n_986);
  xor g829 (n_987, A[16], n_317);
  xor g830 (n_324, n_987, n_318);
  nand g831 (n_988, A[16], n_317);
  nand g832 (n_989, n_318, n_317);
  nand g833 (n_990, A[16], n_318);
  nand g834 (n_340, n_988, n_989, n_990);
  xor g835 (n_991, n_319, n_320);
  xor g836 (n_325, n_991, n_321);
  nand g837 (n_992, n_319, n_320);
  nand g838 (n_993, n_321, n_320);
  nand g839 (n_994, n_319, n_321);
  nand g840 (n_343, n_992, n_993, n_994);
  xor g841 (n_995, n_322, n_323);
  xor g842 (n_327, n_995, n_324);
  nand g843 (n_996, n_322, n_323);
  nand g844 (n_997, n_324, n_323);
  nand g845 (n_998, n_322, n_324);
  nand g846 (n_345, n_996, n_997, n_998);
  xor g847 (n_999, n_325, n_326);
  xor g848 (n_99, n_999, n_327);
  nand g849 (n_1000, n_325, n_326);
  nand g850 (n_1001, n_327, n_326);
  nand g851 (n_1002, n_325, n_327);
  nand g852 (n_50, n_1000, n_1001, n_1002);
  xor g867 (n_1011, n_69, A[13]);
  xor g868 (n_334, n_1011, A[12]);
  xor g873 (n_1015, n_70, n_72);
  xor g874 (n_339, n_1015, n_333);
  nand g876 (n_1017, n_333, n_72);
  nand g877 (n_1018, n_70, n_333);
  nand g878 (n_359, n_770, n_1017, n_1018);
  xor g879 (n_1019, A[21], A[20]);
  xor g880 (n_338, n_1019, A[23]);
  nand g881 (n_1020, A[21], A[20]);
  nand g882 (n_1021, A[23], A[20]);
  nand g883 (n_1022, A[21], A[23]);
  nand g884 (n_358, n_1020, n_1021, n_1022);
  xor g885 (n_1023, A[17], n_334);
  xor g886 (n_341, n_1023, A[16]);
  nand g887 (n_1024, A[17], n_334);
  nand g888 (n_1025, A[16], n_334);
  nand g889 (n_1026, A[17], A[16]);
  nand g890 (n_360, n_1024, n_1025, n_1026);
  xor g891 (n_1027, n_335, n_336);
  xor g892 (n_342, n_1027, n_337);
  nand g893 (n_1028, n_335, n_336);
  nand g894 (n_1029, n_337, n_336);
  nand g895 (n_1030, n_335, n_337);
  nand g896 (n_363, n_1028, n_1029, n_1030);
  xor g897 (n_1031, n_338, n_339);
  xor g898 (n_344, n_1031, n_340);
  nand g899 (n_1032, n_338, n_339);
  nand g900 (n_1033, n_340, n_339);
  nand g901 (n_1034, n_338, n_340);
  nand g902 (n_365, n_1032, n_1033, n_1034);
  xor g903 (n_1035, n_341, n_342);
  xor g904 (n_346, n_1035, n_343);
  nand g905 (n_1036, n_341, n_342);
  nand g906 (n_1037, n_343, n_342);
  nand g907 (n_1038, n_341, n_343);
  nand g908 (n_367, n_1036, n_1037, n_1038);
  xor g909 (n_1039, n_344, n_345);
  xor g910 (n_98, n_1039, n_346);
  nand g911 (n_1040, n_344, n_345);
  nand g912 (n_1041, n_346, n_345);
  nand g913 (n_1042, n_344, n_346);
  nand g914 (n_49, n_1040, n_1041, n_1042);
  xor g917 (n_1043, A[1], n_171);
  nand g922 (n_372, n_625, n_1045, n_1046);
  xor g924 (n_353, n_647, n_178);
  nand g926 (n_1049, n_178, A[6]);
  nand g927 (n_1050, A[5], n_178);
  nand g928 (n_374, n_648, n_1049, n_1050);
  xor g930 (n_355, n_903, n_351);
  nand g932 (n_1053, n_351, A[9]);
  nand g933 (n_1054, A[10], n_351);
  nand g934 (n_375, n_705, n_1053, n_1054);
  xor g936 (n_356, n_791, A[18]);
  nand g938 (n_1057, A[18], A[13]);
  nand g939 (n_1058, A[14], A[18]);
  nand g940 (n_378, n_792, n_1057, n_1058);
  xor g942 (n_357, n_1059, n_353);
  nand g945 (n_1062, n_232, n_353);
  nand g946 (n_379, n_1060, n_1061, n_1062);
  xor g947 (n_1063, A[22], n_234);
  xor g948 (n_361, n_1063, A[21]);
  nand g949 (n_1064, A[22], n_234);
  nand g950 (n_1065, A[21], n_234);
  nand g951 (n_1066, A[22], A[21]);
  nand g952 (n_382, n_1064, n_1065, n_1066);
  xor g953 (n_1067, n_355, n_356);
  xor g954 (n_362, n_1067, A[17]);
  nand g955 (n_1068, n_355, n_356);
  nand g956 (n_1069, A[17], n_356);
  nand g957 (n_1070, n_355, A[17]);
  nand g958 (n_384, n_1068, n_1069, n_1070);
  xor g959 (n_1071, n_357, n_358);
  xor g960 (n_364, n_1071, n_359);
  nand g961 (n_1072, n_357, n_358);
  nand g962 (n_1073, n_359, n_358);
  nand g963 (n_1074, n_357, n_359);
  nand g964 (n_386, n_1072, n_1073, n_1074);
  xor g965 (n_1075, n_360, n_361);
  xor g966 (n_366, n_1075, n_362);
  nand g967 (n_1076, n_360, n_361);
  nand g968 (n_1077, n_362, n_361);
  nand g969 (n_1078, n_360, n_362);
  nand g970 (n_388, n_1076, n_1077, n_1078);
  xor g971 (n_1079, n_363, n_364);
  xor g972 (n_368, n_1079, n_365);
  nand g973 (n_1080, n_363, n_364);
  nand g974 (n_1081, n_365, n_364);
  nand g975 (n_1082, n_363, n_365);
  nand g976 (n_391, n_1080, n_1081, n_1082);
  xor g977 (n_1083, n_366, n_367);
  xor g978 (n_97, n_1083, n_368);
  nand g979 (n_1084, n_366, n_367);
  nand g980 (n_1085, n_368, n_367);
  nand g981 (n_1086, n_366, n_368);
  nand g982 (n_48, n_1084, n_1085, n_1086);
  xor g991 (n_1091, A[6], A[7]);
  xor g992 (n_376, n_1091, n_372);
  nand g993 (n_1092, A[6], A[7]);
  nand g994 (n_1093, n_372, A[7]);
  nand g995 (n_1094, A[6], n_372);
  nand g996 (n_395, n_1092, n_1093, n_1094);
  xor g997 (n_1095, A[10], n_373);
  xor g998 (n_377, n_1095, A[14]);
  nand g999 (n_1096, A[10], n_373);
  nand g1000 (n_1097, A[14], n_373);
  nand g1001 (n_1098, A[10], A[14]);
  nand g1002 (n_397, n_1096, n_1097, n_1098);
  xor g1003 (n_1099, A[11], A[18]);
  xor g1004 (n_380, n_1099, n_374);
  nand g1005 (n_1100, A[11], A[18]);
  nand g1006 (n_1101, n_374, A[18]);
  nand g1007 (n_1102, A[11], n_374);
  nand g1008 (n_399, n_1100, n_1101, n_1102);
  xor g1009 (n_1103, n_375, A[19]);
  xor g1010 (n_381, n_1103, A[15]);
  nand g1011 (n_1104, n_375, A[19]);
  nand g1013 (n_1106, n_375, A[15]);
  nand g1014 (n_400, n_1104, n_948, n_1106);
  xor g1015 (n_1107, n_376, A[22]);
  xor g1016 (n_383, n_1107, n_377);
  nand g1017 (n_1108, n_376, A[22]);
  nand g1018 (n_1109, n_377, A[22]);
  nand g1019 (n_1110, n_376, n_377);
  nand g1020 (n_403, n_1108, n_1109, n_1110);
  xor g1021 (n_1111, A[23], n_378);
  xor g1022 (n_385, n_1111, n_379);
  nand g1023 (n_1112, A[23], n_378);
  nand g1024 (n_1113, n_379, n_378);
  nand g1025 (n_1114, A[23], n_379);
  nand g1026 (n_405, n_1112, n_1113, n_1114);
  xor g1027 (n_1115, n_380, n_381);
  xor g1028 (n_387, n_1115, n_382);
  nand g1029 (n_1116, n_380, n_381);
  nand g1030 (n_1117, n_382, n_381);
  nand g1031 (n_1118, n_380, n_382);
  nand g1032 (n_406, n_1116, n_1117, n_1118);
  xor g1033 (n_1119, n_383, n_384);
  xor g1034 (n_389, n_1119, n_385);
  nand g1035 (n_1120, n_383, n_384);
  nand g1036 (n_1121, n_385, n_384);
  nand g1037 (n_1122, n_383, n_385);
  nand g1038 (n_409, n_1120, n_1121, n_1122);
  xor g1039 (n_1123, n_386, n_387);
  xor g1040 (n_390, n_1123, n_388);
  nand g1041 (n_1124, n_386, n_387);
  nand g1042 (n_1125, n_388, n_387);
  nand g1043 (n_1126, n_386, n_388);
  nand g1044 (n_412, n_1124, n_1125, n_1126);
  xor g1045 (n_1127, n_389, n_390);
  xor g1046 (n_96, n_1127, n_391);
  nand g1047 (n_1128, n_389, n_390);
  nand g1048 (n_1129, n_391, n_390);
  nand g1049 (n_1130, n_389, n_391);
  nand g1050 (n_47, n_1128, n_1129, n_1130);
  xor g1051 (n_1131, A[3], A[4]);
  xor g1052 (n_394, n_1131, A[2]);
  nand g1053 (n_1132, A[3], A[4]);
  nand g1054 (n_1133, A[2], A[4]);
  nand g1056 (n_413, n_1132, n_1133, n_628);
  xor g1057 (n_1135, A[7], n_393);
  xor g1058 (n_396, n_1135, A[8]);
  nand g1059 (n_1136, A[7], n_393);
  nand g1060 (n_1137, A[8], n_393);
  nand g1061 (n_1138, A[7], A[8]);
  nand g1062 (n_415, n_1136, n_1137, n_1138);
  xor g1063 (n_1139, n_394, A[11]);
  xor g1064 (n_398, n_1139, A[12]);
  nand g1065 (n_1140, n_394, A[11]);
  nand g1067 (n_1142, n_394, A[12]);
  nand g1068 (n_417, n_1140, n_973, n_1142);
  xor g1069 (n_1143, n_395, A[19]);
  xor g1070 (n_402, n_1143, n_396);
  nand g1071 (n_1144, n_395, A[19]);
  nand g1072 (n_1145, n_396, A[19]);
  nand g1073 (n_1146, n_395, n_396);
  nand g1074 (n_418, n_1144, n_1145, n_1146);
  xor g1076 (n_401, n_1147, A[23]);
  nand g1078 (n_1149, A[23], A[15]);
  nand g1080 (n_420, n_1148, n_1149, n_1150);
  xor g1081 (n_1151, n_397, A[20]);
  xor g1082 (n_404, n_1151, n_398);
  nand g1083 (n_1152, n_397, A[20]);
  nand g1084 (n_1153, n_398, A[20]);
  nand g1085 (n_1154, n_397, n_398);
  nand g1086 (n_423, n_1152, n_1153, n_1154);
  xor g1087 (n_1155, A[16], n_399);
  xor g1088 (n_407, n_1155, n_400);
  nand g1089 (n_1156, A[16], n_399);
  nand g1090 (n_1157, n_400, n_399);
  nand g1091 (n_1158, A[16], n_400);
  nand g1092 (n_424, n_1156, n_1157, n_1158);
  xor g1093 (n_1159, n_401, n_402);
  xor g1094 (n_408, n_1159, n_403);
  nand g1095 (n_1160, n_401, n_402);
  nand g1096 (n_1161, n_403, n_402);
  nand g1097 (n_1162, n_401, n_403);
  nand g1098 (n_426, n_1160, n_1161, n_1162);
  xor g1099 (n_1163, n_404, n_405);
  xor g1100 (n_410, n_1163, n_406);
  nand g1101 (n_1164, n_404, n_405);
  nand g1102 (n_1165, n_406, n_405);
  nand g1103 (n_1166, n_404, n_406);
  nand g1104 (n_429, n_1164, n_1165, n_1166);
  xor g1105 (n_1167, n_407, n_408);
  xor g1106 (n_411, n_1167, n_409);
  nand g1107 (n_1168, n_407, n_408);
  nand g1108 (n_1169, n_409, n_408);
  nand g1109 (n_1170, n_407, n_409);
  nand g1110 (n_430, n_1168, n_1169, n_1170);
  xor g1111 (n_1171, n_410, n_411);
  xor g1112 (n_95, n_1171, n_412);
  nand g1113 (n_1172, n_410, n_411);
  nand g1114 (n_1173, n_412, n_411);
  nand g1115 (n_1174, n_410, n_412);
  nand g1116 (n_46, n_1172, n_1173, n_1174);
  xor g1117 (n_1175, A[4], A[5]);
  xor g1118 (n_414, n_1175, n_413);
  nand g1119 (n_1176, A[4], A[5]);
  nand g1120 (n_1177, n_413, A[5]);
  nand g1121 (n_1178, A[4], n_413);
  nand g1122 (n_434, n_1176, n_1177, n_1178);
  xor g1123 (n_1179, A[9], A[8]);
  xor g1124 (n_416, n_1179, A[13]);
  nand g1127 (n_1182, A[9], A[13]);
  nand g1128 (n_436, n_761, n_874, n_1182);
  xor g1129 (n_1183, A[12], n_414);
  xor g1130 (n_419, n_1183, n_415);
  nand g1131 (n_1184, A[12], n_414);
  nand g1132 (n_1185, n_415, n_414);
  nand g1133 (n_1186, A[12], n_415);
  nand g1134 (n_438, n_1184, n_1185, n_1186);
  xor g1136 (n_422, n_1187, n_416);
  nand g1138 (n_1189, n_416, A[21]);
  nand g1140 (n_439, n_1188, n_1189, n_1190);
  xor g1141 (n_1191, A[20], n_417);
  xor g1142 (n_421, n_1191, A[17]);
  nand g1143 (n_1192, A[20], n_417);
  nand g1144 (n_1193, A[17], n_417);
  nand g1146 (n_442, n_1192, n_1193, n_918);
  xor g1147 (n_1195, A[16], n_418);
  xor g1148 (n_425, n_1195, n_419);
  nand g1149 (n_1196, A[16], n_418);
  nand g1150 (n_1197, n_419, n_418);
  nand g1151 (n_1198, A[16], n_419);
  nand g1152 (n_443, n_1196, n_1197, n_1198);
  xor g1153 (n_1199, n_420, n_421);
  xor g1154 (n_427, n_1199, n_422);
  nand g1155 (n_1200, n_420, n_421);
  nand g1156 (n_1201, n_422, n_421);
  nand g1157 (n_1202, n_420, n_422);
  nand g1158 (n_445, n_1200, n_1201, n_1202);
  xor g1159 (n_1203, n_423, n_424);
  xor g1160 (n_428, n_1203, n_425);
  nand g1161 (n_1204, n_423, n_424);
  nand g1162 (n_1205, n_425, n_424);
  nand g1163 (n_1206, n_423, n_425);
  nand g1164 (n_448, n_1204, n_1205, n_1206);
  xor g1165 (n_1207, n_426, n_427);
  xor g1166 (n_431, n_1207, n_428);
  nand g1167 (n_1208, n_426, n_427);
  nand g1168 (n_1209, n_428, n_427);
  nand g1169 (n_1210, n_426, n_428);
  nand g1170 (n_450, n_1208, n_1209, n_1210);
  xor g1171 (n_1211, n_429, n_430);
  xor g1172 (n_94, n_1211, n_431);
  nand g1173 (n_1212, n_429, n_430);
  nand g1174 (n_1213, n_431, n_430);
  nand g1175 (n_1214, n_429, n_431);
  nand g1176 (n_45, n_1212, n_1213, n_1214);
  xor g1180 (n_435, n_683, A[10]);
  nand g1183 (n_1218, A[5], A[10]);
  nand g1184 (n_454, n_684, n_705, n_1218);
  xor g1186 (n_437, n_1219, A[13]);
  nand g1190 (n_456, n_1220, n_792, n_1222);
  xor g1191 (n_1223, A[18], n_434);
  xor g1192 (n_440, n_1223, n_435);
  nand g1193 (n_1224, A[18], n_434);
  nand g1194 (n_1225, n_435, n_434);
  nand g1195 (n_1226, A[18], n_435);
  nand g1196 (n_459, n_1224, n_1225, n_1226);
  xor g1197 (n_1227, A[21], A[22]);
  xor g1198 (n_441, n_1227, n_436);
  nand g1200 (n_1229, n_436, A[22]);
  nand g1201 (n_1230, A[21], n_436);
  nand g1202 (n_460, n_1066, n_1229, n_1230);
  xor g1203 (n_1231, A[17], n_437);
  xor g1204 (n_444, n_1231, n_438);
  nand g1205 (n_1232, A[17], n_437);
  nand g1206 (n_1233, n_438, n_437);
  nand g1207 (n_1234, A[17], n_438);
  nand g1208 (n_463, n_1232, n_1233, n_1234);
  xor g1209 (n_1235, n_439, n_440);
  xor g1210 (n_446, n_1235, n_441);
  nand g1211 (n_1236, n_439, n_440);
  nand g1212 (n_1237, n_441, n_440);
  nand g1213 (n_1238, n_439, n_441);
  nand g1214 (n_465, n_1236, n_1237, n_1238);
  xor g1215 (n_1239, n_442, n_443);
  xor g1216 (n_447, n_1239, n_444);
  nand g1217 (n_1240, n_442, n_443);
  nand g1218 (n_1241, n_444, n_443);
  nand g1219 (n_1242, n_442, n_444);
  nand g1220 (n_466, n_1240, n_1241, n_1242);
  xor g1221 (n_1243, n_445, n_446);
  xor g1222 (n_449, n_1243, n_447);
  nand g1223 (n_1244, n_445, n_446);
  nand g1224 (n_1245, n_447, n_446);
  nand g1225 (n_1246, n_445, n_447);
  nand g1226 (n_469, n_1244, n_1245, n_1246);
  xor g1227 (n_1247, n_448, n_449);
  xor g1228 (n_93, n_1247, n_450);
  nand g1229 (n_1248, n_448, n_449);
  nand g1230 (n_1249, n_450, n_449);
  nand g1231 (n_1250, n_448, n_450);
  nand g1232 (n_44, n_1248, n_1249, n_1250);
  xor g1235 (n_1251, A[7], A[10]);
  nand g1240 (n_471, n_722, n_1253, n_1254);
  nand g1243 (n_1256, A[6], A[14]);
  nand g1245 (n_1258, A[6], A[11]);
  nand g1246 (n_473, n_1256, n_744, n_1258);
  xor g1247 (n_1259, A[18], A[19]);
  xor g1248 (n_458, n_1259, A[15]);
  nand g1249 (n_1260, A[18], A[19]);
  nand g1251 (n_1262, A[18], A[15]);
  nand g1252 (n_475, n_1260, n_948, n_1262);
  xor g1253 (n_1263, n_454, A[22]);
  xor g1254 (n_462, n_1263, n_455);
  nand g1255 (n_1264, n_454, A[22]);
  nand g1256 (n_1265, n_455, A[22]);
  nand g1257 (n_1266, n_454, n_455);
  nand g1258 (n_477, n_1264, n_1265, n_1266);
  xor g1259 (n_1267, A[23], n_456);
  xor g1260 (n_461, n_1267, n_457);
  nand g1261 (n_1268, A[23], n_456);
  nand g1262 (n_1269, n_457, n_456);
  nand g1263 (n_1270, A[23], n_457);
  nand g1264 (n_479, n_1268, n_1269, n_1270);
  xor g1265 (n_1271, n_458, n_459);
  xor g1266 (n_464, n_1271, n_460);
  nand g1267 (n_1272, n_458, n_459);
  nand g1268 (n_1273, n_460, n_459);
  nand g1269 (n_1274, n_458, n_460);
  nand g1270 (n_481, n_1272, n_1273, n_1274);
  xor g1271 (n_1275, n_461, n_462);
  xor g1272 (n_467, n_1275, n_463);
  nand g1273 (n_1276, n_461, n_462);
  nand g1274 (n_1277, n_463, n_462);
  nand g1275 (n_1278, n_461, n_463);
  nand g1276 (n_483, n_1276, n_1277, n_1278);
  xor g1277 (n_1279, n_464, n_465);
  xor g1278 (n_468, n_1279, n_466);
  nand g1279 (n_1280, n_464, n_465);
  nand g1280 (n_1281, n_466, n_465);
  nand g1281 (n_1282, n_464, n_466);
  nand g1282 (n_486, n_1280, n_1281, n_1282);
  xor g1283 (n_1283, n_467, n_468);
  xor g1284 (n_92, n_1283, n_469);
  nand g1285 (n_1284, n_467, n_468);
  nand g1286 (n_1285, n_469, n_468);
  nand g1287 (n_1286, n_467, n_469);
  nand g1288 (n_43, n_1284, n_1285, n_1286);
  xor g1289 (n_1287, A[7], A[8]);
  xor g1290 (n_472, n_1287, A[6]);
  nand g1292 (n_1289, A[6], A[8]);
  nand g1294 (n_487, n_1138, n_1289, n_1092);
  xor g1295 (n_1291, A[11], A[12]);
  xor g1296 (n_474, n_1291, A[19]);
  nand g1298 (n_1293, A[19], A[12]);
  nand g1299 (n_1294, A[11], A[19]);
  nand g1300 (n_489, n_973, n_1293, n_1294);
  xor g1302 (n_476, n_1295, A[15]);
  nand g1304 (n_1297, A[15], n_471);
  nand g1306 (n_490, n_1296, n_1297, n_1148);
  xor g1307 (n_1299, A[23], n_472);
  xor g1308 (n_478, n_1299, A[20]);
  nand g1309 (n_1300, A[23], n_472);
  nand g1310 (n_1301, A[20], n_472);
  nand g1312 (n_491, n_1300, n_1301, n_1021);
  xor g1313 (n_1303, n_473, A[16]);
  xor g1314 (n_480, n_1303, n_474);
  nand g1315 (n_1304, n_473, A[16]);
  nand g1316 (n_1305, n_474, A[16]);
  nand g1317 (n_1306, n_473, n_474);
  nand g1318 (n_494, n_1304, n_1305, n_1306);
  xor g1319 (n_1307, n_475, n_476);
  xor g1320 (n_482, n_1307, n_477);
  nand g1321 (n_1308, n_475, n_476);
  nand g1322 (n_1309, n_477, n_476);
  nand g1323 (n_1310, n_475, n_477);
  nand g1324 (n_496, n_1308, n_1309, n_1310);
  xor g1325 (n_1311, n_478, n_479);
  xor g1326 (n_484, n_1311, n_480);
  nand g1327 (n_1312, n_478, n_479);
  nand g1328 (n_1313, n_480, n_479);
  nand g1329 (n_1314, n_478, n_480);
  nand g1330 (n_498, n_1312, n_1313, n_1314);
  xor g1331 (n_1315, n_481, n_482);
  xor g1332 (n_485, n_1315, n_483);
  nand g1333 (n_1316, n_481, n_482);
  nand g1334 (n_1317, n_483, n_482);
  nand g1335 (n_1318, n_481, n_483);
  nand g1336 (n_501, n_1316, n_1317, n_1318);
  xor g1337 (n_1319, n_484, n_485);
  xor g1338 (n_91, n_1319, n_486);
  nand g1339 (n_1320, n_484, n_485);
  nand g1340 (n_1321, n_486, n_485);
  nand g1341 (n_1322, n_484, n_486);
  nand g1342 (n_42, n_1320, n_1321, n_1322);
  xor g1349 (n_1327, A[12], n_487);
  nand g1351 (n_1328, A[12], n_487);
  nand g1354 (n_506, n_1328, n_1329, n_1330);
  xor g1355 (n_1331, A[21], n_416);
  xor g1356 (n_493, n_1331, A[20]);
  nand g1358 (n_1333, A[20], n_416);
  nand g1360 (n_507, n_1189, n_1333, n_1020);
  xor g1361 (n_1335, A[17], A[16]);
  xor g1362 (n_495, n_1335, n_489);
  nand g1364 (n_1337, n_489, A[16]);
  nand g1365 (n_1338, A[17], n_489);
  nand g1366 (n_510, n_1026, n_1337, n_1338);
  xor g1367 (n_1339, n_490, n_491);
  xor g1368 (n_497, n_1339, n_492);
  nand g1369 (n_1340, n_490, n_491);
  nand g1370 (n_1341, n_492, n_491);
  nand g1371 (n_1342, n_490, n_492);
  nand g1372 (n_512, n_1340, n_1341, n_1342);
  xor g1373 (n_1343, n_493, n_494);
  xor g1374 (n_499, n_1343, n_495);
  nand g1375 (n_1344, n_493, n_494);
  nand g1376 (n_1345, n_495, n_494);
  nand g1377 (n_1346, n_493, n_495);
  nand g1378 (n_513, n_1344, n_1345, n_1346);
  xor g1379 (n_1347, n_496, n_497);
  xor g1380 (n_500, n_1347, n_498);
  nand g1381 (n_1348, n_496, n_497);
  nand g1382 (n_1349, n_498, n_497);
  nand g1383 (n_1350, n_496, n_498);
  nand g1384 (n_516, n_1348, n_1349, n_1350);
  xor g1385 (n_1351, n_499, n_500);
  xor g1386 (n_90, n_1351, n_501);
  nand g1387 (n_1352, n_499, n_500);
  nand g1388 (n_1353, n_501, n_500);
  nand g1389 (n_1354, n_499, n_501);
  nand g1390 (n_41, n_1352, n_1353, n_1354);
  xor g1393 (n_1355, A[9], A[14]);
  xor g1394 (n_505, n_1355, A[13]);
  nand g1395 (n_1356, A[9], A[14]);
  nand g1398 (n_520, n_1356, n_792, n_1182);
  xor g1400 (n_508, n_1359, A[21]);
  nand g1403 (n_1362, A[18], A[21]);
  nand g1404 (n_523, n_1360, n_1361, n_1362);
  xor g1405 (n_1363, n_436, A[22]);
  xor g1406 (n_509, n_1363, A[17]);
  nand g1408 (n_1365, A[17], A[22]);
  nand g1409 (n_1366, n_436, A[17]);
  nand g1410 (n_525, n_1229, n_1365, n_1366);
  xor g1411 (n_1367, n_505, n_506);
  xor g1412 (n_511, n_1367, n_507);
  nand g1413 (n_1368, n_505, n_506);
  nand g1414 (n_1369, n_507, n_506);
  nand g1415 (n_1370, n_505, n_507);
  nand g1416 (n_527, n_1368, n_1369, n_1370);
  xor g1417 (n_1371, n_508, n_509);
  xor g1418 (n_514, n_1371, n_510);
  nand g1419 (n_1372, n_508, n_509);
  nand g1420 (n_1373, n_510, n_509);
  nand g1421 (n_1374, n_508, n_510);
  nand g1422 (n_529, n_1372, n_1373, n_1374);
  xor g1423 (n_1375, n_511, n_512);
  xor g1424 (n_515, n_1375, n_513);
  nand g1425 (n_1376, n_511, n_512);
  nand g1426 (n_1377, n_513, n_512);
  nand g1427 (n_1378, n_511, n_513);
  nand g1428 (n_531, n_1376, n_1377, n_1378);
  xor g1429 (n_1379, n_514, n_515);
  xor g1430 (n_89, n_1379, n_516);
  nand g1431 (n_1380, n_514, n_515);
  nand g1432 (n_1381, n_516, n_515);
  nand g1433 (n_1382, n_514, n_516);
  nand g1434 (n_40, n_1380, n_1381, n_1382);
  xor g1438 (n_521, n_743, A[10]);
  nand g1440 (n_1385, A[10], A[11]);
  nand g1442 (n_533, n_744, n_1385, n_1098);
  xor g1444 (n_522, n_1359, A[19]);
  nand g1448 (n_535, n_1360, n_1260, n_1390);
  xor g1449 (n_1391, A[15], n_520);
  xor g1450 (n_524, n_1391, A[23]);
  nand g1451 (n_1392, A[15], n_520);
  nand g1452 (n_1393, A[23], n_520);
  nand g1454 (n_536, n_1392, n_1393, n_1149);
  xor g1455 (n_1395, A[22], n_521);
  xor g1456 (n_526, n_1395, n_522);
  nand g1457 (n_1396, A[22], n_521);
  nand g1458 (n_1397, n_522, n_521);
  nand g1459 (n_1398, A[22], n_522);
  nand g1460 (n_540, n_1396, n_1397, n_1398);
  xor g1461 (n_1399, n_523, n_524);
  xor g1462 (n_528, n_1399, n_525);
  nand g1463 (n_1400, n_523, n_524);
  nand g1464 (n_1401, n_525, n_524);
  nand g1465 (n_1402, n_523, n_525);
  nand g1466 (n_541, n_1400, n_1401, n_1402);
  xor g1467 (n_1403, n_526, n_527);
  xor g1468 (n_530, n_1403, n_528);
  nand g1469 (n_1404, n_526, n_527);
  nand g1470 (n_1405, n_528, n_527);
  nand g1471 (n_1406, n_526, n_528);
  nand g1472 (n_544, n_1404, n_1405, n_1406);
  xor g1473 (n_1407, n_529, n_530);
  xor g1474 (n_88, n_1407, n_531);
  nand g1475 (n_1408, n_529, n_530);
  nand g1476 (n_1409, n_531, n_530);
  nand g1477 (n_1410, n_529, n_531);
  nand g1478 (n_39, n_1408, n_1409, n_1410);
  xor g1480 (n_534, n_1291, A[10]);
  nand g1483 (n_1414, A[12], A[10]);
  nand g1484 (n_545, n_973, n_1385, n_1414);
  xor g1486 (n_537, n_1415, A[15]);
  nand g1490 (n_546, n_1416, n_1148, n_948);
  xor g1491 (n_1419, A[23], A[20]);
  xor g1492 (n_538, n_1419, A[16]);
  nand g1494 (n_1421, A[16], A[20]);
  nand g1495 (n_1422, A[23], A[16]);
  nand g1496 (n_549, n_1021, n_1421, n_1422);
  xor g1497 (n_1423, n_533, n_534);
  xor g1498 (n_539, n_1423, n_535);
  nand g1499 (n_1424, n_533, n_534);
  nand g1500 (n_1425, n_535, n_534);
  nand g1501 (n_1426, n_533, n_535);
  nand g1502 (n_550, n_1424, n_1425, n_1426);
  xor g1503 (n_1427, n_536, n_537);
  xor g1504 (n_542, n_1427, n_538);
  nand g1505 (n_1428, n_536, n_537);
  nand g1506 (n_1429, n_538, n_537);
  nand g1507 (n_1430, n_536, n_538);
  nand g1508 (n_552, n_1428, n_1429, n_1430);
  xor g1509 (n_1431, n_539, n_540);
  xor g1510 (n_543, n_1431, n_541);
  nand g1511 (n_1432, n_539, n_540);
  nand g1512 (n_1433, n_541, n_540);
  nand g1513 (n_1434, n_539, n_541);
  nand g1514 (n_555, n_1432, n_1433, n_1434);
  xor g1515 (n_1435, n_542, n_543);
  xor g1516 (n_87, n_1435, n_544);
  nand g1517 (n_1436, n_542, n_543);
  nand g1518 (n_1437, n_544, n_543);
  nand g1519 (n_1438, n_542, n_544);
  nand g1520 (n_38, n_1436, n_1437, n_1438);
  xor g1521 (n_1439, A[13], A[12]);
  nand g1526 (n_558, n_765, n_1330, n_1442);
  xor g1528 (n_548, n_1019, A[17]);
  nand g1531 (n_1446, A[21], A[17]);
  nand g1532 (n_561, n_1020, n_918, n_1446);
  xor g1533 (n_1447, n_545, A[16]);
  xor g1534 (n_551, n_1447, n_546);
  nand g1535 (n_1448, n_545, A[16]);
  nand g1536 (n_1449, n_546, A[16]);
  nand g1537 (n_1450, n_545, n_546);
  nand g1538 (n_562, n_1448, n_1449, n_1450);
  xor g1539 (n_1451, n_547, n_548);
  xor g1540 (n_553, n_1451, n_549);
  nand g1541 (n_1452, n_547, n_548);
  nand g1542 (n_1453, n_549, n_548);
  nand g1543 (n_1454, n_547, n_549);
  nand g1544 (n_563, n_1452, n_1453, n_1454);
  xor g1545 (n_1455, n_550, n_551);
  xor g1546 (n_554, n_1455, n_552);
  nand g1547 (n_1456, n_550, n_551);
  nand g1548 (n_1457, n_552, n_551);
  nand g1549 (n_1458, n_550, n_552);
  nand g1550 (n_566, n_1456, n_1457, n_1458);
  xor g1551 (n_1459, n_553, n_554);
  xor g1552 (n_86, n_1459, n_555);
  nand g1553 (n_1460, n_553, n_554);
  nand g1554 (n_1461, n_555, n_554);
  nand g1555 (n_1462, n_553, n_555);
  nand g1556 (n_37, n_1460, n_1461, n_1462);
  xor g1559 (n_1463, A[13], A[18]);
  nand g1564 (n_570, n_1057, n_1465, n_1466);
  xor g1566 (n_560, n_1227, A[17]);
  nand g1570 (n_573, n_1066, n_1365, n_1446);
  xor g1571 (n_1471, n_558, n_559);
  xor g1572 (n_564, n_1471, n_560);
  nand g1573 (n_1472, n_558, n_559);
  nand g1574 (n_1473, n_560, n_559);
  nand g1575 (n_1474, n_558, n_560);
  nand g1576 (n_575, n_1472, n_1473, n_1474);
  xor g1577 (n_1475, n_561, n_562);
  xor g1578 (n_565, n_1475, n_563);
  nand g1579 (n_1476, n_561, n_562);
  nand g1580 (n_1477, n_563, n_562);
  nand g1581 (n_1478, n_561, n_563);
  nand g1582 (n_577, n_1476, n_1477, n_1478);
  xor g1583 (n_1479, n_564, n_565);
  xor g1584 (n_85, n_1479, n_566);
  nand g1585 (n_1480, n_564, n_565);
  nand g1586 (n_1481, n_566, n_565);
  nand g1587 (n_1482, n_564, n_566);
  nand g1588 (n_36, n_1480, n_1481, n_1482);
  xor g1592 (n_572, n_1259, A[14]);
  nand g1594 (n_1485, A[14], A[19]);
  nand g1596 (n_579, n_1260, n_1485, n_1058);
  xor g1598 (n_571, n_1487, A[22]);
  nand g1601 (n_1490, A[15], A[22]);
  nand g1602 (n_581, n_1488, n_1489, n_1490);
  xor g1603 (n_1491, A[23], n_570);
  xor g1604 (n_574, n_1491, n_571);
  nand g1605 (n_1492, A[23], n_570);
  nand g1606 (n_1493, n_571, n_570);
  nand g1607 (n_1494, A[23], n_571);
  nand g1608 (n_584, n_1492, n_1493, n_1494);
  xor g1609 (n_1495, n_572, n_573);
  xor g1610 (n_576, n_1495, n_574);
  nand g1611 (n_1496, n_572, n_573);
  nand g1612 (n_1497, n_574, n_573);
  nand g1613 (n_1498, n_572, n_574);
  nand g1614 (n_586, n_1496, n_1497, n_1498);
  xor g1615 (n_1499, n_575, n_576);
  xor g1616 (n_84, n_1499, n_577);
  nand g1617 (n_1500, n_575, n_576);
  nand g1618 (n_1501, n_577, n_576);
  nand g1619 (n_1502, n_575, n_577);
  nand g1620 (n_35, n_1500, n_1501, n_1502);
  xor g1627 (n_1507, A[14], A[23]);
  xor g1628 (n_582, n_1507, A[20]);
  nand g1629 (n_1508, A[14], A[23]);
  nand g1631 (n_1510, A[14], A[20]);
  nand g1632 (n_588, n_1508, n_1021, n_1510);
  xor g1633 (n_1511, A[16], n_579);
  xor g1634 (n_583, n_1511, n_537);
  nand g1635 (n_1512, A[16], n_579);
  nand g1636 (n_1513, n_537, n_579);
  nand g1637 (n_1514, A[16], n_537);
  nand g1638 (n_591, n_1512, n_1513, n_1514);
  xor g1639 (n_1515, n_581, n_582);
  xor g1640 (n_585, n_1515, n_583);
  nand g1641 (n_1516, n_581, n_582);
  nand g1642 (n_1517, n_583, n_582);
  nand g1643 (n_1518, n_581, n_583);
  nand g1644 (n_593, n_1516, n_1517, n_1518);
  xor g1645 (n_1519, n_584, n_585);
  xor g1646 (n_83, n_1519, n_586);
  nand g1647 (n_1520, n_584, n_585);
  nand g1648 (n_1521, n_586, n_585);
  nand g1649 (n_1522, n_584, n_586);
  nand g1650 (n_34, n_1520, n_1521, n_1522);
  xor g1652 (n_589, n_1187, A[20]);
  nand g1656 (n_596, n_1188, n_1020, n_1526);
  xor g1658 (n_590, n_1335, n_546);
  nand g1661 (n_1530, A[17], n_546);
  nand g1662 (n_598, n_1026, n_1449, n_1530);
  xor g1663 (n_1531, n_588, n_589);
  xor g1664 (n_592, n_1531, n_590);
  nand g1665 (n_1532, n_588, n_589);
  nand g1666 (n_1533, n_590, n_589);
  nand g1667 (n_1534, n_588, n_590);
  nand g1668 (n_600, n_1532, n_1533, n_1534);
  xor g1669 (n_1535, n_591, n_592);
  xor g1670 (n_82, n_1535, n_593);
  nand g1671 (n_1536, n_591, n_592);
  nand g1672 (n_1537, n_593, n_592);
  nand g1673 (n_1538, n_591, n_593);
  nand g1674 (n_81, n_1536, n_1537, n_1538);
  xor g1678 (n_597, n_1539, A[22]);
  nand g1682 (n_604, n_1540, n_1541, n_1066);
  xor g1683 (n_1543, A[17], n_596);
  xor g1684 (n_599, n_1543, n_597);
  nand g1685 (n_1544, A[17], n_596);
  nand g1686 (n_1545, n_597, n_596);
  nand g1687 (n_1546, A[17], n_597);
  nand g1688 (n_607, n_1544, n_1545, n_1546);
  xor g1689 (n_1547, n_598, n_599);
  xor g1690 (n_33, n_1547, n_600);
  nand g1691 (n_1548, n_598, n_599);
  nand g1692 (n_1549, n_600, n_599);
  nand g1693 (n_1550, n_598, n_600);
  nand g1694 (n_80, n_1548, n_1549, n_1550);
  xor g1697 (n_1551, A[19], A[22]);
  nand g1699 (n_1552, A[19], A[22]);
  nand g1702 (n_609, n_1552, n_1541, n_1554);
  xor g1703 (n_1555, A[18], A[23]);
  xor g1704 (n_606, n_1555, n_604);
  nand g1705 (n_1556, A[18], A[23]);
  nand g1706 (n_1557, n_604, A[23]);
  nand g1707 (n_1558, A[18], n_604);
  nand g1708 (n_612, n_1556, n_1557, n_1558);
  xor g1709 (n_1559, n_605, n_606);
  xor g1710 (n_32, n_1559, n_607);
  nand g1711 (n_1560, n_605, n_606);
  nand g1712 (n_1561, n_607, n_606);
  nand g1713 (n_1562, n_605, n_607);
  nand g1714 (n_31, n_1560, n_1561, n_1562);
  xor g1716 (n_610, n_1415, A[23]);
  nand g1718 (n_1565, A[23], A[19]);
  nand g1720 (n_613, n_1416, n_1565, n_1150);
  xor g1721 (n_1567, A[18], A[20]);
  xor g1722 (n_611, n_1567, n_609);
  nand g1723 (n_1568, A[18], A[20]);
  nand g1724 (n_1569, n_609, A[20]);
  nand g1725 (n_1570, A[18], n_609);
  nand g1726 (n_615, n_1568, n_1569, n_1570);
  xor g1727 (n_1571, n_610, n_611);
  xor g1728 (n_79, n_1571, n_612);
  nand g1729 (n_1572, n_610, n_611);
  nand g1730 (n_1573, n_612, n_611);
  nand g1731 (n_1574, n_610, n_612);
  nand g1732 (n_30, n_1572, n_1573, n_1574);
  xor g1739 (n_1579, n_613, n_589);
  xor g1740 (n_78, n_1579, n_615);
  nand g1741 (n_1580, n_613, n_589);
  nand g1742 (n_1581, n_615, n_589);
  nand g1743 (n_1582, n_613, n_615);
  nand g1744 (n_77, n_1580, n_1581, n_1582);
  nand g1751 (n_1586, A[22], n_596);
  nand g1752 (n_28, n_1584, n_1585, n_1586);
  xor g1756 (n_76, n_1587, A[21]);
  nand g1760 (n_27, n_1588, n_1589, n_1022);
  xor g1762 (n_75, n_1591, A[22]);
  nand g1764 (n_1593, A[22], A[23]);
  nand g1766 (n_74, n_1150, n_1593, n_1594);
  nor g11 (n_1610, A[0], A[2]);
  nand g12 (n_1605, A[0], A[2]);
  nor g13 (n_1606, A[3], n_118);
  nand g14 (n_1607, A[3], n_118);
  nor g15 (n_1616, A[4], n_117);
  nand g16 (n_1611, A[4], n_117);
  nor g17 (n_1612, n_68, n_116);
  nand g18 (n_1613, n_68, n_116);
  nor g19 (n_1622, n_67, n_115);
  nand g20 (n_1617, n_67, n_115);
  nor g21 (n_1618, n_66, n_114);
  nand g22 (n_1619, n_66, n_114);
  nor g23 (n_1628, n_65, n_113);
  nand g24 (n_1623, n_65, n_113);
  nor g25 (n_1624, n_64, n_112);
  nand g26 (n_1625, n_64, n_112);
  nor g27 (n_1634, n_63, n_111);
  nand g28 (n_1629, n_63, n_111);
  nor g29 (n_1630, n_62, n_110);
  nand g30 (n_1631, n_62, n_110);
  nor g31 (n_1640, n_61, n_109);
  nand g32 (n_1635, n_61, n_109);
  nor g33 (n_1636, n_60, n_108);
  nand g34 (n_1637, n_60, n_108);
  nor g35 (n_1646, n_59, n_107);
  nand g36 (n_1641, n_59, n_107);
  nor g37 (n_1642, n_58, n_106);
  nand g38 (n_1643, n_58, n_106);
  nor g39 (n_1652, n_57, n_105);
  nand g40 (n_1647, n_57, n_105);
  nor g41 (n_1648, n_56, n_104);
  nand g42 (n_1649, n_56, n_104);
  nor g43 (n_1658, n_55, n_103);
  nand g44 (n_1653, n_55, n_103);
  nor g45 (n_1654, n_54, n_102);
  nand g46 (n_1655, n_54, n_102);
  nor g47 (n_1664, n_53, n_101);
  nand g48 (n_1659, n_53, n_101);
  nor g49 (n_1660, n_52, n_100);
  nand g50 (n_1661, n_52, n_100);
  nor g51 (n_1670, n_51, n_99);
  nand g52 (n_1665, n_51, n_99);
  nor g53 (n_1666, n_50, n_98);
  nand g54 (n_1667, n_50, n_98);
  nor g55 (n_1676, n_49, n_97);
  nand g56 (n_1671, n_49, n_97);
  nor g57 (n_1672, n_48, n_96);
  nand g58 (n_1673, n_48, n_96);
  nor g59 (n_1682, n_47, n_95);
  nand g60 (n_1677, n_47, n_95);
  nor g61 (n_1678, n_46, n_94);
  nand g62 (n_1679, n_46, n_94);
  nor g63 (n_1688, n_45, n_93);
  nand g64 (n_1683, n_45, n_93);
  nor g65 (n_1684, n_44, n_92);
  nand g66 (n_1685, n_44, n_92);
  nor g67 (n_1694, n_43, n_91);
  nand g68 (n_1689, n_43, n_91);
  nor g69 (n_1690, n_42, n_90);
  nand g70 (n_1691, n_42, n_90);
  nor g71 (n_1700, n_41, n_89);
  nand g72 (n_1695, n_41, n_89);
  nor g73 (n_1696, n_40, n_88);
  nand g74 (n_1697, n_40, n_88);
  nor g75 (n_1706, n_39, n_87);
  nand g76 (n_1701, n_39, n_87);
  nor g77 (n_1702, n_38, n_86);
  nand g78 (n_1703, n_38, n_86);
  nor g79 (n_1712, n_37, n_85);
  nand g80 (n_1707, n_37, n_85);
  nor g81 (n_1708, n_36, n_84);
  nand g82 (n_1709, n_36, n_84);
  nor g83 (n_1718, n_35, n_83);
  nand g84 (n_1713, n_35, n_83);
  nor g85 (n_1714, n_34, n_82);
  nand g86 (n_1715, n_34, n_82);
  nor g87 (n_1724, n_33, n_81);
  nand g88 (n_1719, n_33, n_81);
  nor g89 (n_1720, n_32, n_80);
  nand g90 (n_1721, n_32, n_80);
  nor g91 (n_1730, n_31, n_79);
  nand g92 (n_1725, n_31, n_79);
  nor g93 (n_1726, n_30, n_78);
  nand g94 (n_1727, n_30, n_78);
  nor g95 (n_1736, n_29, n_77);
  nand g96 (n_1731, n_29, n_77);
  nor g97 (n_1732, n_28, n_76);
  nand g98 (n_1733, n_28, n_76);
  nor g99 (n_1740, n_27, n_75);
  nand g100 (n_1737, n_27, n_75);
  nor g106 (n_1608, n_1605, n_1606);
  nor g110 (n_1614, n_1611, n_1612);
  nor g113 (n_1750, n_1616, n_1612);
  nor g114 (n_1620, n_1617, n_1618);
  nor g117 (n_1752, n_1622, n_1618);
  nor g118 (n_1626, n_1623, n_1624);
  nor g121 (n_1760, n_1628, n_1624);
  nor g122 (n_1632, n_1629, n_1630);
  nor g125 (n_1762, n_1634, n_1630);
  nor g126 (n_1638, n_1635, n_1636);
  nor g129 (n_1770, n_1640, n_1636);
  nor g130 (n_1644, n_1641, n_1642);
  nor g133 (n_1772, n_1646, n_1642);
  nor g134 (n_1650, n_1647, n_1648);
  nor g137 (n_1780, n_1652, n_1648);
  nor g138 (n_1656, n_1653, n_1654);
  nor g141 (n_1782, n_1658, n_1654);
  nor g142 (n_1662, n_1659, n_1660);
  nor g145 (n_1790, n_1664, n_1660);
  nor g146 (n_1668, n_1665, n_1666);
  nor g149 (n_1792, n_1670, n_1666);
  nor g150 (n_1674, n_1671, n_1672);
  nor g153 (n_1800, n_1676, n_1672);
  nor g154 (n_1680, n_1677, n_1678);
  nor g157 (n_1802, n_1682, n_1678);
  nor g158 (n_1686, n_1683, n_1684);
  nor g161 (n_1810, n_1688, n_1684);
  nor g162 (n_1692, n_1689, n_1690);
  nor g165 (n_1812, n_1694, n_1690);
  nor g166 (n_1698, n_1695, n_1696);
  nor g169 (n_1820, n_1700, n_1696);
  nor g170 (n_1704, n_1701, n_1702);
  nor g173 (n_1822, n_1706, n_1702);
  nor g174 (n_1710, n_1707, n_1708);
  nor g177 (n_1830, n_1712, n_1708);
  nor g178 (n_1716, n_1713, n_1714);
  nor g181 (n_1832, n_1718, n_1714);
  nor g182 (n_1722, n_1719, n_1720);
  nor g185 (n_1840, n_1724, n_1720);
  nor g186 (n_1728, n_1725, n_1726);
  nor g189 (n_1842, n_1730, n_1726);
  nor g190 (n_1734, n_1731, n_1732);
  nor g193 (n_1850, n_1736, n_1732);
  nor g203 (n_1748, n_1622, n_1747);
  nand g212 (n_1860, n_1750, n_1752);
  nor g213 (n_1758, n_1634, n_1757);
  nand g222 (n_1867, n_1760, n_1762);
  nor g223 (n_1768, n_1646, n_1767);
  nand g232 (n_1875, n_1770, n_1772);
  nor g233 (n_1778, n_1658, n_1777);
  nand g242 (n_1882, n_1780, n_1782);
  nor g243 (n_1788, n_1670, n_1787);
  nand g252 (n_1890, n_1790, n_1792);
  nor g253 (n_1798, n_1682, n_1797);
  nand g262 (n_1897, n_1800, n_1802);
  nor g263 (n_1808, n_1694, n_1807);
  nand g1776 (n_1905, n_1810, n_1812);
  nor g1777 (n_1818, n_1706, n_1817);
  nand g1786 (n_1912, n_1820, n_1822);
  nor g1787 (n_1828, n_1718, n_1827);
  nand g1796 (n_1920, n_1830, n_1832);
  nor g1797 (n_1838, n_1730, n_1837);
  nand g1806 (n_1927, n_1840, n_1842);
  nor g1807 (n_1848, n_1740, n_1847);
  nand g1814 (n_2131, n_1611, n_1854);
  nand g1816 (n_2133, n_1747, n_1855);
  nand g1819 (n_2136, n_1858, n_1859);
  nand g1822 (n_1935, n_1862, n_1863);
  nor g1823 (n_1865, n_1640, n_1864);
  nor g1826 (n_1945, n_1640, n_1867);
  nor g1832 (n_1873, n_1871, n_1864);
  nor g1835 (n_1951, n_1867, n_1871);
  nor g1836 (n_1877, n_1875, n_1864);
  nor g1839 (n_1954, n_1867, n_1875);
  nor g1840 (n_1880, n_1664, n_1879);
  nor g1843 (n_2034, n_1664, n_1882);
  nor g1849 (n_1888, n_1886, n_1879);
  nor g1852 (n_2040, n_1882, n_1886);
  nor g1853 (n_1892, n_1890, n_1879);
  nor g1856 (n_1960, n_1882, n_1890);
  nor g1857 (n_1895, n_1688, n_1894);
  nor g1860 (n_1973, n_1688, n_1897);
  nor g1866 (n_1903, n_1901, n_1894);
  nor g1869 (n_1983, n_1897, n_1901);
  nor g1870 (n_1907, n_1905, n_1894);
  nor g1873 (n_1988, n_1897, n_1905);
  nor g1874 (n_1910, n_1712, n_1909);
  nor g1877 (n_2086, n_1712, n_1912);
  nor g1883 (n_1918, n_1916, n_1909);
  nor g1886 (n_2092, n_1912, n_1916);
  nor g1887 (n_1922, n_1920, n_1909);
  nor g1890 (n_1996, n_1912, n_1920);
  nor g1891 (n_1925, n_1736, n_1924);
  nor g1894 (n_2009, n_1736, n_1927);
  nor g1900 (n_1933, n_1931, n_1924);
  nor g1903 (n_2019, n_1927, n_1931);
  nand g1906 (n_2140, n_1623, n_1937);
  nand g1907 (n_1938, n_1760, n_1935);
  nand g1908 (n_2142, n_1757, n_1938);
  nand g1911 (n_2145, n_1941, n_1942);
  nand g1914 (n_2148, n_1864, n_1944);
  nand g1915 (n_1947, n_1945, n_1935);
  nand g1916 (n_2151, n_1946, n_1947);
  nand g1917 (n_1950, n_1948, n_1935);
  nand g1918 (n_2153, n_1949, n_1950);
  nand g1919 (n_1953, n_1951, n_1935);
  nand g1920 (n_2156, n_1952, n_1953);
  nand g1921 (n_1956, n_1954, n_1935);
  nand g1922 (n_2024, n_1955, n_1956);
  nor g1923 (n_1958, n_1676, n_1957);
  nand g1932 (n_2048, n_1800, n_1960);
  nor g1933 (n_1967, n_1965, n_1957);
  nor g1938 (n_1970, n_1897, n_1957);
  nand g1947 (n_2060, n_1960, n_1973);
  nand g1952 (n_2064, n_1960, n_1978);
  nand g1957 (n_2068, n_1960, n_1983);
  nand g1962 (n_2072, n_1960, n_1988);
  nor g1963 (n_1994, n_1724, n_1993);
  nand g1972 (n_2100, n_1840, n_1996);
  nor g1973 (n_2003, n_2001, n_1993);
  nor g1978 (n_2006, n_1927, n_1993);
  nand g1987 (n_2112, n_1996, n_2009);
  nand g1992 (n_2116, n_1996, n_2014);
  nand g1997 (n_2120, n_1996, n_2019);
  nand g2000 (n_2160, n_1647, n_2026);
  nand g2001 (n_2027, n_1780, n_2024);
  nand g2002 (n_2162, n_1777, n_2027);
  nand g2005 (n_2165, n_2030, n_2031);
  nand g2008 (n_2168, n_1879, n_2033);
  nand g2009 (n_2036, n_2034, n_2024);
  nand g2010 (n_2171, n_2035, n_2036);
  nand g2011 (n_2039, n_2037, n_2024);
  nand g2012 (n_2173, n_2038, n_2039);
  nand g2013 (n_2042, n_2040, n_2024);
  nand g2014 (n_2176, n_2041, n_2042);
  nand g2015 (n_2043, n_1960, n_2024);
  nand g2016 (n_2178, n_1957, n_2043);
  nand g2019 (n_2181, n_2046, n_2047);
  nand g2022 (n_2183, n_2050, n_2051);
  nand g2025 (n_2186, n_2054, n_2055);
  nand g2028 (n_2189, n_2058, n_2059);
  nand g2031 (n_2192, n_2062, n_2063);
  nand g2034 (n_2194, n_2066, n_2067);
  nand g2037 (n_2197, n_2070, n_2071);
  nand g2040 (n_2076, n_2074, n_2075);
  nand g2043 (n_2201, n_1695, n_2078);
  nand g2044 (n_2079, n_1820, n_2076);
  nand g2045 (n_2203, n_1817, n_2079);
  nand g2048 (n_2206, n_2082, n_2083);
  nand g2051 (n_2209, n_1909, n_2085);
  nand g2052 (n_2088, n_2086, n_2076);
  nand g2053 (n_2212, n_2087, n_2088);
  nand g2054 (n_2091, n_2089, n_2076);
  nand g2055 (n_2214, n_2090, n_2091);
  nand g2056 (n_2094, n_2092, n_2076);
  nand g2057 (n_2217, n_2093, n_2094);
  nand g2058 (n_2095, n_1996, n_2076);
  nand g2059 (n_2219, n_1993, n_2095);
  nand g2062 (n_2222, n_2098, n_2099);
  nand g2065 (n_2224, n_2102, n_2103);
  nand g2068 (n_2227, n_2106, n_2107);
  nand g2071 (n_2230, n_2110, n_2111);
  nand g2074 (n_2233, n_2114, n_2115);
  nand g2077 (n_2235, n_2118, n_2119);
  nand g2080 (n_2238, n_2122, n_2123);
  xnor g2092 (Z[5], n_2131, n_2132);
  xnor g2094 (Z[6], n_2133, n_2134);
  xnor g2097 (Z[7], n_2136, n_2137);
  xnor g2099 (Z[8], n_1935, n_2138);
  xnor g2102 (Z[9], n_2140, n_2141);
  xnor g2104 (Z[10], n_2142, n_2143);
  xnor g2107 (Z[11], n_2145, n_2146);
  xnor g2110 (Z[12], n_2148, n_2149);
  xnor g2113 (Z[13], n_2151, n_2152);
  xnor g2115 (Z[14], n_2153, n_2154);
  xnor g2118 (Z[15], n_2156, n_2157);
  xnor g2120 (Z[16], n_2024, n_2158);
  xnor g2123 (Z[17], n_2160, n_2161);
  xnor g2125 (Z[18], n_2162, n_2163);
  xnor g2128 (Z[19], n_2165, n_2166);
  xnor g2131 (Z[20], n_2168, n_2169);
  xnor g2134 (Z[21], n_2171, n_2172);
  xnor g2136 (Z[22], n_2173, n_2174);
  xnor g2139 (Z[23], n_2176, n_2177);
  xnor g2141 (Z[24], n_2178, n_2179);
  xnor g2144 (Z[25], n_2181, n_2182);
  xnor g2146 (Z[26], n_2183, n_2184);
  xnor g2149 (Z[27], n_2186, n_2187);
  xnor g2152 (Z[28], n_2189, n_2190);
  xnor g2155 (Z[29], n_2192, n_2193);
  xnor g2157 (Z[30], n_2194, n_2195);
  xnor g2160 (Z[31], n_2197, n_2198);
  xnor g2162 (Z[32], n_2076, n_2199);
  xnor g2165 (Z[33], n_2201, n_2202);
  xnor g2167 (Z[34], n_2203, n_2204);
  xnor g2170 (Z[35], n_2206, n_2207);
  xnor g2173 (Z[36], n_2209, n_2210);
  xnor g2176 (Z[37], n_2212, n_2213);
  xnor g2178 (Z[38], n_2214, n_2215);
  xnor g2181 (Z[39], n_2217, n_2218);
  xnor g2183 (Z[40], n_2219, n_2220);
  xnor g2186 (Z[41], n_2222, n_2223);
  xnor g2188 (Z[42], n_2224, n_2225);
  xnor g2191 (Z[43], n_2227, n_2228);
  xnor g2194 (Z[44], n_2230, n_2231);
  xnor g2197 (Z[45], n_2233, n_2234);
  xnor g2199 (Z[46], n_2235, n_2236);
  xnor g2202 (Z[47], n_2238, n_2239);
  or g2212 (n_1045, A[2], wc);
  not gc (wc, n_171);
  or g2213 (n_1046, wc0, A[2]);
  not gc0 (wc0, A[1]);
  or g2214 (n_1090, A[2], wc1);
  not gc1 (wc1, A[3]);
  xnor g2215 (n_1147, A[24], A[15]);
  or g2216 (n_1148, wc2, A[24]);
  not gc2 (wc2, A[15]);
  or g2217 (n_1150, wc3, A[24]);
  not gc3 (wc3, A[23]);
  xnor g2218 (n_1187, A[24], A[21]);
  or g2219 (n_1188, wc4, A[24]);
  not gc4 (wc4, A[21]);
  xnor g2220 (n_1219, A[14], A[6]);
  or g2221 (n_1220, A[6], wc5);
  not gc5 (wc5, A[14]);
  or g2222 (n_1222, A[6], wc6);
  not gc6 (wc6, A[13]);
  xnor g2223 (n_455, n_1251, A[6]);
  or g2224 (n_1253, A[6], wc7);
  not gc7 (wc7, A[10]);
  or g2225 (n_1254, A[6], wc8);
  not gc8 (wc8, A[7]);
  or g2227 (n_1330, wc9, A[24]);
  not gc9 (wc9, A[12]);
  xnor g2228 (n_1359, A[18], A[10]);
  or g2229 (n_1360, A[10], wc10);
  not gc10 (wc10, A[18]);
  or g2230 (n_1361, A[10], wc11);
  not gc11 (wc11, A[21]);
  or g2231 (n_1390, A[10], wc12);
  not gc12 (wc12, A[19]);
  xnor g2232 (n_1415, A[24], A[19]);
  or g2233 (n_1416, wc13, A[24]);
  not gc13 (wc13, A[19]);
  xnor g2234 (n_547, n_1439, A[24]);
  or g2235 (n_1442, wc14, A[24]);
  not gc14 (wc14, A[13]);
  xnor g2236 (n_559, n_1463, A[14]);
  or g2237 (n_1465, A[14], wc15);
  not gc15 (wc15, A[18]);
  or g2238 (n_1466, wc16, A[14]);
  not gc16 (wc16, A[13]);
  xnor g2239 (n_1487, A[15], A[14]);
  or g2240 (n_1488, A[14], wc17);
  not gc17 (wc17, A[15]);
  or g2241 (n_1489, A[14], wc18);
  not gc18 (wc18, A[22]);
  or g2242 (n_1526, wc19, A[24]);
  not gc19 (wc19, A[20]);
  xnor g2243 (n_1539, A[21], A[18]);
  or g2244 (n_1540, A[18], wc20);
  not gc20 (wc20, A[21]);
  or g2245 (n_1541, A[18], wc21);
  not gc21 (wc21, A[22]);
  xnor g2246 (n_605, n_1551, A[18]);
  or g2247 (n_1554, A[18], wc22);
  not gc22 (wc22, A[19]);
  or g2249 (n_1584, A[21], wc23);
  not gc23 (wc23, A[22]);
  xnor g2250 (n_1587, A[23], A[22]);
  or g2251 (n_1588, A[22], wc24);
  not gc24 (wc24, A[23]);
  or g2252 (n_1589, wc25, A[22]);
  not gc25 (wc25, A[21]);
  xnor g2253 (n_1591, A[24], A[23]);
  or g2254 (n_1594, wc26, A[24]);
  not gc26 (wc26, A[22]);
  xnor g2255 (n_351, n_1043, A[2]);
  xnor g2256 (n_1059, n_232, A[24]);
  or g2257 (n_1060, A[24], wc27);
  not gc27 (wc27, n_232);
  xnor g2258 (n_373, n_627, A[2]);
  nand g2259 (n_393, n_628, n_1090);
  or g2260 (n_1190, A[24], wc28);
  not gc28 (wc28, n_416);
  xnor g2261 (n_457, n_1219, A[11]);
  or g2263 (n_2125, wc29, n_1610);
  not gc29 (wc29, n_1605);
  xnor g2264 (n_1295, n_471, A[24]);
  or g2265 (n_1296, A[24], wc30);
  not gc30 (wc30, n_471);
  or g2266 (n_1329, A[24], wc31);
  not gc31 (wc31, n_487);
  xnor g2267 (n_29, n_1227, n_596);
  or g2268 (n_1585, A[21], wc32);
  not gc32 (wc32, n_596);
  and g2269 (n_1745, wc33, n_1607);
  not gc33 (wc33, n_1608);
  or g2270 (n_2128, wc34, n_1606);
  not gc34 (wc34, n_1607);
  or g2271 (n_1061, A[24], wc35);
  not gc35 (wc35, n_353);
  xnor g2272 (n_492, n_1327, A[24]);
  and g2273 (n_1738, wc36, n_74);
  not gc36 (wc36, A[24]);
  or g2274 (n_1739, wc37, n_74);
  not gc37 (wc37, A[24]);
  not g2275 (Z[2], n_2125);
  or g2276 (n_2129, wc38, n_1616);
  not gc38 (wc38, n_1611);
  and g2277 (n_1747, wc39, n_1613);
  not gc39 (wc39, n_1614);
  or g2280 (n_1856, wc40, n_1622);
  not gc40 (wc40, n_1750);
  or g2281 (n_2132, wc41, n_1612);
  not gc41 (wc41, n_1613);
  or g2282 (n_2134, wc42, n_1622);
  not gc42 (wc42, n_1617);
  or g2283 (n_2236, wc43, n_1740);
  not gc43 (wc43, n_1737);
  and g2284 (n_1754, wc44, n_1619);
  not gc44 (wc44, n_1620);
  or g2285 (n_1854, n_1616, n_1745);
  or g2286 (n_1855, n_1745, wc45);
  not gc45 (wc45, n_1750);
  xor g2287 (Z[3], n_1605, n_2128);
  xor g2288 (Z[4], n_1745, n_2129);
  or g2289 (n_2137, wc46, n_1618);
  not gc46 (wc46, n_1619);
  or g2290 (n_2239, wc47, n_1738);
  not gc47 (wc47, n_1739);
  and g2291 (n_1858, wc48, n_1617);
  not gc48 (wc48, n_1748);
  and g2292 (n_1755, wc49, n_1752);
  not gc49 (wc49, n_1747);
  or g2293 (n_1859, n_1745, n_1856);
  or g2294 (n_2138, wc50, n_1628);
  not gc50 (wc50, n_1623);
  or g2295 (n_2234, wc51, n_1732);
  not gc51 (wc51, n_1733);
  and g2296 (n_1757, wc52, n_1625);
  not gc52 (wc52, n_1626);
  and g2297 (n_1862, wc53, n_1754);
  not gc53 (wc53, n_1755);
  or g2298 (n_1863, n_1860, n_1745);
  or g2299 (n_2141, wc54, n_1624);
  not gc54 (wc54, n_1625);
  and g2300 (n_1764, wc55, n_1631);
  not gc55 (wc55, n_1632);
  and g2301 (n_1844, wc56, n_1727);
  not gc56 (wc56, n_1728);
  and g2302 (n_1847, wc57, n_1733);
  not gc57 (wc57, n_1734);
  or g2303 (n_1939, wc58, n_1634);
  not gc58 (wc58, n_1760);
  or g2304 (n_1931, wc59, n_1740);
  not gc59 (wc59, n_1850);
  or g2305 (n_2143, wc60, n_1634);
  not gc60 (wc60, n_1629);
  or g2306 (n_2146, wc61, n_1630);
  not gc61 (wc61, n_1631);
  or g2307 (n_2149, wc62, n_1640);
  not gc62 (wc62, n_1635);
  or g2308 (n_2225, wc63, n_1730);
  not gc63 (wc63, n_1725);
  or g2309 (n_2228, wc64, n_1726);
  not gc64 (wc64, n_1727);
  or g2310 (n_2231, wc65, n_1736);
  not gc65 (wc65, n_1731);
  and g2311 (n_1941, wc66, n_1629);
  not gc66 (wc66, n_1758);
  and g2312 (n_1765, wc67, n_1762);
  not gc67 (wc67, n_1757);
  or g2313 (n_1937, wc68, n_1628);
  not gc68 (wc68, n_1935);
  or g2314 (n_2223, wc69, n_1720);
  not gc69 (wc69, n_1721);
  and g2315 (n_1767, wc70, n_1637);
  not gc70 (wc70, n_1638);
  and g2316 (n_1774, wc71, n_1643);
  not gc71 (wc71, n_1644);
  and g2317 (n_1834, wc72, n_1715);
  not gc72 (wc72, n_1716);
  and g2318 (n_1837, wc73, n_1721);
  not gc73 (wc73, n_1722);
  and g2319 (n_1864, wc74, n_1764);
  not gc74 (wc74, n_1765);
  or g2320 (n_1871, wc75, n_1646);
  not gc75 (wc75, n_1770);
  or g2321 (n_2001, wc76, n_1730);
  not gc76 (wc76, n_1840);
  and g2322 (n_1932, wc77, n_1737);
  not gc77 (wc77, n_1848);
  or g2323 (n_1942, n_1939, wc78);
  not gc78 (wc78, n_1935);
  or g2324 (n_1944, wc79, n_1867);
  not gc79 (wc79, n_1935);
  or g2325 (n_2152, wc80, n_1636);
  not gc80 (wc80, n_1637);
  or g2326 (n_2154, wc81, n_1646);
  not gc81 (wc81, n_1641);
  or g2327 (n_2157, wc82, n_1642);
  not gc82 (wc82, n_1643);
  or g2328 (n_2158, wc83, n_1652);
  not gc83 (wc83, n_1647);
  or g2329 (n_2215, wc84, n_1718);
  not gc84 (wc84, n_1713);
  or g2330 (n_2218, wc85, n_1714);
  not gc85 (wc85, n_1715);
  or g2331 (n_2220, wc86, n_1724);
  not gc86 (wc86, n_1719);
  and g2332 (n_1777, wc87, n_1649);
  not gc87 (wc87, n_1650);
  and g2333 (n_1827, wc88, n_1709);
  not gc88 (wc88, n_1710);
  and g2334 (n_1775, wc89, n_1772);
  not gc89 (wc89, n_1767);
  or g2335 (n_1916, wc90, n_1718);
  not gc90 (wc90, n_1830);
  and g2336 (n_1845, wc91, n_1842);
  not gc91 (wc91, n_1837);
  and g2337 (n_1869, wc92, n_1770);
  not gc92 (wc92, n_1864);
  and g2338 (n_1948, wc93, n_1770);
  not gc93 (wc93, n_1867);
  and g2339 (n_2014, wc94, n_1850);
  not gc94 (wc94, n_1927);
  or g2340 (n_2161, wc95, n_1648);
  not gc95 (wc95, n_1649);
  or g2341 (n_2210, wc96, n_1712);
  not gc96 (wc96, n_1707);
  or g2342 (n_2213, wc97, n_1708);
  not gc97 (wc97, n_1709);
  and g2343 (n_1784, wc98, n_1655);
  not gc98 (wc98, n_1656);
  and g2344 (n_1824, wc99, n_1703);
  not gc99 (wc99, n_1704);
  and g2345 (n_1872, wc100, n_1641);
  not gc100 (wc100, n_1768);
  and g2346 (n_1876, wc101, n_1774);
  not gc101 (wc101, n_1775);
  or g2347 (n_2028, wc102, n_1658);
  not gc102 (wc102, n_1780);
  and g2348 (n_1835, wc103, n_1832);
  not gc103 (wc103, n_1827);
  and g2349 (n_2002, wc104, n_1725);
  not gc104 (wc104, n_1838);
  and g2350 (n_1924, wc105, n_1844);
  not gc105 (wc105, n_1845);
  and g2351 (n_1946, wc106, n_1635);
  not gc106 (wc106, n_1865);
  and g2352 (n_1949, wc107, n_1767);
  not gc107 (wc107, n_1869);
  or g2353 (n_2163, wc108, n_1658);
  not gc108 (wc108, n_1653);
  or g2354 (n_2166, wc109, n_1654);
  not gc109 (wc109, n_1655);
  or g2355 (n_2202, wc110, n_1696);
  not gc110 (wc110, n_1697);
  or g2356 (n_2204, wc111, n_1706);
  not gc111 (wc111, n_1701);
  or g2357 (n_2207, wc112, n_1702);
  not gc112 (wc112, n_1703);
  and g2358 (n_2030, wc113, n_1653);
  not gc113 (wc113, n_1778);
  and g2359 (n_1785, wc114, n_1782);
  not gc114 (wc114, n_1777);
  and g2360 (n_1917, wc115, n_1713);
  not gc115 (wc115, n_1828);
  and g2361 (n_1921, wc116, n_1834);
  not gc116 (wc116, n_1835);
  and g2362 (n_1929, wc117, n_1850);
  not gc117 (wc117, n_1924);
  and g2363 (n_1787, wc118, n_1661);
  not gc118 (wc118, n_1662);
  and g2364 (n_1794, wc119, n_1667);
  not gc119 (wc119, n_1668);
  and g2365 (n_1879, wc120, n_1784);
  not gc120 (wc120, n_1785);
  or g2366 (n_1886, wc121, n_1670);
  not gc121 (wc121, n_1790);
  and g2367 (n_1952, n_1872, wc122);
  not gc122 (wc122, n_1873);
  and g2368 (n_1955, n_1876, wc123);
  not gc123 (wc123, n_1877);
  and g2369 (n_2011, wc124, n_1731);
  not gc124 (wc124, n_1925);
  and g2370 (n_2016, wc125, n_1847);
  not gc125 (wc125, n_1929);
  and g2371 (n_2021, n_1932, wc126);
  not gc126 (wc126, n_1933);
  or g2372 (n_2169, wc127, n_1664);
  not gc127 (wc127, n_1659);
  or g2373 (n_2172, wc128, n_1660);
  not gc128 (wc128, n_1661);
  or g2374 (n_2174, wc129, n_1670);
  not gc129 (wc129, n_1665);
  or g2375 (n_2177, wc130, n_1666);
  not gc130 (wc130, n_1667);
  or g2376 (n_2179, wc131, n_1676);
  not gc131 (wc131, n_1671);
  or g2377 (n_2187, wc132, n_1678);
  not gc132 (wc132, n_1679);
  and g2378 (n_1797, wc133, n_1673);
  not gc133 (wc133, n_1674);
  and g2379 (n_1795, wc134, n_1792);
  not gc134 (wc134, n_1787);
  and g2380 (n_1884, wc135, n_1790);
  not gc135 (wc135, n_1879);
  and g2381 (n_2037, wc136, n_1790);
  not gc136 (wc136, n_1882);
  or g2382 (n_2182, wc137, n_1672);
  not gc137 (wc137, n_1673);
  or g2383 (n_2190, wc138, n_1688);
  not gc138 (wc138, n_1683);
  and g2384 (n_1804, wc139, n_1679);
  not gc139 (wc139, n_1680);
  and g2385 (n_1807, wc140, n_1685);
  not gc140 (wc140, n_1686);
  and g2386 (n_1814, wc141, n_1691);
  not gc141 (wc141, n_1692);
  and g2387 (n_1817, wc142, n_1697);
  not gc142 (wc142, n_1698);
  and g2388 (n_1887, wc143, n_1665);
  not gc143 (wc143, n_1788);
  and g2389 (n_1891, wc144, n_1794);
  not gc144 (wc144, n_1795);
  or g2390 (n_1965, wc145, n_1682);
  not gc145 (wc145, n_1800);
  or g2391 (n_1901, wc146, n_1694);
  not gc146 (wc146, n_1810);
  or g2392 (n_2080, wc147, n_1706);
  not gc147 (wc147, n_1820);
  and g2393 (n_2035, wc148, n_1659);
  not gc148 (wc148, n_1880);
  and g2394 (n_2038, wc149, n_1787);
  not gc149 (wc149, n_1884);
  or g2395 (n_2044, wc150, n_1676);
  not gc150 (wc150, n_1960);
  or g2396 (n_2026, wc151, n_1652);
  not gc151 (wc151, n_2024);
  or g2397 (n_2031, n_2028, wc152);
  not gc152 (wc152, n_2024);
  or g2398 (n_2033, wc153, n_1882);
  not gc153 (wc153, n_2024);
  or g2399 (n_2184, wc154, n_1682);
  not gc154 (wc154, n_1677);
  or g2400 (n_2193, wc155, n_1684);
  not gc155 (wc155, n_1685);
  or g2401 (n_2195, wc156, n_1694);
  not gc156 (wc156, n_1689);
  or g2402 (n_2198, wc157, n_1690);
  not gc157 (wc157, n_1691);
  or g2403 (n_2199, wc158, n_1700);
  not gc158 (wc158, n_1695);
  and g2404 (n_1966, wc159, n_1677);
  not gc159 (wc159, n_1798);
  and g2405 (n_1805, wc160, n_1802);
  not gc160 (wc160, n_1797);
  and g2406 (n_1815, wc161, n_1812);
  not gc161 (wc161, n_1807);
  and g2407 (n_1825, wc162, n_1822);
  not gc162 (wc162, n_1817);
  and g2408 (n_1978, wc163, n_1810);
  not gc163 (wc163, n_1897);
  and g2409 (n_2089, wc164, n_1830);
  not gc164 (wc164, n_1912);
  and g2410 (n_1894, wc165, n_1804);
  not gc165 (wc165, n_1805);
  and g2411 (n_1902, wc166, n_1689);
  not gc166 (wc166, n_1808);
  and g2412 (n_1906, wc167, n_1814);
  not gc167 (wc167, n_1815);
  and g2413 (n_2082, wc168, n_1701);
  not gc168 (wc168, n_1818);
  and g2414 (n_1909, wc169, n_1824);
  not gc169 (wc169, n_1825);
  and g2415 (n_2041, n_1887, wc170);
  not gc170 (wc170, n_1888);
  and g2416 (n_1957, n_1891, wc171);
  not gc171 (wc171, n_1892);
  or g2417 (n_2052, n_1965, wc172);
  not gc172 (wc172, n_1960);
  or g2418 (n_2056, wc173, n_1897);
  not gc173 (wc173, n_1960);
  or g2419 (n_2096, wc174, n_1724);
  not gc174 (wc174, n_1996);
  or g2420 (n_2104, n_2001, wc175);
  not gc175 (wc175, n_1996);
  or g2421 (n_2108, wc176, n_1927);
  not gc176 (wc176, n_1996);
  or g2422 (n_2047, n_2044, wc177);
  not gc177 (wc177, n_2024);
  or g2423 (n_2051, n_2048, wc178);
  not gc178 (wc178, n_2024);
  and g2424 (n_1899, wc179, n_1810);
  not gc179 (wc179, n_1894);
  and g2425 (n_1914, wc180, n_1830);
  not gc180 (wc180, n_1909);
  and g2426 (n_1963, wc181, n_1800);
  not gc181 (wc181, n_1957);
  and g2427 (n_1976, wc182, n_1973);
  not gc182 (wc182, n_1957);
  and g2428 (n_1981, wc183, n_1978);
  not gc183 (wc183, n_1957);
  and g2429 (n_1986, wc184, n_1983);
  not gc184 (wc184, n_1957);
  and g2430 (n_1991, wc185, n_1988);
  not gc185 (wc185, n_1957);
  and g2431 (n_1975, wc186, n_1683);
  not gc186 (wc186, n_1895);
  and g2432 (n_1980, wc187, n_1807);
  not gc187 (wc187, n_1899);
  and g2433 (n_1985, n_1902, wc188);
  not gc188 (wc188, n_1903);
  and g2434 (n_1990, n_1906, wc189);
  not gc189 (wc189, n_1907);
  and g2435 (n_2087, wc190, n_1707);
  not gc190 (wc190, n_1910);
  and g2436 (n_2090, wc191, n_1827);
  not gc191 (wc191, n_1914);
  and g2437 (n_2093, n_1917, wc192);
  not gc192 (wc192, n_1918);
  and g2438 (n_1993, n_1921, wc193);
  not gc193 (wc193, n_1922);
  and g2439 (n_2046, wc194, n_1671);
  not gc194 (wc194, n_1958);
  and g2440 (n_2050, wc195, n_1797);
  not gc195 (wc195, n_1963);
  and g2441 (n_2054, n_1966, wc196);
  not gc196 (wc196, n_1967);
  and g2442 (n_2058, n_1894, wc197);
  not gc197 (wc197, n_1970);
  or g2443 (n_2055, n_2052, wc198);
  not gc198 (wc198, n_2024);
  or g2444 (n_2059, n_2056, wc199);
  not gc199 (wc199, n_2024);
  or g2445 (n_2063, n_2060, wc200);
  not gc200 (wc200, n_2024);
  or g2446 (n_2067, n_2064, wc201);
  not gc201 (wc201, n_2024);
  or g2447 (n_2071, n_2068, wc202);
  not gc202 (wc202, n_2024);
  or g2448 (n_2075, n_2072, wc203);
  not gc203 (wc203, n_2024);
  and g2449 (n_1999, wc204, n_1840);
  not gc204 (wc204, n_1993);
  and g2450 (n_2012, wc205, n_2009);
  not gc205 (wc205, n_1993);
  and g2451 (n_2017, wc206, n_2014);
  not gc206 (wc206, n_1993);
  and g2452 (n_2022, wc207, n_2019);
  not gc207 (wc207, n_1993);
  and g2453 (n_2062, n_1975, wc208);
  not gc208 (wc208, n_1976);
  and g2454 (n_2066, n_1980, wc209);
  not gc209 (wc209, n_1981);
  and g2455 (n_2070, n_1985, wc210);
  not gc210 (wc210, n_1986);
  and g2456 (n_2074, n_1990, wc211);
  not gc211 (wc211, n_1991);
  and g2457 (n_2098, wc212, n_1719);
  not gc212 (wc212, n_1994);
  and g2458 (n_2102, wc213, n_1837);
  not gc213 (wc213, n_1999);
  and g2459 (n_2106, n_2002, wc214);
  not gc214 (wc214, n_2003);
  and g2460 (n_2110, n_1924, wc215);
  not gc215 (wc215, n_2006);
  and g2461 (n_2114, wc216, n_2011);
  not gc216 (wc216, n_2012);
  and g2462 (n_2118, wc217, n_2016);
  not gc217 (wc217, n_2017);
  and g2463 (n_2122, wc218, n_2021);
  not gc218 (wc218, n_2022);
  or g2464 (n_2078, wc219, n_1700);
  not gc219 (wc219, n_2076);
  or g2465 (n_2083, n_2080, wc220);
  not gc220 (wc220, n_2076);
  or g2466 (n_2085, wc221, n_1912);
  not gc221 (wc221, n_2076);
  or g2467 (n_2099, n_2096, wc222);
  not gc222 (wc222, n_2076);
  or g2468 (n_2103, wc223, n_2100);
  not gc223 (wc223, n_2076);
  or g2469 (n_2107, n_2104, wc224);
  not gc224 (wc224, n_2076);
  or g2470 (n_2111, n_2108, wc225);
  not gc225 (wc225, n_2076);
  or g2471 (n_2115, wc226, n_2112);
  not gc226 (wc226, n_2076);
  or g2472 (n_2119, wc227, n_2116);
  not gc227 (wc227, n_2076);
  or g2473 (n_2123, wc228, n_2120);
  not gc228 (wc228, n_2076);
endmodule

module mult_signed_const_4952_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_4952_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_5219_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_176;
  wire n_178, n_179, n_180, n_183, n_184, n_187, n_188, n_189;
  wire n_196, n_200, n_201, n_202, n_203, n_204, n_207, n_209;
  wire n_210, n_211, n_212, n_217, n_218, n_219, n_220, n_221;
  wire n_223, n_224, n_225, n_226, n_227, n_233, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_244, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_257, n_259, n_260, n_261;
  wire n_262, n_267, n_270, n_272, n_273, n_274, n_275, n_276;
  wire n_277, n_282, n_283, n_284, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_298, n_300, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_317;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_334, n_335, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_349, n_351, n_353, n_354, n_355;
  wire n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_366, n_367, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477;
  wire n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485;
  wire n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539;
  wire n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_588, n_589, n_590, n_591, n_592, n_596, n_597;
  wire n_598, n_599, n_603, n_604, n_605, n_606, n_609, n_610;
  wire n_611, n_614, n_622, n_623, n_624, n_625, n_626, n_627;
  wire n_628, n_629, n_630, n_631, n_632, n_633, n_634, n_635;
  wire n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_646;
  wire n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_658;
  wire n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_668;
  wire n_669, n_670, n_671, n_672, n_673, n_674, n_675, n_676;
  wire n_677, n_684, n_685, n_686, n_687, n_688, n_689, n_690;
  wire n_691, n_692, n_693, n_698, n_699, n_701, n_702, n_703;
  wire n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711;
  wire n_712, n_713, n_722, n_723, n_724, n_725, n_726, n_727;
  wire n_728, n_729, n_730, n_731, n_732, n_733, n_738, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_752, n_753, n_764, n_765, n_766, n_767, n_768;
  wire n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776;
  wire n_777, n_788, n_789, n_790, n_791, n_792, n_793, n_794;
  wire n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802;
  wire n_803, n_804, n_805, n_814, n_815, n_818, n_819, n_820;
  wire n_821, n_822, n_823, n_824, n_825, n_826, n_827, n_828;
  wire n_829, n_830, n_831, n_832, n_833, n_846, n_847, n_848;
  wire n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856;
  wire n_857, n_858, n_859, n_860, n_861, n_868, n_869, n_870;
  wire n_871, n_872, n_873, n_878, n_879, n_880, n_881, n_882;
  wire n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890;
  wire n_891, n_892, n_893, n_904, n_906, n_907, n_908, n_909;
  wire n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917;
  wire n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925;
  wire n_926, n_927, n_928, n_929, n_942, n_943, n_944, n_948;
  wire n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956;
  wire n_957, n_958, n_959, n_960, n_961, n_962, n_963, n_964;
  wire n_965, n_982, n_983, n_984, n_986, n_987, n_988, n_989;
  wire n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997;
  wire n_998, n_999, n_1000, n_1001, n_1013, n_1014, n_1015, n_1016;
  wire n_1018, n_1019, n_1020, n_1022, n_1023, n_1025, n_1026, n_1027;
  wire n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035;
  wire n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1044;
  wire n_1045, n_1046, n_1047, n_1049, n_1050, n_1051, n_1052, n_1054;
  wire n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062;
  wire n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070;
  wire n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078;
  wire n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086;
  wire n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094;
  wire n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102;
  wire n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110;
  wire n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118;
  wire n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126;
  wire n_1127, n_1128, n_1129, n_1132, n_1133, n_1134, n_1135, n_1136;
  wire n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1144, n_1145;
  wire n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153;
  wire n_1154, n_1155, n_1156, n_1158, n_1159, n_1160, n_1161, n_1162;
  wire n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170;
  wire n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178;
  wire n_1179, n_1180, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187;
  wire n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195;
  wire n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205;
  wire n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213;
  wire n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221;
  wire n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229;
  wire n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237;
  wire n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
  wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1252, n_1253, n_1254;
  wire n_1255, n_1256, n_1257, n_1258, n_1259, n_1261, n_1262, n_1263;
  wire n_1264, n_1265, n_1266, n_1268, n_1269, n_1270, n_1271, n_1272;
  wire n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281;
  wire n_1282, n_1283, n_1284, n_1285, n_1286, n_1288, n_1290, n_1291;
  wire n_1292, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300;
  wire n_1301, n_1302, n_1303, n_1305, n_1306, n_1307, n_1308, n_1309;
  wire n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317;
  wire n_1318, n_1319, n_1320, n_1321, n_1325, n_1326, n_1327, n_1328;
  wire n_1329, n_1330, n_1331, n_1333, n_1334, n_1335, n_1337, n_1338;
  wire n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346;
  wire n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1355;
  wire n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363;
  wire n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372;
  wire n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380;
  wire n_1381, n_1385, n_1386, n_1388, n_1389, n_1390, n_1391, n_1393;
  wire n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403;
  wire n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1412, n_1414;
  wire n_1415, n_1416, n_1417, n_1418, n_1419, n_1421, n_1422, n_1423;
  wire n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431;
  wire n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1440;
  wire n_1441, n_1442, n_1445, n_1446, n_1448, n_1449, n_1450, n_1451;
  wire n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1468;
  wire n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476;
  wire n_1477, n_1478, n_1479, n_1480, n_1481, n_1485, n_1488, n_1489;
  wire n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
  wire n_1498, n_1499, n_1500, n_1501, n_1504, n_1506, n_1507, n_1508;
  wire n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519;
  wire n_1520, n_1521, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533;
  wire n_1534, n_1535, n_1536, n_1537, n_1541, n_1542, n_1543, n_1544;
  wire n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1553, n_1555;
  wire n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1566, n_1567;
  wire n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1578, n_1580;
  wire n_1581, n_1583, n_1584, n_1585, n_1587, n_1588, n_1589, n_1590;
  wire n_1591, n_1593, n_1604, n_1605, n_1606, n_1607, n_1609, n_1610;
  wire n_1611, n_1612, n_1613, n_1615, n_1616, n_1617, n_1618, n_1619;
  wire n_1621, n_1622, n_1623, n_1624, n_1625, n_1627, n_1628, n_1629;
  wire n_1630, n_1631, n_1633, n_1634, n_1635, n_1636, n_1637, n_1639;
  wire n_1640, n_1641, n_1642, n_1643, n_1645, n_1646, n_1647, n_1648;
  wire n_1649, n_1651, n_1652, n_1653, n_1654, n_1655, n_1657, n_1658;
  wire n_1659, n_1660, n_1661, n_1663, n_1664, n_1665, n_1666, n_1667;
  wire n_1669, n_1670, n_1671, n_1672, n_1673, n_1675, n_1676, n_1677;
  wire n_1678, n_1679, n_1681, n_1682, n_1683, n_1684, n_1685, n_1687;
  wire n_1688, n_1689, n_1690, n_1691, n_1693, n_1694, n_1695, n_1696;
  wire n_1697, n_1699, n_1700, n_1701, n_1702, n_1703, n_1705, n_1706;
  wire n_1707, n_1708, n_1709, n_1711, n_1712, n_1713, n_1714, n_1715;
  wire n_1717, n_1718, n_1719, n_1720, n_1721, n_1723, n_1724, n_1725;
  wire n_1726, n_1727, n_1729, n_1730, n_1731, n_1732, n_1733, n_1735;
  wire n_1736, n_1737, n_1738, n_1739, n_1744, n_1746, n_1747, n_1749;
  wire n_1751, n_1753, n_1754, n_1756, n_1757, n_1759, n_1761, n_1763;
  wire n_1764, n_1766, n_1767, n_1769, n_1771, n_1773, n_1774, n_1776;
  wire n_1777, n_1779, n_1781, n_1783, n_1784, n_1786, n_1787, n_1789;
  wire n_1791, n_1793, n_1794, n_1796, n_1797, n_1799, n_1801, n_1803;
  wire n_1804, n_1806, n_1807, n_1809, n_1811, n_1813, n_1814, n_1816;
  wire n_1817, n_1819, n_1821, n_1823, n_1824, n_1826, n_1827, n_1829;
  wire n_1831, n_1833, n_1834, n_1836, n_1837, n_1839, n_1841, n_1843;
  wire n_1844, n_1846, n_1847, n_1849, n_1853, n_1854, n_1855, n_1857;
  wire n_1858, n_1859, n_1861, n_1862, n_1863, n_1864, n_1866, n_1868;
  wire n_1870, n_1871, n_1872, n_1874, n_1875, n_1876, n_1878, n_1879;
  wire n_1881, n_1883, n_1885, n_1886, n_1887, n_1889, n_1890, n_1891;
  wire n_1893, n_1894, n_1896, n_1898, n_1900, n_1901, n_1902, n_1904;
  wire n_1905, n_1906, n_1908, n_1909, n_1911, n_1913, n_1915, n_1916;
  wire n_1917, n_1919, n_1920, n_1921, n_1923, n_1924, n_1926, n_1928;
  wire n_1930, n_1931, n_1932, n_1934, n_1936, n_1937, n_1938, n_1940;
  wire n_1941, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949;
  wire n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957;
  wire n_1959, n_1962, n_1964, n_1965, n_1966, n_1969, n_1972, n_1974;
  wire n_1975, n_1977, n_1979, n_1980, n_1982, n_1984, n_1985, n_1987;
  wire n_1989, n_1990, n_1992, n_1993, n_1995, n_1998, n_2000, n_2001;
  wire n_2002, n_2005, n_2008, n_2010, n_2011, n_2013, n_2015, n_2016;
  wire n_2018, n_2020, n_2021, n_2023, n_2025, n_2026, n_2027, n_2029;
  wire n_2030, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038;
  wire n_2039, n_2040, n_2041, n_2042, n_2043, n_2045, n_2046, n_2047;
  wire n_2049, n_2050, n_2051, n_2053, n_2054, n_2055, n_2057, n_2058;
  wire n_2059, n_2061, n_2062, n_2063, n_2065, n_2066, n_2067, n_2069;
  wire n_2070, n_2071, n_2073, n_2074, n_2075, n_2077, n_2078, n_2079;
  wire n_2081, n_2082, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089;
  wire n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2097, n_2098;
  wire n_2099, n_2101, n_2102, n_2103, n_2105, n_2106, n_2107, n_2109;
  wire n_2110, n_2111, n_2113, n_2114, n_2115, n_2117, n_2118, n_2119;
  wire n_2121, n_2122, n_2124, n_2127, n_2128, n_2130, n_2131, n_2132;
  wire n_2133, n_2135, n_2136, n_2137, n_2139, n_2140, n_2141, n_2142;
  wire n_2144, n_2145, n_2147, n_2148, n_2150, n_2151, n_2152, n_2153;
  wire n_2155, n_2156, n_2157, n_2159, n_2160, n_2161, n_2162, n_2164;
  wire n_2165, n_2167, n_2168, n_2170, n_2171, n_2172, n_2173, n_2175;
  wire n_2176, n_2177, n_2178, n_2180, n_2181, n_2182, n_2183, n_2185;
  wire n_2186, n_2188, n_2189, n_2191, n_2192, n_2193, n_2194, n_2196;
  wire n_2197, n_2198, n_2200, n_2201, n_2202, n_2203, n_2205, n_2206;
  wire n_2208, n_2209, n_2211, n_2212, n_2213, n_2214, n_2216, n_2217;
  wire n_2218, n_2219, n_2221, n_2222, n_2223, n_2224, n_2226, n_2227;
  wire n_2229, n_2230, n_2232, n_2233, n_2234, n_2235, n_2237, n_2238;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], n_171);
  xor g270 (n_117, n_622, A[2]);
  nand g3 (n_623, A[1], n_171);
  nand g271 (n_624, A[2], n_171);
  nand g272 (n_625, A[1], A[2]);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, A[4]);
  xor g288 (n_176, n_634, n_69);
  nand g289 (n_635, n_68, A[4]);
  nand g290 (n_636, n_69, A[4]);
  nand g291 (n_637, n_68, n_69);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_176);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_176);
  nand g296 (n_640, A[7], n_176);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g299 (n_642, A[1], A[2]);
  xor g300 (n_178, n_642, n_171);
  xor g305 (n_646, n_178, A[5]);
  xor g306 (n_180, n_646, A[6]);
  nand g307 (n_647, n_178, A[5]);
  nand g308 (n_648, A[6], A[5]);
  nand g309 (n_649, n_178, A[6]);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, n_179, n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, n_179, n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, n_179, A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_188, n_659, n_660, n_661);
  xor g329 (n_662, n_183, n_184);
  xor g330 (n_112, n_662, A[9]);
  nand g331 (n_663, n_183, n_184);
  nand g332 (n_664, A[9], n_184);
  nand g333 (n_665, n_183, A[9]);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_187, n_630, n_67);
  nand g340 (n_668, n_67, n_173);
  nand g341 (n_669, A[4], n_67);
  nand g342 (n_71, n_631, n_668, n_669);
  xor g343 (n_670, A[7], n_187);
  xor g344 (n_189, n_670, A[8]);
  nand g345 (n_671, A[7], n_187);
  nand g346 (n_672, A[8], n_187);
  nand g347 (n_673, A[7], A[8]);
  nand g348 (n_73, n_671, n_672, n_673);
  xor g349 (n_674, A[10], n_188);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, A[10], n_188);
  nand g352 (n_676, n_189, n_188);
  nand g353 (n_677, A[10], n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_72, n_638, n_71);
  nand g366 (n_684, n_71, n_176);
  nand g367 (n_685, A[5], n_71);
  nand g368 (n_201, n_639, n_684, n_685);
  xor g369 (n_686, A[8], A[9]);
  xor g370 (n_196, n_686, A[11]);
  nand g371 (n_687, A[8], A[9]);
  nand g372 (n_688, A[11], A[9]);
  nand g373 (n_689, A[8], A[11]);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, n_73, n_72);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, n_73, n_72);
  nand g378 (n_692, n_196, n_72);
  nand g379 (n_693, n_73, n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g387 (n_698, n_117, A[5]);
  xor g388 (n_200, n_698, A[6]);
  nand g389 (n_699, n_117, A[5]);
  nand g391 (n_701, n_117, A[6]);
  nand g392 (n_207, n_699, n_648, n_701);
  xor g393 (n_702, n_179, n_200);
  xor g394 (n_202, n_702, A[10]);
  nand g395 (n_703, n_179, n_200);
  nand g396 (n_704, A[10], n_200);
  nand g397 (n_705, n_179, A[10]);
  nand g398 (n_209, n_703, n_704, n_705);
  xor g399 (n_706, A[9], A[12]);
  xor g400 (n_204, n_706, n_201);
  nand g401 (n_707, A[9], A[12]);
  nand g402 (n_708, n_201, A[12]);
  nand g403 (n_709, A[9], n_201);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, n_202, n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, n_202, n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, n_202, n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g423 (n_722, n_207, A[10]);
  xor g424 (n_210, n_722, n_184);
  nand g425 (n_723, n_207, A[10]);
  nand g426 (n_724, n_184, A[10]);
  nand g427 (n_725, n_207, n_184);
  nand g428 (n_217, n_723, n_724, n_725);
  xor g429 (n_726, A[11], A[13]);
  xor g430 (n_212, n_726, n_209);
  nand g431 (n_727, A[11], A[13]);
  nand g432 (n_728, n_209, A[13]);
  nand g433 (n_729, A[11], n_209);
  nand g434 (n_220, n_727, n_728, n_729);
  xor g435 (n_730, n_210, n_211);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, n_210, n_211);
  nand g438 (n_732, n_212, n_211);
  nand g439 (n_733, n_210, n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_218, n_738, n_187);
  xor g455 (n_742, n_188, A[11]);
  xor g456 (n_219, n_742, A[12]);
  nand g457 (n_743, n_188, A[11]);
  nand g458 (n_744, A[12], A[11]);
  nand g459 (n_745, n_188, A[12]);
  nand g460 (n_224, n_743, n_744, n_745);
  xor g461 (n_746, A[14], n_217);
  xor g462 (n_221, n_746, n_218);
  nand g463 (n_747, A[14], n_217);
  nand g464 (n_748, n_218, n_217);
  nand g465 (n_749, A[14], n_218);
  nand g466 (n_225, n_747, n_748, n_749);
  xor g467 (n_750, n_219, n_220);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, n_219, n_220);
  nand g470 (n_752, n_221, n_220);
  nand g471 (n_753, n_219, n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g488 (n_223, n_686, n_72);
  nand g490 (n_764, n_72, A[9]);
  nand g491 (n_765, A[8], n_72);
  nand g492 (n_234, n_687, n_764, n_765);
  xor g493 (n_766, A[12], n_73);
  xor g494 (n_226, n_766, A[13]);
  nand g495 (n_767, A[12], n_73);
  nand g496 (n_768, A[13], n_73);
  nand g497 (n_769, A[12], A[13]);
  nand g498 (n_236, n_767, n_768, n_769);
  xor g499 (n_770, A[15], n_223);
  xor g500 (n_227, n_770, n_224);
  nand g501 (n_771, A[15], n_223);
  nand g502 (n_772, n_224, n_223);
  nand g503 (n_773, A[15], n_224);
  nand g504 (n_238, n_771, n_772, n_773);
  xor g505 (n_774, n_225, n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, n_225, n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, n_225, n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g524 (n_233, n_650, A[9]);
  nand g526 (n_788, A[9], n_180);
  nand g527 (n_789, n_179, A[9]);
  nand g528 (n_244, n_651, n_788, n_789);
  xor g529 (n_790, A[10], n_201);
  xor g530 (n_235, n_790, A[13]);
  nand g531 (n_791, A[10], n_201);
  nand g532 (n_792, A[13], n_201);
  nand g533 (n_793, A[10], A[13]);
  nand g534 (n_246, n_791, n_792, n_793);
  xor g535 (n_794, A[14], n_233);
  xor g536 (n_237, n_794, n_234);
  nand g537 (n_795, A[14], n_233);
  nand g538 (n_796, n_234, n_233);
  nand g539 (n_797, A[14], n_234);
  nand g540 (n_248, n_795, n_796, n_797);
  xor g541 (n_798, A[16], n_235);
  xor g542 (n_239, n_798, n_236);
  nand g543 (n_799, A[16], n_235);
  nand g544 (n_800, n_236, n_235);
  nand g545 (n_801, A[16], n_236);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, n_237, n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, n_237, n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, n_237, n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g565 (n_814, n_183, A[10]);
  xor g566 (n_245, n_814, n_184);
  nand g567 (n_815, n_183, A[10]);
  nand g570 (n_257, n_815, n_724, n_663);
  xor g571 (n_818, A[11], A[14]);
  xor g572 (n_247, n_818, n_244);
  nand g573 (n_819, A[11], A[14]);
  nand g574 (n_820, n_244, A[14]);
  nand g575 (n_821, A[11], n_244);
  nand g576 (n_259, n_819, n_820, n_821);
  xor g577 (n_822, A[15], n_245);
  xor g578 (n_249, n_822, n_246);
  nand g579 (n_823, A[15], n_245);
  nand g580 (n_824, n_246, n_245);
  nand g581 (n_825, A[15], n_246);
  nand g582 (n_261, n_823, n_824, n_825);
  xor g583 (n_826, n_247, A[17]);
  xor g584 (n_251, n_826, n_248);
  nand g585 (n_827, n_247, A[17]);
  nand g586 (n_828, n_248, A[17]);
  nand g587 (n_829, n_247, n_248);
  nand g588 (n_118, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g615 (n_846, n_218, n_257);
  xor g616 (n_260, n_846, A[15]);
  nand g617 (n_847, n_218, n_257);
  nand g618 (n_848, A[15], n_257);
  nand g619 (n_849, n_218, A[15]);
  nand g620 (n_272, n_847, n_848, n_849);
  xor g621 (n_850, n_219, n_259);
  xor g622 (n_262, n_850, A[16]);
  nand g623 (n_851, n_219, n_259);
  nand g624 (n_852, A[16], n_259);
  nand g625 (n_853, n_219, A[16]);
  nand g626 (n_273, n_851, n_852, n_853);
  xor g627 (n_854, n_260, A[18]);
  xor g628 (n_119, n_854, n_261);
  nand g629 (n_855, n_260, A[18]);
  nand g630 (n_856, n_261, A[18]);
  nand g631 (n_857, n_260, n_261);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_262, n_118);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_262, n_118);
  nand g636 (n_860, n_119, n_118);
  nand g637 (n_861, n_262, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g648 (n_267, n_638, A[8]);
  nand g650 (n_868, A[8], n_176);
  nand g651 (n_869, A[5], A[8]);
  nand g652 (n_282, n_639, n_868, n_869);
  xor g653 (n_870, n_71, A[9]);
  xor g654 (n_270, n_870, n_267);
  nand g655 (n_871, n_71, A[9]);
  nand g656 (n_872, n_267, A[9]);
  nand g657 (n_873, n_71, n_267);
  nand g658 (n_284, n_871, n_872, n_873);
  xor g665 (n_878, n_224, n_270);
  xor g666 (n_274, n_878, A[16]);
  nand g667 (n_879, n_224, n_270);
  nand g668 (n_880, A[16], n_270);
  nand g669 (n_881, n_224, A[16]);
  nand g670 (n_288, n_879, n_880, n_881);
  xor g671 (n_882, n_226, A[17]);
  xor g672 (n_275, n_882, n_272);
  nand g673 (n_883, n_226, A[17]);
  nand g674 (n_884, n_272, A[17]);
  nand g675 (n_885, n_226, n_272);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, A[19], n_273);
  xor g678 (n_277, n_886, n_274);
  nand g679 (n_887, A[19], n_273);
  nand g680 (n_888, n_274, n_273);
  nand g681 (n_889, A[19], n_274);
  nand g682 (n_291, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g702 (n_283, n_650, A[10]);
  nand g704 (n_904, A[10], n_180);
  nand g706 (n_298, n_651, n_904, n_705);
  xor g707 (n_906, A[9], n_282);
  xor g708 (n_286, n_906, A[13]);
  nand g709 (n_907, A[9], n_282);
  nand g710 (n_908, A[13], n_282);
  nand g711 (n_909, A[9], A[13]);
  nand g712 (n_300, n_907, n_908, n_909);
  xor g713 (n_910, n_283, A[14]);
  xor g714 (n_287, n_910, n_284);
  nand g715 (n_911, n_283, A[14]);
  nand g716 (n_912, n_284, A[14]);
  nand g717 (n_913, n_283, n_284);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, n_236, n_286);
  xor g720 (n_289, n_914, A[18]);
  nand g721 (n_915, n_236, n_286);
  nand g722 (n_916, A[18], n_286);
  nand g723 (n_917, n_236, A[18]);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, A[17], n_287);
  xor g726 (n_292, n_918, A[20]);
  nand g727 (n_919, A[17], n_287);
  nand g728 (n_920, A[20], n_287);
  nand g729 (n_921, A[17], A[20]);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, n_288, n_289);
  xor g732 (n_293, n_922, n_290);
  nand g733 (n_923, n_288, n_289);
  nand g734 (n_924, n_290, n_289);
  nand g735 (n_925, n_288, n_290);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g761 (n_942, A[11], n_298);
  xor g762 (n_301, n_942, A[14]);
  nand g763 (n_943, A[11], n_298);
  nand g764 (n_944, A[14], n_298);
  nand g766 (n_317, n_943, n_944, n_819);
  xor g768 (n_303, n_822, n_300);
  nand g770 (n_948, n_300, n_245);
  nand g771 (n_949, A[15], n_300);
  nand g772 (n_319, n_823, n_948, n_949);
  xor g773 (n_950, A[19], n_301);
  xor g774 (n_305, n_950, A[18]);
  nand g775 (n_951, A[19], n_301);
  nand g776 (n_952, A[18], n_301);
  nand g777 (n_953, A[19], A[18]);
  nand g778 (n_320, n_951, n_952, n_953);
  xor g779 (n_954, n_302, A[21]);
  xor g780 (n_307, n_954, n_303);
  nand g781 (n_955, n_302, A[21]);
  nand g782 (n_956, n_303, A[21]);
  nand g783 (n_957, n_302, n_303);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, n_304, n_305);
  xor g786 (n_309, n_958, n_306);
  nand g787 (n_959, n_304, n_305);
  nand g788 (n_960, n_306, n_305);
  nand g789 (n_961, n_304, n_306);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g823 (n_982, n_219, n_317);
  xor g824 (n_321, n_982, A[16]);
  nand g825 (n_983, n_219, n_317);
  nand g826 (n_984, A[16], n_317);
  nand g828 (n_337, n_983, n_984, n_853);
  xor g829 (n_986, A[19], n_260);
  xor g830 (n_322, n_986, A[20]);
  nand g831 (n_987, A[19], n_260);
  nand g832 (n_988, A[20], n_260);
  nand g833 (n_989, A[19], A[20]);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, A[22], n_319);
  xor g836 (n_324, n_990, n_320);
  nand g837 (n_991, A[22], n_319);
  nand g838 (n_992, n_320, n_319);
  nand g839 (n_993, A[22], n_320);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, n_321, n_322);
  xor g842 (n_326, n_994, n_323);
  nand g843 (n_995, n_321, n_322);
  nand g844 (n_996, n_323, n_322);
  nand g845 (n_997, n_321, n_323);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, n_324, n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, n_324, n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, n_324, n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g868 (n_334, n_870, A[12]);
  nand g871 (n_1013, n_71, A[12]);
  nand g872 (n_354, n_871, n_707, n_1013);
  xor g873 (n_1014, n_73, n_267);
  xor g874 (n_335, n_1014, A[13]);
  nand g875 (n_1015, n_73, n_267);
  nand g876 (n_1016, A[13], n_267);
  nand g878 (n_356, n_1015, n_1016, n_768);
  xor g879 (n_1018, n_224, n_334);
  xor g880 (n_338, n_1018, A[16]);
  nand g881 (n_1019, n_224, n_334);
  nand g882 (n_1020, A[16], n_334);
  nand g884 (n_358, n_1019, n_1020, n_881);
  xor g885 (n_1022, n_335, A[17]);
  xor g886 (n_339, n_1022, n_272);
  nand g887 (n_1023, n_335, A[17]);
  nand g889 (n_1025, n_335, n_272);
  nand g890 (n_359, n_1023, n_884, n_1025);
  xor g891 (n_1026, A[21], A[20]);
  xor g892 (n_341, n_1026, n_337);
  nand g893 (n_1027, A[21], A[20]);
  nand g894 (n_1028, n_337, A[20]);
  nand g895 (n_1029, A[21], n_337);
  nand g896 (n_361, n_1027, n_1028, n_1029);
  xor g897 (n_1030, A[23], n_338);
  xor g898 (n_343, n_1030, n_339);
  nand g899 (n_1031, A[23], n_338);
  nand g900 (n_1032, n_339, n_338);
  nand g901 (n_1033, A[23], n_339);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, n_340, n_341);
  xor g904 (n_345, n_1034, n_342);
  nand g905 (n_1035, n_340, n_341);
  nand g906 (n_1036, n_342, n_341);
  nand g907 (n_1037, n_340, n_342);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, n_343, n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, n_343, n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, n_343, n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  xor g917 (n_1042, A[2], n_171);
  nand g922 (n_371, n_624, n_1044, n_1045);
  xor g923 (n_1046, n_349, A[5]);
  xor g924 (n_351, n_1046, A[6]);
  nand g925 (n_1047, n_349, A[5]);
  nand g927 (n_1049, n_349, A[6]);
  nand g928 (n_373, n_1047, n_648, n_1049);
  xor g929 (n_1050, n_179, n_351);
  xor g930 (n_353, n_1050, A[9]);
  nand g931 (n_1051, n_179, n_351);
  nand g932 (n_1052, A[9], n_351);
  nand g934 (n_375, n_1051, n_1052, n_789);
  xor g935 (n_1054, A[10], n_282);
  xor g936 (n_355, n_1054, A[14]);
  nand g937 (n_1055, A[10], n_282);
  nand g938 (n_1056, A[14], n_282);
  nand g939 (n_1057, A[10], A[14]);
  nand g940 (n_377, n_1055, n_1056, n_1057);
  xor g941 (n_1058, n_353, A[13]);
  xor g942 (n_357, n_1058, n_354);
  nand g943 (n_1059, n_353, A[13]);
  nand g944 (n_1060, n_354, A[13]);
  nand g945 (n_1061, n_353, n_354);
  nand g946 (n_380, n_1059, n_1060, n_1061);
  xor g947 (n_1062, n_355, n_356);
  xor g948 (n_360, n_1062, A[17]);
  nand g949 (n_1063, n_355, n_356);
  nand g950 (n_1064, A[17], n_356);
  nand g951 (n_1065, n_355, A[17]);
  nand g952 (n_381, n_1063, n_1064, n_1065);
  xor g953 (n_1066, A[18], n_357);
  nand g955 (n_1067, A[18], n_357);
  nand g958 (n_384, n_1067, n_1068, n_1069);
  xor g959 (n_1070, A[21], A[22]);
  xor g960 (n_362, n_1070, n_358);
  nand g961 (n_1071, A[21], A[22]);
  nand g962 (n_1072, n_358, A[22]);
  nand g963 (n_1073, A[21], n_358);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, n_359, n_360);
  xor g966 (n_365, n_1074, n_361);
  nand g967 (n_1075, n_359, n_360);
  nand g968 (n_1076, n_361, n_360);
  nand g969 (n_1077, n_359, n_361);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g971 (n_1078, n_362, n_363);
  xor g972 (n_367, n_1078, n_364);
  nand g973 (n_1079, n_362, n_363);
  nand g974 (n_1080, n_364, n_363);
  nand g975 (n_1081, n_362, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  xor g985 (n_1086, A[1], A[3]);
  nand g987 (n_1087, A[1], A[3]);
  nand g990 (n_392, n_1087, n_1088, n_1089);
  xor g991 (n_1090, n_371, A[6]);
  xor g992 (n_374, n_1090, n_372);
  nand g993 (n_1091, n_371, A[6]);
  nand g994 (n_1092, n_372, A[6]);
  nand g995 (n_1093, n_371, n_372);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, A[10]);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, A[10], n_373);
  nand g1001 (n_1097, A[7], A[10]);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, n_374, A[11]);
  xor g1004 (n_378, n_1098, n_375);
  nand g1005 (n_1099, n_374, A[11]);
  nand g1006 (n_1100, n_375, A[11]);
  nand g1007 (n_1101, n_374, n_375);
  nand g1008 (n_398, n_1099, n_1100, n_1101);
  xor g1009 (n_1102, n_376, A[14]);
  xor g1010 (n_379, n_1102, A[15]);
  nand g1011 (n_1103, n_376, A[14]);
  nand g1012 (n_1104, A[15], A[14]);
  nand g1013 (n_1105, n_376, A[15]);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, n_377, n_378);
  xor g1016 (n_382, n_1106, A[19]);
  nand g1017 (n_1107, n_377, n_378);
  nand g1018 (n_1108, A[19], n_378);
  nand g1019 (n_1109, n_377, A[19]);
  nand g1020 (n_403, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, A[18], n_379);
  xor g1022 (n_383, n_1110, n_380);
  nand g1023 (n_1111, A[18], n_379);
  nand g1024 (n_1112, n_380, n_379);
  nand g1025 (n_1113, A[18], n_380);
  nand g1026 (n_404, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, A[22], A[23]);
  xor g1028 (n_386, n_1114, n_381);
  nand g1029 (n_1115, A[22], A[23]);
  nand g1030 (n_1116, n_381, A[23]);
  nand g1031 (n_1117, A[22], n_381);
  nand g1032 (n_407, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_382, n_383);
  xor g1034 (n_388, n_1118, n_384);
  nand g1035 (n_1119, n_382, n_383);
  nand g1036 (n_1120, n_384, n_383);
  nand g1037 (n_1121, n_382, n_384);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, n_385, n_386);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, n_385, n_386);
  nand g1042 (n_1124, n_387, n_386);
  nand g1043 (n_1125, n_385, n_387);
  nand g1044 (n_411, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1052 (n_393, n_626, A[4]);
  nand g1054 (n_1132, A[4], A[2]);
  nand g1055 (n_1133, A[3], A[4]);
  nand g1056 (n_412, n_627, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, A[11], A[12]);
  xor g1070 (n_399, n_1142, n_396);
  nand g1072 (n_1144, n_396, A[12]);
  nand g1073 (n_1145, A[11], n_396);
  nand g1074 (n_418, n_744, n_1144, n_1145);
  xor g1075 (n_1146, n_397, A[15]);
  xor g1076 (n_401, n_1146, n_398);
  nand g1077 (n_1147, n_397, A[15]);
  nand g1078 (n_1148, n_398, A[15]);
  nand g1079 (n_1149, n_397, n_398);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, n_399, A[16]);
  xor g1082 (n_402, n_1150, n_400);
  nand g1083 (n_1151, n_399, A[16]);
  nand g1084 (n_1152, n_400, A[16]);
  nand g1085 (n_1153, n_399, n_400);
  nand g1086 (n_422, n_1151, n_1152, n_1153);
  xor g1088 (n_405, n_1154, A[20]);
  nand g1092 (n_423, n_1155, n_1156, n_989);
  xor g1093 (n_1158, n_401, A[23]);
  xor g1094 (n_406, n_1158, n_402);
  nand g1095 (n_1159, n_401, A[23]);
  nand g1096 (n_1160, n_402, A[23]);
  nand g1097 (n_1161, n_401, n_402);
  nand g1098 (n_426, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_403, n_404);
  xor g1100 (n_409, n_1162, n_405);
  nand g1101 (n_1163, n_403, n_404);
  nand g1102 (n_1164, n_405, n_404);
  nand g1103 (n_1165, n_403, n_405);
  nand g1104 (n_427, n_1163, n_1164, n_1165);
  xor g1105 (n_1166, n_406, n_407);
  xor g1106 (n_410, n_1166, n_408);
  nand g1107 (n_1167, n_406, n_407);
  nand g1108 (n_1168, n_408, n_407);
  nand g1109 (n_1169, n_406, n_408);
  nand g1110 (n_429, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1123 (n_1178, A[8], n_413);
  xor g1124 (n_415, n_1178, A[9]);
  nand g1125 (n_1179, A[8], n_413);
  nand g1126 (n_1180, A[9], n_413);
  nand g1128 (n_435, n_1179, n_1180, n_687);
  xor g1129 (n_1182, n_414, A[12]);
  xor g1130 (n_417, n_1182, n_415);
  nand g1131 (n_1183, n_414, A[12]);
  nand g1132 (n_1184, n_415, A[12]);
  nand g1133 (n_1185, n_414, n_415);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, A[13], n_416);
  xor g1136 (n_420, n_1186, n_417);
  nand g1137 (n_1187, A[13], n_416);
  nand g1138 (n_1188, n_417, n_416);
  nand g1139 (n_1189, A[13], n_417);
  nand g1140 (n_439, n_1187, n_1188, n_1189);
  xor g1141 (n_1190, A[16], n_418);
  xor g1142 (n_421, n_1190, A[17]);
  nand g1143 (n_1191, A[16], n_418);
  nand g1144 (n_1192, A[17], n_418);
  nand g1145 (n_1193, A[16], A[17]);
  nand g1146 (n_440, n_1191, n_1192, n_1193);
  xor g1148 (n_424, n_1194, A[20]);
  nand g1152 (n_442, n_1195, n_1156, n_1027);
  xor g1153 (n_1198, n_419, n_420);
  xor g1154 (n_425, n_1198, n_421);
  nand g1155 (n_1199, n_419, n_420);
  nand g1156 (n_1200, n_421, n_420);
  nand g1157 (n_1201, n_419, n_421);
  nand g1158 (n_444, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_422, n_423);
  xor g1160 (n_428, n_1202, n_424);
  nand g1161 (n_1203, n_422, n_423);
  nand g1162 (n_1204, n_424, n_423);
  nand g1163 (n_1205, n_422, n_424);
  nand g1164 (n_447, n_1203, n_1204, n_1205);
  xor g1165 (n_1206, n_425, n_426);
  xor g1166 (n_430, n_1206, n_427);
  nand g1167 (n_1207, n_425, n_426);
  nand g1168 (n_1208, n_427, n_426);
  nand g1169 (n_1209, n_425, n_427);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, n_433);
  nand g1183 (n_1217, A[6], n_433);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, A[9], A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, A[9], A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, A[9], n_434);
  nand g1190 (n_456, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, A[14], n_435);
  xor g1192 (n_438, n_1222, A[13]);
  nand g1193 (n_1223, A[14], n_435);
  nand g1194 (n_1224, A[13], n_435);
  nand g1195 (n_1225, A[14], A[13]);
  nand g1196 (n_457, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, n_436, n_437);
  xor g1198 (n_441, n_1226, A[18]);
  nand g1199 (n_1227, n_436, n_437);
  nand g1200 (n_1228, A[18], n_437);
  nand g1201 (n_1229, n_436, A[18]);
  nand g1202 (n_460, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, A[17], n_438);
  xor g1204 (n_443, n_1230, A[21]);
  nand g1205 (n_1231, A[17], n_438);
  nand g1206 (n_1232, A[21], n_438);
  nand g1207 (n_1233, A[17], A[21]);
  nand g1208 (n_462, n_1231, n_1232, n_1233);
  xor g1209 (n_1234, A[22], n_439);
  xor g1210 (n_445, n_1234, n_440);
  nand g1211 (n_1235, A[22], n_439);
  nand g1212 (n_1236, n_440, n_439);
  nand g1213 (n_1237, A[22], n_440);
  nand g1214 (n_463, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_441, n_442);
  xor g1216 (n_446, n_1238, n_443);
  nand g1217 (n_1239, n_441, n_442);
  nand g1218 (n_1240, n_443, n_442);
  nand g1219 (n_1241, n_441, n_443);
  nand g1220 (n_465, n_1239, n_1240, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[7], A[5]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], A[11]);
  xor g1242 (n_455, n_1254, n_453);
  nand g1243 (n_1255, A[10], A[11]);
  nand g1244 (n_1256, n_453, A[11]);
  nand g1245 (n_1257, A[10], n_453);
  nand g1246 (n_472, n_1255, n_1256, n_1257);
  xor g1247 (n_1258, n_454, A[14]);
  xor g1248 (n_458, n_1258, A[15]);
  nand g1249 (n_1259, n_454, A[14]);
  nand g1251 (n_1261, n_454, A[15]);
  nand g1252 (n_474, n_1259, n_1104, n_1261);
  xor g1253 (n_1262, n_455, n_456);
  xor g1254 (n_459, n_1262, n_457);
  nand g1255 (n_1263, n_455, n_456);
  nand g1256 (n_1264, n_457, n_456);
  nand g1257 (n_1265, n_455, n_457);
  nand g1258 (n_476, n_1263, n_1264, n_1265);
  xor g1259 (n_1266, A[19], A[18]);
  xor g1260 (n_461, n_1266, n_458);
  nand g1262 (n_1268, n_458, A[18]);
  nand g1263 (n_1269, A[19], n_458);
  nand g1264 (n_478, n_953, n_1268, n_1269);
  xor g1265 (n_1270, A[22], n_459);
  xor g1266 (n_464, n_1270, A[23]);
  nand g1267 (n_1271, A[22], n_459);
  nand g1268 (n_1272, A[23], n_459);
  nand g1270 (n_479, n_1271, n_1272, n_1115);
  xor g1271 (n_1274, n_460, n_461);
  xor g1272 (n_466, n_1274, n_462);
  nand g1273 (n_1275, n_460, n_461);
  nand g1274 (n_1276, n_462, n_461);
  nand g1275 (n_1277, n_460, n_462);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1277 (n_1278, n_463, n_464);
  xor g1278 (n_467, n_1278, n_465);
  nand g1279 (n_1279, n_463, n_464);
  nand g1280 (n_1280, n_465, n_464);
  nand g1281 (n_1281, n_463, n_465);
  nand g1282 (n_485, n_1279, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1289 (n_1286, A[7], A[6]);
  xor g1290 (n_471, n_1286, A[8]);
  nand g1292 (n_1288, A[8], A[6]);
  nand g1294 (n_486, n_661, n_1288, n_673);
  xor g1295 (n_1290, A[11], n_470);
  xor g1296 (n_473, n_1290, A[12]);
  nand g1297 (n_1291, A[11], n_470);
  nand g1298 (n_1292, A[12], n_470);
  nand g1300 (n_487, n_1291, n_1292, n_744);
  xor g1301 (n_1294, n_471, A[15]);
  xor g1302 (n_475, n_1294, n_472);
  nand g1303 (n_1295, n_471, A[15]);
  nand g1304 (n_1296, n_472, A[15]);
  nand g1305 (n_1297, n_471, n_472);
  nand g1306 (n_489, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, n_473, A[16]);
  xor g1308 (n_477, n_1298, A[19]);
  nand g1309 (n_1299, n_473, A[16]);
  nand g1310 (n_1300, A[19], A[16]);
  nand g1311 (n_1301, n_473, A[19]);
  nand g1312 (n_492, n_1299, n_1300, n_1301);
  xor g1314 (n_480, n_1302, A[20]);
  nand g1317 (n_1305, n_474, A[20]);
  nand g1318 (n_493, n_1303, n_1156, n_1305);
  xor g1319 (n_1306, n_475, n_476);
  xor g1320 (n_481, n_1306, A[23]);
  nand g1321 (n_1307, n_475, n_476);
  nand g1322 (n_1308, A[23], n_476);
  nand g1323 (n_1309, n_475, A[23]);
  nand g1324 (n_494, n_1307, n_1308, n_1309);
  xor g1325 (n_1310, n_477, n_478);
  xor g1326 (n_483, n_1310, n_479);
  nand g1327 (n_1311, n_477, n_478);
  nand g1328 (n_1312, n_479, n_478);
  nand g1329 (n_1313, n_477, n_479);
  nand g1330 (n_497, n_1311, n_1312, n_1313);
  xor g1331 (n_1314, n_480, n_481);
  xor g1332 (n_484, n_1314, n_482);
  nand g1333 (n_1315, n_480, n_481);
  nand g1334 (n_1316, n_482, n_481);
  nand g1335 (n_1317, n_480, n_482);
  nand g1336 (n_499, n_1315, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1344 (n_488, n_686, A[12]);
  nand g1347 (n_1325, A[8], A[12]);
  nand g1348 (n_503, n_687, n_707, n_1325);
  xor g1349 (n_1326, n_486, A[13]);
  xor g1350 (n_490, n_1326, n_487);
  nand g1351 (n_1327, n_486, A[13]);
  nand g1352 (n_1328, n_487, A[13]);
  nand g1353 (n_1329, n_486, n_487);
  nand g1354 (n_505, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, n_488, A[16]);
  xor g1356 (n_491, n_1330, A[17]);
  nand g1357 (n_1331, n_488, A[16]);
  nand g1359 (n_1333, n_488, A[17]);
  nand g1360 (n_507, n_1331, n_1193, n_1333);
  xor g1362 (n_495, n_1334, A[20]);
  nand g1365 (n_1337, n_489, A[20]);
  nand g1366 (n_509, n_1335, n_1156, n_1337);
  xor g1367 (n_1338, n_490, A[21]);
  xor g1368 (n_496, n_1338, n_491);
  nand g1369 (n_1339, n_490, A[21]);
  nand g1370 (n_1340, n_491, A[21]);
  nand g1371 (n_1341, n_490, n_491);
  nand g1372 (n_511, n_1339, n_1340, n_1341);
  xor g1373 (n_1342, n_492, n_493);
  xor g1374 (n_498, n_1342, n_494);
  nand g1375 (n_1343, n_492, n_493);
  nand g1376 (n_1344, n_494, n_493);
  nand g1377 (n_1345, n_492, n_494);
  nand g1378 (n_513, n_1343, n_1344, n_1345);
  xor g1379 (n_1346, n_495, n_496);
  xor g1380 (n_500, n_1346, n_497);
  nand g1381 (n_1347, n_495, n_496);
  nand g1382 (n_1348, n_497, n_496);
  nand g1383 (n_1349, n_495, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  nand g1397 (n_1357, A[9], A[14]);
  nand g1398 (n_519, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], n_503);
  xor g1400 (n_506, n_1358, n_504);
  nand g1401 (n_1359, A[13], n_503);
  nand g1402 (n_1360, n_504, n_503);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_522, n_1359, n_1360, n_1361);
  xor g1405 (n_1362, A[18], A[17]);
  xor g1406 (n_508, n_1362, A[21]);
  nand g1407 (n_1363, A[18], A[17]);
  nand g1409 (n_1365, A[18], A[21]);
  nand g1410 (n_523, n_1363, n_1233, n_1365);
  xor g1411 (n_1366, n_505, A[22]);
  xor g1412 (n_510, n_1366, n_506);
  nand g1413 (n_1367, n_505, A[22]);
  nand g1414 (n_1368, n_506, A[22]);
  nand g1415 (n_1369, n_505, n_506);
  nand g1416 (n_525, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_507, n_508);
  xor g1418 (n_512, n_1370, n_509);
  nand g1419 (n_1371, n_507, n_508);
  nand g1420 (n_1372, n_509, n_508);
  nand g1421 (n_1373, n_507, n_509);
  nand g1422 (n_527, n_1371, n_1372, n_1373);
  xor g1423 (n_1374, n_510, n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, n_510, n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, n_510, n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1443 (n_1386, A[14], A[15]);
  xor g1444 (n_521, n_1386, n_519);
  nand g1446 (n_1388, n_519, A[15]);
  nand g1447 (n_1389, A[14], n_519);
  nand g1448 (n_534, n_1104, n_1388, n_1389);
  xor g1449 (n_1390, n_520, A[19]);
  xor g1450 (n_524, n_1390, A[18]);
  nand g1451 (n_1391, n_520, A[19]);
  nand g1453 (n_1393, n_520, A[18]);
  nand g1454 (n_536, n_1391, n_953, n_1393);
  xor g1456 (n_526, n_1114, n_521);
  nand g1458 (n_1396, n_521, A[23]);
  nand g1459 (n_1397, A[22], n_521);
  nand g1460 (n_538, n_1115, n_1396, n_1397);
  xor g1461 (n_1398, n_522, n_523);
  xor g1462 (n_528, n_1398, n_524);
  nand g1463 (n_1399, n_522, n_523);
  nand g1464 (n_1400, n_524, n_523);
  nand g1465 (n_1401, n_522, n_524);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1467 (n_1402, n_525, n_526);
  xor g1468 (n_529, n_1402, n_527);
  nand g1469 (n_1403, n_525, n_526);
  nand g1470 (n_1404, n_527, n_526);
  nand g1471 (n_1405, n_525, n_527);
  nand g1472 (n_543, n_1403, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1480 (n_533, n_1142, A[10]);
  nand g1482 (n_1412, A[10], A[12]);
  nand g1484 (n_544, n_744, n_1412, n_1255);
  xor g1485 (n_1414, A[15], n_532);
  xor g1486 (n_535, n_1414, A[16]);
  nand g1487 (n_1415, A[15], n_532);
  nand g1488 (n_1416, A[16], n_532);
  nand g1489 (n_1417, A[15], A[16]);
  nand g1490 (n_546, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, n_533, A[19]);
  nand g1493 (n_1419, n_533, A[19]);
  nand g1496 (n_547, n_1419, n_1155, n_1421);
  xor g1497 (n_1422, A[20], A[23]);
  xor g1498 (n_539, n_1422, n_534);
  nand g1499 (n_1423, A[20], A[23]);
  nand g1500 (n_1424, n_534, A[23]);
  nand g1501 (n_1425, A[20], n_534);
  nand g1502 (n_550, n_1423, n_1424, n_1425);
  xor g1503 (n_1426, n_535, n_536);
  xor g1504 (n_541, n_1426, n_537);
  nand g1505 (n_1427, n_535, n_536);
  nand g1506 (n_1428, n_537, n_536);
  nand g1507 (n_1429, n_535, n_537);
  nand g1508 (n_551, n_1427, n_1428, n_1429);
  xor g1509 (n_1430, n_538, n_539);
  xor g1510 (n_542, n_1430, n_540);
  nand g1511 (n_1431, n_538, n_539);
  nand g1512 (n_1432, n_540, n_539);
  nand g1513 (n_1433, n_538, n_540);
  nand g1514 (n_554, n_1431, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1521 (n_1438, A[12], A[13]);
  xor g1522 (n_545, n_1438, n_544);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_769, n_1440, n_1441);
  xor g1527 (n_1442, A[16], A[17]);
  xor g1528 (n_548, n_1442, A[21]);
  nand g1531 (n_1445, A[16], A[21]);
  nand g1532 (n_560, n_1193, n_1233, n_1445);
  xor g1534 (n_549, n_1446, n_545);
  nand g1536 (n_1448, n_545, A[20]);
  nand g1538 (n_559, n_1156, n_1448, n_1449);
  xor g1539 (n_1450, n_546, n_547);
  xor g1540 (n_552, n_1450, n_548);
  nand g1541 (n_1451, n_546, n_547);
  nand g1542 (n_1452, n_548, n_547);
  nand g1543 (n_1453, n_546, n_548);
  nand g1544 (n_563, n_1451, n_1452, n_1453);
  xor g1545 (n_1454, n_549, n_550);
  xor g1546 (n_553, n_1454, n_551);
  nand g1547 (n_1455, n_549, n_550);
  nand g1548 (n_1456, n_551, n_550);
  nand g1549 (n_1457, n_549, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  xor g1560 (n_558, n_1462, A[18]);
  nand g1563 (n_1465, A[13], A[18]);
  nand g1564 (n_570, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, A[17], A[21]);
  xor g1566 (n_561, n_1466, n_557);
  nand g1568 (n_1468, n_557, A[21]);
  nand g1569 (n_1469, A[17], n_557);
  nand g1570 (n_572, n_1233, n_1468, n_1469);
  xor g1571 (n_1470, A[22], n_558);
  xor g1572 (n_562, n_1470, n_559);
  nand g1573 (n_1471, A[22], n_558);
  nand g1574 (n_1472, n_559, n_558);
  nand g1575 (n_1473, A[22], n_559);
  nand g1576 (n_574, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, n_560, n_561);
  xor g1578 (n_564, n_1474, n_562);
  nand g1579 (n_1475, n_560, n_561);
  nand g1580 (n_1476, n_562, n_561);
  nand g1581 (n_1477, n_560, n_562);
  nand g1582 (n_576, n_1475, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  xor g1598 (n_571, n_1266, A[22]);
  nand g1600 (n_1488, A[22], A[18]);
  nand g1601 (n_1489, A[19], A[22]);
  nand g1602 (n_580, n_953, n_1488, n_1489);
  xor g1603 (n_1490, A[23], n_569);
  xor g1604 (n_573, n_1490, n_570);
  nand g1605 (n_1491, A[23], n_569);
  nand g1606 (n_1492, n_570, n_569);
  nand g1607 (n_1493, A[23], n_570);
  nand g1608 (n_583, n_1491, n_1492, n_1493);
  xor g1609 (n_1494, n_571, n_572);
  xor g1610 (n_575, n_1494, n_573);
  nand g1611 (n_1495, n_571, n_572);
  nand g1612 (n_1496, n_573, n_572);
  nand g1613 (n_1497, n_571, n_573);
  nand g1614 (n_585, n_1495, n_1496, n_1497);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1622 (n_579, n_1386, A[16]);
  nand g1624 (n_1504, A[16], A[14]);
  nand g1626 (n_586, n_1104, n_1504, n_1417);
  xor g1627 (n_1506, A[19], n_578);
  nand g1629 (n_1507, A[19], n_578);
  nand g1632 (n_588, n_1507, n_1508, n_1155);
  xor g1634 (n_582, n_1422, n_579);
  nand g1636 (n_1512, n_579, A[23]);
  nand g1637 (n_1513, A[20], n_579);
  nand g1638 (n_589, n_1423, n_1512, n_1513);
  xor g1639 (n_1514, n_580, n_581);
  xor g1640 (n_584, n_1514, n_582);
  nand g1641 (n_1515, n_580, n_581);
  nand g1642 (n_1516, n_582, n_581);
  nand g1643 (n_1517, n_580, n_582);
  nand g1644 (n_592, n_1515, n_1516, n_1517);
  xor g1645 (n_1518, n_583, n_584);
  xor g1646 (n_83, n_1518, n_585);
  nand g1647 (n_1519, n_583, n_584);
  nand g1648 (n_1520, n_585, n_584);
  nand g1649 (n_1521, n_583, n_585);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1658 (n_590, n_1446, n_586);
  nand g1660 (n_1528, n_586, A[20]);
  nand g1662 (n_596, n_1156, n_1528, n_1529);
  xor g1663 (n_1530, n_548, n_588);
  xor g1664 (n_591, n_1530, n_589);
  nand g1665 (n_1531, n_548, n_588);
  nand g1666 (n_1532, n_589, n_588);
  nand g1667 (n_1533, n_548, n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_33, n_1535, n_1536, n_1537);
  xor g1678 (n_597, n_1466, A[22]);
  nand g1681 (n_1541, A[17], A[22]);
  nand g1682 (n_603, n_1233, n_1071, n_1541);
  xor g1684 (n_598, n_1542, n_596);
  nand g1686 (n_1544, n_596, n_560);
  nand g1688 (n_606, n_1543, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_81, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[18], A[22]);
  xor g1698 (n_604, n_1550, A[23]);
  nand g1701 (n_1553, A[18], A[23]);
  nand g1702 (n_609, n_1488, n_1115, n_1553);
  nand g1706 (n_1556, n_603, A[18]);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, n_604, n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, n_604, n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, n_604, n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1721 (n_1566, A[23], A[19]);
  xor g1722 (n_611, n_1566, n_405);
  nand g1723 (n_1567, A[23], A[19]);
  nand g1724 (n_1568, n_405, A[19]);
  nand g1725 (n_1569, A[23], n_405);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1727 (n_1570, n_609, n_610);
  xor g1728 (n_79, n_1570, n_611);
  nand g1729 (n_1571, n_609, n_610);
  nand g1730 (n_1572, n_611, n_610);
  nand g1731 (n_1573, n_609, n_611);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1739 (n_1578, n_423, n_424);
  xor g1740 (n_78, n_1578, n_614);
  nand g1742 (n_1580, n_614, n_424);
  nand g1743 (n_1581, n_423, n_614);
  nand g1744 (n_77, n_1204, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_442);
  nand g1752 (n_28, n_1583, n_1584, n_1585);
  nand g1759 (n_1589, A[23], A[21]);
  nand g1760 (n_27, n_1587, n_1588, n_1589);
  xor g1762 (n_75, n_1590, A[22]);
  nand g1766 (n_74, n_1591, n_1115, n_1593);
  nor g11 (n_1609, A[0], A[2]);
  nand g12 (n_1604, A[0], A[2]);
  nor g13 (n_1605, n_68, A[3]);
  nand g14 (n_1606, n_68, A[3]);
  nor g15 (n_1615, A[4], n_117);
  nand g16 (n_1610, A[4], n_117);
  nor g17 (n_1611, A[5], n_116);
  nand g18 (n_1612, A[5], n_116);
  nor g19 (n_1621, n_67, n_115);
  nand g20 (n_1616, n_67, n_115);
  nor g21 (n_1617, n_66, n_114);
  nand g22 (n_1618, n_66, n_114);
  nor g23 (n_1627, n_65, n_113);
  nand g24 (n_1622, n_65, n_113);
  nor g25 (n_1623, n_64, n_112);
  nand g26 (n_1624, n_64, n_112);
  nor g27 (n_1633, n_63, n_111);
  nand g28 (n_1628, n_63, n_111);
  nor g29 (n_1629, n_62, n_110);
  nand g30 (n_1630, n_62, n_110);
  nor g31 (n_1639, n_61, n_109);
  nand g32 (n_1634, n_61, n_109);
  nor g33 (n_1635, n_60, n_108);
  nand g34 (n_1636, n_60, n_108);
  nor g35 (n_1645, n_59, n_107);
  nand g36 (n_1640, n_59, n_107);
  nor g37 (n_1641, n_58, n_106);
  nand g38 (n_1642, n_58, n_106);
  nor g39 (n_1651, n_57, n_105);
  nand g40 (n_1646, n_57, n_105);
  nor g41 (n_1647, n_56, n_104);
  nand g42 (n_1648, n_56, n_104);
  nor g43 (n_1657, n_55, n_103);
  nand g44 (n_1652, n_55, n_103);
  nor g45 (n_1653, n_54, n_102);
  nand g46 (n_1654, n_54, n_102);
  nor g47 (n_1663, n_53, n_101);
  nand g48 (n_1658, n_53, n_101);
  nor g49 (n_1659, n_52, n_100);
  nand g50 (n_1660, n_52, n_100);
  nor g51 (n_1669, n_51, n_99);
  nand g52 (n_1664, n_51, n_99);
  nor g53 (n_1665, n_50, n_98);
  nand g54 (n_1666, n_50, n_98);
  nor g55 (n_1675, n_49, n_97);
  nand g56 (n_1670, n_49, n_97);
  nor g57 (n_1671, n_48, n_96);
  nand g58 (n_1672, n_48, n_96);
  nor g59 (n_1681, n_47, n_95);
  nand g60 (n_1676, n_47, n_95);
  nor g61 (n_1677, n_46, n_94);
  nand g62 (n_1678, n_46, n_94);
  nor g63 (n_1687, n_45, n_93);
  nand g64 (n_1682, n_45, n_93);
  nor g65 (n_1683, n_44, n_92);
  nand g66 (n_1684, n_44, n_92);
  nor g67 (n_1693, n_43, n_91);
  nand g68 (n_1688, n_43, n_91);
  nor g69 (n_1689, n_42, n_90);
  nand g70 (n_1690, n_42, n_90);
  nor g71 (n_1699, n_41, n_89);
  nand g72 (n_1694, n_41, n_89);
  nor g73 (n_1695, n_40, n_88);
  nand g74 (n_1696, n_40, n_88);
  nor g75 (n_1705, n_39, n_87);
  nand g76 (n_1700, n_39, n_87);
  nor g77 (n_1701, n_38, n_86);
  nand g78 (n_1702, n_38, n_86);
  nor g79 (n_1711, n_37, n_85);
  nand g80 (n_1706, n_37, n_85);
  nor g81 (n_1707, n_36, n_84);
  nand g82 (n_1708, n_36, n_84);
  nor g83 (n_1717, n_35, n_83);
  nand g84 (n_1712, n_35, n_83);
  nor g85 (n_1713, n_34, n_82);
  nand g86 (n_1714, n_34, n_82);
  nor g87 (n_1723, n_33, n_81);
  nand g88 (n_1718, n_33, n_81);
  nor g89 (n_1719, n_32, n_80);
  nand g90 (n_1720, n_32, n_80);
  nor g91 (n_1729, n_31, n_79);
  nand g92 (n_1724, n_31, n_79);
  nor g93 (n_1725, n_30, n_78);
  nand g94 (n_1726, n_30, n_78);
  nor g95 (n_1735, n_29, n_77);
  nand g96 (n_1730, n_29, n_77);
  nor g97 (n_1731, n_28, n_76);
  nand g98 (n_1732, n_28, n_76);
  nor g99 (n_1739, n_27, n_75);
  nand g100 (n_1736, n_27, n_75);
  nor g106 (n_1607, n_1604, n_1605);
  nor g110 (n_1613, n_1610, n_1611);
  nor g113 (n_1749, n_1615, n_1611);
  nor g114 (n_1619, n_1616, n_1617);
  nor g117 (n_1751, n_1621, n_1617);
  nor g118 (n_1625, n_1622, n_1623);
  nor g121 (n_1759, n_1627, n_1623);
  nor g122 (n_1631, n_1628, n_1629);
  nor g125 (n_1761, n_1633, n_1629);
  nor g126 (n_1637, n_1634, n_1635);
  nor g129 (n_1769, n_1639, n_1635);
  nor g130 (n_1643, n_1640, n_1641);
  nor g133 (n_1771, n_1645, n_1641);
  nor g134 (n_1649, n_1646, n_1647);
  nor g137 (n_1779, n_1651, n_1647);
  nor g138 (n_1655, n_1652, n_1653);
  nor g141 (n_1781, n_1657, n_1653);
  nor g142 (n_1661, n_1658, n_1659);
  nor g145 (n_1789, n_1663, n_1659);
  nor g146 (n_1667, n_1664, n_1665);
  nor g149 (n_1791, n_1669, n_1665);
  nor g150 (n_1673, n_1670, n_1671);
  nor g153 (n_1799, n_1675, n_1671);
  nor g154 (n_1679, n_1676, n_1677);
  nor g157 (n_1801, n_1681, n_1677);
  nor g158 (n_1685, n_1682, n_1683);
  nor g161 (n_1809, n_1687, n_1683);
  nor g162 (n_1691, n_1688, n_1689);
  nor g165 (n_1811, n_1693, n_1689);
  nor g166 (n_1697, n_1694, n_1695);
  nor g169 (n_1819, n_1699, n_1695);
  nor g170 (n_1703, n_1700, n_1701);
  nor g173 (n_1821, n_1705, n_1701);
  nor g174 (n_1709, n_1706, n_1707);
  nor g177 (n_1829, n_1711, n_1707);
  nor g178 (n_1715, n_1712, n_1713);
  nor g181 (n_1831, n_1717, n_1713);
  nor g182 (n_1721, n_1718, n_1719);
  nor g185 (n_1839, n_1723, n_1719);
  nor g186 (n_1727, n_1724, n_1725);
  nor g189 (n_1841, n_1729, n_1725);
  nor g190 (n_1733, n_1730, n_1731);
  nor g193 (n_1849, n_1735, n_1731);
  nor g203 (n_1747, n_1621, n_1746);
  nand g212 (n_1859, n_1749, n_1751);
  nor g213 (n_1757, n_1633, n_1756);
  nand g222 (n_1866, n_1759, n_1761);
  nor g223 (n_1767, n_1645, n_1766);
  nand g232 (n_1874, n_1769, n_1771);
  nor g233 (n_1777, n_1657, n_1776);
  nand g242 (n_1881, n_1779, n_1781);
  nor g243 (n_1787, n_1669, n_1786);
  nand g252 (n_1889, n_1789, n_1791);
  nor g253 (n_1797, n_1681, n_1796);
  nand g262 (n_1896, n_1799, n_1801);
  nor g263 (n_1807, n_1693, n_1806);
  nand g1776 (n_1904, n_1809, n_1811);
  nor g1777 (n_1817, n_1705, n_1816);
  nand g1786 (n_1911, n_1819, n_1821);
  nor g1787 (n_1827, n_1717, n_1826);
  nand g1796 (n_1919, n_1829, n_1831);
  nor g1797 (n_1837, n_1729, n_1836);
  nand g1806 (n_1926, n_1839, n_1841);
  nor g1807 (n_1847, n_1739, n_1846);
  nand g1814 (n_2130, n_1610, n_1853);
  nand g1816 (n_2132, n_1746, n_1854);
  nand g1819 (n_2135, n_1857, n_1858);
  nand g1822 (n_1934, n_1861, n_1862);
  nor g1823 (n_1864, n_1639, n_1863);
  nor g1826 (n_1944, n_1639, n_1866);
  nor g1832 (n_1872, n_1870, n_1863);
  nor g1835 (n_1950, n_1866, n_1870);
  nor g1836 (n_1876, n_1874, n_1863);
  nor g1839 (n_1953, n_1866, n_1874);
  nor g1840 (n_1879, n_1663, n_1878);
  nor g1843 (n_2033, n_1663, n_1881);
  nor g1849 (n_1887, n_1885, n_1878);
  nor g1852 (n_2039, n_1881, n_1885);
  nor g1853 (n_1891, n_1889, n_1878);
  nor g1856 (n_1959, n_1881, n_1889);
  nor g1857 (n_1894, n_1687, n_1893);
  nor g1860 (n_1972, n_1687, n_1896);
  nor g1866 (n_1902, n_1900, n_1893);
  nor g1869 (n_1982, n_1896, n_1900);
  nor g1870 (n_1906, n_1904, n_1893);
  nor g1873 (n_1987, n_1896, n_1904);
  nor g1874 (n_1909, n_1711, n_1908);
  nor g1877 (n_2085, n_1711, n_1911);
  nor g1883 (n_1917, n_1915, n_1908);
  nor g1886 (n_2091, n_1911, n_1915);
  nor g1887 (n_1921, n_1919, n_1908);
  nor g1890 (n_1995, n_1911, n_1919);
  nor g1891 (n_1924, n_1735, n_1923);
  nor g1894 (n_2008, n_1735, n_1926);
  nor g1900 (n_1932, n_1930, n_1923);
  nor g1903 (n_2018, n_1926, n_1930);
  nand g1906 (n_2139, n_1622, n_1936);
  nand g1907 (n_1937, n_1759, n_1934);
  nand g1908 (n_2141, n_1756, n_1937);
  nand g1911 (n_2144, n_1940, n_1941);
  nand g1914 (n_2147, n_1863, n_1943);
  nand g1915 (n_1946, n_1944, n_1934);
  nand g1916 (n_2150, n_1945, n_1946);
  nand g1917 (n_1949, n_1947, n_1934);
  nand g1918 (n_2152, n_1948, n_1949);
  nand g1919 (n_1952, n_1950, n_1934);
  nand g1920 (n_2155, n_1951, n_1952);
  nand g1921 (n_1955, n_1953, n_1934);
  nand g1922 (n_2023, n_1954, n_1955);
  nor g1923 (n_1957, n_1675, n_1956);
  nand g1932 (n_2047, n_1799, n_1959);
  nor g1933 (n_1966, n_1964, n_1956);
  nor g1938 (n_1969, n_1896, n_1956);
  nand g1947 (n_2059, n_1959, n_1972);
  nand g1952 (n_2063, n_1959, n_1977);
  nand g1957 (n_2067, n_1959, n_1982);
  nand g1962 (n_2071, n_1959, n_1987);
  nor g1963 (n_1993, n_1723, n_1992);
  nand g1972 (n_2099, n_1839, n_1995);
  nor g1973 (n_2002, n_2000, n_1992);
  nor g1978 (n_2005, n_1926, n_1992);
  nand g1987 (n_2111, n_1995, n_2008);
  nand g1992 (n_2115, n_1995, n_2013);
  nand g1997 (n_2119, n_1995, n_2018);
  nand g2000 (n_2159, n_1646, n_2025);
  nand g2001 (n_2026, n_1779, n_2023);
  nand g2002 (n_2161, n_1776, n_2026);
  nand g2005 (n_2164, n_2029, n_2030);
  nand g2008 (n_2167, n_1878, n_2032);
  nand g2009 (n_2035, n_2033, n_2023);
  nand g2010 (n_2170, n_2034, n_2035);
  nand g2011 (n_2038, n_2036, n_2023);
  nand g2012 (n_2172, n_2037, n_2038);
  nand g2013 (n_2041, n_2039, n_2023);
  nand g2014 (n_2175, n_2040, n_2041);
  nand g2015 (n_2042, n_1959, n_2023);
  nand g2016 (n_2177, n_1956, n_2042);
  nand g2019 (n_2180, n_2045, n_2046);
  nand g2022 (n_2182, n_2049, n_2050);
  nand g2025 (n_2185, n_2053, n_2054);
  nand g2028 (n_2188, n_2057, n_2058);
  nand g2031 (n_2191, n_2061, n_2062);
  nand g2034 (n_2193, n_2065, n_2066);
  nand g2037 (n_2196, n_2069, n_2070);
  nand g2040 (n_2075, n_2073, n_2074);
  nand g2043 (n_2200, n_1694, n_2077);
  nand g2044 (n_2078, n_1819, n_2075);
  nand g2045 (n_2202, n_1816, n_2078);
  nand g2048 (n_2205, n_2081, n_2082);
  nand g2051 (n_2208, n_1908, n_2084);
  nand g2052 (n_2087, n_2085, n_2075);
  nand g2053 (n_2211, n_2086, n_2087);
  nand g2054 (n_2090, n_2088, n_2075);
  nand g2055 (n_2213, n_2089, n_2090);
  nand g2056 (n_2093, n_2091, n_2075);
  nand g2057 (n_2216, n_2092, n_2093);
  nand g2058 (n_2094, n_1995, n_2075);
  nand g2059 (n_2218, n_1992, n_2094);
  nand g2062 (n_2221, n_2097, n_2098);
  nand g2065 (n_2223, n_2101, n_2102);
  nand g2068 (n_2226, n_2105, n_2106);
  nand g2071 (n_2229, n_2109, n_2110);
  nand g2074 (n_2232, n_2113, n_2114);
  nand g2077 (n_2234, n_2117, n_2118);
  nand g2080 (n_2237, n_2121, n_2122);
  xnor g2092 (Z[5], n_2130, n_2131);
  xnor g2094 (Z[6], n_2132, n_2133);
  xnor g2097 (Z[7], n_2135, n_2136);
  xnor g2099 (Z[8], n_1934, n_2137);
  xnor g2102 (Z[9], n_2139, n_2140);
  xnor g2104 (Z[10], n_2141, n_2142);
  xnor g2107 (Z[11], n_2144, n_2145);
  xnor g2110 (Z[12], n_2147, n_2148);
  xnor g2113 (Z[13], n_2150, n_2151);
  xnor g2115 (Z[14], n_2152, n_2153);
  xnor g2118 (Z[15], n_2155, n_2156);
  xnor g2120 (Z[16], n_2023, n_2157);
  xnor g2123 (Z[17], n_2159, n_2160);
  xnor g2125 (Z[18], n_2161, n_2162);
  xnor g2128 (Z[19], n_2164, n_2165);
  xnor g2131 (Z[20], n_2167, n_2168);
  xnor g2134 (Z[21], n_2170, n_2171);
  xnor g2136 (Z[22], n_2172, n_2173);
  xnor g2139 (Z[23], n_2175, n_2176);
  xnor g2141 (Z[24], n_2177, n_2178);
  xnor g2144 (Z[25], n_2180, n_2181);
  xnor g2146 (Z[26], n_2182, n_2183);
  xnor g2149 (Z[27], n_2185, n_2186);
  xnor g2152 (Z[28], n_2188, n_2189);
  xnor g2155 (Z[29], n_2191, n_2192);
  xnor g2157 (Z[30], n_2193, n_2194);
  xnor g2160 (Z[31], n_2196, n_2197);
  xnor g2162 (Z[32], n_2075, n_2198);
  xnor g2165 (Z[33], n_2200, n_2201);
  xnor g2167 (Z[34], n_2202, n_2203);
  xnor g2170 (Z[35], n_2205, n_2206);
  xnor g2173 (Z[36], n_2208, n_2209);
  xnor g2176 (Z[37], n_2211, n_2212);
  xnor g2178 (Z[38], n_2213, n_2214);
  xnor g2181 (Z[39], n_2216, n_2217);
  xnor g2183 (Z[40], n_2218, n_2219);
  xnor g2186 (Z[41], n_2221, n_2222);
  xnor g2188 (Z[42], n_2223, n_2224);
  xnor g2191 (Z[43], n_2226, n_2227);
  xnor g2194 (Z[44], n_2229, n_2230);
  xnor g2197 (Z[45], n_2232, n_2233);
  xnor g2199 (Z[46], n_2234, n_2235);
  xnor g2202 (Z[47], n_2237, n_2238);
  or g2214 (n_1044, A[1], wc);
  not gc (wc, n_171);
  or g2215 (n_1045, A[1], wc0);
  not gc0 (wc0, A[2]);
  or g2216 (n_1069, wc1, A[24]);
  not gc1 (wc1, A[18]);
  or g2217 (n_1088, A[2], wc2);
  not gc2 (wc2, A[3]);
  or g2218 (n_1089, wc3, A[2]);
  not gc3 (wc3, A[1]);
  xnor g2219 (n_1154, A[24], A[19]);
  or g2220 (n_1155, wc4, A[24]);
  not gc4 (wc4, A[19]);
  or g2221 (n_1156, wc5, A[24]);
  not gc5 (wc5, A[20]);
  xnor g2222 (n_1194, A[24], A[21]);
  or g2223 (n_1195, wc6, A[24]);
  not gc6 (wc6, A[21]);
  xnor g2224 (n_1214, A[6], A[5]);
  or g2225 (n_1215, A[5], wc7);
  not gc7 (wc7, A[6]);
  or g2226 (n_1252, wc8, A[6]);
  not gc8 (wc8, A[5]);
  or g2227 (n_1253, A[6], wc9);
  not gc9 (wc9, A[7]);
  or g2229 (n_1355, wc10, A[10]);
  not gc10 (wc10, A[9]);
  or g2230 (n_1356, A[10], wc11);
  not gc11 (wc11, A[14]);
  or g2231 (n_1385, A[10], wc12);
  not gc12 (wc12, A[11]);
  xnor g2232 (n_1446, A[24], A[20]);
  xnor g2233 (n_1462, A[14], A[13]);
  or g2234 (n_1463, wc13, A[14]);
  not gc13 (wc13, A[13]);
  or g2235 (n_1464, A[14], wc14);
  not gc14 (wc14, A[18]);
  or g2236 (n_1485, A[14], wc15);
  not gc15 (wc15, A[15]);
  or g2238 (n_1555, wc16, A[19]);
  not gc16 (wc16, A[18]);
  or g2240 (n_1583, A[21], wc17);
  not gc17 (wc17, A[22]);
  or g2242 (n_1587, A[22], wc18);
  not gc18 (wc18, A[23]);
  or g2243 (n_1588, wc19, A[22]);
  not gc19 (wc19, A[21]);
  xnor g2244 (n_1590, A[24], A[23]);
  or g2245 (n_1591, wc20, A[24]);
  not gc20 (wc20, A[23]);
  or g2246 (n_1593, wc21, A[24]);
  not gc21 (wc21, A[22]);
  xnor g2247 (n_349, n_1042, A[1]);
  xnor g2248 (n_372, n_1086, A[2]);
  xnor g2249 (n_453, n_1250, A[6]);
  xnor g2250 (n_504, n_1218, A[14]);
  xnor g2251 (n_520, n_1254, A[10]);
  nand g2252 (n_532, n_1255, n_1385);
  or g2253 (n_1421, A[24], wc22);
  not gc22 (wc22, n_533);
  xnor g2254 (n_569, n_1386, A[14]);
  nand g2255 (n_578, n_1104, n_1485);
  xnor g2256 (n_1542, n_560, A[18]);
  or g2257 (n_1543, A[18], wc23);
  not gc23 (wc23, n_560);
  xnor g2258 (n_605, n_1266, n_603);
  or g2259 (n_1557, A[19], wc24);
  not gc24 (wc24, n_603);
  xnor g2260 (n_76, n_1114, A[21]);
  or g2262 (n_2124, wc25, n_1609);
  not gc25 (wc25, n_1604);
  xnor g2263 (n_537, n_1418, A[24]);
  or g2264 (n_1508, A[24], wc26);
  not gc26 (wc26, n_578);
  or g2265 (n_1529, A[24], wc27);
  not gc27 (wc27, n_586);
  xnor g2266 (n_29, n_1070, n_442);
  or g2267 (n_1584, A[21], wc28);
  not gc28 (wc28, n_442);
  and g2268 (n_1744, wc29, n_1606);
  not gc29 (wc29, n_1607);
  or g2269 (n_2127, wc30, n_1605);
  not gc30 (wc30, n_1606);
  or g2270 (n_1449, A[24], wc31);
  not gc31 (wc31, n_545);
  xnor g2271 (n_581, n_1506, A[24]);
  and g2272 (n_1737, wc32, n_74);
  not gc32 (wc32, A[24]);
  or g2273 (n_1738, wc33, n_74);
  not gc33 (wc33, A[24]);
  not g2274 (Z[2], n_2124);
  or g2275 (n_1216, A[5], wc34);
  not gc34 (wc34, n_433);
  or g2276 (n_1545, A[18], wc35);
  not gc35 (wc35, n_596);
  or g2279 (n_2128, wc36, n_1615);
  not gc36 (wc36, n_1610);
  or g2280 (n_2235, wc37, n_1739);
  not gc37 (wc37, n_1736);
  and g2281 (n_1746, wc38, n_1612);
  not gc38 (wc38, n_1613);
  or g2282 (n_1853, n_1615, n_1744);
  or g2283 (n_1854, n_1744, wc39);
  not gc39 (wc39, n_1749);
  xor g2284 (Z[3], n_1604, n_2127);
  xor g2285 (Z[4], n_1744, n_2128);
  or g2286 (n_2131, wc40, n_1611);
  not gc40 (wc40, n_1612);
  or g2287 (n_2238, wc41, n_1737);
  not gc41 (wc41, n_1738);
  xnor g2288 (n_1334, n_489, A[24]);
  or g2289 (n_1335, A[24], wc42);
  not gc42 (wc42, n_489);
  and g2290 (n_1753, wc43, n_1618);
  not gc43 (wc43, n_1619);
  or g2291 (n_1855, wc44, n_1621);
  not gc44 (wc44, n_1749);
  or g2292 (n_2133, wc45, n_1621);
  not gc45 (wc45, n_1616);
  or g2293 (n_2136, wc46, n_1617);
  not gc46 (wc46, n_1618);
  or g2294 (n_2233, wc47, n_1731);
  not gc47 (wc47, n_1732);
  and g2295 (n_1857, wc48, n_1616);
  not gc48 (wc48, n_1747);
  and g2296 (n_1754, wc49, n_1751);
  not gc49 (wc49, n_1746);
  or g2297 (n_2137, wc50, n_1627);
  not gc50 (wc50, n_1622);
  or g2298 (n_2227, wc51, n_1725);
  not gc51 (wc51, n_1726);
  xnor g2299 (n_1302, n_474, A[24]);
  or g2300 (n_1303, A[24], wc52);
  not gc52 (wc52, n_474);
  and g2301 (n_1846, wc53, n_1732);
  not gc53 (wc53, n_1733);
  and g2302 (n_1861, wc54, n_1753);
  not gc54 (wc54, n_1754);
  or g2303 (n_1930, wc55, n_1739);
  not gc55 (wc55, n_1849);
  or g2304 (n_1858, n_1744, n_1855);
  or g2305 (n_1862, n_1859, n_1744);
  or g2306 (n_2230, wc56, n_1735);
  not gc56 (wc56, n_1730);
  or g2307 (n_1068, A[24], wc57);
  not gc57 (wc57, n_357);
  and g2308 (n_1756, wc58, n_1624);
  not gc58 (wc58, n_1625);
  or g2309 (n_2140, wc59, n_1623);
  not gc59 (wc59, n_1624);
  xnor g2310 (n_363, n_1066, A[24]);
  and g2311 (n_1836, wc60, n_1720);
  not gc60 (wc60, n_1721);
  and g2312 (n_1843, wc61, n_1726);
  not gc61 (wc61, n_1727);
  or g2313 (n_1938, wc62, n_1633);
  not gc62 (wc62, n_1759);
  or g2314 (n_2000, wc63, n_1729);
  not gc63 (wc63, n_1839);
  and g2315 (n_1931, wc64, n_1736);
  not gc64 (wc64, n_1847);
  or g2316 (n_1936, wc65, n_1627);
  not gc65 (wc65, n_1934);
  or g2317 (n_2142, wc66, n_1633);
  not gc66 (wc66, n_1628);
  or g2318 (n_2219, wc67, n_1723);
  not gc67 (wc67, n_1718);
  or g2319 (n_2222, wc68, n_1719);
  not gc68 (wc68, n_1720);
  or g2320 (n_2224, wc69, n_1729);
  not gc69 (wc69, n_1724);
  and g2321 (n_1763, wc70, n_1630);
  not gc70 (wc70, n_1631);
  and g2322 (n_1940, wc71, n_1628);
  not gc71 (wc71, n_1757);
  and g2323 (n_1844, wc72, n_1841);
  not gc72 (wc72, n_1836);
  and g2324 (n_2013, wc73, n_1849);
  not gc73 (wc73, n_1926);
  or g2325 (n_2145, wc74, n_1629);
  not gc74 (wc74, n_1630);
  and g2326 (n_1826, wc75, n_1708);
  not gc75 (wc75, n_1709);
  and g2327 (n_1833, wc76, n_1714);
  not gc76 (wc76, n_1715);
  and g2328 (n_1764, wc77, n_1761);
  not gc77 (wc77, n_1756);
  or g2329 (n_1915, wc78, n_1717);
  not gc78 (wc78, n_1829);
  and g2330 (n_2001, wc79, n_1724);
  not gc79 (wc79, n_1837);
  and g2331 (n_1923, wc80, n_1843);
  not gc80 (wc80, n_1844);
  or g2332 (n_1941, n_1938, wc81);
  not gc81 (wc81, n_1934);
  or g2333 (n_2148, wc82, n_1639);
  not gc82 (wc82, n_1634);
  or g2334 (n_2209, wc83, n_1711);
  not gc83 (wc83, n_1706);
  or g2335 (n_2212, wc84, n_1707);
  not gc84 (wc84, n_1708);
  or g2336 (n_2214, wc85, n_1717);
  not gc85 (wc85, n_1712);
  or g2337 (n_2217, wc86, n_1713);
  not gc86 (wc86, n_1714);
  and g2338 (n_1863, wc87, n_1763);
  not gc87 (wc87, n_1764);
  and g2339 (n_1834, wc88, n_1831);
  not gc88 (wc88, n_1826);
  and g2340 (n_1928, wc89, n_1849);
  not gc89 (wc89, n_1923);
  or g2341 (n_1943, wc90, n_1866);
  not gc90 (wc90, n_1934);
  or g2342 (n_2156, wc91, n_1641);
  not gc91 (wc91, n_1642);
  and g2343 (n_1766, wc92, n_1636);
  not gc92 (wc92, n_1637);
  and g2344 (n_1773, wc93, n_1642);
  not gc93 (wc93, n_1643);
  or g2345 (n_1870, wc94, n_1645);
  not gc94 (wc94, n_1769);
  and g2346 (n_1916, wc95, n_1712);
  not gc95 (wc95, n_1827);
  and g2347 (n_1920, wc96, n_1833);
  not gc96 (wc96, n_1834);
  and g2348 (n_2010, wc97, n_1730);
  not gc97 (wc97, n_1924);
  and g2349 (n_2015, wc98, n_1846);
  not gc98 (wc98, n_1928);
  and g2350 (n_2020, n_1931, wc99);
  not gc99 (wc99, n_1932);
  or g2351 (n_2151, wc100, n_1635);
  not gc100 (wc100, n_1636);
  or g2352 (n_2153, wc101, n_1645);
  not gc101 (wc101, n_1640);
  and g2353 (n_1774, wc102, n_1771);
  not gc102 (wc102, n_1766);
  and g2354 (n_1945, wc103, n_1634);
  not gc103 (wc103, n_1864);
  and g2355 (n_1868, wc104, n_1769);
  not gc104 (wc104, n_1863);
  and g2356 (n_1947, wc105, n_1769);
  not gc105 (wc105, n_1866);
  or g2357 (n_2157, wc106, n_1651);
  not gc106 (wc106, n_1646);
  or g2358 (n_2203, wc107, n_1705);
  not gc107 (wc107, n_1700);
  and g2359 (n_1776, wc108, n_1648);
  not gc108 (wc108, n_1649);
  and g2360 (n_1823, wc109, n_1702);
  not gc109 (wc109, n_1703);
  and g2361 (n_1871, wc110, n_1640);
  not gc110 (wc110, n_1767);
  and g2362 (n_1875, wc111, n_1773);
  not gc111 (wc111, n_1774);
  and g2363 (n_1948, wc112, n_1766);
  not gc112 (wc112, n_1868);
  or g2364 (n_2160, wc113, n_1647);
  not gc113 (wc113, n_1648);
  or g2365 (n_2206, wc114, n_1701);
  not gc114 (wc114, n_1702);
  or g2366 (n_2027, wc115, n_1657);
  not gc115 (wc115, n_1779);
  or g2367 (n_2162, wc116, n_1657);
  not gc116 (wc116, n_1652);
  or g2368 (n_2171, wc117, n_1659);
  not gc117 (wc117, n_1660);
  or g2369 (n_2173, wc118, n_1669);
  not gc118 (wc118, n_1664);
  and g2370 (n_1783, wc119, n_1654);
  not gc119 (wc119, n_1655);
  and g2371 (n_1786, wc120, n_1660);
  not gc120 (wc120, n_1661);
  and g2372 (n_1793, wc121, n_1666);
  not gc121 (wc121, n_1667);
  and g2373 (n_1813, wc122, n_1690);
  not gc122 (wc122, n_1691);
  and g2374 (n_2029, wc123, n_1652);
  not gc123 (wc123, n_1777);
  or g2375 (n_1885, wc124, n_1669);
  not gc124 (wc124, n_1789);
  and g2376 (n_1951, n_1871, wc125);
  not gc125 (wc125, n_1872);
  and g2377 (n_1954, n_1875, wc126);
  not gc126 (wc126, n_1876);
  or g2378 (n_2165, wc127, n_1653);
  not gc127 (wc127, n_1654);
  or g2379 (n_2168, wc128, n_1663);
  not gc128 (wc128, n_1658);
  or g2380 (n_2176, wc129, n_1665);
  not gc129 (wc129, n_1666);
  or g2381 (n_2178, wc130, n_1675);
  not gc130 (wc130, n_1670);
  or g2382 (n_2194, wc131, n_1693);
  not gc131 (wc131, n_1688);
  or g2383 (n_2197, wc132, n_1689);
  not gc132 (wc132, n_1690);
  or g2384 (n_2198, wc133, n_1699);
  not gc133 (wc133, n_1694);
  and g2385 (n_1796, wc134, n_1672);
  not gc134 (wc134, n_1673);
  and g2386 (n_1803, wc135, n_1678);
  not gc135 (wc135, n_1679);
  and g2387 (n_1816, wc136, n_1696);
  not gc136 (wc136, n_1697);
  and g2388 (n_1784, wc137, n_1781);
  not gc137 (wc137, n_1776);
  and g2389 (n_1794, wc138, n_1791);
  not gc138 (wc138, n_1786);
  or g2390 (n_1964, wc139, n_1681);
  not gc139 (wc139, n_1799);
  or g2391 (n_2079, wc140, n_1705);
  not gc140 (wc140, n_1819);
  and g2392 (n_2036, wc141, n_1789);
  not gc141 (wc141, n_1881);
  or g2393 (n_2181, wc142, n_1671);
  not gc142 (wc142, n_1672);
  or g2394 (n_2183, wc143, n_1681);
  not gc143 (wc143, n_1676);
  or g2395 (n_2186, wc144, n_1677);
  not gc144 (wc144, n_1678);
  or g2396 (n_2189, wc145, n_1687);
  not gc145 (wc145, n_1682);
  or g2397 (n_2201, wc146, n_1695);
  not gc146 (wc146, n_1696);
  and g2398 (n_1806, wc147, n_1684);
  not gc147 (wc147, n_1685);
  and g2399 (n_1878, wc148, n_1783);
  not gc148 (wc148, n_1784);
  and g2400 (n_1886, wc149, n_1664);
  not gc149 (wc149, n_1787);
  and g2401 (n_1890, wc150, n_1793);
  not gc150 (wc150, n_1794);
  and g2402 (n_1804, wc151, n_1801);
  not gc151 (wc151, n_1796);
  or g2403 (n_1900, wc152, n_1693);
  not gc152 (wc152, n_1809);
  and g2404 (n_1824, wc153, n_1821);
  not gc153 (wc153, n_1816);
  and g2405 (n_2088, wc154, n_1829);
  not gc154 (wc154, n_1911);
  or g2406 (n_2043, wc155, n_1675);
  not gc155 (wc155, n_1959);
  or g2407 (n_2025, wc156, n_1651);
  not gc156 (wc156, n_2023);
  or g2408 (n_2030, n_2027, wc157);
  not gc157 (wc157, n_2023);
  or g2409 (n_2032, wc158, n_1881);
  not gc158 (wc158, n_2023);
  or g2410 (n_2192, wc159, n_1683);
  not gc159 (wc159, n_1684);
  and g2411 (n_1965, wc160, n_1676);
  not gc160 (wc160, n_1797);
  and g2412 (n_1893, wc161, n_1803);
  not gc161 (wc161, n_1804);
  and g2413 (n_1814, wc162, n_1811);
  not gc162 (wc162, n_1806);
  and g2414 (n_2081, wc163, n_1700);
  not gc163 (wc163, n_1817);
  and g2415 (n_1908, wc164, n_1823);
  not gc164 (wc164, n_1824);
  and g2416 (n_1883, wc165, n_1789);
  not gc165 (wc165, n_1878);
  and g2417 (n_1977, wc166, n_1809);
  not gc166 (wc166, n_1896);
  or g2418 (n_2051, n_1964, wc167);
  not gc167 (wc167, n_1959);
  or g2419 (n_2055, wc168, n_1896);
  not gc168 (wc168, n_1959);
  or g2420 (n_2095, wc169, n_1723);
  not gc169 (wc169, n_1995);
  or g2421 (n_2103, n_2000, wc170);
  not gc170 (wc170, n_1995);
  or g2422 (n_2107, wc171, n_1926);
  not gc171 (wc171, n_1995);
  and g2423 (n_1901, wc172, n_1688);
  not gc172 (wc172, n_1807);
  and g2424 (n_1905, wc173, n_1813);
  not gc173 (wc173, n_1814);
  and g2425 (n_2034, wc174, n_1658);
  not gc174 (wc174, n_1879);
  and g2426 (n_2037, wc175, n_1786);
  not gc175 (wc175, n_1883);
  and g2427 (n_2040, n_1886, wc176);
  not gc176 (wc176, n_1887);
  and g2428 (n_1956, n_1890, wc177);
  not gc177 (wc177, n_1891);
  and g2429 (n_1898, wc178, n_1809);
  not gc178 (wc178, n_1893);
  and g2430 (n_1913, wc179, n_1829);
  not gc179 (wc179, n_1908);
  or g2431 (n_2046, n_2043, wc180);
  not gc180 (wc180, n_2023);
  or g2432 (n_2050, n_2047, wc181);
  not gc181 (wc181, n_2023);
  and g2433 (n_1974, wc182, n_1682);
  not gc182 (wc182, n_1894);
  and g2434 (n_1979, wc183, n_1806);
  not gc183 (wc183, n_1898);
  and g2435 (n_2086, wc184, n_1706);
  not gc184 (wc184, n_1909);
  and g2436 (n_2089, wc185, n_1826);
  not gc185 (wc185, n_1913);
  and g2437 (n_2092, n_1916, wc186);
  not gc186 (wc186, n_1917);
  and g2438 (n_1992, n_1920, wc187);
  not gc187 (wc187, n_1921);
  and g2439 (n_1962, wc188, n_1799);
  not gc188 (wc188, n_1956);
  and g2440 (n_1975, wc189, n_1972);
  not gc189 (wc189, n_1956);
  and g2441 (n_1980, wc190, n_1977);
  not gc190 (wc190, n_1956);
  and g2442 (n_1985, wc191, n_1982);
  not gc191 (wc191, n_1956);
  and g2443 (n_1990, wc192, n_1987);
  not gc192 (wc192, n_1956);
  or g2444 (n_2054, n_2051, wc193);
  not gc193 (wc193, n_2023);
  or g2445 (n_2058, n_2055, wc194);
  not gc194 (wc194, n_2023);
  or g2446 (n_2062, n_2059, wc195);
  not gc195 (wc195, n_2023);
  and g2447 (n_1984, n_1901, wc196);
  not gc196 (wc196, n_1902);
  and g2448 (n_1989, n_1905, wc197);
  not gc197 (wc197, n_1906);
  and g2449 (n_2045, wc198, n_1670);
  not gc198 (wc198, n_1957);
  and g2450 (n_2049, wc199, n_1796);
  not gc199 (wc199, n_1962);
  and g2451 (n_2053, n_1965, wc200);
  not gc200 (wc200, n_1966);
  and g2452 (n_2057, n_1893, wc201);
  not gc201 (wc201, n_1969);
  and g2453 (n_1998, wc202, n_1839);
  not gc202 (wc202, n_1992);
  and g2454 (n_2011, wc203, n_2008);
  not gc203 (wc203, n_1992);
  and g2455 (n_2016, wc204, n_2013);
  not gc204 (wc204, n_1992);
  and g2456 (n_2021, wc205, n_2018);
  not gc205 (wc205, n_1992);
  or g2457 (n_2066, n_2063, wc206);
  not gc206 (wc206, n_2023);
  or g2458 (n_2070, n_2067, wc207);
  not gc207 (wc207, n_2023);
  or g2459 (n_2074, n_2071, wc208);
  not gc208 (wc208, n_2023);
  and g2460 (n_2061, wc209, n_1974);
  not gc209 (wc209, n_1975);
  and g2461 (n_2065, wc210, n_1979);
  not gc210 (wc210, n_1980);
  and g2462 (n_2097, wc211, n_1718);
  not gc211 (wc211, n_1993);
  and g2463 (n_2101, wc212, n_1836);
  not gc212 (wc212, n_1998);
  and g2464 (n_2105, n_2001, wc213);
  not gc213 (wc213, n_2002);
  and g2465 (n_2109, n_1923, wc214);
  not gc214 (wc214, n_2005);
  and g2466 (n_2113, wc215, n_2010);
  not gc215 (wc215, n_2011);
  and g2467 (n_2117, wc216, n_2015);
  not gc216 (wc216, n_2016);
  and g2468 (n_2121, wc217, n_2020);
  not gc217 (wc217, n_2021);
  and g2469 (n_2069, n_1984, wc218);
  not gc218 (wc218, n_1985);
  and g2470 (n_2073, n_1989, wc219);
  not gc219 (wc219, n_1990);
  or g2471 (n_2077, wc220, n_1699);
  not gc220 (wc220, n_2075);
  or g2472 (n_2082, n_2079, wc221);
  not gc221 (wc221, n_2075);
  or g2473 (n_2084, wc222, n_1911);
  not gc222 (wc222, n_2075);
  or g2474 (n_2098, n_2095, wc223);
  not gc223 (wc223, n_2075);
  or g2475 (n_2102, wc224, n_2099);
  not gc224 (wc224, n_2075);
  or g2476 (n_2106, n_2103, wc225);
  not gc225 (wc225, n_2075);
  or g2477 (n_2110, n_2107, wc226);
  not gc226 (wc226, n_2075);
  or g2478 (n_2114, wc227, n_2111);
  not gc227 (wc227, n_2075);
  or g2479 (n_2118, wc228, n_2115);
  not gc228 (wc228, n_2075);
  or g2480 (n_2122, wc229, n_2119);
  not gc229 (wc229, n_2075);
endmodule

module mult_signed_const_5219_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_5219_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_5486_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_171, n_172, n_173, n_176, n_179;
  wire n_180, n_183, n_184, n_187, n_188, n_189, n_193, n_195;
  wire n_196, n_201, n_202, n_203, n_204, n_208, n_209, n_210;
  wire n_211, n_212, n_215, n_217, n_218, n_219, n_220, n_221;
  wire n_223, n_224, n_225, n_226, n_227, n_228, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_245, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_257, n_259, n_260;
  wire n_261, n_262, n_263, n_269, n_270, n_272, n_273, n_274;
  wire n_275, n_276, n_277, n_278, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_300, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_315, n_317, n_318, n_319, n_320, n_321, n_322, n_323;
  wire n_324, n_325, n_326, n_327, n_333, n_334, n_336, n_337;
  wire n_338, n_339, n_340, n_341, n_342, n_343, n_344, n_345;
  wire n_346, n_350, n_352, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_372, n_373, n_374, n_375, n_377, n_378, n_379, n_380;
  wire n_381, n_382, n_383, n_384, n_385, n_386, n_387, n_388;
  wire n_389, n_390, n_391, n_393, n_394, n_395, n_396, n_397;
  wire n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405;
  wire n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413;
  wire n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421;
  wire n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429;
  wire n_430, n_431, n_434, n_435, n_436, n_437, n_438, n_439;
  wire n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447;
  wire n_448, n_449, n_450, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_471, n_472, n_473, n_474, n_475;
  wire n_476, n_477, n_479, n_480, n_481, n_482, n_483, n_484;
  wire n_485, n_486, n_487, n_488, n_489, n_491, n_492, n_493;
  wire n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_521, n_522, n_523, n_524;
  wire n_525, n_526, n_527, n_528, n_529, n_530, n_531, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_546, n_547, n_548, n_549, n_550, n_551;
  wire n_552, n_553, n_554, n_555, n_558, n_559, n_561, n_562;
  wire n_563, n_564, n_565, n_566, n_571, n_572, n_573, n_574;
  wire n_575, n_576, n_577, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_590, n_591, n_592, n_593, n_596;
  wire n_597, n_598, n_599, n_600, n_604, n_606, n_607, n_609;
  wire n_611, n_612, n_613, n_614, n_615, n_618, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_642, n_647, n_648, n_649, n_650, n_651, n_652;
  wire n_653, n_654, n_659, n_660, n_661, n_662, n_663, n_664;
  wire n_665, n_666, n_669, n_670, n_671, n_672, n_673, n_674;
  wire n_675, n_676, n_677, n_678, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_691, n_692, n_693, n_694, n_703, n_704;
  wire n_705, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_714, n_719, n_723, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_734, n_737, n_738;
  wire n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746;
  wire n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_754;
  wire n_765, n_766, n_767, n_768, n_769, n_770, n_771, n_772;
  wire n_773, n_774, n_775, n_776, n_777, n_778, n_787, n_788;
  wire n_789, n_791, n_792, n_793, n_794, n_795, n_796, n_797;
  wire n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805;
  wire n_806, n_815, n_819, n_820, n_821, n_822, n_823, n_824;
  wire n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832;
  wire n_833, n_834, n_841, n_842, n_843, n_844, n_845, n_846;
  wire n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854;
  wire n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862;
  wire n_875, n_876, n_877, n_878, n_879, n_880, n_881, n_882;
  wire n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890;
  wire n_891, n_892, n_893, n_894, n_907, n_910, n_911, n_912;
  wire n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920;
  wire n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928;
  wire n_929, n_930, n_939, n_945, n_946, n_947, n_948, n_949;
  wire n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957;
  wire n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965;
  wire n_966, n_974, n_975, n_976, n_977, n_978, n_979, n_980;
  wire n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988;
  wire n_989, n_990, n_991, n_992, n_993, n_994, n_995, n_996;
  wire n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1017, n_1018;
  wire n_1019, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027;
  wire n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035;
  wire n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043;
  wire n_1045, n_1046, n_1047, n_1048, n_1049, n_1055, n_1056, n_1058;
  wire n_1059, n_1060, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067;
  wire n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075;
  wire n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083;
  wire n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091;
  wire n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099;
  wire n_1100, n_1101, n_1103, n_1104, n_1106, n_1107, n_1108, n_1109;
  wire n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117;
  wire n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125;
  wire n_1126, n_1127, n_1128, n_1129, n_1130, n_1133, n_1134, n_1135;
  wire n_1136, n_1137, n_1138, n_1139, n_1141, n_1143, n_1144, n_1145;
  wire n_1146, n_1147, n_1148, n_1150, n_1151, n_1152, n_1153, n_1154;
  wire n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162;
  wire n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170;
  wire n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178;
  wire n_1179, n_1180, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188;
  wire n_1191, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199;
  wire n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207;
  wire n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215;
  wire n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223;
  wire n_1224, n_1226, n_1227, n_1228, n_1229, n_1231, n_1232, n_1233;
  wire n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241;
  wire n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249;
  wire n_1250, n_1251, n_1253, n_1254, n_1258, n_1259, n_1261, n_1262;
  wire n_1263, n_1264, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271;
  wire n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279;
  wire n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1289;
  wire n_1291, n_1299, n_1300, n_1302, n_1303, n_1304, n_1305, n_1306;
  wire n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314;
  wire n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322;
  wire n_1323, n_1327, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335;
  wire n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343;
  wire n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351;
  wire n_1352, n_1353, n_1354, n_1355, n_1359, n_1360, n_1361, n_1363;
  wire n_1364, n_1365, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372;
  wire n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380;
  wire n_1381, n_1382, n_1383, n_1387, n_1388, n_1389, n_1391, n_1392;
  wire n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401;
  wire n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409;
  wire n_1410, n_1416, n_1417, n_1419, n_1422, n_1423, n_1424, n_1425;
  wire n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433;
  wire n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1442, n_1446;
  wire n_1447, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455;
  wire n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1467;
  wire n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476;
  wire n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1487, n_1488;
  wire n_1489, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497;
  wire n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1506;
  wire n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518;
  wire n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1527, n_1529;
  wire n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537;
  wire n_1538, n_1539, n_1540, n_1542, n_1543, n_1544, n_1545, n_1546;
  wire n_1547, n_1548, n_1549, n_1550, n_1556, n_1557, n_1558, n_1559;
  wire n_1560, n_1561, n_1562, n_1563, n_1564, n_1567, n_1568, n_1569;
  wire n_1570, n_1571, n_1572, n_1573, n_1574, n_1579, n_1580, n_1581;
  wire n_1582, n_1584, n_1585, n_1586, n_1588, n_1589, n_1590, n_1605;
  wire n_1606, n_1607, n_1608, n_1610, n_1611, n_1612, n_1613, n_1614;
  wire n_1616, n_1617, n_1618, n_1619, n_1620, n_1622, n_1623, n_1624;
  wire n_1625, n_1626, n_1628, n_1629, n_1630, n_1631, n_1632, n_1634;
  wire n_1635, n_1636, n_1637, n_1638, n_1640, n_1641, n_1642, n_1643;
  wire n_1644, n_1646, n_1647, n_1648, n_1649, n_1650, n_1652, n_1653;
  wire n_1654, n_1655, n_1656, n_1658, n_1659, n_1660, n_1661, n_1662;
  wire n_1664, n_1665, n_1666, n_1667, n_1668, n_1670, n_1671, n_1672;
  wire n_1673, n_1674, n_1676, n_1677, n_1678, n_1679, n_1680, n_1682;
  wire n_1683, n_1684, n_1685, n_1686, n_1688, n_1689, n_1690, n_1691;
  wire n_1692, n_1694, n_1695, n_1696, n_1697, n_1698, n_1700, n_1701;
  wire n_1702, n_1703, n_1704, n_1706, n_1707, n_1708, n_1709, n_1710;
  wire n_1712, n_1713, n_1714, n_1715, n_1716, n_1718, n_1719, n_1720;
  wire n_1721, n_1722, n_1724, n_1725, n_1726, n_1727, n_1728, n_1730;
  wire n_1731, n_1732, n_1733, n_1734, n_1736, n_1737, n_1738, n_1739;
  wire n_1740, n_1745, n_1747, n_1748, n_1750, n_1752, n_1754, n_1755;
  wire n_1757, n_1758, n_1760, n_1762, n_1764, n_1765, n_1767, n_1768;
  wire n_1770, n_1772, n_1774, n_1775, n_1777, n_1778, n_1780, n_1782;
  wire n_1784, n_1785, n_1787, n_1788, n_1790, n_1792, n_1794, n_1795;
  wire n_1797, n_1798, n_1800, n_1802, n_1804, n_1805, n_1807, n_1808;
  wire n_1810, n_1812, n_1814, n_1815, n_1817, n_1818, n_1820, n_1822;
  wire n_1824, n_1825, n_1827, n_1828, n_1830, n_1832, n_1834, n_1835;
  wire n_1837, n_1838, n_1840, n_1842, n_1844, n_1845, n_1847, n_1848;
  wire n_1850, n_1854, n_1855, n_1856, n_1858, n_1859, n_1860, n_1862;
  wire n_1863, n_1864, n_1865, n_1867, n_1869, n_1871, n_1872, n_1873;
  wire n_1875, n_1876, n_1877, n_1879, n_1880, n_1882, n_1884, n_1886;
  wire n_1887, n_1888, n_1890, n_1891, n_1892, n_1894, n_1895, n_1897;
  wire n_1899, n_1901, n_1902, n_1903, n_1905, n_1906, n_1907, n_1909;
  wire n_1910, n_1912, n_1914, n_1916, n_1917, n_1918, n_1920, n_1921;
  wire n_1922, n_1924, n_1925, n_1927, n_1929, n_1931, n_1932, n_1933;
  wire n_1935, n_1937, n_1938, n_1939, n_1941, n_1942, n_1944, n_1945;
  wire n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953;
  wire n_1954, n_1955, n_1956, n_1957, n_1958, n_1960, n_1963, n_1965;
  wire n_1966, n_1967, n_1970, n_1973, n_1975, n_1976, n_1978, n_1980;
  wire n_1981, n_1983, n_1985, n_1986, n_1988, n_1990, n_1991, n_1993;
  wire n_1994, n_1996, n_1999, n_2001, n_2002, n_2003, n_2006, n_2009;
  wire n_2011, n_2012, n_2014, n_2016, n_2017, n_2019, n_2021, n_2022;
  wire n_2024, n_2026, n_2027, n_2028, n_2030, n_2031, n_2033, n_2034;
  wire n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042;
  wire n_2043, n_2044, n_2046, n_2047, n_2048, n_2050, n_2051, n_2052;
  wire n_2054, n_2055, n_2056, n_2058, n_2059, n_2060, n_2062, n_2063;
  wire n_2064, n_2066, n_2067, n_2068, n_2070, n_2071, n_2072, n_2074;
  wire n_2075, n_2076, n_2078, n_2079, n_2080, n_2082, n_2083, n_2085;
  wire n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093;
  wire n_2094, n_2095, n_2096, n_2098, n_2099, n_2100, n_2102, n_2103;
  wire n_2104, n_2106, n_2107, n_2108, n_2110, n_2111, n_2112, n_2114;
  wire n_2115, n_2116, n_2118, n_2119, n_2120, n_2122, n_2123, n_2125;
  wire n_2128, n_2129, n_2131, n_2132, n_2133, n_2134, n_2136, n_2137;
  wire n_2138, n_2140, n_2141, n_2142, n_2143, n_2145, n_2146, n_2148;
  wire n_2149, n_2151, n_2152, n_2153, n_2154, n_2156, n_2157, n_2158;
  wire n_2160, n_2161, n_2162, n_2163, n_2165, n_2166, n_2168, n_2169;
  wire n_2171, n_2172, n_2173, n_2174, n_2176, n_2177, n_2178, n_2179;
  wire n_2181, n_2182, n_2183, n_2184, n_2186, n_2187, n_2189, n_2190;
  wire n_2192, n_2193, n_2194, n_2195, n_2197, n_2198, n_2199, n_2201;
  wire n_2202, n_2203, n_2204, n_2206, n_2207, n_2209, n_2210, n_2212;
  wire n_2213, n_2214, n_2215, n_2217, n_2218, n_2219, n_2220, n_2222;
  wire n_2223, n_2224, n_2225, n_2227, n_2228, n_2230, n_2231, n_2233;
  wire n_2234, n_2235, n_2236, n_2238, n_2239;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_623, A[1], A[2]);
  xor g270 (n_117, n_623, n_171);
  nand g3 (n_624, A[1], A[2]);
  nand g271 (n_625, n_171, A[2]);
  nand g272 (n_626, A[1], n_171);
  nand g273 (n_172, n_624, n_625, n_626);
  xor g274 (n_627, A[2], A[3]);
  xor g275 (n_116, n_627, n_172);
  nand g276 (n_628, A[2], A[3]);
  nand g4 (n_629, n_172, A[3]);
  nand g277 (n_630, A[2], n_172);
  nand g278 (n_67, n_628, n_629, n_630);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_631, A[4], n_173);
  xor g282 (n_115, n_631, A[6]);
  nand g283 (n_632, A[4], n_173);
  nand g284 (n_633, A[6], n_173);
  nand g5 (n_634, A[4], A[6]);
  nand g6 (n_66, n_632, n_633, n_634);
  xor g287 (n_635, n_68, A[4]);
  xor g288 (n_176, n_635, n_69);
  nand g289 (n_636, n_68, A[4]);
  nand g290 (n_637, n_69, A[4]);
  nand g291 (n_638, n_68, n_69);
  nand g292 (n_179, n_636, n_637, n_638);
  xor g293 (n_639, A[5], n_176);
  xor g294 (n_114, n_639, A[7]);
  nand g295 (n_640, A[5], n_176);
  nand g296 (n_641, A[7], n_176);
  nand g297 (n_642, A[5], A[7]);
  nand g298 (n_65, n_640, n_641, n_642);
  xor g305 (n_647, n_117, A[5]);
  xor g306 (n_180, n_647, A[6]);
  nand g307 (n_648, n_117, A[5]);
  nand g308 (n_649, A[6], A[5]);
  nand g309 (n_650, n_117, A[6]);
  nand g310 (n_183, n_648, n_649, n_650);
  xor g311 (n_651, n_179, A[8]);
  xor g312 (n_113, n_651, n_180);
  nand g313 (n_652, n_179, A[8]);
  nand g314 (n_653, n_180, A[8]);
  nand g315 (n_654, n_179, n_180);
  nand g316 (n_64, n_652, n_653, n_654);
  xor g323 (n_659, A[6], n_116);
  xor g324 (n_184, n_659, A[7]);
  nand g325 (n_660, A[6], n_116);
  nand g326 (n_661, A[7], n_116);
  nand g327 (n_662, A[6], A[7]);
  nand g328 (n_187, n_660, n_661, n_662);
  xor g329 (n_663, A[9], n_183);
  xor g330 (n_112, n_663, n_184);
  nand g331 (n_664, A[9], n_183);
  nand g332 (n_665, n_184, n_183);
  nand g333 (n_666, A[9], n_184);
  nand g334 (n_63, n_664, n_665, n_666);
  xor g338 (n_188, n_631, A[7]);
  nand g340 (n_669, A[7], n_173);
  nand g341 (n_670, A[4], A[7]);
  nand g342 (n_193, n_632, n_669, n_670);
  xor g343 (n_671, n_67, A[8]);
  xor g344 (n_189, n_671, A[10]);
  nand g345 (n_672, n_67, A[8]);
  nand g346 (n_673, A[10], A[8]);
  nand g347 (n_674, n_67, A[10]);
  nand g348 (n_195, n_672, n_673, n_674);
  xor g349 (n_675, n_187, n_188);
  xor g350 (n_111, n_675, n_189);
  nand g351 (n_676, n_187, n_188);
  nand g352 (n_677, n_189, n_188);
  nand g353 (n_678, n_187, n_189);
  nand g354 (n_62, n_676, n_677, n_678);
  xor g364 (n_73, n_639, A[8]);
  nand g366 (n_685, A[8], n_176);
  nand g367 (n_686, A[5], A[8]);
  nand g368 (n_201, n_640, n_685, n_686);
  xor g369 (n_687, A[9], A[11]);
  xor g370 (n_196, n_687, n_193);
  nand g371 (n_688, A[9], A[11]);
  nand g372 (n_689, n_193, A[11]);
  nand g373 (n_690, A[9], n_193);
  nand g374 (n_202, n_688, n_689, n_690);
  xor g375 (n_691, n_73, n_195);
  xor g376 (n_110, n_691, n_196);
  nand g377 (n_692, n_73, n_195);
  nand g378 (n_693, n_196, n_195);
  nand g379 (n_694, n_73, n_196);
  nand g380 (n_61, n_692, n_693, n_694);
  xor g393 (n_703, n_179, A[10]);
  xor g394 (n_203, n_703, n_180);
  nand g395 (n_704, n_179, A[10]);
  nand g396 (n_705, n_180, A[10]);
  nand g398 (n_209, n_704, n_705, n_654);
  xor g399 (n_707, A[12], A[9]);
  xor g400 (n_204, n_707, n_201);
  nand g401 (n_708, A[12], A[9]);
  nand g402 (n_709, n_201, A[9]);
  nand g403 (n_710, A[12], n_201);
  nand g404 (n_211, n_708, n_709, n_710);
  xor g405 (n_711, n_202, n_203);
  xor g406 (n_109, n_711, n_204);
  nand g407 (n_712, n_202, n_203);
  nand g408 (n_713, n_204, n_203);
  nand g409 (n_714, n_202, n_204);
  nand g410 (n_60, n_712, n_713, n_714);
  xor g417 (n_719, A[6], A[7]);
  xor g418 (n_208, n_719, n_116);
  xor g423 (n_723, n_183, A[11]);
  xor g424 (n_210, n_723, A[10]);
  nand g425 (n_724, n_183, A[11]);
  nand g426 (n_725, A[10], A[11]);
  nand g427 (n_726, n_183, A[10]);
  nand g428 (n_217, n_724, n_725, n_726);
  xor g429 (n_727, A[13], n_208);
  xor g430 (n_212, n_727, n_209);
  nand g431 (n_728, A[13], n_208);
  nand g432 (n_729, n_209, n_208);
  nand g433 (n_730, A[13], n_209);
  nand g434 (n_220, n_728, n_729, n_730);
  xor g435 (n_731, n_210, n_211);
  xor g436 (n_108, n_731, n_212);
  nand g437 (n_732, n_210, n_211);
  nand g438 (n_733, n_212, n_211);
  nand g439 (n_734, n_210, n_212);
  nand g440 (n_59, n_732, n_733, n_734);
  xor g444 (n_215, n_631, n_67);
  nand g446 (n_737, n_67, n_173);
  nand g447 (n_738, A[4], n_67);
  nand g448 (n_71, n_632, n_737, n_738);
  xor g449 (n_739, A[7], A[8]);
  xor g450 (n_218, n_739, A[12]);
  nand g451 (n_740, A[7], A[8]);
  nand g452 (n_741, A[12], A[8]);
  nand g453 (n_742, A[7], A[12]);
  nand g454 (n_223, n_740, n_741, n_742);
  xor g455 (n_743, A[11], A[14]);
  xor g456 (n_219, n_743, n_215);
  nand g457 (n_744, A[11], A[14]);
  nand g458 (n_745, n_215, A[14]);
  nand g459 (n_746, A[11], n_215);
  nand g460 (n_225, n_744, n_745, n_746);
  xor g461 (n_747, n_187, n_217);
  xor g462 (n_221, n_747, n_218);
  nand g463 (n_748, n_187, n_217);
  nand g464 (n_749, n_218, n_217);
  nand g465 (n_750, n_187, n_218);
  nand g466 (n_227, n_748, n_749, n_750);
  xor g467 (n_751, n_219, n_220);
  xor g468 (n_107, n_751, n_221);
  nand g469 (n_752, n_219, n_220);
  nand g470 (n_753, n_221, n_220);
  nand g471 (n_754, n_219, n_221);
  nand g472 (n_58, n_752, n_753, n_754);
  xor g488 (n_224, n_707, A[13]);
  nand g490 (n_765, A[13], A[9]);
  nand g491 (n_766, A[12], A[13]);
  nand g492 (n_235, n_708, n_765, n_766);
  xor g493 (n_767, n_71, A[15]);
  xor g494 (n_226, n_767, n_73);
  nand g495 (n_768, n_71, A[15]);
  nand g496 (n_769, n_73, A[15]);
  nand g497 (n_770, n_71, n_73);
  nand g498 (n_236, n_768, n_769, n_770);
  xor g499 (n_771, n_223, n_224);
  xor g500 (n_228, n_771, n_225);
  nand g501 (n_772, n_223, n_224);
  nand g502 (n_773, n_225, n_224);
  nand g503 (n_774, n_223, n_225);
  nand g504 (n_238, n_772, n_773, n_774);
  xor g505 (n_775, n_226, n_227);
  xor g506 (n_106, n_775, n_228);
  nand g507 (n_776, n_226, n_227);
  nand g508 (n_777, n_228, n_227);
  nand g509 (n_778, n_226, n_228);
  nand g510 (n_57, n_776, n_777, n_778);
  xor g523 (n_787, n_179, A[9]);
  xor g524 (n_234, n_787, A[10]);
  nand g525 (n_788, n_179, A[9]);
  nand g526 (n_789, A[10], A[9]);
  nand g528 (n_245, n_788, n_789, n_704);
  xor g529 (n_791, n_180, A[13]);
  xor g530 (n_237, n_791, A[14]);
  nand g531 (n_792, n_180, A[13]);
  nand g532 (n_793, A[14], A[13]);
  nand g533 (n_794, n_180, A[14]);
  nand g534 (n_246, n_792, n_793, n_794);
  xor g535 (n_795, n_201, A[16]);
  xor g536 (n_239, n_795, n_234);
  nand g537 (n_796, n_201, A[16]);
  nand g538 (n_797, n_234, A[16]);
  nand g539 (n_798, n_201, n_234);
  nand g540 (n_249, n_796, n_797, n_798);
  xor g541 (n_799, n_235, n_236);
  xor g542 (n_240, n_799, n_237);
  nand g543 (n_800, n_235, n_236);
  nand g544 (n_801, n_237, n_236);
  nand g545 (n_802, n_235, n_237);
  nand g546 (n_251, n_800, n_801, n_802);
  xor g547 (n_803, n_238, n_239);
  xor g548 (n_105, n_803, n_240);
  nand g549 (n_804, n_238, n_239);
  nand g550 (n_805, n_240, n_239);
  nand g551 (n_806, n_238, n_240);
  nand g552 (n_56, n_804, n_805, n_806);
  xor g565 (n_815, A[10], n_183);
  xor g566 (n_247, n_815, A[11]);
  xor g571 (n_819, A[15], A[14]);
  xor g572 (n_248, n_819, A[17]);
  nand g573 (n_820, A[15], A[14]);
  nand g574 (n_821, A[17], A[14]);
  nand g575 (n_822, A[15], A[17]);
  nand g576 (n_260, n_820, n_821, n_822);
  xor g577 (n_823, n_208, n_245);
  xor g578 (n_250, n_823, n_246);
  nand g579 (n_824, n_208, n_245);
  nand g580 (n_825, n_246, n_245);
  nand g581 (n_826, n_208, n_246);
  nand g582 (n_262, n_824, n_825, n_826);
  xor g583 (n_827, n_247, n_248);
  xor g584 (n_252, n_827, n_249);
  nand g585 (n_828, n_247, n_248);
  nand g586 (n_829, n_249, n_248);
  nand g587 (n_830, n_247, n_249);
  nand g588 (n_119, n_828, n_829, n_830);
  xor g589 (n_831, n_250, n_251);
  xor g590 (n_104, n_831, n_252);
  nand g591 (n_832, n_250, n_251);
  nand g592 (n_833, n_252, n_251);
  nand g593 (n_834, n_250, n_252);
  nand g594 (n_55, n_832, n_833, n_834);
  xor g604 (n_257, n_671, A[11]);
  nand g606 (n_841, A[11], A[8]);
  nand g607 (n_842, n_67, A[11]);
  nand g608 (n_269, n_672, n_841, n_842);
  xor g609 (n_843, A[12], A[15]);
  xor g610 (n_259, n_843, n_187);
  nand g611 (n_844, A[12], A[15]);
  nand g612 (n_845, n_187, A[15]);
  nand g613 (n_846, A[12], n_187);
  nand g614 (n_270, n_844, n_845, n_846);
  xor g615 (n_847, n_188, A[16]);
  xor g616 (n_261, n_847, A[18]);
  nand g617 (n_848, n_188, A[16]);
  nand g618 (n_849, A[18], A[16]);
  nand g619 (n_850, n_188, A[18]);
  nand g620 (n_272, n_848, n_849, n_850);
  xor g621 (n_851, n_257, n_217);
  xor g622 (n_263, n_851, n_259);
  nand g623 (n_852, n_257, n_217);
  nand g624 (n_853, n_259, n_217);
  nand g625 (n_854, n_257, n_259);
  nand g626 (n_275, n_852, n_853, n_854);
  xor g627 (n_855, n_260, n_261);
  xor g628 (n_118, n_855, n_262);
  nand g629 (n_856, n_260, n_261);
  nand g630 (n_857, n_262, n_261);
  nand g631 (n_858, n_260, n_262);
  nand g632 (n_277, n_856, n_857, n_858);
  xor g633 (n_859, n_263, n_118);
  xor g634 (n_103, n_859, n_119);
  nand g635 (n_860, n_263, n_118);
  nand g636 (n_861, n_119, n_118);
  nand g637 (n_862, n_263, n_119);
  nand g638 (n_54, n_860, n_861, n_862);
  xor g659 (n_875, n_193, A[17]);
  xor g660 (n_274, n_875, A[19]);
  nand g661 (n_876, n_193, A[17]);
  nand g662 (n_877, A[19], A[17]);
  nand g663 (n_878, n_193, A[19]);
  nand g664 (n_287, n_876, n_877, n_878);
  xor g665 (n_879, A[16], n_73);
  xor g666 (n_273, n_879, n_269);
  nand g667 (n_880, A[16], n_73);
  nand g668 (n_881, n_269, n_73);
  nand g669 (n_882, A[16], n_269);
  nand g670 (n_288, n_880, n_881, n_882);
  xor g671 (n_883, n_270, n_224);
  xor g672 (n_276, n_883, n_272);
  nand g673 (n_884, n_270, n_224);
  nand g674 (n_885, n_272, n_224);
  nand g675 (n_886, n_270, n_272);
  nand g676 (n_290, n_884, n_885, n_886);
  xor g677 (n_887, n_273, n_274);
  xor g678 (n_278, n_887, n_275);
  nand g679 (n_888, n_273, n_274);
  nand g680 (n_889, n_275, n_274);
  nand g681 (n_890, n_273, n_275);
  nand g682 (n_293, n_888, n_889, n_890);
  xor g683 (n_891, n_276, n_277);
  xor g684 (n_102, n_891, n_278);
  nand g685 (n_892, n_276, n_277);
  nand g686 (n_893, n_278, n_277);
  nand g687 (n_894, n_276, n_278);
  nand g688 (n_53, n_892, n_893, n_894);
  xor g707 (n_907, A[9], A[13]);
  xor g708 (n_286, n_907, A[14]);
  nand g711 (n_910, A[9], A[14]);
  nand g712 (n_300, n_765, n_793, n_910);
  xor g713 (n_911, A[18], A[20]);
  xor g714 (n_289, n_911, A[17]);
  nand g715 (n_912, A[18], A[20]);
  nand g716 (n_913, A[17], A[20]);
  nand g717 (n_914, A[18], A[17]);
  nand g718 (n_302, n_912, n_913, n_914);
  xor g719 (n_915, n_201, n_203);
  xor g720 (n_291, n_915, n_235);
  nand g721 (n_916, n_201, n_203);
  nand g722 (n_917, n_235, n_203);
  nand g723 (n_918, n_201, n_235);
  nand g724 (n_305, n_916, n_917, n_918);
  xor g725 (n_919, n_286, n_287);
  xor g726 (n_292, n_919, n_288);
  nand g727 (n_920, n_286, n_287);
  nand g728 (n_921, n_288, n_287);
  nand g729 (n_922, n_286, n_288);
  nand g730 (n_307, n_920, n_921, n_922);
  xor g731 (n_923, n_289, n_290);
  xor g732 (n_294, n_923, n_291);
  nand g733 (n_924, n_289, n_290);
  nand g734 (n_925, n_291, n_290);
  nand g735 (n_926, n_289, n_291);
  nand g736 (n_309, n_924, n_925, n_926);
  xor g737 (n_927, n_292, n_293);
  xor g738 (n_101, n_927, n_294);
  nand g739 (n_928, n_292, n_293);
  nand g740 (n_929, n_294, n_293);
  nand g741 (n_930, n_292, n_294);
  nand g742 (n_52, n_928, n_929, n_930);
  xor g755 (n_939, A[11], A[10]);
  xor g756 (n_301, n_939, n_183);
  xor g762 (n_303, n_819, n_208);
  nand g764 (n_945, n_208, A[15]);
  nand g765 (n_946, A[14], n_208);
  nand g766 (n_318, n_820, n_945, n_946);
  xor g767 (n_947, A[19], A[18]);
  xor g768 (n_304, n_947, A[21]);
  nand g769 (n_948, A[19], A[18]);
  nand g770 (n_949, A[21], A[18]);
  nand g771 (n_950, A[19], A[21]);
  nand g772 (n_320, n_948, n_949, n_950);
  xor g773 (n_951, n_209, n_300);
  xor g774 (n_306, n_951, n_301);
  nand g775 (n_952, n_209, n_300);
  nand g776 (n_953, n_301, n_300);
  nand g777 (n_954, n_209, n_301);
  nand g778 (n_322, n_952, n_953, n_954);
  xor g779 (n_955, n_302, n_303);
  xor g780 (n_308, n_955, n_304);
  nand g781 (n_956, n_302, n_303);
  nand g782 (n_957, n_304, n_303);
  nand g783 (n_958, n_302, n_304);
  nand g784 (n_323, n_956, n_957, n_958);
  xor g785 (n_959, n_305, n_306);
  xor g786 (n_310, n_959, n_307);
  nand g787 (n_960, n_305, n_306);
  nand g788 (n_961, n_307, n_306);
  nand g789 (n_962, n_305, n_307);
  nand g790 (n_326, n_960, n_961, n_962);
  xor g791 (n_963, n_308, n_309);
  xor g792 (n_100, n_963, n_310);
  nand g793 (n_964, n_308, n_309);
  nand g794 (n_965, n_310, n_309);
  nand g795 (n_966, n_308, n_310);
  nand g796 (n_51, n_964, n_965, n_966);
  xor g806 (n_315, n_671, A[12]);
  nand g809 (n_974, n_67, A[12]);
  nand g810 (n_333, n_672, n_741, n_974);
  xor g811 (n_975, A[11], n_188);
  xor g812 (n_317, n_975, A[15]);
  nand g813 (n_976, A[11], n_188);
  nand g814 (n_977, A[15], n_188);
  nand g815 (n_978, A[11], A[15]);
  nand g816 (n_334, n_976, n_977, n_978);
  xor g817 (n_979, n_187, A[20]);
  xor g818 (n_319, n_979, A[16]);
  nand g819 (n_980, n_187, A[20]);
  nand g820 (n_981, A[16], A[20]);
  nand g821 (n_982, n_187, A[16]);
  nand g822 (n_336, n_980, n_981, n_982);
  xor g823 (n_983, A[19], n_315);
  xor g824 (n_321, n_983, A[22]);
  nand g825 (n_984, A[19], n_315);
  nand g826 (n_985, A[22], n_315);
  nand g827 (n_986, A[19], A[22]);
  nand g828 (n_337, n_984, n_985, n_986);
  xor g829 (n_987, n_217, n_317);
  xor g830 (n_324, n_987, n_318);
  nand g831 (n_988, n_217, n_317);
  nand g832 (n_989, n_318, n_317);
  nand g833 (n_990, n_217, n_318);
  nand g834 (n_341, n_988, n_989, n_990);
  xor g835 (n_991, n_319, n_320);
  xor g836 (n_325, n_991, n_321);
  nand g837 (n_992, n_319, n_320);
  nand g838 (n_993, n_321, n_320);
  nand g839 (n_994, n_319, n_321);
  nand g840 (n_343, n_992, n_993, n_994);
  xor g841 (n_995, n_322, n_323);
  xor g842 (n_327, n_995, n_324);
  nand g843 (n_996, n_322, n_323);
  nand g844 (n_997, n_324, n_323);
  nand g845 (n_998, n_322, n_324);
  nand g846 (n_345, n_996, n_997, n_998);
  xor g847 (n_999, n_325, n_326);
  xor g848 (n_99, n_999, n_327);
  nand g849 (n_1000, n_325, n_326);
  nand g850 (n_1001, n_327, n_326);
  nand g851 (n_1002, n_325, n_327);
  nand g852 (n_50, n_1000, n_1001, n_1002);
  xor g874 (n_339, n_875, n_73);
  nand g876 (n_1017, n_73, A[17]);
  nand g877 (n_1018, n_193, n_73);
  nand g878 (n_357, n_876, n_1017, n_1018);
  xor g879 (n_1019, A[16], A[20]);
  xor g880 (n_338, n_1019, A[21]);
  nand g882 (n_1021, A[21], A[20]);
  nand g883 (n_1022, A[16], A[21]);
  nand g884 (n_358, n_981, n_1021, n_1022);
  xor g885 (n_1023, A[23], n_333);
  xor g886 (n_340, n_1023, n_334);
  nand g887 (n_1024, A[23], n_333);
  nand g888 (n_1025, n_334, n_333);
  nand g889 (n_1026, A[23], n_334);
  nand g890 (n_360, n_1024, n_1025, n_1026);
  xor g891 (n_1027, n_224, n_336);
  xor g892 (n_342, n_1027, n_337);
  nand g893 (n_1028, n_224, n_336);
  nand g894 (n_1029, n_337, n_336);
  nand g895 (n_1030, n_224, n_337);
  nand g896 (n_363, n_1028, n_1029, n_1030);
  xor g897 (n_1031, n_338, n_339);
  xor g898 (n_344, n_1031, n_340);
  nand g899 (n_1032, n_338, n_339);
  nand g900 (n_1033, n_340, n_339);
  nand g901 (n_1034, n_338, n_340);
  nand g902 (n_364, n_1032, n_1033, n_1034);
  xor g903 (n_1035, n_341, n_342);
  xor g904 (n_346, n_1035, n_343);
  nand g905 (n_1036, n_341, n_342);
  nand g906 (n_1037, n_343, n_342);
  nand g907 (n_1038, n_341, n_343);
  nand g908 (n_367, n_1036, n_1037, n_1038);
  xor g909 (n_1039, n_344, n_345);
  xor g910 (n_98, n_1039, n_346);
  nand g911 (n_1040, n_344, n_345);
  nand g912 (n_1041, n_346, n_345);
  nand g913 (n_1042, n_344, n_346);
  nand g914 (n_49, n_1040, n_1041, n_1042);
  xor g917 (n_1043, A[2], n_171);
  nand g922 (n_372, n_625, n_1045, n_1046);
  xor g923 (n_1047, A[5], n_350);
  xor g924 (n_352, n_1047, A[6]);
  nand g925 (n_1048, A[5], n_350);
  nand g926 (n_1049, A[6], n_350);
  nand g928 (n_374, n_1048, n_1049, n_649);
  xor g935 (n_1055, n_352, A[14]);
  xor g936 (n_356, n_1055, A[13]);
  nand g937 (n_1056, n_352, A[14]);
  nand g939 (n_1058, n_352, A[13]);
  nand g940 (n_378, n_1056, n_793, n_1058);
  xor g941 (n_1059, n_201, A[18]);
  xor g942 (n_359, n_1059, A[17]);
  nand g943 (n_1060, n_201, A[18]);
  nand g945 (n_1062, n_201, A[17]);
  nand g946 (n_380, n_1060, n_914, n_1062);
  xor g948 (n_361, n_1063, A[21]);
  nand g950 (n_1065, A[21], A[22]);
  nand g952 (n_381, n_1064, n_1065, n_1066);
  xor g953 (n_1067, n_235, n_234);
  xor g954 (n_362, n_1067, n_356);
  nand g955 (n_1068, n_235, n_234);
  nand g956 (n_1069, n_356, n_234);
  nand g957 (n_1070, n_235, n_356);
  nand g958 (n_384, n_1068, n_1069, n_1070);
  xor g959 (n_1071, n_357, n_358);
  xor g960 (n_365, n_1071, n_359);
  nand g961 (n_1072, n_357, n_358);
  nand g962 (n_1073, n_359, n_358);
  nand g963 (n_1074, n_357, n_359);
  nand g964 (n_386, n_1072, n_1073, n_1074);
  xor g965 (n_1075, n_360, n_361);
  xor g966 (n_366, n_1075, n_362);
  nand g967 (n_1076, n_360, n_361);
  nand g968 (n_1077, n_362, n_361);
  nand g969 (n_1078, n_360, n_362);
  nand g970 (n_388, n_1076, n_1077, n_1078);
  xor g971 (n_1079, n_363, n_364);
  xor g972 (n_368, n_1079, n_365);
  nand g973 (n_1080, n_363, n_364);
  nand g974 (n_1081, n_365, n_364);
  nand g975 (n_1082, n_363, n_365);
  nand g976 (n_390, n_1080, n_1081, n_1082);
  xor g977 (n_1083, n_366, n_367);
  xor g978 (n_97, n_1083, n_368);
  nand g979 (n_1084, n_366, n_367);
  nand g980 (n_1085, n_368, n_367);
  nand g981 (n_1086, n_366, n_368);
  nand g982 (n_48, n_1084, n_1085, n_1086);
  xor g985 (n_1087, A[1], A[3]);
  nand g987 (n_1088, A[1], A[3]);
  nand g990 (n_393, n_1088, n_1089, n_1090);
  xor g991 (n_1091, n_372, A[6]);
  xor g992 (n_375, n_1091, n_373);
  nand g993 (n_1092, n_372, A[6]);
  nand g994 (n_1093, n_373, A[6]);
  nand g995 (n_1094, n_372, n_373);
  nand g996 (n_395, n_1092, n_1093, n_1094);
  xor g997 (n_1095, A[7], A[10]);
  xor g998 (n_377, n_1095, n_374);
  nand g999 (n_1096, A[7], A[10]);
  nand g1000 (n_1097, n_374, A[10]);
  nand g1001 (n_1098, A[7], n_374);
  nand g1002 (n_397, n_1096, n_1097, n_1098);
  xor g1003 (n_1099, A[11], n_375);
  xor g1004 (n_379, n_1099, A[15]);
  nand g1005 (n_1100, A[11], n_375);
  nand g1006 (n_1101, A[15], n_375);
  nand g1008 (n_399, n_1100, n_1101, n_978);
  xor g1009 (n_1103, A[14], A[18]);
  xor g1010 (n_382, n_1103, A[19]);
  nand g1011 (n_1104, A[14], A[18]);
  nand g1013 (n_1106, A[14], A[19]);
  nand g1014 (n_401, n_1104, n_948, n_1106);
  xor g1015 (n_1107, A[22], A[23]);
  xor g1016 (n_383, n_1107, n_245);
  nand g1017 (n_1108, A[22], A[23]);
  nand g1018 (n_1109, n_245, A[23]);
  nand g1019 (n_1110, A[22], n_245);
  nand g1020 (n_402, n_1108, n_1109, n_1110);
  xor g1021 (n_1111, n_377, n_378);
  xor g1022 (n_385, n_1111, n_379);
  nand g1023 (n_1112, n_377, n_378);
  nand g1024 (n_1113, n_379, n_378);
  nand g1025 (n_1114, n_377, n_379);
  nand g1026 (n_406, n_1112, n_1113, n_1114);
  xor g1027 (n_1115, n_380, n_381);
  xor g1028 (n_387, n_1115, n_382);
  nand g1029 (n_1116, n_380, n_381);
  nand g1030 (n_1117, n_382, n_381);
  nand g1031 (n_1118, n_380, n_382);
  nand g1032 (n_407, n_1116, n_1117, n_1118);
  xor g1033 (n_1119, n_383, n_384);
  xor g1034 (n_389, n_1119, n_385);
  nand g1035 (n_1120, n_383, n_384);
  nand g1036 (n_1121, n_385, n_384);
  nand g1037 (n_1122, n_383, n_385);
  nand g1038 (n_409, n_1120, n_1121, n_1122);
  xor g1039 (n_1123, n_386, n_387);
  xor g1040 (n_391, n_1123, n_388);
  nand g1041 (n_1124, n_386, n_387);
  nand g1042 (n_1125, n_388, n_387);
  nand g1043 (n_1126, n_386, n_388);
  nand g1044 (n_412, n_1124, n_1125, n_1126);
  xor g1045 (n_1127, n_389, n_390);
  xor g1046 (n_96, n_1127, n_391);
  nand g1047 (n_1128, n_389, n_390);
  nand g1048 (n_1129, n_391, n_390);
  nand g1049 (n_1130, n_389, n_391);
  nand g1050 (n_47, n_1128, n_1129, n_1130);
  xor g1052 (n_394, n_627, A[4]);
  nand g1054 (n_1133, A[4], A[2]);
  nand g1055 (n_1134, A[3], A[4]);
  nand g1056 (n_413, n_628, n_1133, n_1134);
  xor g1057 (n_1135, n_393, n_394);
  xor g1058 (n_396, n_1135, A[7]);
  nand g1059 (n_1136, n_393, n_394);
  nand g1060 (n_1137, A[7], n_394);
  nand g1061 (n_1138, n_393, A[7]);
  nand g1062 (n_415, n_1136, n_1137, n_1138);
  xor g1063 (n_1139, A[8], A[11]);
  xor g1064 (n_398, n_1139, A[12]);
  nand g1066 (n_1141, A[12], A[11]);
  nand g1068 (n_416, n_841, n_1141, n_741);
  xor g1069 (n_1143, n_395, n_396);
  xor g1070 (n_400, n_1143, A[15]);
  nand g1071 (n_1144, n_395, n_396);
  nand g1072 (n_1145, A[15], n_396);
  nand g1073 (n_1146, n_395, A[15]);
  nand g1074 (n_418, n_1144, n_1145, n_1146);
  xor g1075 (n_1147, A[19], A[16]);
  xor g1076 (n_403, n_1147, A[20]);
  nand g1077 (n_1148, A[19], A[16]);
  nand g1079 (n_1150, A[19], A[20]);
  nand g1080 (n_419, n_1148, n_981, n_1150);
  xor g1082 (n_404, n_1151, n_397);
  nand g1084 (n_1153, n_397, A[23]);
  nand g1086 (n_422, n_1152, n_1153, n_1154);
  xor g1087 (n_1155, n_398, n_399);
  xor g1088 (n_405, n_1155, n_400);
  nand g1089 (n_1156, n_398, n_399);
  nand g1090 (n_1157, n_400, n_399);
  nand g1091 (n_1158, n_398, n_400);
  nand g1092 (n_424, n_1156, n_1157, n_1158);
  xor g1093 (n_1159, n_401, n_402);
  xor g1094 (n_408, n_1159, n_403);
  nand g1095 (n_1160, n_401, n_402);
  nand g1096 (n_1161, n_403, n_402);
  nand g1097 (n_1162, n_401, n_403);
  nand g1098 (n_426, n_1160, n_1161, n_1162);
  xor g1099 (n_1163, n_404, n_405);
  xor g1100 (n_410, n_1163, n_406);
  nand g1101 (n_1164, n_404, n_405);
  nand g1102 (n_1165, n_406, n_405);
  nand g1103 (n_1166, n_404, n_406);
  nand g1104 (n_428, n_1164, n_1165, n_1166);
  xor g1105 (n_1167, n_407, n_408);
  xor g1106 (n_411, n_1167, n_409);
  nand g1107 (n_1168, n_407, n_408);
  nand g1108 (n_1169, n_409, n_408);
  nand g1109 (n_1170, n_407, n_409);
  nand g1110 (n_431, n_1168, n_1169, n_1170);
  xor g1111 (n_1171, n_410, n_411);
  xor g1112 (n_95, n_1171, n_412);
  nand g1113 (n_1172, n_410, n_411);
  nand g1114 (n_1173, n_412, n_411);
  nand g1115 (n_1174, n_410, n_412);
  nand g1116 (n_46, n_1172, n_1173, n_1174);
  xor g1117 (n_1175, A[4], A[5]);
  xor g1118 (n_414, n_1175, n_413);
  nand g1119 (n_1176, A[4], A[5]);
  nand g1120 (n_1177, n_413, A[5]);
  nand g1121 (n_1178, A[4], n_413);
  nand g1122 (n_434, n_1176, n_1177, n_1178);
  xor g1123 (n_1179, A[8], A[9]);
  xor g1124 (n_417, n_1179, A[12]);
  nand g1125 (n_1180, A[8], A[9]);
  nand g1128 (n_436, n_1180, n_708, n_741);
  xor g1129 (n_1183, n_414, A[13]);
  xor g1130 (n_420, n_1183, n_415);
  nand g1131 (n_1184, n_414, A[13]);
  nand g1132 (n_1185, n_415, A[13]);
  nand g1133 (n_1186, n_414, n_415);
  nand g1134 (n_438, n_1184, n_1185, n_1186);
  xor g1135 (n_1187, A[17], A[16]);
  xor g1136 (n_421, n_1187, A[20]);
  nand g1137 (n_1188, A[17], A[16]);
  nand g1140 (n_439, n_1188, n_981, n_913);
  xor g1142 (n_423, n_1191, n_416);
  nand g1144 (n_1193, n_416, A[21]);
  nand g1146 (n_441, n_1066, n_1193, n_1194);
  xor g1147 (n_1195, n_417, n_418);
  xor g1148 (n_425, n_1195, n_419);
  nand g1149 (n_1196, n_417, n_418);
  nand g1150 (n_1197, n_419, n_418);
  nand g1151 (n_1198, n_417, n_419);
  nand g1152 (n_443, n_1196, n_1197, n_1198);
  xor g1153 (n_1199, n_420, n_421);
  xor g1154 (n_427, n_1199, n_422);
  nand g1155 (n_1200, n_420, n_421);
  nand g1156 (n_1201, n_422, n_421);
  nand g1157 (n_1202, n_420, n_422);
  nand g1158 (n_445, n_1200, n_1201, n_1202);
  xor g1159 (n_1203, n_423, n_424);
  xor g1160 (n_429, n_1203, n_425);
  nand g1161 (n_1204, n_423, n_424);
  nand g1162 (n_1205, n_425, n_424);
  nand g1163 (n_1206, n_423, n_425);
  nand g1164 (n_447, n_1204, n_1205, n_1206);
  xor g1165 (n_1207, n_426, n_427);
  xor g1166 (n_430, n_1207, n_428);
  nand g1167 (n_1208, n_426, n_427);
  nand g1168 (n_1209, n_428, n_427);
  nand g1169 (n_1210, n_426, n_428);
  nand g1170 (n_450, n_1208, n_1209, n_1210);
  xor g1171 (n_1211, n_429, n_430);
  xor g1172 (n_94, n_1211, n_431);
  nand g1173 (n_1212, n_429, n_430);
  nand g1174 (n_1213, n_431, n_430);
  nand g1175 (n_1214, n_429, n_431);
  nand g1176 (n_45, n_1212, n_1213, n_1214);
  xor g1180 (n_435, n_1215, A[9]);
  nand g1183 (n_1218, A[6], A[9]);
  nand g1184 (n_455, n_1216, n_1217, n_1218);
  xor g1185 (n_1219, A[10], n_434);
  xor g1186 (n_437, n_1219, A[14]);
  nand g1187 (n_1220, A[10], n_434);
  nand g1188 (n_1221, A[14], n_434);
  nand g1189 (n_1222, A[10], A[14]);
  nand g1190 (n_457, n_1220, n_1221, n_1222);
  xor g1191 (n_1223, A[13], A[18]);
  xor g1192 (n_440, n_1223, A[17]);
  nand g1193 (n_1224, A[13], A[18]);
  nand g1195 (n_1226, A[13], A[17]);
  nand g1196 (n_458, n_1224, n_914, n_1226);
  xor g1197 (n_1227, A[21], n_435);
  xor g1198 (n_442, n_1227, A[22]);
  nand g1199 (n_1228, A[21], n_435);
  nand g1200 (n_1229, A[22], n_435);
  nand g1202 (n_460, n_1228, n_1229, n_1065);
  xor g1203 (n_1231, n_436, n_437);
  xor g1204 (n_444, n_1231, n_438);
  nand g1205 (n_1232, n_436, n_437);
  nand g1206 (n_1233, n_438, n_437);
  nand g1207 (n_1234, n_436, n_438);
  nand g1208 (n_462, n_1232, n_1233, n_1234);
  xor g1209 (n_1235, n_439, n_440);
  xor g1210 (n_446, n_1235, n_441);
  nand g1211 (n_1236, n_439, n_440);
  nand g1212 (n_1237, n_441, n_440);
  nand g1213 (n_1238, n_439, n_441);
  nand g1214 (n_464, n_1236, n_1237, n_1238);
  xor g1215 (n_1239, n_442, n_443);
  xor g1216 (n_448, n_1239, n_444);
  nand g1217 (n_1240, n_442, n_443);
  nand g1218 (n_1241, n_444, n_443);
  nand g1219 (n_1242, n_442, n_444);
  nand g1220 (n_466, n_1240, n_1241, n_1242);
  xor g1221 (n_1243, n_445, n_446);
  xor g1222 (n_449, n_1243, n_447);
  nand g1223 (n_1244, n_445, n_446);
  nand g1224 (n_1245, n_447, n_446);
  nand g1225 (n_1246, n_445, n_447);
  nand g1226 (n_469, n_1244, n_1245, n_1246);
  xor g1227 (n_1247, n_448, n_449);
  xor g1228 (n_93, n_1247, n_450);
  nand g1229 (n_1248, n_448, n_449);
  nand g1230 (n_1249, n_450, n_449);
  nand g1231 (n_1250, n_448, n_450);
  nand g1232 (n_44, n_1248, n_1249, n_1250);
  xor g1235 (n_1251, A[7], A[5]);
  nand g1240 (n_471, n_642, n_1253, n_1254);
  xor g1242 (n_456, n_939, A[15]);
  nand g1245 (n_1258, A[10], A[15]);
  nand g1246 (n_474, n_725, n_978, n_1258);
  xor g1247 (n_1259, A[14], A[19]);
  xor g1248 (n_459, n_1259, n_454);
  nand g1250 (n_1261, n_454, A[19]);
  nand g1251 (n_1262, A[14], n_454);
  nand g1252 (n_475, n_1106, n_1261, n_1262);
  xor g1253 (n_1263, A[18], A[22]);
  xor g1254 (n_461, n_1263, A[23]);
  nand g1255 (n_1264, A[18], A[22]);
  nand g1257 (n_1266, A[18], A[23]);
  nand g1258 (n_477, n_1264, n_1108, n_1266);
  xor g1259 (n_1267, n_455, n_456);
  xor g1260 (n_463, n_1267, n_457);
  nand g1261 (n_1268, n_455, n_456);
  nand g1262 (n_1269, n_457, n_456);
  nand g1263 (n_1270, n_455, n_457);
  nand g1264 (n_479, n_1268, n_1269, n_1270);
  xor g1265 (n_1271, n_458, n_459);
  xor g1266 (n_465, n_1271, n_460);
  nand g1267 (n_1272, n_458, n_459);
  nand g1268 (n_1273, n_460, n_459);
  nand g1269 (n_1274, n_458, n_460);
  nand g1270 (n_481, n_1272, n_1273, n_1274);
  xor g1271 (n_1275, n_461, n_462);
  xor g1272 (n_467, n_1275, n_463);
  nand g1273 (n_1276, n_461, n_462);
  nand g1274 (n_1277, n_463, n_462);
  nand g1275 (n_1278, n_461, n_463);
  nand g1276 (n_484, n_1276, n_1277, n_1278);
  xor g1277 (n_1279, n_464, n_465);
  xor g1278 (n_468, n_1279, n_466);
  nand g1279 (n_1280, n_464, n_465);
  nand g1280 (n_1281, n_466, n_465);
  nand g1281 (n_1282, n_464, n_466);
  nand g1282 (n_486, n_1280, n_1281, n_1282);
  xor g1283 (n_1283, n_467, n_468);
  xor g1284 (n_92, n_1283, n_469);
  nand g1285 (n_1284, n_467, n_468);
  nand g1286 (n_1285, n_469, n_468);
  nand g1287 (n_1286, n_467, n_469);
  nand g1288 (n_43, n_1284, n_1285, n_1286);
  xor g1290 (n_472, n_739, A[6]);
  nand g1292 (n_1289, A[6], A[8]);
  nand g1294 (n_487, n_740, n_1289, n_662);
  xor g1295 (n_1291, A[11], A[12]);
  xor g1296 (n_473, n_1291, A[15]);
  nand g1300 (n_489, n_1141, n_844, n_978);
  xor g1308 (n_476, n_1299, A[23]);
  nand g1311 (n_1302, n_471, A[23]);
  nand g1312 (n_492, n_1300, n_1152, n_1302);
  xor g1313 (n_1303, n_472, n_473);
  xor g1314 (n_480, n_1303, n_474);
  nand g1315 (n_1304, n_472, n_473);
  nand g1316 (n_1305, n_474, n_473);
  nand g1317 (n_1306, n_472, n_474);
  nand g1318 (n_494, n_1304, n_1305, n_1306);
  xor g1319 (n_1307, n_475, n_476);
  xor g1320 (n_482, n_1307, n_477);
  nand g1321 (n_1308, n_475, n_476);
  nand g1322 (n_1309, n_477, n_476);
  nand g1323 (n_1310, n_475, n_477);
  nand g1324 (n_496, n_1308, n_1309, n_1310);
  xor g1325 (n_1311, n_403, n_479);
  xor g1326 (n_483, n_1311, n_480);
  nand g1327 (n_1312, n_403, n_479);
  nand g1328 (n_1313, n_480, n_479);
  nand g1329 (n_1314, n_403, n_480);
  nand g1330 (n_499, n_1312, n_1313, n_1314);
  xor g1331 (n_1315, n_481, n_482);
  xor g1332 (n_485, n_1315, n_483);
  nand g1333 (n_1316, n_481, n_482);
  nand g1334 (n_1317, n_483, n_482);
  nand g1335 (n_1318, n_481, n_483);
  nand g1336 (n_501, n_1316, n_1317, n_1318);
  xor g1337 (n_1319, n_484, n_485);
  xor g1338 (n_91, n_1319, n_486);
  nand g1339 (n_1320, n_484, n_485);
  nand g1340 (n_1321, n_486, n_485);
  nand g1341 (n_1322, n_484, n_486);
  nand g1342 (n_42, n_1320, n_1321, n_1322);
  xor g1343 (n_1323, A[8], A[12]);
  xor g1344 (n_488, n_1323, A[9]);
  xor g1349 (n_1327, A[13], A[17]);
  xor g1350 (n_493, n_1327, A[16]);
  nand g1353 (n_1330, A[13], A[16]);
  nand g1354 (n_505, n_1226, n_1188, n_1330);
  xor g1355 (n_1331, n_487, A[20]);
  nand g1357 (n_1332, n_487, A[20]);
  nand g1360 (n_506, n_1332, n_1333, n_1334);
  xor g1361 (n_1335, A[21], n_488);
  xor g1362 (n_495, n_1335, n_489);
  nand g1363 (n_1336, A[21], n_488);
  nand g1364 (n_1337, n_489, n_488);
  nand g1365 (n_1338, A[21], n_489);
  nand g1366 (n_509, n_1336, n_1337, n_1338);
  xor g1367 (n_1339, n_419, n_491);
  xor g1368 (n_497, n_1339, n_492);
  nand g1369 (n_1340, n_419, n_491);
  nand g1370 (n_1341, n_492, n_491);
  nand g1371 (n_1342, n_419, n_492);
  nand g1372 (n_512, n_1340, n_1341, n_1342);
  xor g1373 (n_1343, n_493, n_494);
  xor g1374 (n_498, n_1343, n_495);
  nand g1375 (n_1344, n_493, n_494);
  nand g1376 (n_1345, n_495, n_494);
  nand g1377 (n_1346, n_493, n_495);
  nand g1378 (n_513, n_1344, n_1345, n_1346);
  xor g1379 (n_1347, n_496, n_497);
  xor g1380 (n_500, n_1347, n_498);
  nand g1381 (n_1348, n_496, n_497);
  nand g1382 (n_1349, n_498, n_497);
  nand g1383 (n_1350, n_496, n_498);
  nand g1384 (n_516, n_1348, n_1349, n_1350);
  xor g1385 (n_1351, n_499, n_500);
  xor g1386 (n_90, n_1351, n_501);
  nand g1387 (n_1352, n_499, n_500);
  nand g1388 (n_1353, n_501, n_500);
  nand g1389 (n_1354, n_499, n_501);
  nand g1390 (n_41, n_1352, n_1353, n_1354);
  xor g1393 (n_1355, A[9], A[14]);
  xor g1394 (n_507, n_1355, A[13]);
  xor g1400 (n_508, n_1359, A[17]);
  nand g1404 (n_521, n_1360, n_1361, n_914);
  xor g1405 (n_1363, A[21], n_436);
  xor g1406 (n_510, n_1363, A[22]);
  nand g1407 (n_1364, A[21], n_436);
  nand g1408 (n_1365, A[22], n_436);
  nand g1410 (n_524, n_1364, n_1365, n_1065);
  xor g1411 (n_1367, n_505, n_506);
  xor g1412 (n_511, n_1367, n_507);
  nand g1413 (n_1368, n_505, n_506);
  nand g1414 (n_1369, n_507, n_506);
  nand g1415 (n_1370, n_505, n_507);
  nand g1416 (n_526, n_1368, n_1369, n_1370);
  xor g1417 (n_1371, n_508, n_509);
  xor g1418 (n_514, n_1371, n_510);
  nand g1419 (n_1372, n_508, n_509);
  nand g1420 (n_1373, n_510, n_509);
  nand g1421 (n_1374, n_508, n_510);
  nand g1422 (n_528, n_1372, n_1373, n_1374);
  xor g1423 (n_1375, n_511, n_512);
  xor g1424 (n_515, n_1375, n_513);
  nand g1425 (n_1376, n_511, n_512);
  nand g1426 (n_1377, n_513, n_512);
  nand g1427 (n_1378, n_511, n_513);
  nand g1428 (n_531, n_1376, n_1377, n_1378);
  xor g1429 (n_1379, n_514, n_515);
  xor g1430 (n_89, n_1379, n_516);
  nand g1431 (n_1380, n_514, n_515);
  nand g1432 (n_1381, n_516, n_515);
  nand g1433 (n_1382, n_514, n_516);
  nand g1434 (n_40, n_1380, n_1381, n_1382);
  xor g1437 (n_1383, A[10], A[15]);
  xor g1438 (n_522, n_1383, A[14]);
  nand g1442 (n_534, n_1258, n_820, n_1222);
  xor g1444 (n_523, n_1387, A[18]);
  nand g1448 (n_535, n_1388, n_1389, n_948);
  xor g1449 (n_1391, A[10], A[22]);
  xor g1450 (n_525, n_1391, A[23]);
  nand g1451 (n_1392, A[10], A[22]);
  nand g1453 (n_1394, A[10], A[23]);
  nand g1454 (n_538, n_1392, n_1108, n_1394);
  xor g1455 (n_1395, n_300, n_521);
  xor g1456 (n_527, n_1395, n_522);
  nand g1457 (n_1396, n_300, n_521);
  nand g1458 (n_1397, n_522, n_521);
  nand g1459 (n_1398, n_300, n_522);
  nand g1460 (n_539, n_1396, n_1397, n_1398);
  xor g1461 (n_1399, n_523, n_524);
  xor g1462 (n_529, n_1399, n_525);
  nand g1463 (n_1400, n_523, n_524);
  nand g1464 (n_1401, n_525, n_524);
  nand g1465 (n_1402, n_523, n_525);
  nand g1466 (n_542, n_1400, n_1401, n_1402);
  xor g1467 (n_1403, n_526, n_527);
  xor g1468 (n_530, n_1403, n_528);
  nand g1469 (n_1404, n_526, n_527);
  nand g1470 (n_1405, n_528, n_527);
  nand g1471 (n_1406, n_526, n_528);
  nand g1472 (n_544, n_1404, n_1405, n_1406);
  xor g1473 (n_1407, n_529, n_530);
  xor g1474 (n_88, n_1407, n_531);
  nand g1475 (n_1408, n_529, n_530);
  nand g1476 (n_1409, n_531, n_530);
  nand g1477 (n_1410, n_529, n_531);
  nand g1478 (n_39, n_1408, n_1409, n_1410);
  nand g1487 (n_1416, A[19], A[11]);
  nand g1488 (n_1417, A[16], A[11]);
  nand g1490 (n_546, n_1416, n_1417, n_1148);
  xor g1492 (n_536, n_1419, A[23]);
  nand g1495 (n_1422, A[20], A[23]);
  nand g1496 (n_549, n_1333, n_1152, n_1422);
  xor g1497 (n_1423, n_473, n_534);
  xor g1498 (n_540, n_1423, n_535);
  nand g1499 (n_1424, n_473, n_534);
  nand g1500 (n_1425, n_535, n_534);
  nand g1501 (n_1426, n_473, n_535);
  nand g1502 (n_551, n_1424, n_1425, n_1426);
  xor g1503 (n_1427, n_536, n_537);
  xor g1504 (n_541, n_1427, n_538);
  nand g1505 (n_1428, n_536, n_537);
  nand g1506 (n_1429, n_538, n_537);
  nand g1507 (n_1430, n_536, n_538);
  nand g1508 (n_552, n_1428, n_1429, n_1430);
  xor g1509 (n_1431, n_539, n_540);
  xor g1510 (n_543, n_1431, n_541);
  nand g1511 (n_1432, n_539, n_540);
  nand g1512 (n_1433, n_541, n_540);
  nand g1513 (n_1434, n_539, n_541);
  nand g1514 (n_555, n_1432, n_1433, n_1434);
  xor g1515 (n_1435, n_542, n_543);
  xor g1516 (n_87, n_1435, n_544);
  nand g1517 (n_1436, n_542, n_543);
  nand g1518 (n_1437, n_544, n_543);
  nand g1519 (n_1438, n_542, n_544);
  nand g1520 (n_38, n_1436, n_1437, n_1438);
  xor g1521 (n_1439, A[12], A[13]);
  xor g1522 (n_547, n_1439, A[17]);
  nand g1525 (n_1442, A[12], A[17]);
  nand g1526 (n_558, n_766, n_1226, n_1442);
  nand g1532 (n_559, n_981, n_1333, n_1446);
  xor g1533 (n_1447, A[21], n_489);
  xor g1534 (n_550, n_1447, n_546);
  nand g1536 (n_1449, n_546, n_489);
  nand g1537 (n_1450, A[21], n_546);
  nand g1538 (n_562, n_1338, n_1449, n_1450);
  xor g1539 (n_1451, n_547, n_548);
  xor g1540 (n_553, n_1451, n_549);
  nand g1541 (n_1452, n_547, n_548);
  nand g1542 (n_1453, n_549, n_548);
  nand g1543 (n_1454, n_547, n_549);
  nand g1544 (n_563, n_1452, n_1453, n_1454);
  xor g1545 (n_1455, n_550, n_551);
  xor g1546 (n_554, n_1455, n_552);
  nand g1547 (n_1456, n_550, n_551);
  nand g1548 (n_1457, n_552, n_551);
  nand g1549 (n_1458, n_550, n_552);
  nand g1550 (n_566, n_1456, n_1457, n_1458);
  xor g1551 (n_1459, n_553, n_554);
  xor g1552 (n_86, n_1459, n_555);
  nand g1553 (n_1460, n_553, n_554);
  nand g1554 (n_1461, n_555, n_554);
  nand g1555 (n_1462, n_553, n_555);
  nand g1556 (n_37, n_1460, n_1461, n_1462);
  xor g1565 (n_1467, A[21], A[22]);
  nand g1570 (n_572, n_1065, n_1469, n_1470);
  xor g1571 (n_1471, n_558, n_559);
  xor g1572 (n_564, n_1471, n_440);
  nand g1573 (n_1472, n_558, n_559);
  nand g1574 (n_1473, n_440, n_559);
  nand g1575 (n_1474, n_558, n_440);
  nand g1576 (n_575, n_1472, n_1473, n_1474);
  xor g1577 (n_1475, n_561, n_562);
  xor g1578 (n_565, n_1475, n_563);
  nand g1579 (n_1476, n_561, n_562);
  nand g1580 (n_1477, n_563, n_562);
  nand g1581 (n_1478, n_561, n_563);
  nand g1582 (n_577, n_1476, n_1477, n_1478);
  xor g1583 (n_1479, n_564, n_565);
  xor g1584 (n_85, n_1479, n_566);
  nand g1585 (n_1480, n_564, n_565);
  nand g1586 (n_1481, n_566, n_565);
  nand g1587 (n_1482, n_564, n_566);
  nand g1588 (n_36, n_1480, n_1481, n_1482);
  xor g1592 (n_571, n_1259, A[18]);
  xor g1597 (n_1487, A[22], A[14]);
  xor g1598 (n_573, n_1487, A[23]);
  nand g1599 (n_1488, A[22], A[14]);
  nand g1600 (n_1489, A[23], A[14]);
  nand g1602 (n_581, n_1488, n_1489, n_1108);
  xor g1604 (n_574, n_1491, n_571);
  nand g1606 (n_1493, n_571, n_458);
  nand g1608 (n_584, n_1492, n_1493, n_1494);
  xor g1609 (n_1495, n_572, n_573);
  xor g1610 (n_576, n_1495, n_574);
  nand g1611 (n_1496, n_572, n_573);
  nand g1612 (n_1497, n_574, n_573);
  nand g1613 (n_1498, n_572, n_574);
  nand g1614 (n_586, n_1496, n_1497, n_1498);
  xor g1615 (n_1499, n_575, n_576);
  xor g1616 (n_84, n_1499, n_577);
  nand g1617 (n_1500, n_575, n_576);
  nand g1618 (n_1501, n_577, n_576);
  nand g1619 (n_1502, n_575, n_577);
  nand g1620 (n_35, n_1500, n_1501, n_1502);
  xor g1621 (n_1503, A[15], A[19]);
  xor g1622 (n_582, n_1503, A[16]);
  nand g1623 (n_1504, A[15], A[19]);
  nand g1625 (n_1506, A[15], A[16]);
  nand g1626 (n_587, n_1504, n_1148, n_1506);
  xor g1633 (n_1511, A[15], n_401);
  xor g1634 (n_583, n_1511, n_536);
  nand g1635 (n_1512, A[15], n_401);
  nand g1636 (n_1513, n_536, n_401);
  nand g1637 (n_1514, A[15], n_536);
  nand g1638 (n_591, n_1512, n_1513, n_1514);
  xor g1639 (n_1515, n_581, n_582);
  xor g1640 (n_585, n_1515, n_583);
  nand g1641 (n_1516, n_581, n_582);
  nand g1642 (n_1517, n_583, n_582);
  nand g1643 (n_1518, n_581, n_583);
  nand g1644 (n_593, n_1516, n_1517, n_1518);
  xor g1645 (n_1519, n_584, n_585);
  xor g1646 (n_83, n_1519, n_586);
  nand g1647 (n_1520, n_584, n_585);
  nand g1648 (n_1521, n_586, n_585);
  nand g1649 (n_1522, n_584, n_586);
  nand g1650 (n_34, n_1520, n_1521, n_1522);
  xor g1652 (n_588, n_1523, A[16]);
  nand g1656 (n_596, n_1524, n_1188, n_1446);
  xor g1657 (n_1527, A[20], A[21]);
  xor g1658 (n_590, n_1527, n_587);
  nand g1660 (n_1529, n_587, A[21]);
  nand g1661 (n_1530, A[20], n_587);
  nand g1662 (n_598, n_1021, n_1529, n_1530);
  xor g1663 (n_1531, n_588, n_549);
  xor g1664 (n_592, n_1531, n_590);
  nand g1665 (n_1532, n_588, n_549);
  nand g1666 (n_1533, n_590, n_549);
  nand g1667 (n_1534, n_588, n_590);
  nand g1668 (n_600, n_1532, n_1533, n_1534);
  xor g1669 (n_1535, n_591, n_592);
  xor g1670 (n_82, n_1535, n_593);
  nand g1671 (n_1536, n_591, n_592);
  nand g1672 (n_1537, n_593, n_592);
  nand g1673 (n_1538, n_591, n_593);
  nand g1674 (n_81, n_1536, n_1537, n_1538);
  xor g1677 (n_1539, A[17], A[21]);
  xor g1678 (n_597, n_1539, A[22]);
  nand g1679 (n_1540, A[17], A[21]);
  nand g1681 (n_1542, A[17], A[22]);
  nand g1682 (n_604, n_1540, n_1065, n_1542);
  xor g1684 (n_599, n_1543, n_597);
  nand g1686 (n_1545, n_597, n_596);
  nand g1688 (n_607, n_1544, n_1545, n_1546);
  xor g1689 (n_1547, n_598, n_599);
  xor g1690 (n_33, n_1547, n_600);
  nand g1691 (n_1548, n_598, n_599);
  nand g1692 (n_1549, n_600, n_599);
  nand g1693 (n_1550, n_598, n_600);
  nand g1694 (n_80, n_1548, n_1549, n_1550);
  nand g1706 (n_1557, n_604, A[18]);
  nand g1708 (n_612, n_1556, n_1557, n_1558);
  xor g1709 (n_1559, n_461, n_606);
  xor g1710 (n_32, n_1559, n_607);
  nand g1711 (n_1560, n_461, n_606);
  nand g1712 (n_1561, n_607, n_606);
  nand g1713 (n_1562, n_461, n_607);
  nand g1714 (n_31, n_1560, n_1561, n_1562);
  xor g1716 (n_609, n_1563, A[20]);
  nand g1720 (n_613, n_1564, n_1150, n_1333);
  xor g1721 (n_1567, A[23], A[19]);
  xor g1722 (n_611, n_1567, n_609);
  nand g1723 (n_1568, A[23], A[19]);
  nand g1724 (n_1569, n_609, A[19]);
  nand g1725 (n_1570, A[23], n_609);
  nand g1726 (n_615, n_1568, n_1569, n_1570);
  xor g1727 (n_1571, n_477, n_611);
  xor g1728 (n_79, n_1571, n_612);
  nand g1729 (n_1572, n_477, n_611);
  nand g1730 (n_1573, n_612, n_611);
  nand g1731 (n_1574, n_477, n_612);
  nand g1732 (n_30, n_1572, n_1573, n_1574);
  xor g1734 (n_614, n_1419, A[21]);
  nand g1738 (n_618, n_1333, n_1021, n_1066);
  xor g1739 (n_1579, n_613, n_614);
  xor g1740 (n_78, n_1579, n_615);
  nand g1741 (n_1580, n_613, n_614);
  nand g1742 (n_1581, n_615, n_614);
  nand g1743 (n_1582, n_613, n_615);
  nand g1744 (n_77, n_1580, n_1581, n_1582);
  nand g1751 (n_1586, A[22], n_618);
  nand g1752 (n_28, n_1584, n_1585, n_1586);
  nand g1759 (n_1590, A[23], A[21]);
  nand g1760 (n_27, n_1588, n_1589, n_1590);
  xor g1762 (n_75, n_1151, A[22]);
  nand g1766 (n_74, n_1152, n_1108, n_1064);
  nor g11 (n_1610, A[0], A[2]);
  nand g12 (n_1605, A[0], A[2]);
  nor g13 (n_1606, n_68, A[3]);
  nand g14 (n_1607, n_68, A[3]);
  nor g15 (n_1616, A[4], n_117);
  nand g16 (n_1611, A[4], n_117);
  nor g17 (n_1612, A[5], n_116);
  nand g18 (n_1613, A[5], n_116);
  nor g19 (n_1622, n_67, n_115);
  nand g20 (n_1617, n_67, n_115);
  nor g21 (n_1618, n_66, n_114);
  nand g22 (n_1619, n_66, n_114);
  nor g23 (n_1628, n_65, n_113);
  nand g24 (n_1623, n_65, n_113);
  nor g25 (n_1624, n_64, n_112);
  nand g26 (n_1625, n_64, n_112);
  nor g27 (n_1634, n_63, n_111);
  nand g28 (n_1629, n_63, n_111);
  nor g29 (n_1630, n_62, n_110);
  nand g30 (n_1631, n_62, n_110);
  nor g31 (n_1640, n_61, n_109);
  nand g32 (n_1635, n_61, n_109);
  nor g33 (n_1636, n_60, n_108);
  nand g34 (n_1637, n_60, n_108);
  nor g35 (n_1646, n_59, n_107);
  nand g36 (n_1641, n_59, n_107);
  nor g37 (n_1642, n_58, n_106);
  nand g38 (n_1643, n_58, n_106);
  nor g39 (n_1652, n_57, n_105);
  nand g40 (n_1647, n_57, n_105);
  nor g41 (n_1648, n_56, n_104);
  nand g42 (n_1649, n_56, n_104);
  nor g43 (n_1658, n_55, n_103);
  nand g44 (n_1653, n_55, n_103);
  nor g45 (n_1654, n_54, n_102);
  nand g46 (n_1655, n_54, n_102);
  nor g47 (n_1664, n_53, n_101);
  nand g48 (n_1659, n_53, n_101);
  nor g49 (n_1660, n_52, n_100);
  nand g50 (n_1661, n_52, n_100);
  nor g51 (n_1670, n_51, n_99);
  nand g52 (n_1665, n_51, n_99);
  nor g53 (n_1666, n_50, n_98);
  nand g54 (n_1667, n_50, n_98);
  nor g55 (n_1676, n_49, n_97);
  nand g56 (n_1671, n_49, n_97);
  nor g57 (n_1672, n_48, n_96);
  nand g58 (n_1673, n_48, n_96);
  nor g59 (n_1682, n_47, n_95);
  nand g60 (n_1677, n_47, n_95);
  nor g61 (n_1678, n_46, n_94);
  nand g62 (n_1679, n_46, n_94);
  nor g63 (n_1688, n_45, n_93);
  nand g64 (n_1683, n_45, n_93);
  nor g65 (n_1684, n_44, n_92);
  nand g66 (n_1685, n_44, n_92);
  nor g67 (n_1694, n_43, n_91);
  nand g68 (n_1689, n_43, n_91);
  nor g69 (n_1690, n_42, n_90);
  nand g70 (n_1691, n_42, n_90);
  nor g71 (n_1700, n_41, n_89);
  nand g72 (n_1695, n_41, n_89);
  nor g73 (n_1696, n_40, n_88);
  nand g74 (n_1697, n_40, n_88);
  nor g75 (n_1706, n_39, n_87);
  nand g76 (n_1701, n_39, n_87);
  nor g77 (n_1702, n_38, n_86);
  nand g78 (n_1703, n_38, n_86);
  nor g79 (n_1712, n_37, n_85);
  nand g80 (n_1707, n_37, n_85);
  nor g81 (n_1708, n_36, n_84);
  nand g82 (n_1709, n_36, n_84);
  nor g83 (n_1718, n_35, n_83);
  nand g84 (n_1713, n_35, n_83);
  nor g85 (n_1714, n_34, n_82);
  nand g86 (n_1715, n_34, n_82);
  nor g87 (n_1724, n_33, n_81);
  nand g88 (n_1719, n_33, n_81);
  nor g89 (n_1720, n_32, n_80);
  nand g90 (n_1721, n_32, n_80);
  nor g91 (n_1730, n_31, n_79);
  nand g92 (n_1725, n_31, n_79);
  nor g93 (n_1726, n_30, n_78);
  nand g94 (n_1727, n_30, n_78);
  nor g95 (n_1736, n_29, n_77);
  nand g96 (n_1731, n_29, n_77);
  nor g97 (n_1732, n_28, n_76);
  nand g98 (n_1733, n_28, n_76);
  nor g99 (n_1740, n_27, n_75);
  nand g100 (n_1737, n_27, n_75);
  nor g106 (n_1608, n_1605, n_1606);
  nor g110 (n_1614, n_1611, n_1612);
  nor g113 (n_1750, n_1616, n_1612);
  nor g114 (n_1620, n_1617, n_1618);
  nor g117 (n_1752, n_1622, n_1618);
  nor g118 (n_1626, n_1623, n_1624);
  nor g121 (n_1760, n_1628, n_1624);
  nor g122 (n_1632, n_1629, n_1630);
  nor g125 (n_1762, n_1634, n_1630);
  nor g126 (n_1638, n_1635, n_1636);
  nor g129 (n_1770, n_1640, n_1636);
  nor g130 (n_1644, n_1641, n_1642);
  nor g133 (n_1772, n_1646, n_1642);
  nor g134 (n_1650, n_1647, n_1648);
  nor g137 (n_1780, n_1652, n_1648);
  nor g138 (n_1656, n_1653, n_1654);
  nor g141 (n_1782, n_1658, n_1654);
  nor g142 (n_1662, n_1659, n_1660);
  nor g145 (n_1790, n_1664, n_1660);
  nor g146 (n_1668, n_1665, n_1666);
  nor g149 (n_1792, n_1670, n_1666);
  nor g150 (n_1674, n_1671, n_1672);
  nor g153 (n_1800, n_1676, n_1672);
  nor g154 (n_1680, n_1677, n_1678);
  nor g157 (n_1802, n_1682, n_1678);
  nor g158 (n_1686, n_1683, n_1684);
  nor g161 (n_1810, n_1688, n_1684);
  nor g162 (n_1692, n_1689, n_1690);
  nor g165 (n_1812, n_1694, n_1690);
  nor g166 (n_1698, n_1695, n_1696);
  nor g169 (n_1820, n_1700, n_1696);
  nor g170 (n_1704, n_1701, n_1702);
  nor g173 (n_1822, n_1706, n_1702);
  nor g174 (n_1710, n_1707, n_1708);
  nor g177 (n_1830, n_1712, n_1708);
  nor g178 (n_1716, n_1713, n_1714);
  nor g181 (n_1832, n_1718, n_1714);
  nor g182 (n_1722, n_1719, n_1720);
  nor g185 (n_1840, n_1724, n_1720);
  nor g186 (n_1728, n_1725, n_1726);
  nor g189 (n_1842, n_1730, n_1726);
  nor g190 (n_1734, n_1731, n_1732);
  nor g193 (n_1850, n_1736, n_1732);
  nor g203 (n_1748, n_1622, n_1747);
  nand g212 (n_1860, n_1750, n_1752);
  nor g213 (n_1758, n_1634, n_1757);
  nand g222 (n_1867, n_1760, n_1762);
  nor g223 (n_1768, n_1646, n_1767);
  nand g232 (n_1875, n_1770, n_1772);
  nor g233 (n_1778, n_1658, n_1777);
  nand g242 (n_1882, n_1780, n_1782);
  nor g243 (n_1788, n_1670, n_1787);
  nand g252 (n_1890, n_1790, n_1792);
  nor g253 (n_1798, n_1682, n_1797);
  nand g262 (n_1897, n_1800, n_1802);
  nor g263 (n_1808, n_1694, n_1807);
  nand g1776 (n_1905, n_1810, n_1812);
  nor g1777 (n_1818, n_1706, n_1817);
  nand g1786 (n_1912, n_1820, n_1822);
  nor g1787 (n_1828, n_1718, n_1827);
  nand g1796 (n_1920, n_1830, n_1832);
  nor g1797 (n_1838, n_1730, n_1837);
  nand g1806 (n_1927, n_1840, n_1842);
  nor g1807 (n_1848, n_1740, n_1847);
  nand g1814 (n_2131, n_1611, n_1854);
  nand g1816 (n_2133, n_1747, n_1855);
  nand g1819 (n_2136, n_1858, n_1859);
  nand g1822 (n_1935, n_1862, n_1863);
  nor g1823 (n_1865, n_1640, n_1864);
  nor g1826 (n_1945, n_1640, n_1867);
  nor g1832 (n_1873, n_1871, n_1864);
  nor g1835 (n_1951, n_1867, n_1871);
  nor g1836 (n_1877, n_1875, n_1864);
  nor g1839 (n_1954, n_1867, n_1875);
  nor g1840 (n_1880, n_1664, n_1879);
  nor g1843 (n_2034, n_1664, n_1882);
  nor g1849 (n_1888, n_1886, n_1879);
  nor g1852 (n_2040, n_1882, n_1886);
  nor g1853 (n_1892, n_1890, n_1879);
  nor g1856 (n_1960, n_1882, n_1890);
  nor g1857 (n_1895, n_1688, n_1894);
  nor g1860 (n_1973, n_1688, n_1897);
  nor g1866 (n_1903, n_1901, n_1894);
  nor g1869 (n_1983, n_1897, n_1901);
  nor g1870 (n_1907, n_1905, n_1894);
  nor g1873 (n_1988, n_1897, n_1905);
  nor g1874 (n_1910, n_1712, n_1909);
  nor g1877 (n_2086, n_1712, n_1912);
  nor g1883 (n_1918, n_1916, n_1909);
  nor g1886 (n_2092, n_1912, n_1916);
  nor g1887 (n_1922, n_1920, n_1909);
  nor g1890 (n_1996, n_1912, n_1920);
  nor g1891 (n_1925, n_1736, n_1924);
  nor g1894 (n_2009, n_1736, n_1927);
  nor g1900 (n_1933, n_1931, n_1924);
  nor g1903 (n_2019, n_1927, n_1931);
  nand g1906 (n_2140, n_1623, n_1937);
  nand g1907 (n_1938, n_1760, n_1935);
  nand g1908 (n_2142, n_1757, n_1938);
  nand g1911 (n_2145, n_1941, n_1942);
  nand g1914 (n_2148, n_1864, n_1944);
  nand g1915 (n_1947, n_1945, n_1935);
  nand g1916 (n_2151, n_1946, n_1947);
  nand g1917 (n_1950, n_1948, n_1935);
  nand g1918 (n_2153, n_1949, n_1950);
  nand g1919 (n_1953, n_1951, n_1935);
  nand g1920 (n_2156, n_1952, n_1953);
  nand g1921 (n_1956, n_1954, n_1935);
  nand g1922 (n_2024, n_1955, n_1956);
  nor g1923 (n_1958, n_1676, n_1957);
  nand g1932 (n_2048, n_1800, n_1960);
  nor g1933 (n_1967, n_1965, n_1957);
  nor g1938 (n_1970, n_1897, n_1957);
  nand g1947 (n_2060, n_1960, n_1973);
  nand g1952 (n_2064, n_1960, n_1978);
  nand g1957 (n_2068, n_1960, n_1983);
  nand g1962 (n_2072, n_1960, n_1988);
  nor g1963 (n_1994, n_1724, n_1993);
  nand g1972 (n_2100, n_1840, n_1996);
  nor g1973 (n_2003, n_2001, n_1993);
  nor g1978 (n_2006, n_1927, n_1993);
  nand g1987 (n_2112, n_1996, n_2009);
  nand g1992 (n_2116, n_1996, n_2014);
  nand g1997 (n_2120, n_1996, n_2019);
  nand g2000 (n_2160, n_1647, n_2026);
  nand g2001 (n_2027, n_1780, n_2024);
  nand g2002 (n_2162, n_1777, n_2027);
  nand g2005 (n_2165, n_2030, n_2031);
  nand g2008 (n_2168, n_1879, n_2033);
  nand g2009 (n_2036, n_2034, n_2024);
  nand g2010 (n_2171, n_2035, n_2036);
  nand g2011 (n_2039, n_2037, n_2024);
  nand g2012 (n_2173, n_2038, n_2039);
  nand g2013 (n_2042, n_2040, n_2024);
  nand g2014 (n_2176, n_2041, n_2042);
  nand g2015 (n_2043, n_1960, n_2024);
  nand g2016 (n_2178, n_1957, n_2043);
  nand g2019 (n_2181, n_2046, n_2047);
  nand g2022 (n_2183, n_2050, n_2051);
  nand g2025 (n_2186, n_2054, n_2055);
  nand g2028 (n_2189, n_2058, n_2059);
  nand g2031 (n_2192, n_2062, n_2063);
  nand g2034 (n_2194, n_2066, n_2067);
  nand g2037 (n_2197, n_2070, n_2071);
  nand g2040 (n_2076, n_2074, n_2075);
  nand g2043 (n_2201, n_1695, n_2078);
  nand g2044 (n_2079, n_1820, n_2076);
  nand g2045 (n_2203, n_1817, n_2079);
  nand g2048 (n_2206, n_2082, n_2083);
  nand g2051 (n_2209, n_1909, n_2085);
  nand g2052 (n_2088, n_2086, n_2076);
  nand g2053 (n_2212, n_2087, n_2088);
  nand g2054 (n_2091, n_2089, n_2076);
  nand g2055 (n_2214, n_2090, n_2091);
  nand g2056 (n_2094, n_2092, n_2076);
  nand g2057 (n_2217, n_2093, n_2094);
  nand g2058 (n_2095, n_1996, n_2076);
  nand g2059 (n_2219, n_1993, n_2095);
  nand g2062 (n_2222, n_2098, n_2099);
  nand g2065 (n_2224, n_2102, n_2103);
  nand g2068 (n_2227, n_2106, n_2107);
  nand g2071 (n_2230, n_2110, n_2111);
  nand g2074 (n_2233, n_2114, n_2115);
  nand g2077 (n_2235, n_2118, n_2119);
  nand g2080 (n_2238, n_2122, n_2123);
  xnor g2092 (Z[5], n_2131, n_2132);
  xnor g2094 (Z[6], n_2133, n_2134);
  xnor g2097 (Z[7], n_2136, n_2137);
  xnor g2099 (Z[8], n_1935, n_2138);
  xnor g2102 (Z[9], n_2140, n_2141);
  xnor g2104 (Z[10], n_2142, n_2143);
  xnor g2107 (Z[11], n_2145, n_2146);
  xnor g2110 (Z[12], n_2148, n_2149);
  xnor g2113 (Z[13], n_2151, n_2152);
  xnor g2115 (Z[14], n_2153, n_2154);
  xnor g2118 (Z[15], n_2156, n_2157);
  xnor g2120 (Z[16], n_2024, n_2158);
  xnor g2123 (Z[17], n_2160, n_2161);
  xnor g2125 (Z[18], n_2162, n_2163);
  xnor g2128 (Z[19], n_2165, n_2166);
  xnor g2131 (Z[20], n_2168, n_2169);
  xnor g2134 (Z[21], n_2171, n_2172);
  xnor g2136 (Z[22], n_2173, n_2174);
  xnor g2139 (Z[23], n_2176, n_2177);
  xnor g2141 (Z[24], n_2178, n_2179);
  xnor g2144 (Z[25], n_2181, n_2182);
  xnor g2146 (Z[26], n_2183, n_2184);
  xnor g2149 (Z[27], n_2186, n_2187);
  xnor g2152 (Z[28], n_2189, n_2190);
  xnor g2155 (Z[29], n_2192, n_2193);
  xnor g2157 (Z[30], n_2194, n_2195);
  xnor g2160 (Z[31], n_2197, n_2198);
  xnor g2162 (Z[32], n_2076, n_2199);
  xnor g2165 (Z[33], n_2201, n_2202);
  xnor g2167 (Z[34], n_2203, n_2204);
  xnor g2170 (Z[35], n_2206, n_2207);
  xnor g2173 (Z[36], n_2209, n_2210);
  xnor g2176 (Z[37], n_2212, n_2213);
  xnor g2178 (Z[38], n_2214, n_2215);
  xnor g2181 (Z[39], n_2217, n_2218);
  xnor g2183 (Z[40], n_2219, n_2220);
  xnor g2186 (Z[41], n_2222, n_2223);
  xnor g2188 (Z[42], n_2224, n_2225);
  xnor g2191 (Z[43], n_2227, n_2228);
  xnor g2194 (Z[44], n_2230, n_2231);
  xnor g2197 (Z[45], n_2233, n_2234);
  xnor g2199 (Z[46], n_2235, n_2236);
  xnor g2202 (Z[47], n_2238, n_2239);
  or g2216 (n_1045, A[1], wc);
  not gc (wc, n_171);
  or g2217 (n_1046, A[1], wc0);
  not gc0 (wc0, A[2]);
  xnor g2218 (n_1063, A[24], A[22]);
  or g2219 (n_1064, wc1, A[24]);
  not gc1 (wc1, A[22]);
  or g2220 (n_1066, wc2, A[24]);
  not gc2 (wc2, A[21]);
  or g2221 (n_1089, A[2], wc3);
  not gc3 (wc3, A[3]);
  or g2222 (n_1090, wc4, A[2]);
  not gc4 (wc4, A[1]);
  xnor g2223 (n_1151, A[24], A[23]);
  or g2224 (n_1152, wc5, A[24]);
  not gc5 (wc5, A[23]);
  xnor g2225 (n_1191, A[24], A[21]);
  xnor g2226 (n_1215, A[6], A[5]);
  or g2227 (n_1216, A[5], wc6);
  not gc6 (wc6, A[6]);
  or g2228 (n_1217, A[5], wc7);
  not gc7 (wc7, A[9]);
  or g2229 (n_1253, wc8, A[6]);
  not gc8 (wc8, A[5]);
  or g2230 (n_1254, A[6], wc9);
  not gc9 (wc9, A[7]);
  or g2231 (n_1333, wc10, A[24]);
  not gc10 (wc10, A[20]);
  xnor g2232 (n_1359, A[18], A[10]);
  or g2233 (n_1360, A[10], wc11);
  not gc11 (wc11, A[18]);
  or g2234 (n_1361, A[10], wc12);
  not gc12 (wc12, A[17]);
  xnor g2235 (n_1387, A[19], A[11]);
  or g2236 (n_1388, A[11], wc13);
  not gc13 (wc13, A[19]);
  or g2237 (n_1389, A[11], wc14);
  not gc14 (wc14, A[18]);
  xnor g2239 (n_1419, A[24], A[20]);
  xnor g2240 (n_548, n_1019, A[24]);
  or g2241 (n_1446, wc15, A[24]);
  not gc15 (wc15, A[16]);
  xnor g2242 (n_561, n_1467, A[14]);
  or g2243 (n_1469, A[14], wc16);
  not gc16 (wc16, A[22]);
  or g2244 (n_1470, A[14], wc17);
  not gc17 (wc17, A[21]);
  xnor g2245 (n_1523, A[24], A[17]);
  or g2246 (n_1524, wc18, A[24]);
  not gc18 (wc18, A[17]);
  or g2248 (n_1556, wc19, A[19]);
  not gc19 (wc19, A[18]);
  xnor g2249 (n_1563, A[24], A[19]);
  or g2250 (n_1564, wc20, A[24]);
  not gc20 (wc20, A[19]);
  or g2252 (n_1584, A[21], wc21);
  not gc21 (wc21, A[22]);
  or g2254 (n_1588, A[22], wc22);
  not gc22 (wc22, A[23]);
  or g2255 (n_1589, wc23, A[22]);
  not gc23 (wc23, A[21]);
  xnor g2256 (n_350, n_1043, A[1]);
  xnor g2257 (n_373, n_1087, A[2]);
  or g2258 (n_1194, A[24], wc24);
  not gc24 (wc24, n_416);
  xnor g2259 (n_454, n_1251, A[6]);
  xnor g2260 (n_537, n_1387, A[16]);
  xnor g2261 (n_1491, n_458, A[15]);
  or g2262 (n_1492, A[15], wc25);
  not gc25 (wc25, n_458);
  or g2263 (n_1494, A[15], wc26);
  not gc26 (wc26, n_571);
  or g2264 (n_1546, A[18], wc27);
  not gc27 (wc27, n_597);
  xnor g2265 (n_606, n_947, n_604);
  or g2266 (n_1558, A[19], wc28);
  not gc28 (wc28, n_604);
  xnor g2267 (n_76, n_1107, A[21]);
  or g2269 (n_2125, wc29, n_1610);
  not gc29 (wc29, n_1605);
  xnor g2270 (n_1299, n_471, A[24]);
  or g2271 (n_1300, A[24], wc30);
  not gc30 (wc30, n_471);
  or g2272 (n_1334, A[24], wc31);
  not gc31 (wc31, n_487);
  xnor g2273 (n_1543, n_596, A[18]);
  or g2274 (n_1544, A[18], wc32);
  not gc32 (wc32, n_596);
  xnor g2275 (n_29, n_1467, n_618);
  or g2276 (n_1585, A[21], wc33);
  not gc33 (wc33, n_618);
  and g2277 (n_1745, wc34, n_1607);
  not gc34 (wc34, n_1608);
  or g2278 (n_2128, wc35, n_1606);
  not gc35 (wc35, n_1607);
  xnor g2279 (n_491, n_1331, A[24]);
  and g2280 (n_1738, wc36, n_74);
  not gc36 (wc36, A[24]);
  or g2281 (n_1739, wc37, n_74);
  not gc37 (wc37, A[24]);
  not g2282 (Z[2], n_2125);
  or g2283 (n_2129, wc38, n_1616);
  not gc38 (wc38, n_1611);
  or g2286 (n_2236, wc39, n_1740);
  not gc39 (wc39, n_1737);
  and g2287 (n_1747, wc40, n_1613);
  not gc40 (wc40, n_1614);
  or g2288 (n_1854, n_1616, n_1745);
  or g2289 (n_1855, n_1745, wc41);
  not gc41 (wc41, n_1750);
  xor g2290 (Z[3], n_1605, n_2128);
  xor g2291 (Z[4], n_1745, n_2129);
  or g2292 (n_2132, wc42, n_1612);
  not gc42 (wc42, n_1613);
  or g2293 (n_2239, wc43, n_1738);
  not gc43 (wc43, n_1739);
  or g2294 (n_1154, A[24], wc44);
  not gc44 (wc44, n_397);
  and g2295 (n_1754, wc45, n_1619);
  not gc45 (wc45, n_1620);
  or g2296 (n_1856, wc46, n_1622);
  not gc46 (wc46, n_1750);
  or g2297 (n_2134, wc47, n_1622);
  not gc47 (wc47, n_1617);
  or g2298 (n_2137, wc48, n_1618);
  not gc48 (wc48, n_1619);
  or g2299 (n_2138, wc49, n_1628);
  not gc49 (wc49, n_1623);
  or g2300 (n_2234, wc50, n_1732);
  not gc50 (wc50, n_1733);
  and g2301 (n_1858, wc51, n_1617);
  not gc51 (wc51, n_1748);
  and g2302 (n_1755, wc52, n_1752);
  not gc52 (wc52, n_1747);
  or g2303 (n_2228, wc53, n_1726);
  not gc53 (wc53, n_1727);
  and g2304 (n_1757, wc54, n_1625);
  not gc54 (wc54, n_1626);
  and g2305 (n_1844, wc55, n_1727);
  not gc55 (wc55, n_1728);
  and g2306 (n_1847, wc56, n_1733);
  not gc56 (wc56, n_1734);
  and g2307 (n_1862, wc57, n_1754);
  not gc57 (wc57, n_1755);
  or g2308 (n_1931, wc58, n_1740);
  not gc58 (wc58, n_1850);
  or g2309 (n_1859, n_1745, n_1856);
  or g2310 (n_1863, n_1860, n_1745);
  or g2311 (n_2141, wc59, n_1624);
  not gc59 (wc59, n_1625);
  or g2312 (n_2223, wc60, n_1720);
  not gc60 (wc60, n_1721);
  or g2313 (n_2225, wc61, n_1730);
  not gc61 (wc61, n_1725);
  or g2314 (n_2231, wc62, n_1736);
  not gc62 (wc62, n_1731);
  and g2315 (n_1837, wc63, n_1721);
  not gc63 (wc63, n_1722);
  or g2316 (n_1939, wc64, n_1634);
  not gc64 (wc64, n_1760);
  or g2317 (n_2001, wc65, n_1730);
  not gc65 (wc65, n_1840);
  or g2318 (n_2143, wc66, n_1634);
  not gc66 (wc66, n_1629);
  or g2319 (n_2218, wc67, n_1714);
  not gc67 (wc67, n_1715);
  or g2320 (n_2220, wc68, n_1724);
  not gc68 (wc68, n_1719);
  and g2321 (n_1764, wc69, n_1631);
  not gc69 (wc69, n_1632);
  and g2322 (n_1767, wc70, n_1637);
  not gc70 (wc70, n_1638);
  and g2323 (n_1827, wc71, n_1709);
  not gc71 (wc71, n_1710);
  and g2324 (n_1834, wc72, n_1715);
  not gc72 (wc72, n_1716);
  and g2325 (n_1941, wc73, n_1629);
  not gc73 (wc73, n_1758);
  or g2326 (n_1916, wc74, n_1718);
  not gc74 (wc74, n_1830);
  and g2327 (n_1845, wc75, n_1842);
  not gc75 (wc75, n_1837);
  and g2328 (n_1932, wc76, n_1737);
  not gc76 (wc76, n_1848);
  and g2329 (n_2014, wc77, n_1850);
  not gc77 (wc77, n_1927);
  or g2330 (n_1937, wc78, n_1628);
  not gc78 (wc78, n_1935);
  or g2331 (n_2146, wc79, n_1630);
  not gc79 (wc79, n_1631);
  or g2332 (n_2149, wc80, n_1640);
  not gc80 (wc80, n_1635);
  or g2333 (n_2152, wc81, n_1636);
  not gc81 (wc81, n_1637);
  or g2334 (n_2210, wc82, n_1712);
  not gc82 (wc82, n_1707);
  or g2335 (n_2213, wc83, n_1708);
  not gc83 (wc83, n_1709);
  or g2336 (n_2215, wc84, n_1718);
  not gc84 (wc84, n_1713);
  and g2337 (n_1765, wc85, n_1762);
  not gc85 (wc85, n_1757);
  or g2338 (n_1871, wc86, n_1646);
  not gc86 (wc86, n_1770);
  and g2339 (n_1835, wc87, n_1832);
  not gc87 (wc87, n_1827);
  and g2340 (n_2002, wc88, n_1725);
  not gc88 (wc88, n_1838);
  and g2341 (n_1924, wc89, n_1844);
  not gc89 (wc89, n_1845);
  and g2342 (n_1948, wc90, n_1770);
  not gc90 (wc90, n_1867);
  or g2343 (n_1942, n_1939, wc91);
  not gc91 (wc91, n_1935);
  or g2344 (n_2154, wc92, n_1646);
  not gc92 (wc92, n_1641);
  and g2345 (n_1774, wc93, n_1643);
  not gc93 (wc93, n_1644);
  and g2346 (n_1824, wc94, n_1703);
  not gc94 (wc94, n_1704);
  and g2347 (n_1864, wc95, n_1764);
  not gc95 (wc95, n_1765);
  and g2348 (n_1872, wc96, n_1641);
  not gc96 (wc96, n_1768);
  and g2349 (n_1917, wc97, n_1713);
  not gc97 (wc97, n_1828);
  and g2350 (n_1921, wc98, n_1834);
  not gc98 (wc98, n_1835);
  and g2351 (n_1929, wc99, n_1850);
  not gc99 (wc99, n_1924);
  or g2352 (n_1944, wc100, n_1867);
  not gc100 (wc100, n_1935);
  or g2353 (n_2157, wc101, n_1642);
  not gc101 (wc101, n_1643);
  or g2354 (n_2202, wc102, n_1696);
  not gc102 (wc102, n_1697);
  or g2355 (n_2204, wc103, n_1706);
  not gc103 (wc103, n_1701);
  or g2356 (n_2207, wc104, n_1702);
  not gc104 (wc104, n_1703);
  and g2357 (n_1775, wc105, n_1772);
  not gc105 (wc105, n_1767);
  and g2358 (n_1869, wc106, n_1770);
  not gc106 (wc106, n_1864);
  and g2359 (n_2011, wc107, n_1731);
  not gc107 (wc107, n_1925);
  and g2360 (n_2016, wc108, n_1847);
  not gc108 (wc108, n_1929);
  and g2361 (n_2021, n_1932, wc109);
  not gc109 (wc109, n_1933);
  or g2362 (n_2158, wc110, n_1652);
  not gc110 (wc110, n_1647);
  or g2363 (n_2166, wc111, n_1654);
  not gc111 (wc111, n_1655);
  and g2364 (n_1777, wc112, n_1649);
  not gc112 (wc112, n_1650);
  and g2365 (n_1784, wc113, n_1655);
  not gc113 (wc113, n_1656);
  and g2366 (n_1876, wc114, n_1774);
  not gc114 (wc114, n_1775);
  or g2367 (n_2028, wc115, n_1658);
  not gc115 (wc115, n_1780);
  and g2368 (n_1946, wc116, n_1635);
  not gc116 (wc116, n_1865);
  and g2369 (n_1949, wc117, n_1767);
  not gc117 (wc117, n_1869);
  and g2370 (n_1952, n_1872, wc118);
  not gc118 (wc118, n_1873);
  or g2371 (n_2161, wc119, n_1648);
  not gc119 (wc119, n_1649);
  or g2372 (n_2163, wc120, n_1658);
  not gc120 (wc120, n_1653);
  or g2373 (n_2169, wc121, n_1664);
  not gc121 (wc121, n_1659);
  and g2374 (n_1787, wc122, n_1661);
  not gc122 (wc122, n_1662);
  and g2375 (n_1785, wc123, n_1782);
  not gc123 (wc123, n_1777);
  or g2376 (n_2172, wc124, n_1660);
  not gc124 (wc124, n_1661);
  and g2377 (n_1794, wc125, n_1667);
  not gc125 (wc125, n_1668);
  and g2378 (n_1797, wc126, n_1673);
  not gc126 (wc126, n_1674);
  and g2379 (n_1804, wc127, n_1679);
  not gc127 (wc127, n_1680);
  and g2380 (n_1807, wc128, n_1685);
  not gc128 (wc128, n_1686);
  and g2381 (n_1814, wc129, n_1691);
  not gc129 (wc129, n_1692);
  and g2382 (n_1817, wc130, n_1697);
  not gc130 (wc130, n_1698);
  and g2383 (n_2030, wc131, n_1653);
  not gc131 (wc131, n_1778);
  and g2384 (n_1879, wc132, n_1784);
  not gc132 (wc132, n_1785);
  or g2385 (n_1886, wc133, n_1670);
  not gc133 (wc133, n_1790);
  or g2386 (n_1965, wc134, n_1682);
  not gc134 (wc134, n_1800);
  or g2387 (n_1901, wc135, n_1694);
  not gc135 (wc135, n_1810);
  or g2388 (n_2080, wc136, n_1706);
  not gc136 (wc136, n_1820);
  and g2389 (n_1955, n_1876, wc137);
  not gc137 (wc137, n_1877);
  and g2390 (n_2037, wc138, n_1790);
  not gc138 (wc138, n_1882);
  or g2391 (n_2174, wc139, n_1670);
  not gc139 (wc139, n_1665);
  or g2392 (n_2177, wc140, n_1666);
  not gc140 (wc140, n_1667);
  or g2393 (n_2179, wc141, n_1676);
  not gc141 (wc141, n_1671);
  or g2394 (n_2182, wc142, n_1672);
  not gc142 (wc142, n_1673);
  or g2395 (n_2184, wc143, n_1682);
  not gc143 (wc143, n_1677);
  or g2396 (n_2187, wc144, n_1678);
  not gc144 (wc144, n_1679);
  or g2397 (n_2190, wc145, n_1688);
  not gc145 (wc145, n_1683);
  or g2398 (n_2193, wc146, n_1684);
  not gc146 (wc146, n_1685);
  or g2399 (n_2195, wc147, n_1694);
  not gc147 (wc147, n_1689);
  or g2400 (n_2198, wc148, n_1690);
  not gc148 (wc148, n_1691);
  or g2401 (n_2199, wc149, n_1700);
  not gc149 (wc149, n_1695);
  and g2402 (n_1887, wc150, n_1665);
  not gc150 (wc150, n_1788);
  and g2403 (n_1795, wc151, n_1792);
  not gc151 (wc151, n_1787);
  and g2404 (n_1805, wc152, n_1802);
  not gc152 (wc152, n_1797);
  and g2405 (n_1815, wc153, n_1812);
  not gc153 (wc153, n_1807);
  and g2406 (n_1825, wc154, n_1822);
  not gc154 (wc154, n_1817);
  and g2407 (n_1884, wc155, n_1790);
  not gc155 (wc155, n_1879);
  and g2408 (n_1978, wc156, n_1810);
  not gc156 (wc156, n_1897);
  and g2409 (n_2089, wc157, n_1830);
  not gc157 (wc157, n_1912);
  and g2410 (n_1891, wc158, n_1794);
  not gc158 (wc158, n_1795);
  and g2411 (n_1966, wc159, n_1677);
  not gc159 (wc159, n_1798);
  and g2412 (n_1894, wc160, n_1804);
  not gc160 (wc160, n_1805);
  and g2413 (n_1902, wc161, n_1689);
  not gc161 (wc161, n_1808);
  and g2414 (n_1906, wc162, n_1814);
  not gc162 (wc162, n_1815);
  and g2415 (n_2082, wc163, n_1701);
  not gc163 (wc163, n_1818);
  and g2416 (n_1909, wc164, n_1824);
  not gc164 (wc164, n_1825);
  and g2417 (n_2035, wc165, n_1659);
  not gc165 (wc165, n_1880);
  and g2418 (n_2038, wc166, n_1787);
  not gc166 (wc166, n_1884);
  or g2419 (n_2044, wc167, n_1676);
  not gc167 (wc167, n_1960);
  or g2420 (n_2052, n_1965, wc168);
  not gc168 (wc168, n_1960);
  or g2421 (n_2056, wc169, n_1897);
  not gc169 (wc169, n_1960);
  or g2422 (n_2096, wc170, n_1724);
  not gc170 (wc170, n_1996);
  or g2423 (n_2104, n_2001, wc171);
  not gc171 (wc171, n_1996);
  or g2424 (n_2108, wc172, n_1927);
  not gc172 (wc172, n_1996);
  or g2425 (n_2026, wc173, n_1652);
  not gc173 (wc173, n_2024);
  or g2426 (n_2031, n_2028, wc174);
  not gc174 (wc174, n_2024);
  or g2427 (n_2033, wc175, n_1882);
  not gc175 (wc175, n_2024);
  and g2428 (n_2041, n_1887, wc176);
  not gc176 (wc176, n_1888);
  and g2429 (n_1899, wc177, n_1810);
  not gc177 (wc177, n_1894);
  and g2430 (n_1914, wc178, n_1830);
  not gc178 (wc178, n_1909);
  and g2431 (n_1957, n_1891, wc179);
  not gc179 (wc179, n_1892);
  and g2432 (n_1975, wc180, n_1683);
  not gc180 (wc180, n_1895);
  and g2433 (n_1980, wc181, n_1807);
  not gc181 (wc181, n_1899);
  and g2434 (n_1985, n_1902, wc182);
  not gc182 (wc182, n_1903);
  and g2435 (n_1990, n_1906, wc183);
  not gc183 (wc183, n_1907);
  and g2436 (n_2087, wc184, n_1707);
  not gc184 (wc184, n_1910);
  and g2437 (n_2090, wc185, n_1827);
  not gc185 (wc185, n_1914);
  and g2438 (n_2093, n_1917, wc186);
  not gc186 (wc186, n_1918);
  and g2439 (n_1993, n_1921, wc187);
  not gc187 (wc187, n_1922);
  or g2440 (n_2047, n_2044, wc188);
  not gc188 (wc188, n_2024);
  or g2441 (n_2051, n_2048, wc189);
  not gc189 (wc189, n_2024);
  or g2442 (n_2055, n_2052, wc190);
  not gc190 (wc190, n_2024);
  or g2443 (n_2059, n_2056, wc191);
  not gc191 (wc191, n_2024);
  or g2444 (n_2063, n_2060, wc192);
  not gc192 (wc192, n_2024);
  or g2445 (n_2067, n_2064, wc193);
  not gc193 (wc193, n_2024);
  or g2446 (n_2071, n_2068, wc194);
  not gc194 (wc194, n_2024);
  or g2447 (n_2075, n_2072, wc195);
  not gc195 (wc195, n_2024);
  and g2448 (n_1963, wc196, n_1800);
  not gc196 (wc196, n_1957);
  and g2449 (n_1976, wc197, n_1973);
  not gc197 (wc197, n_1957);
  and g2450 (n_1981, wc198, n_1978);
  not gc198 (wc198, n_1957);
  and g2451 (n_1986, wc199, n_1983);
  not gc199 (wc199, n_1957);
  and g2452 (n_1991, wc200, n_1988);
  not gc200 (wc200, n_1957);
  and g2453 (n_1999, wc201, n_1840);
  not gc201 (wc201, n_1993);
  and g2454 (n_2012, wc202, n_2009);
  not gc202 (wc202, n_1993);
  and g2455 (n_2017, wc203, n_2014);
  not gc203 (wc203, n_1993);
  and g2456 (n_2022, wc204, n_2019);
  not gc204 (wc204, n_1993);
  and g2457 (n_2046, wc205, n_1671);
  not gc205 (wc205, n_1958);
  and g2458 (n_2050, wc206, n_1797);
  not gc206 (wc206, n_1963);
  and g2459 (n_2054, n_1966, wc207);
  not gc207 (wc207, n_1967);
  and g2460 (n_2058, n_1894, wc208);
  not gc208 (wc208, n_1970);
  and g2461 (n_2062, wc209, n_1975);
  not gc209 (wc209, n_1976);
  and g2462 (n_2066, wc210, n_1980);
  not gc210 (wc210, n_1981);
  and g2463 (n_2070, wc211, n_1985);
  not gc211 (wc211, n_1986);
  and g2464 (n_2074, wc212, n_1990);
  not gc212 (wc212, n_1991);
  and g2465 (n_2098, wc213, n_1719);
  not gc213 (wc213, n_1994);
  and g2466 (n_2102, wc214, n_1837);
  not gc214 (wc214, n_1999);
  and g2467 (n_2106, n_2002, wc215);
  not gc215 (wc215, n_2003);
  and g2468 (n_2110, n_1924, wc216);
  not gc216 (wc216, n_2006);
  and g2469 (n_2114, wc217, n_2011);
  not gc217 (wc217, n_2012);
  and g2470 (n_2118, wc218, n_2016);
  not gc218 (wc218, n_2017);
  and g2471 (n_2122, wc219, n_2021);
  not gc219 (wc219, n_2022);
  or g2472 (n_2078, wc220, n_1700);
  not gc220 (wc220, n_2076);
  or g2473 (n_2083, n_2080, wc221);
  not gc221 (wc221, n_2076);
  or g2474 (n_2085, wc222, n_1912);
  not gc222 (wc222, n_2076);
  or g2475 (n_2099, n_2096, wc223);
  not gc223 (wc223, n_2076);
  or g2476 (n_2103, wc224, n_2100);
  not gc224 (wc224, n_2076);
  or g2477 (n_2107, n_2104, wc225);
  not gc225 (wc225, n_2076);
  or g2478 (n_2111, n_2108, wc226);
  not gc226 (wc226, n_2076);
  or g2479 (n_2115, wc227, n_2112);
  not gc227 (wc227, n_2076);
  or g2480 (n_2119, wc228, n_2116);
  not gc228 (wc228, n_2076);
  or g2481 (n_2123, wc229, n_2120);
  not gc229 (wc229, n_2076);
endmodule

module mult_signed_const_5486_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_5486_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_5753_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_171, n_172, n_173, n_176, n_178;
  wire n_179, n_180, n_183, n_184, n_187, n_188, n_189, n_193;
  wire n_195, n_196, n_200, n_201, n_202, n_203, n_204, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_215, n_217, n_218;
  wire n_219, n_220, n_221, n_223, n_224, n_225, n_226, n_227;
  wire n_228, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252;
  wire n_257, n_258, n_260, n_261, n_262, n_263, n_266, n_268;
  wire n_269, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_278, n_281, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_299, n_300;
  wire n_301, n_302, n_303, n_304, n_305, n_306, n_307, n_308;
  wire n_309, n_310, n_315, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_333, n_334;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_350, n_352, n_354, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_431, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_498, n_499, n_500, n_501, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_516, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_530, n_531, n_533, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550;
  wire n_551, n_552, n_553, n_554, n_555, n_558, n_559, n_560;
  wire n_561, n_562, n_563, n_564, n_565, n_566, n_570, n_571;
  wire n_572, n_573, n_574, n_575, n_576, n_577, n_579, n_580;
  wire n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_589;
  wire n_590, n_591, n_592, n_593, n_597, n_599, n_600, n_605;
  wire n_606, n_607, n_609, n_610, n_611, n_612, n_613, n_615;
  wire n_623, n_624, n_625, n_626, n_627, n_628, n_629, n_630;
  wire n_631, n_632, n_633, n_634, n_635, n_636, n_637, n_638;
  wire n_639, n_640, n_641, n_642, n_643, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_654, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_666, n_669, n_670, n_671;
  wire n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_685;
  wire n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693;
  wire n_694, n_699, n_700, n_701, n_703, n_704, n_705, n_706;
  wire n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714;
  wire n_719, n_723, n_724, n_725, n_726, n_727, n_728, n_729;
  wire n_730, n_731, n_732, n_733, n_734, n_737, n_738, n_739;
  wire n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747;
  wire n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_763;
  wire n_764, n_765, n_767, n_768, n_769, n_770, n_771, n_772;
  wire n_773, n_774, n_775, n_776, n_777, n_778, n_789, n_790;
  wire n_791, n_792, n_793, n_794, n_795, n_796, n_797, n_798;
  wire n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_806;
  wire n_815, n_816, n_818, n_819, n_820, n_821, n_822, n_823;
  wire n_824, n_825, n_826, n_827, n_828, n_829, n_830, n_831;
  wire n_832, n_833, n_834, n_841, n_842, n_847, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_865, n_866, n_867;
  wire n_868, n_869, n_870, n_873, n_875, n_876, n_877, n_878;
  wire n_879, n_880, n_881, n_882, n_883, n_884, n_885, n_886;
  wire n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_894;
  wire n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910;
  wire n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918;
  wire n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926;
  wire n_927, n_928, n_929, n_930, n_939, n_945, n_946, n_947;
  wire n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955;
  wire n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963;
  wire n_964, n_965, n_966, n_973, n_974, n_975, n_976, n_978;
  wire n_979, n_980, n_982, n_983, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1017;
  wire n_1018, n_1019, n_1020, n_1022, n_1023, n_1024, n_1025, n_1026;
  wire n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034;
  wire n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042;
  wire n_1043, n_1045, n_1046, n_1047, n_1048, n_1049, n_1051, n_1052;
  wire n_1053, n_1054, n_1055, n_1057, n_1058, n_1059, n_1060, n_1061;
  wire n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069;
  wire n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077;
  wire n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085;
  wire n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093;
  wire n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101;
  wire n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109;
  wire n_1110, n_1111, n_1112, n_1113, n_1115, n_1116, n_1117, n_1118;
  wire n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126;
  wire n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1135;
  wire n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1143, n_1144;
  wire n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152;
  wire n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160;
  wire n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168;
  wire n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1177;
  wire n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185;
  wire n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193;
  wire n_1194, n_1195, n_1196, n_1199, n_1200, n_1201, n_1202, n_1203;
  wire n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211;
  wire n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219;
  wire n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227;
  wire n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235;
  wire n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243;
  wire n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251;
  wire n_1253, n_1254, n_1255, n_1257, n_1258, n_1259, n_1260, n_1261;
  wire n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270;
  wire n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278;
  wire n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286;
  wire n_1289, n_1291, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298;
  wire n_1299, n_1300, n_1302, n_1303, n_1304, n_1306, n_1307, n_1308;
  wire n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316;
  wire n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1326;
  wire n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1334, n_1335;
  wire n_1336, n_1337, n_1338, n_1341, n_1342, n_1343, n_1344, n_1345;
  wire n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353;
  wire n_1354, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362;
  wire n_1363, n_1364, n_1365, n_1367, n_1368, n_1369, n_1370, n_1371;
  wire n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379;
  wire n_1380, n_1381, n_1382, n_1385, n_1387, n_1389, n_1390, n_1391;
  wire n_1393, n_1394, n_1395, n_1396, n_1397, n_1399, n_1400, n_1401;
  wire n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409;
  wire n_1410, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421;
  wire n_1422, n_1423, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430;
  wire n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438;
  wire n_1439, n_1441, n_1442, n_1446, n_1447, n_1449, n_1450, n_1451;
  wire n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1460, n_1461, n_1462, n_1464, n_1465, n_1467, n_1470, n_1471;
  wire n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479;
  wire n_1480, n_1481, n_1482, n_1486, n_1489, n_1491, n_1492, n_1493;
  wire n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501;
  wire n_1502, n_1505, n_1507, n_1508, n_1509, n_1513, n_1514, n_1515;
  wire n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1529;
  wire n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537;
  wire n_1538, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1551, n_1554, n_1556, n_1557, n_1558, n_1559, n_1560;
  wire n_1561, n_1562, n_1563, n_1566, n_1567, n_1568, n_1569, n_1570;
  wire n_1571, n_1572, n_1573, n_1574, n_1579, n_1580, n_1581, n_1582;
  wire n_1584, n_1585, n_1586, n_1588, n_1589, n_1591, n_1592, n_1594;
  wire n_1605, n_1606, n_1607, n_1608, n_1610, n_1611, n_1612, n_1613;
  wire n_1614, n_1616, n_1617, n_1618, n_1619, n_1620, n_1622, n_1623;
  wire n_1624, n_1625, n_1626, n_1628, n_1629, n_1630, n_1631, n_1632;
  wire n_1634, n_1635, n_1636, n_1637, n_1638, n_1640, n_1641, n_1642;
  wire n_1643, n_1644, n_1646, n_1647, n_1648, n_1649, n_1650, n_1652;
  wire n_1653, n_1654, n_1655, n_1656, n_1658, n_1659, n_1660, n_1661;
  wire n_1662, n_1664, n_1665, n_1666, n_1667, n_1668, n_1670, n_1671;
  wire n_1672, n_1673, n_1674, n_1676, n_1677, n_1678, n_1679, n_1680;
  wire n_1682, n_1683, n_1684, n_1685, n_1686, n_1688, n_1689, n_1690;
  wire n_1691, n_1692, n_1694, n_1695, n_1696, n_1697, n_1698, n_1700;
  wire n_1701, n_1702, n_1703, n_1704, n_1706, n_1707, n_1708, n_1709;
  wire n_1710, n_1712, n_1713, n_1714, n_1715, n_1716, n_1718, n_1719;
  wire n_1720, n_1721, n_1722, n_1724, n_1725, n_1726, n_1727, n_1728;
  wire n_1730, n_1731, n_1732, n_1733, n_1734, n_1736, n_1737, n_1738;
  wire n_1739, n_1740, n_1745, n_1747, n_1748, n_1750, n_1752, n_1754;
  wire n_1755, n_1757, n_1758, n_1760, n_1762, n_1764, n_1765, n_1767;
  wire n_1768, n_1770, n_1772, n_1774, n_1775, n_1777, n_1778, n_1780;
  wire n_1782, n_1784, n_1785, n_1787, n_1788, n_1790, n_1792, n_1794;
  wire n_1795, n_1797, n_1798, n_1800, n_1802, n_1804, n_1805, n_1807;
  wire n_1808, n_1810, n_1812, n_1814, n_1815, n_1817, n_1818, n_1820;
  wire n_1822, n_1824, n_1825, n_1827, n_1828, n_1830, n_1832, n_1834;
  wire n_1835, n_1837, n_1838, n_1840, n_1842, n_1844, n_1845, n_1847;
  wire n_1848, n_1850, n_1854, n_1855, n_1856, n_1858, n_1859, n_1860;
  wire n_1862, n_1863, n_1864, n_1865, n_1867, n_1869, n_1871, n_1872;
  wire n_1873, n_1875, n_1876, n_1877, n_1879, n_1880, n_1882, n_1884;
  wire n_1886, n_1887, n_1888, n_1890, n_1891, n_1892, n_1894, n_1895;
  wire n_1897, n_1899, n_1901, n_1902, n_1903, n_1905, n_1906, n_1907;
  wire n_1909, n_1910, n_1912, n_1914, n_1916, n_1917, n_1918, n_1920;
  wire n_1921, n_1922, n_1924, n_1925, n_1927, n_1929, n_1931, n_1932;
  wire n_1933, n_1935, n_1937, n_1938, n_1939, n_1941, n_1942, n_1944;
  wire n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952;
  wire n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1960, n_1963;
  wire n_1965, n_1966, n_1967, n_1970, n_1973, n_1975, n_1976, n_1978;
  wire n_1980, n_1981, n_1983, n_1985, n_1986, n_1988, n_1990, n_1991;
  wire n_1993, n_1994, n_1996, n_1999, n_2001, n_2002, n_2003, n_2006;
  wire n_2009, n_2011, n_2012, n_2014, n_2016, n_2017, n_2019, n_2021;
  wire n_2022, n_2024, n_2026, n_2027, n_2028, n_2030, n_2031, n_2033;
  wire n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041;
  wire n_2042, n_2043, n_2044, n_2046, n_2047, n_2048, n_2050, n_2051;
  wire n_2052, n_2054, n_2055, n_2056, n_2058, n_2059, n_2060, n_2062;
  wire n_2063, n_2064, n_2066, n_2067, n_2068, n_2070, n_2071, n_2072;
  wire n_2074, n_2075, n_2076, n_2078, n_2079, n_2080, n_2082, n_2083;
  wire n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092;
  wire n_2093, n_2094, n_2095, n_2096, n_2098, n_2099, n_2100, n_2102;
  wire n_2103, n_2104, n_2106, n_2107, n_2108, n_2110, n_2111, n_2112;
  wire n_2114, n_2115, n_2116, n_2118, n_2119, n_2120, n_2122, n_2123;
  wire n_2125, n_2128, n_2129, n_2131, n_2132, n_2133, n_2134, n_2136;
  wire n_2137, n_2138, n_2140, n_2141, n_2142, n_2143, n_2145, n_2146;
  wire n_2148, n_2149, n_2151, n_2152, n_2153, n_2154, n_2156, n_2157;
  wire n_2158, n_2160, n_2161, n_2162, n_2163, n_2165, n_2166, n_2168;
  wire n_2169, n_2171, n_2172, n_2173, n_2174, n_2176, n_2177, n_2178;
  wire n_2179, n_2181, n_2182, n_2183, n_2184, n_2186, n_2187, n_2189;
  wire n_2190, n_2192, n_2193, n_2194, n_2195, n_2197, n_2198, n_2199;
  wire n_2201, n_2202, n_2203, n_2204, n_2206, n_2207, n_2209, n_2210;
  wire n_2212, n_2213, n_2214, n_2215, n_2217, n_2218, n_2219, n_2220;
  wire n_2222, n_2223, n_2224, n_2225, n_2227, n_2228, n_2230, n_2231;
  wire n_2233, n_2234, n_2235, n_2236, n_2238, n_2239;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_623, A[1], n_171);
  xor g270 (n_117, n_623, A[2]);
  nand g3 (n_624, A[1], n_171);
  nand g271 (n_625, A[2], n_171);
  nand g272 (n_626, A[1], A[2]);
  nand g273 (n_172, n_624, n_625, n_626);
  xor g274 (n_627, A[2], A[3]);
  xor g275 (n_116, n_627, n_172);
  nand g276 (n_628, A[2], A[3]);
  nand g4 (n_629, n_172, A[3]);
  nand g277 (n_630, A[2], n_172);
  nand g278 (n_67, n_628, n_629, n_630);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_631, A[4], n_173);
  xor g282 (n_115, n_631, A[6]);
  nand g283 (n_632, A[4], n_173);
  nand g284 (n_633, A[6], n_173);
  nand g5 (n_634, A[4], A[6]);
  nand g6 (n_66, n_632, n_633, n_634);
  xor g287 (n_635, n_68, A[4]);
  xor g288 (n_176, n_635, n_69);
  nand g289 (n_636, n_68, A[4]);
  nand g290 (n_637, n_69, A[4]);
  nand g291 (n_638, n_68, n_69);
  nand g292 (n_179, n_636, n_637, n_638);
  xor g293 (n_639, A[5], n_176);
  xor g294 (n_114, n_639, A[7]);
  nand g295 (n_640, A[5], n_176);
  nand g296 (n_641, A[7], n_176);
  nand g297 (n_642, A[5], A[7]);
  nand g298 (n_65, n_640, n_641, n_642);
  xor g299 (n_643, A[1], A[2]);
  xor g300 (n_178, n_643, n_171);
  xor g305 (n_647, A[5], n_178);
  xor g306 (n_180, n_647, A[6]);
  nand g307 (n_648, A[5], n_178);
  nand g308 (n_649, A[6], n_178);
  nand g309 (n_650, A[5], A[6]);
  nand g310 (n_183, n_648, n_649, n_650);
  xor g311 (n_651, n_179, n_180);
  xor g312 (n_113, n_651, A[8]);
  nand g313 (n_652, n_179, n_180);
  nand g314 (n_653, A[8], n_180);
  nand g315 (n_654, n_179, A[8]);
  nand g316 (n_64, n_652, n_653, n_654);
  xor g323 (n_659, A[6], n_116);
  xor g324 (n_184, n_659, A[7]);
  nand g325 (n_660, A[6], n_116);
  nand g326 (n_661, A[7], n_116);
  nand g327 (n_662, A[6], A[7]);
  nand g328 (n_187, n_660, n_661, n_662);
  xor g329 (n_663, n_183, A[9]);
  xor g330 (n_112, n_663, n_184);
  nand g331 (n_664, n_183, A[9]);
  nand g332 (n_665, n_184, A[9]);
  nand g333 (n_666, n_183, n_184);
  nand g334 (n_63, n_664, n_665, n_666);
  xor g338 (n_188, n_631, A[7]);
  nand g340 (n_669, A[7], n_173);
  nand g341 (n_670, A[4], A[7]);
  nand g342 (n_193, n_632, n_669, n_670);
  xor g343 (n_671, n_67, A[8]);
  xor g344 (n_189, n_671, n_187);
  nand g345 (n_672, n_67, A[8]);
  nand g346 (n_673, n_187, A[8]);
  nand g347 (n_674, n_67, n_187);
  nand g348 (n_195, n_672, n_673, n_674);
  xor g349 (n_675, A[10], n_188);
  xor g350 (n_111, n_675, n_189);
  nand g351 (n_676, A[10], n_188);
  nand g352 (n_677, n_189, n_188);
  nand g353 (n_678, A[10], n_189);
  nand g354 (n_62, n_676, n_677, n_678);
  xor g364 (n_72, n_639, A[8]);
  nand g366 (n_685, A[8], n_176);
  nand g367 (n_686, A[5], A[8]);
  nand g368 (n_201, n_640, n_685, n_686);
  xor g369 (n_687, A[9], n_193);
  xor g370 (n_196, n_687, A[11]);
  nand g371 (n_688, A[9], n_193);
  nand g372 (n_689, A[11], n_193);
  nand g373 (n_690, A[9], A[11]);
  nand g374 (n_202, n_688, n_689, n_690);
  xor g375 (n_691, n_72, n_195);
  xor g376 (n_110, n_691, n_196);
  nand g377 (n_692, n_72, n_195);
  nand g378 (n_693, n_196, n_195);
  nand g379 (n_694, n_72, n_196);
  nand g380 (n_61, n_692, n_693, n_694);
  xor g387 (n_699, A[5], n_117);
  xor g388 (n_200, n_699, A[6]);
  nand g389 (n_700, A[5], n_117);
  nand g390 (n_701, A[6], n_117);
  nand g392 (n_207, n_700, n_701, n_650);
  xor g393 (n_703, n_179, n_200);
  xor g394 (n_203, n_703, A[10]);
  nand g395 (n_704, n_179, n_200);
  nand g396 (n_705, A[10], n_200);
  nand g397 (n_706, n_179, A[10]);
  nand g398 (n_209, n_704, n_705, n_706);
  xor g399 (n_707, A[9], A[12]);
  xor g400 (n_204, n_707, n_201);
  nand g401 (n_708, A[9], A[12]);
  nand g402 (n_709, n_201, A[12]);
  nand g403 (n_710, A[9], n_201);
  nand g404 (n_211, n_708, n_709, n_710);
  xor g405 (n_711, n_202, n_203);
  xor g406 (n_109, n_711, n_204);
  nand g407 (n_712, n_202, n_203);
  nand g408 (n_713, n_204, n_203);
  nand g409 (n_714, n_202, n_204);
  nand g410 (n_60, n_712, n_713, n_714);
  xor g417 (n_719, A[6], A[7]);
  xor g418 (n_208, n_719, n_116);
  xor g423 (n_723, n_207, A[11]);
  xor g424 (n_210, n_723, A[10]);
  nand g425 (n_724, n_207, A[11]);
  nand g426 (n_725, A[10], A[11]);
  nand g427 (n_726, n_207, A[10]);
  nand g428 (n_217, n_724, n_725, n_726);
  xor g429 (n_727, n_208, A[13]);
  xor g430 (n_212, n_727, n_209);
  nand g431 (n_728, n_208, A[13]);
  nand g432 (n_729, n_209, A[13]);
  nand g433 (n_730, n_208, n_209);
  nand g434 (n_220, n_728, n_729, n_730);
  xor g435 (n_731, n_210, n_211);
  xor g436 (n_108, n_731, n_212);
  nand g437 (n_732, n_210, n_211);
  nand g438 (n_733, n_212, n_211);
  nand g439 (n_734, n_210, n_212);
  nand g440 (n_59, n_732, n_733, n_734);
  xor g444 (n_215, n_631, n_67);
  nand g446 (n_737, n_67, n_173);
  nand g447 (n_738, A[4], n_67);
  nand g448 (n_71, n_632, n_737, n_738);
  xor g449 (n_739, A[7], A[8]);
  xor g450 (n_218, n_739, n_215);
  nand g451 (n_740, A[7], A[8]);
  nand g452 (n_741, n_215, A[8]);
  nand g453 (n_742, A[7], n_215);
  nand g454 (n_223, n_740, n_741, n_742);
  xor g455 (n_743, A[11], n_187);
  xor g456 (n_219, n_743, A[12]);
  nand g457 (n_744, A[11], n_187);
  nand g458 (n_745, A[12], n_187);
  nand g459 (n_746, A[11], A[12]);
  nand g460 (n_225, n_744, n_745, n_746);
  xor g461 (n_747, A[14], n_217);
  xor g462 (n_221, n_747, n_218);
  nand g463 (n_748, A[14], n_217);
  nand g464 (n_749, n_218, n_217);
  nand g465 (n_750, A[14], n_218);
  nand g466 (n_227, n_748, n_749, n_750);
  xor g467 (n_751, n_219, n_220);
  xor g468 (n_107, n_751, n_221);
  nand g469 (n_752, n_219, n_220);
  nand g470 (n_753, n_221, n_220);
  nand g471 (n_754, n_219, n_221);
  nand g472 (n_58, n_752, n_753, n_754);
  xor g487 (n_763, A[9], n_71);
  xor g488 (n_224, n_763, A[12]);
  nand g489 (n_764, A[9], n_71);
  nand g490 (n_765, A[12], n_71);
  nand g492 (n_235, n_764, n_765, n_708);
  xor g493 (n_767, n_72, A[13]);
  xor g494 (n_226, n_767, A[15]);
  nand g495 (n_768, n_72, A[13]);
  nand g496 (n_769, A[15], A[13]);
  nand g497 (n_770, n_72, A[15]);
  nand g498 (n_237, n_768, n_769, n_770);
  xor g499 (n_771, n_223, n_224);
  xor g500 (n_228, n_771, n_225);
  nand g501 (n_772, n_223, n_224);
  nand g502 (n_773, n_225, n_224);
  nand g503 (n_774, n_223, n_225);
  nand g504 (n_239, n_772, n_773, n_774);
  xor g505 (n_775, n_226, n_227);
  xor g506 (n_106, n_775, n_228);
  nand g507 (n_776, n_226, n_227);
  nand g508 (n_777, n_228, n_227);
  nand g509 (n_778, n_226, n_228);
  nand g510 (n_57, n_776, n_777, n_778);
  xor g524 (n_234, n_651, A[9]);
  nand g526 (n_789, A[9], n_180);
  nand g527 (n_790, n_179, A[9]);
  nand g528 (n_245, n_652, n_789, n_790);
  xor g529 (n_791, A[10], n_201);
  xor g530 (n_236, n_791, A[14]);
  nand g531 (n_792, A[10], n_201);
  nand g532 (n_793, A[14], n_201);
  nand g533 (n_794, A[10], A[14]);
  nand g534 (n_247, n_792, n_793, n_794);
  xor g535 (n_795, A[13], n_234);
  xor g536 (n_238, n_795, n_235);
  nand g537 (n_796, A[13], n_234);
  nand g538 (n_797, n_235, n_234);
  nand g539 (n_798, A[13], n_235);
  nand g540 (n_249, n_796, n_797, n_798);
  xor g541 (n_799, A[16], n_236);
  xor g542 (n_240, n_799, n_237);
  nand g543 (n_800, A[16], n_236);
  nand g544 (n_801, n_237, n_236);
  nand g545 (n_802, A[16], n_237);
  nand g546 (n_251, n_800, n_801, n_802);
  xor g547 (n_803, n_238, n_239);
  xor g548 (n_105, n_803, n_240);
  nand g549 (n_804, n_238, n_239);
  nand g550 (n_805, n_240, n_239);
  nand g551 (n_806, n_238, n_240);
  nand g552 (n_56, n_804, n_805, n_806);
  xor g565 (n_815, n_183, A[10]);
  xor g566 (n_246, n_815, A[11]);
  nand g567 (n_816, n_183, A[10]);
  nand g569 (n_818, n_183, A[11]);
  nand g570 (n_258, n_816, n_725, n_818);
  xor g571 (n_819, n_208, A[14]);
  xor g572 (n_248, n_819, n_245);
  nand g573 (n_820, n_208, A[14]);
  nand g574 (n_821, n_245, A[14]);
  nand g575 (n_822, n_208, n_245);
  nand g576 (n_260, n_820, n_821, n_822);
  xor g577 (n_823, A[15], n_246);
  xor g578 (n_250, n_823, n_247);
  nand g579 (n_824, A[15], n_246);
  nand g580 (n_825, n_247, n_246);
  nand g581 (n_826, A[15], n_247);
  nand g582 (n_262, n_824, n_825, n_826);
  xor g583 (n_827, n_248, A[17]);
  xor g584 (n_252, n_827, n_249);
  nand g585 (n_828, n_248, A[17]);
  nand g586 (n_829, n_249, A[17]);
  nand g587 (n_830, n_248, n_249);
  nand g588 (n_118, n_828, n_829, n_830);
  xor g589 (n_831, n_250, n_251);
  xor g590 (n_104, n_831, n_252);
  nand g591 (n_832, n_250, n_251);
  nand g592 (n_833, n_252, n_251);
  nand g593 (n_834, n_250, n_252);
  nand g594 (n_55, n_832, n_833, n_834);
  xor g604 (n_257, n_671, n_188);
  nand g606 (n_841, n_188, A[8]);
  nand g607 (n_842, n_67, n_188);
  nand g608 (n_269, n_672, n_841, n_842);
  xor g615 (n_847, A[15], n_257);
  xor g616 (n_261, n_847, n_258);
  nand g617 (n_848, A[15], n_257);
  nand g618 (n_849, n_258, n_257);
  nand g619 (n_850, A[15], n_258);
  nand g620 (n_273, n_848, n_849, n_850);
  xor g621 (n_851, n_219, A[16]);
  xor g622 (n_263, n_851, A[18]);
  nand g623 (n_852, n_219, A[16]);
  nand g624 (n_853, A[18], A[16]);
  nand g625 (n_854, n_219, A[18]);
  nand g626 (n_275, n_852, n_853, n_854);
  xor g627 (n_855, n_260, n_261);
  xor g628 (n_119, n_855, n_262);
  nand g629 (n_856, n_260, n_261);
  nand g630 (n_857, n_262, n_261);
  nand g631 (n_858, n_260, n_262);
  nand g632 (n_277, n_856, n_857, n_858);
  xor g633 (n_859, n_263, n_118);
  xor g634 (n_103, n_859, n_119);
  nand g635 (n_860, n_263, n_118);
  nand g636 (n_861, n_119, n_118);
  nand g637 (n_862, n_263, n_119);
  nand g638 (n_54, n_860, n_861, n_862);
  xor g642 (n_266, n_635, A[5]);
  nand g644 (n_865, A[5], A[4]);
  nand g645 (n_866, n_68, A[5]);
  nand g646 (n_281, n_636, n_865, n_866);
  xor g647 (n_867, n_69, n_266);
  xor g648 (n_268, n_867, A[8]);
  nand g649 (n_868, n_69, n_266);
  nand g650 (n_869, A[8], n_266);
  nand g651 (n_870, n_69, A[8]);
  nand g652 (n_283, n_868, n_869, n_870);
  xor g654 (n_271, n_687, A[12]);
  nand g656 (n_873, A[12], n_193);
  nand g658 (n_285, n_688, n_873, n_708);
  xor g659 (n_875, A[13], n_268);
  xor g660 (n_272, n_875, n_269);
  nand g661 (n_876, A[13], n_268);
  nand g662 (n_877, n_269, n_268);
  nand g663 (n_878, A[13], n_269);
  nand g664 (n_286, n_876, n_877, n_878);
  xor g665 (n_879, n_225, n_271);
  xor g666 (n_274, n_879, A[16]);
  nand g667 (n_880, n_225, n_271);
  nand g668 (n_881, A[16], n_271);
  nand g669 (n_882, n_225, A[16]);
  nand g670 (n_289, n_880, n_881, n_882);
  xor g671 (n_883, A[19], A[17]);
  xor g672 (n_276, n_883, n_272);
  nand g673 (n_884, A[19], A[17]);
  nand g674 (n_885, n_272, A[17]);
  nand g675 (n_886, A[19], n_272);
  nand g676 (n_290, n_884, n_885, n_886);
  xor g677 (n_887, n_273, n_274);
  xor g678 (n_278, n_887, n_275);
  nand g679 (n_888, n_273, n_274);
  nand g680 (n_889, n_275, n_274);
  nand g681 (n_890, n_273, n_275);
  nand g682 (n_293, n_888, n_889, n_890);
  xor g683 (n_891, n_276, n_277);
  xor g684 (n_102, n_891, n_278);
  nand g685 (n_892, n_276, n_277);
  nand g686 (n_893, n_278, n_277);
  nand g687 (n_894, n_276, n_278);
  nand g688 (n_53, n_892, n_893, n_894);
  xor g701 (n_903, n_281, n_180);
  xor g702 (n_284, n_903, A[10]);
  nand g703 (n_904, n_281, n_180);
  nand g704 (n_905, A[10], n_180);
  nand g705 (n_906, n_281, A[10]);
  nand g706 (n_299, n_904, n_905, n_906);
  xor g707 (n_907, A[9], A[13]);
  xor g708 (n_287, n_907, n_283);
  nand g709 (n_908, A[9], A[13]);
  nand g710 (n_909, n_283, A[13]);
  nand g711 (n_910, A[9], n_283);
  nand g712 (n_301, n_908, n_909, n_910);
  xor g713 (n_911, A[14], n_284);
  xor g714 (n_288, n_911, n_285);
  nand g715 (n_912, A[14], n_284);
  nand g716 (n_913, n_285, n_284);
  nand g717 (n_914, A[14], n_285);
  nand g718 (n_303, n_912, n_913, n_914);
  xor g719 (n_915, n_286, A[18]);
  xor g720 (n_291, n_915, A[17]);
  nand g721 (n_916, n_286, A[18]);
  nand g722 (n_917, A[17], A[18]);
  nand g723 (n_918, n_286, A[17]);
  nand g724 (n_305, n_916, n_917, n_918);
  xor g725 (n_919, n_287, A[20]);
  xor g726 (n_292, n_919, n_288);
  nand g727 (n_920, n_287, A[20]);
  nand g728 (n_921, n_288, A[20]);
  nand g729 (n_922, n_287, n_288);
  nand g730 (n_306, n_920, n_921, n_922);
  xor g731 (n_923, n_289, n_290);
  xor g732 (n_294, n_923, n_291);
  nand g733 (n_924, n_289, n_290);
  nand g734 (n_925, n_291, n_290);
  nand g735 (n_926, n_289, n_291);
  nand g736 (n_309, n_924, n_925, n_926);
  xor g737 (n_927, n_292, n_293);
  xor g738 (n_101, n_927, n_294);
  nand g739 (n_928, n_292, n_293);
  nand g740 (n_929, n_294, n_293);
  nand g741 (n_930, n_292, n_294);
  nand g742 (n_52, n_928, n_929, n_930);
  xor g755 (n_939, n_183, A[11]);
  xor g756 (n_300, n_939, A[10]);
  xor g762 (n_302, n_819, A[15]);
  nand g764 (n_945, A[15], A[14]);
  nand g765 (n_946, n_208, A[15]);
  nand g766 (n_318, n_820, n_945, n_946);
  xor g767 (n_947, n_299, n_300);
  xor g768 (n_304, n_947, n_301);
  nand g769 (n_948, n_299, n_300);
  nand g770 (n_949, n_301, n_300);
  nand g771 (n_950, n_299, n_301);
  nand g772 (n_320, n_948, n_949, n_950);
  xor g773 (n_951, A[19], n_302);
  xor g774 (n_307, n_951, A[18]);
  nand g775 (n_952, A[19], n_302);
  nand g776 (n_953, A[18], n_302);
  nand g777 (n_954, A[19], A[18]);
  nand g778 (n_321, n_952, n_953, n_954);
  xor g779 (n_955, A[21], n_303);
  xor g780 (n_308, n_955, n_304);
  nand g781 (n_956, A[21], n_303);
  nand g782 (n_957, n_304, n_303);
  nand g783 (n_958, A[21], n_304);
  nand g784 (n_324, n_956, n_957, n_958);
  xor g785 (n_959, n_305, n_306);
  xor g786 (n_310, n_959, n_307);
  nand g787 (n_960, n_305, n_306);
  nand g788 (n_961, n_307, n_306);
  nand g789 (n_962, n_305, n_307);
  nand g790 (n_326, n_960, n_961, n_962);
  xor g791 (n_963, n_308, n_309);
  xor g792 (n_100, n_963, n_310);
  nand g793 (n_964, n_308, n_309);
  nand g794 (n_965, n_310, n_309);
  nand g795 (n_966, n_308, n_310);
  nand g796 (n_51, n_964, n_965, n_966);
  xor g806 (n_315, n_671, A[11]);
  nand g808 (n_973, A[11], A[8]);
  nand g809 (n_974, n_67, A[11]);
  nand g810 (n_333, n_672, n_973, n_974);
  xor g811 (n_975, n_188, n_187);
  xor g812 (n_317, n_975, A[12]);
  nand g813 (n_976, n_188, n_187);
  nand g815 (n_978, n_188, A[12]);
  nand g816 (n_334, n_976, n_745, n_978);
  xor g817 (n_979, n_315, n_258);
  xor g818 (n_319, n_979, A[15]);
  nand g819 (n_980, n_315, n_258);
  nand g821 (n_982, n_315, A[15]);
  nand g822 (n_336, n_980, n_850, n_982);
  xor g823 (n_983, n_317, A[16]);
  xor g824 (n_322, n_983, n_318);
  nand g825 (n_984, n_317, A[16]);
  nand g826 (n_985, n_318, A[16]);
  nand g827 (n_986, n_317, n_318);
  nand g828 (n_339, n_984, n_985, n_986);
  xor g829 (n_987, A[19], n_319);
  xor g830 (n_323, n_987, A[22]);
  nand g831 (n_988, A[19], n_319);
  nand g832 (n_989, A[22], n_319);
  nand g833 (n_990, A[19], A[22]);
  nand g834 (n_340, n_988, n_989, n_990);
  xor g835 (n_991, A[20], n_320);
  xor g836 (n_325, n_991, n_321);
  nand g837 (n_992, A[20], n_320);
  nand g838 (n_993, n_321, n_320);
  nand g839 (n_994, A[20], n_321);
  nand g840 (n_343, n_992, n_993, n_994);
  xor g841 (n_995, n_322, n_323);
  xor g842 (n_327, n_995, n_324);
  nand g843 (n_996, n_322, n_323);
  nand g844 (n_997, n_324, n_323);
  nand g845 (n_998, n_322, n_324);
  nand g846 (n_345, n_996, n_997, n_998);
  xor g847 (n_999, n_325, n_326);
  xor g848 (n_99, n_999, n_327);
  nand g849 (n_1000, n_325, n_326);
  nand g850 (n_1001, n_327, n_326);
  nand g851 (n_1002, n_325, n_327);
  nand g852 (n_50, n_1000, n_1001, n_1002);
  xor g874 (n_337, n_875, n_333);
  nand g876 (n_1017, n_333, A[13]);
  nand g877 (n_1018, n_268, n_333);
  nand g878 (n_357, n_876, n_1017, n_1018);
  xor g879 (n_1019, n_334, n_271);
  xor g880 (n_338, n_1019, A[16]);
  nand g881 (n_1020, n_334, n_271);
  nand g883 (n_1022, n_334, A[16]);
  nand g884 (n_359, n_1020, n_881, n_1022);
  xor g885 (n_1023, n_336, A[17]);
  xor g886 (n_341, n_1023, n_337);
  nand g887 (n_1024, n_336, A[17]);
  nand g888 (n_1025, n_337, A[17]);
  nand g889 (n_1026, n_336, n_337);
  nand g890 (n_360, n_1024, n_1025, n_1026);
  xor g891 (n_1027, A[21], A[20]);
  xor g892 (n_342, n_1027, A[23]);
  nand g893 (n_1028, A[21], A[20]);
  nand g894 (n_1029, A[23], A[20]);
  nand g895 (n_1030, A[21], A[23]);
  nand g896 (n_362, n_1028, n_1029, n_1030);
  xor g897 (n_1031, n_338, n_339);
  xor g898 (n_344, n_1031, n_340);
  nand g899 (n_1032, n_338, n_339);
  nand g900 (n_1033, n_340, n_339);
  nand g901 (n_1034, n_338, n_340);
  nand g902 (n_365, n_1032, n_1033, n_1034);
  xor g903 (n_1035, n_341, n_342);
  xor g904 (n_346, n_1035, n_343);
  nand g905 (n_1036, n_341, n_342);
  nand g906 (n_1037, n_343, n_342);
  nand g907 (n_1038, n_341, n_343);
  nand g908 (n_367, n_1036, n_1037, n_1038);
  xor g909 (n_1039, n_344, n_345);
  xor g910 (n_98, n_1039, n_346);
  nand g911 (n_1040, n_344, n_345);
  nand g912 (n_1041, n_346, n_345);
  nand g913 (n_1042, n_344, n_346);
  nand g914 (n_49, n_1040, n_1041, n_1042);
  xor g917 (n_1043, A[2], n_171);
  nand g922 (n_372, n_625, n_1045, n_1046);
  xor g923 (n_1047, A[5], n_350);
  xor g924 (n_352, n_1047, A[6]);
  nand g925 (n_1048, A[5], n_350);
  nand g926 (n_1049, A[6], n_350);
  nand g928 (n_374, n_1048, n_1049, n_650);
  xor g929 (n_1051, n_281, n_352);
  xor g930 (n_354, n_1051, A[9]);
  nand g931 (n_1052, n_281, n_352);
  nand g932 (n_1053, A[9], n_352);
  nand g933 (n_1054, n_281, A[9]);
  nand g934 (n_376, n_1052, n_1053, n_1054);
  xor g935 (n_1055, A[10], A[14]);
  xor g936 (n_356, n_1055, n_283);
  nand g938 (n_1057, n_283, A[14]);
  nand g939 (n_1058, A[10], n_283);
  nand g940 (n_378, n_794, n_1057, n_1058);
  xor g941 (n_1059, A[13], n_354);
  xor g942 (n_358, n_1059, n_285);
  nand g943 (n_1060, A[13], n_354);
  nand g944 (n_1061, n_285, n_354);
  nand g945 (n_1062, A[13], n_285);
  nand g946 (n_380, n_1060, n_1061, n_1062);
  xor g947 (n_1063, n_356, A[17]);
  xor g948 (n_361, n_1063, n_357);
  nand g949 (n_1064, n_356, A[17]);
  nand g950 (n_1065, n_357, A[17]);
  nand g951 (n_1066, n_356, n_357);
  nand g952 (n_382, n_1064, n_1065, n_1066);
  xor g953 (n_1067, A[18], n_358);
  nand g955 (n_1068, A[18], n_358);
  nand g958 (n_384, n_1068, n_1069, n_1070);
  xor g959 (n_1071, A[21], A[22]);
  xor g960 (n_363, n_1071, n_359);
  nand g961 (n_1072, A[21], A[22]);
  nand g962 (n_1073, n_359, A[22]);
  nand g963 (n_1074, A[21], n_359);
  nand g964 (n_386, n_1072, n_1073, n_1074);
  xor g965 (n_1075, n_360, n_361);
  xor g966 (n_366, n_1075, n_362);
  nand g967 (n_1076, n_360, n_361);
  nand g968 (n_1077, n_362, n_361);
  nand g969 (n_1078, n_360, n_362);
  nand g970 (n_389, n_1076, n_1077, n_1078);
  xor g971 (n_1079, n_363, n_364);
  xor g972 (n_368, n_1079, n_365);
  nand g973 (n_1080, n_363, n_364);
  nand g974 (n_1081, n_365, n_364);
  nand g975 (n_1082, n_363, n_365);
  nand g976 (n_390, n_1080, n_1081, n_1082);
  xor g977 (n_1083, n_366, n_367);
  xor g978 (n_97, n_1083, n_368);
  nand g979 (n_1084, n_366, n_367);
  nand g980 (n_1085, n_368, n_367);
  nand g981 (n_1086, n_366, n_368);
  nand g982 (n_48, n_1084, n_1085, n_1086);
  xor g985 (n_1087, A[1], A[3]);
  nand g987 (n_1088, A[1], A[3]);
  nand g990 (n_393, n_1088, n_1089, n_1090);
  xor g991 (n_1091, n_372, A[6]);
  xor g992 (n_375, n_1091, n_373);
  nand g993 (n_1092, n_372, A[6]);
  nand g994 (n_1093, n_373, A[6]);
  nand g995 (n_1094, n_372, n_373);
  nand g996 (n_395, n_1092, n_1093, n_1094);
  xor g997 (n_1095, A[7], n_374);
  xor g998 (n_377, n_1095, A[10]);
  nand g999 (n_1096, A[7], n_374);
  nand g1000 (n_1097, A[10], n_374);
  nand g1001 (n_1098, A[7], A[10]);
  nand g1002 (n_397, n_1096, n_1097, n_1098);
  xor g1003 (n_1099, A[11], n_375);
  xor g1004 (n_379, n_1099, A[14]);
  nand g1005 (n_1100, A[11], n_375);
  nand g1006 (n_1101, A[14], n_375);
  nand g1007 (n_1102, A[11], A[14]);
  nand g1008 (n_399, n_1100, n_1101, n_1102);
  xor g1009 (n_1103, n_376, n_377);
  xor g1010 (n_381, n_1103, A[15]);
  nand g1011 (n_1104, n_376, n_377);
  nand g1012 (n_1105, A[15], n_377);
  nand g1013 (n_1106, n_376, A[15]);
  nand g1014 (n_401, n_1104, n_1105, n_1106);
  xor g1015 (n_1107, n_378, n_379);
  xor g1016 (n_383, n_1107, A[18]);
  nand g1017 (n_1108, n_378, n_379);
  nand g1018 (n_1109, A[18], n_379);
  nand g1019 (n_1110, n_378, A[18]);
  nand g1020 (n_403, n_1108, n_1109, n_1110);
  xor g1021 (n_1111, A[19], n_380);
  xor g1022 (n_385, n_1111, A[22]);
  nand g1023 (n_1112, A[19], n_380);
  nand g1024 (n_1113, A[22], n_380);
  nand g1026 (n_405, n_1112, n_1113, n_990);
  xor g1027 (n_1115, n_381, A[23]);
  xor g1028 (n_387, n_1115, n_382);
  nand g1029 (n_1116, n_381, A[23]);
  nand g1030 (n_1117, n_382, A[23]);
  nand g1031 (n_1118, n_381, n_382);
  nand g1032 (n_408, n_1116, n_1117, n_1118);
  xor g1033 (n_1119, n_383, n_384);
  xor g1034 (n_388, n_1119, n_385);
  nand g1035 (n_1120, n_383, n_384);
  nand g1036 (n_1121, n_385, n_384);
  nand g1037 (n_1122, n_383, n_385);
  nand g1038 (n_409, n_1120, n_1121, n_1122);
  xor g1039 (n_1123, n_386, n_387);
  xor g1040 (n_391, n_1123, n_388);
  nand g1041 (n_1124, n_386, n_387);
  nand g1042 (n_1125, n_388, n_387);
  nand g1043 (n_1126, n_386, n_388);
  nand g1044 (n_412, n_1124, n_1125, n_1126);
  xor g1045 (n_1127, n_389, n_390);
  xor g1046 (n_96, n_1127, n_391);
  nand g1047 (n_1128, n_389, n_390);
  nand g1048 (n_1129, n_391, n_390);
  nand g1049 (n_1130, n_389, n_391);
  nand g1050 (n_47, n_1128, n_1129, n_1130);
  xor g1051 (n_1131, A[3], A[4]);
  xor g1052 (n_394, n_1131, A[2]);
  nand g1053 (n_1132, A[3], A[4]);
  nand g1054 (n_1133, A[2], A[4]);
  nand g1056 (n_413, n_1132, n_1133, n_628);
  xor g1057 (n_1135, n_393, A[7]);
  xor g1058 (n_396, n_1135, n_394);
  nand g1059 (n_1136, n_393, A[7]);
  nand g1060 (n_1137, n_394, A[7]);
  nand g1061 (n_1138, n_393, n_394);
  nand g1062 (n_415, n_1136, n_1137, n_1138);
  xor g1063 (n_1139, A[8], n_395);
  xor g1064 (n_398, n_1139, A[11]);
  nand g1065 (n_1140, A[8], n_395);
  nand g1066 (n_1141, A[11], n_395);
  nand g1068 (n_417, n_1140, n_1141, n_973);
  xor g1069 (n_1143, A[12], n_396);
  xor g1070 (n_400, n_1143, n_397);
  nand g1071 (n_1144, A[12], n_396);
  nand g1072 (n_1145, n_397, n_396);
  nand g1073 (n_1146, A[12], n_397);
  nand g1074 (n_419, n_1144, n_1145, n_1146);
  xor g1075 (n_1147, n_398, A[15]);
  xor g1076 (n_402, n_1147, n_399);
  nand g1077 (n_1148, n_398, A[15]);
  nand g1078 (n_1149, n_399, A[15]);
  nand g1079 (n_1150, n_398, n_399);
  nand g1080 (n_420, n_1148, n_1149, n_1150);
  xor g1081 (n_1151, A[16], A[19]);
  xor g1082 (n_404, n_1151, n_400);
  nand g1083 (n_1152, A[16], A[19]);
  nand g1084 (n_1153, n_400, A[19]);
  nand g1085 (n_1154, A[16], n_400);
  nand g1086 (n_422, n_1152, n_1153, n_1154);
  xor g1088 (n_406, n_1155, A[20]);
  nand g1091 (n_1158, n_401, A[20]);
  nand g1092 (n_423, n_1156, n_1157, n_1158);
  xor g1093 (n_1159, n_402, A[23]);
  xor g1094 (n_407, n_1159, n_403);
  nand g1095 (n_1160, n_402, A[23]);
  nand g1096 (n_1161, n_403, A[23]);
  nand g1097 (n_1162, n_402, n_403);
  nand g1098 (n_426, n_1160, n_1161, n_1162);
  xor g1099 (n_1163, n_404, n_405);
  xor g1100 (n_410, n_1163, n_406);
  nand g1101 (n_1164, n_404, n_405);
  nand g1102 (n_1165, n_406, n_405);
  nand g1103 (n_1166, n_404, n_406);
  nand g1104 (n_428, n_1164, n_1165, n_1166);
  xor g1105 (n_1167, n_407, n_408);
  xor g1106 (n_411, n_1167, n_409);
  nand g1107 (n_1168, n_407, n_408);
  nand g1108 (n_1169, n_409, n_408);
  nand g1109 (n_1170, n_407, n_409);
  nand g1110 (n_431, n_1168, n_1169, n_1170);
  xor g1111 (n_1171, n_410, n_411);
  xor g1112 (n_95, n_1171, n_412);
  nand g1113 (n_1172, n_410, n_411);
  nand g1114 (n_1173, n_412, n_411);
  nand g1115 (n_1174, n_410, n_412);
  nand g1116 (n_46, n_1172, n_1173, n_1174);
  xor g1117 (n_1175, A[4], A[5]);
  xor g1118 (n_414, n_1175, n_413);
  nand g1120 (n_1177, n_413, A[5]);
  nand g1121 (n_1178, A[4], n_413);
  nand g1122 (n_434, n_865, n_1177, n_1178);
  xor g1123 (n_1179, A[8], n_414);
  xor g1124 (n_416, n_1179, A[9]);
  nand g1125 (n_1180, A[8], n_414);
  nand g1126 (n_1181, A[9], n_414);
  nand g1127 (n_1182, A[8], A[9]);
  nand g1128 (n_436, n_1180, n_1181, n_1182);
  xor g1129 (n_1183, n_415, A[12]);
  xor g1130 (n_418, n_1183, A[13]);
  nand g1131 (n_1184, n_415, A[12]);
  nand g1132 (n_1185, A[13], A[12]);
  nand g1133 (n_1186, n_415, A[13]);
  nand g1134 (n_438, n_1184, n_1185, n_1186);
  xor g1135 (n_1187, n_416, n_417);
  xor g1136 (n_421, n_1187, n_418);
  nand g1137 (n_1188, n_416, n_417);
  nand g1138 (n_1189, n_418, n_417);
  nand g1139 (n_1190, n_416, n_418);
  nand g1140 (n_440, n_1188, n_1189, n_1190);
  xor g1141 (n_1191, A[16], A[17]);
  xor g1142 (n_424, n_1191, n_419);
  nand g1143 (n_1192, A[16], A[17]);
  nand g1144 (n_1193, n_419, A[17]);
  nand g1145 (n_1194, A[16], n_419);
  nand g1146 (n_441, n_1192, n_1193, n_1194);
  xor g1148 (n_425, n_1195, A[20]);
  nand g1152 (n_443, n_1196, n_1157, n_1028);
  xor g1153 (n_1199, n_420, n_421);
  xor g1154 (n_427, n_1199, n_422);
  nand g1155 (n_1200, n_420, n_421);
  nand g1156 (n_1201, n_422, n_421);
  nand g1157 (n_1202, n_420, n_422);
  nand g1158 (n_445, n_1200, n_1201, n_1202);
  xor g1159 (n_1203, n_423, n_424);
  xor g1160 (n_429, n_1203, n_425);
  nand g1161 (n_1204, n_423, n_424);
  nand g1162 (n_1205, n_425, n_424);
  nand g1163 (n_1206, n_423, n_425);
  nand g1164 (n_448, n_1204, n_1205, n_1206);
  xor g1165 (n_1207, n_426, n_427);
  xor g1166 (n_430, n_1207, n_428);
  nand g1167 (n_1208, n_426, n_427);
  nand g1168 (n_1209, n_428, n_427);
  nand g1169 (n_1210, n_426, n_428);
  nand g1170 (n_450, n_1208, n_1209, n_1210);
  xor g1171 (n_1211, n_429, n_430);
  xor g1172 (n_94, n_1211, n_431);
  nand g1173 (n_1212, n_429, n_430);
  nand g1174 (n_1213, n_431, n_430);
  nand g1175 (n_1214, n_429, n_431);
  nand g1176 (n_45, n_1212, n_1213, n_1214);
  xor g1180 (n_435, n_1215, n_434);
  nand g1183 (n_1218, A[6], n_434);
  nand g1184 (n_455, n_1216, n_1217, n_1218);
  xor g1185 (n_1219, A[9], A[10]);
  xor g1186 (n_437, n_1219, n_435);
  nand g1187 (n_1220, A[9], A[10]);
  nand g1188 (n_1221, n_435, A[10]);
  nand g1189 (n_1222, A[9], n_435);
  nand g1190 (n_457, n_1220, n_1221, n_1222);
  xor g1191 (n_1223, A[14], A[13]);
  xor g1192 (n_439, n_1223, n_436);
  nand g1193 (n_1224, A[14], A[13]);
  nand g1194 (n_1225, n_436, A[13]);
  nand g1195 (n_1226, A[14], n_436);
  nand g1196 (n_459, n_1224, n_1225, n_1226);
  xor g1197 (n_1227, n_437, n_438);
  xor g1198 (n_442, n_1227, A[18]);
  nand g1199 (n_1228, n_437, n_438);
  nand g1200 (n_1229, A[18], n_438);
  nand g1201 (n_1230, n_437, A[18]);
  nand g1202 (n_460, n_1228, n_1229, n_1230);
  xor g1203 (n_1231, A[17], n_439);
  xor g1204 (n_444, n_1231, A[21]);
  nand g1205 (n_1232, A[17], n_439);
  nand g1206 (n_1233, A[21], n_439);
  nand g1207 (n_1234, A[17], A[21]);
  nand g1208 (n_462, n_1232, n_1233, n_1234);
  xor g1209 (n_1235, A[22], n_440);
  xor g1210 (n_446, n_1235, n_441);
  nand g1211 (n_1236, A[22], n_440);
  nand g1212 (n_1237, n_441, n_440);
  nand g1213 (n_1238, A[22], n_441);
  nand g1214 (n_464, n_1236, n_1237, n_1238);
  xor g1215 (n_1239, n_442, n_443);
  xor g1216 (n_447, n_1239, n_444);
  nand g1217 (n_1240, n_442, n_443);
  nand g1218 (n_1241, n_444, n_443);
  nand g1219 (n_1242, n_442, n_444);
  nand g1220 (n_466, n_1240, n_1241, n_1242);
  xor g1221 (n_1243, n_445, n_446);
  xor g1222 (n_449, n_1243, n_447);
  nand g1223 (n_1244, n_445, n_446);
  nand g1224 (n_1245, n_447, n_446);
  nand g1225 (n_1246, n_445, n_447);
  nand g1226 (n_469, n_1244, n_1245, n_1246);
  xor g1227 (n_1247, n_448, n_449);
  xor g1228 (n_93, n_1247, n_450);
  nand g1229 (n_1248, n_448, n_449);
  nand g1230 (n_1249, n_450, n_449);
  nand g1231 (n_1250, n_448, n_450);
  nand g1232 (n_44, n_1248, n_1249, n_1250);
  xor g1235 (n_1251, A[5], A[7]);
  nand g1240 (n_471, n_642, n_1253, n_1254);
  xor g1241 (n_1255, A[10], A[11]);
  xor g1242 (n_456, n_1255, n_454);
  nand g1244 (n_1257, n_454, A[11]);
  nand g1245 (n_1258, A[10], n_454);
  nand g1246 (n_473, n_725, n_1257, n_1258);
  xor g1247 (n_1259, A[14], n_455);
  xor g1248 (n_458, n_1259, A[15]);
  nand g1249 (n_1260, A[14], n_455);
  nand g1250 (n_1261, A[15], n_455);
  nand g1252 (n_475, n_1260, n_1261, n_945);
  xor g1253 (n_1263, n_456, n_457);
  xor g1254 (n_461, n_1263, A[19]);
  nand g1255 (n_1264, n_456, n_457);
  nand g1256 (n_1265, A[19], n_457);
  nand g1257 (n_1266, n_456, A[19]);
  nand g1258 (n_478, n_1264, n_1265, n_1266);
  xor g1259 (n_1267, A[18], n_458);
  xor g1260 (n_463, n_1267, n_459);
  nand g1261 (n_1268, A[18], n_458);
  nand g1262 (n_1269, n_459, n_458);
  nand g1263 (n_1270, A[18], n_459);
  nand g1264 (n_479, n_1268, n_1269, n_1270);
  xor g1265 (n_1271, A[22], A[23]);
  xor g1266 (n_465, n_1271, n_460);
  nand g1267 (n_1272, A[22], A[23]);
  nand g1268 (n_1273, n_460, A[23]);
  nand g1269 (n_1274, A[22], n_460);
  nand g1270 (n_481, n_1272, n_1273, n_1274);
  xor g1271 (n_1275, n_461, n_462);
  xor g1272 (n_467, n_1275, n_463);
  nand g1273 (n_1276, n_461, n_462);
  nand g1274 (n_1277, n_463, n_462);
  nand g1275 (n_1278, n_461, n_463);
  nand g1276 (n_483, n_1276, n_1277, n_1278);
  xor g1277 (n_1279, n_464, n_465);
  xor g1278 (n_468, n_1279, n_466);
  nand g1279 (n_1280, n_464, n_465);
  nand g1280 (n_1281, n_466, n_465);
  nand g1281 (n_1282, n_464, n_466);
  nand g1282 (n_486, n_1280, n_1281, n_1282);
  xor g1283 (n_1283, n_467, n_468);
  xor g1284 (n_92, n_1283, n_469);
  nand g1285 (n_1284, n_467, n_468);
  nand g1286 (n_1285, n_469, n_468);
  nand g1287 (n_1286, n_467, n_469);
  nand g1288 (n_43, n_1284, n_1285, n_1286);
  xor g1290 (n_472, n_719, A[8]);
  nand g1292 (n_1289, A[8], A[6]);
  nand g1294 (n_487, n_662, n_1289, n_740);
  xor g1295 (n_1291, A[11], A[12]);
  xor g1296 (n_474, n_1291, n_471);
  nand g1298 (n_1293, n_471, A[12]);
  nand g1299 (n_1294, A[11], n_471);
  nand g1300 (n_488, n_746, n_1293, n_1294);
  xor g1301 (n_1295, n_472, A[15]);
  xor g1302 (n_476, n_1295, n_473);
  nand g1303 (n_1296, n_472, A[15]);
  nand g1304 (n_1297, n_473, A[15]);
  nand g1305 (n_1298, n_472, n_473);
  nand g1306 (n_490, n_1296, n_1297, n_1298);
  xor g1307 (n_1299, n_474, A[16]);
  xor g1308 (n_477, n_1299, A[19]);
  nand g1309 (n_1300, n_474, A[16]);
  nand g1311 (n_1302, n_474, A[19]);
  nand g1312 (n_493, n_1300, n_1152, n_1302);
  xor g1314 (n_480, n_1303, A[20]);
  nand g1317 (n_1306, n_475, A[20]);
  nand g1318 (n_494, n_1304, n_1157, n_1306);
  xor g1319 (n_1307, n_476, A[23]);
  xor g1320 (n_482, n_1307, n_477);
  nand g1321 (n_1308, n_476, A[23]);
  nand g1322 (n_1309, n_477, A[23]);
  nand g1323 (n_1310, n_476, n_477);
  nand g1324 (n_497, n_1308, n_1309, n_1310);
  xor g1325 (n_1311, n_478, n_479);
  xor g1326 (n_484, n_1311, n_480);
  nand g1327 (n_1312, n_478, n_479);
  nand g1328 (n_1313, n_480, n_479);
  nand g1329 (n_1314, n_478, n_480);
  nand g1330 (n_499, n_1312, n_1313, n_1314);
  xor g1331 (n_1315, n_481, n_482);
  xor g1332 (n_485, n_1315, n_483);
  nand g1333 (n_1316, n_481, n_482);
  nand g1334 (n_1317, n_483, n_482);
  nand g1335 (n_1318, n_481, n_483);
  nand g1336 (n_500, n_1316, n_1317, n_1318);
  xor g1337 (n_1319, n_484, n_485);
  xor g1338 (n_91, n_1319, n_486);
  nand g1339 (n_1320, n_484, n_485);
  nand g1340 (n_1321, n_486, n_485);
  nand g1341 (n_1322, n_484, n_486);
  nand g1342 (n_42, n_1320, n_1321, n_1322);
  xor g1343 (n_1323, A[8], A[9]);
  xor g1344 (n_489, n_1323, A[12]);
  nand g1347 (n_1326, A[8], A[12]);
  nand g1348 (n_504, n_1182, n_708, n_1326);
  xor g1349 (n_1327, n_487, A[13]);
  xor g1350 (n_491, n_1327, n_488);
  nand g1351 (n_1328, n_487, A[13]);
  nand g1352 (n_1329, n_488, A[13]);
  nand g1353 (n_1330, n_487, n_488);
  nand g1354 (n_506, n_1328, n_1329, n_1330);
  xor g1355 (n_1331, n_489, A[16]);
  xor g1356 (n_492, n_1331, A[17]);
  nand g1357 (n_1332, n_489, A[16]);
  nand g1359 (n_1334, n_489, A[17]);
  nand g1360 (n_507, n_1332, n_1192, n_1334);
  xor g1362 (n_495, n_1335, n_491);
  nand g1365 (n_1338, n_490, n_491);
  nand g1366 (n_509, n_1336, n_1337, n_1338);
  xor g1368 (n_496, n_1027, n_492);
  nand g1370 (n_1341, n_492, A[21]);
  nand g1371 (n_1342, A[20], n_492);
  nand g1372 (n_511, n_1028, n_1341, n_1342);
  xor g1373 (n_1343, n_493, n_494);
  xor g1374 (n_498, n_1343, n_495);
  nand g1375 (n_1344, n_493, n_494);
  nand g1376 (n_1345, n_495, n_494);
  nand g1377 (n_1346, n_493, n_495);
  nand g1378 (n_514, n_1344, n_1345, n_1346);
  xor g1379 (n_1347, n_496, n_497);
  xor g1380 (n_501, n_1347, n_498);
  nand g1381 (n_1348, n_496, n_497);
  nand g1382 (n_1349, n_498, n_497);
  nand g1383 (n_1350, n_496, n_498);
  nand g1384 (n_516, n_1348, n_1349, n_1350);
  xor g1385 (n_1351, n_499, n_500);
  xor g1386 (n_90, n_1351, n_501);
  nand g1387 (n_1352, n_499, n_500);
  nand g1388 (n_1353, n_501, n_500);
  nand g1389 (n_1354, n_499, n_501);
  nand g1390 (n_41, n_1352, n_1353, n_1354);
  nand g1397 (n_1358, A[9], A[14]);
  nand g1398 (n_520, n_1356, n_1357, n_1358);
  xor g1399 (n_1359, A[13], n_504);
  xor g1400 (n_508, n_1359, A[18]);
  nand g1401 (n_1360, A[13], n_504);
  nand g1402 (n_1361, A[18], n_504);
  nand g1403 (n_1362, A[13], A[18]);
  nand g1404 (n_523, n_1360, n_1361, n_1362);
  xor g1405 (n_1363, A[17], n_505);
  xor g1406 (n_510, n_1363, A[21]);
  nand g1407 (n_1364, A[17], n_505);
  nand g1408 (n_1365, A[21], n_505);
  nand g1410 (n_524, n_1364, n_1365, n_1234);
  xor g1411 (n_1367, n_506, A[22]);
  xor g1412 (n_512, n_1367, n_507);
  nand g1413 (n_1368, n_506, A[22]);
  nand g1414 (n_1369, n_507, A[22]);
  nand g1415 (n_1370, n_506, n_507);
  nand g1416 (n_527, n_1368, n_1369, n_1370);
  xor g1417 (n_1371, n_508, n_509);
  xor g1418 (n_513, n_1371, n_510);
  nand g1419 (n_1372, n_508, n_509);
  nand g1420 (n_1373, n_510, n_509);
  nand g1421 (n_1374, n_508, n_510);
  nand g1422 (n_528, n_1372, n_1373, n_1374);
  xor g1423 (n_1375, n_511, n_512);
  xor g1424 (n_515, n_1375, n_513);
  nand g1425 (n_1376, n_511, n_512);
  nand g1426 (n_1377, n_513, n_512);
  nand g1427 (n_1378, n_511, n_513);
  nand g1428 (n_531, n_1376, n_1377, n_1378);
  xor g1429 (n_1379, n_514, n_515);
  xor g1430 (n_89, n_1379, n_516);
  nand g1431 (n_1380, n_514, n_515);
  nand g1432 (n_1381, n_516, n_515);
  nand g1433 (n_1382, n_514, n_516);
  nand g1434 (n_40, n_1380, n_1381, n_1382);
  xor g1443 (n_1387, A[14], A[15]);
  xor g1444 (n_522, n_1387, n_520);
  nand g1446 (n_1389, n_520, A[15]);
  nand g1447 (n_1390, A[14], n_520);
  nand g1448 (n_535, n_945, n_1389, n_1390);
  xor g1449 (n_1391, A[19], A[18]);
  nand g1454 (n_537, n_954, n_1393, n_1394);
  xor g1455 (n_1395, A[22], n_522);
  xor g1456 (n_526, n_1395, A[23]);
  nand g1457 (n_1396, A[22], n_522);
  nand g1458 (n_1397, A[23], n_522);
  nand g1460 (n_539, n_1396, n_1397, n_1272);
  xor g1461 (n_1399, n_523, n_524);
  xor g1462 (n_529, n_1399, n_525);
  nand g1463 (n_1400, n_523, n_524);
  nand g1464 (n_1401, n_525, n_524);
  nand g1465 (n_1402, n_523, n_525);
  nand g1466 (n_541, n_1400, n_1401, n_1402);
  xor g1467 (n_1403, n_526, n_527);
  xor g1468 (n_530, n_1403, n_528);
  nand g1469 (n_1404, n_526, n_527);
  nand g1470 (n_1405, n_528, n_527);
  nand g1471 (n_1406, n_526, n_528);
  nand g1472 (n_544, n_1404, n_1405, n_1406);
  xor g1473 (n_1407, n_529, n_530);
  xor g1474 (n_88, n_1407, n_531);
  nand g1475 (n_1408, n_529, n_530);
  nand g1476 (n_1409, n_531, n_530);
  nand g1477 (n_1410, n_529, n_531);
  nand g1478 (n_39, n_1408, n_1409, n_1410);
  xor g1480 (n_534, n_1291, A[11]);
  xor g1485 (n_1415, A[15], n_533);
  xor g1486 (n_536, n_1415, A[16]);
  nand g1487 (n_1416, A[15], n_533);
  nand g1488 (n_1417, A[16], n_533);
  nand g1489 (n_1418, A[15], A[16]);
  nand g1490 (n_546, n_1416, n_1417, n_1418);
  xor g1491 (n_1419, n_534, A[19]);
  nand g1493 (n_1420, n_534, A[19]);
  nand g1496 (n_548, n_1420, n_1421, n_1422);
  xor g1497 (n_1423, A[20], A[23]);
  xor g1498 (n_540, n_1423, n_535);
  nand g1500 (n_1425, n_535, A[23]);
  nand g1501 (n_1426, A[20], n_535);
  nand g1502 (n_551, n_1029, n_1425, n_1426);
  xor g1503 (n_1427, n_536, n_537);
  xor g1504 (n_542, n_1427, n_538);
  nand g1505 (n_1428, n_536, n_537);
  nand g1506 (n_1429, n_538, n_537);
  nand g1507 (n_1430, n_536, n_538);
  nand g1508 (n_552, n_1428, n_1429, n_1430);
  xor g1509 (n_1431, n_539, n_540);
  xor g1510 (n_543, n_1431, n_541);
  nand g1511 (n_1432, n_539, n_540);
  nand g1512 (n_1433, n_541, n_540);
  nand g1513 (n_1434, n_539, n_541);
  nand g1514 (n_555, n_1432, n_1433, n_1434);
  xor g1515 (n_1435, n_542, n_543);
  xor g1516 (n_87, n_1435, n_544);
  nand g1517 (n_1436, n_542, n_543);
  nand g1518 (n_1437, n_544, n_543);
  nand g1519 (n_1438, n_542, n_544);
  nand g1520 (n_38, n_1436, n_1437, n_1438);
  xor g1521 (n_1439, A[12], A[13]);
  xor g1522 (n_547, n_1439, n_545);
  nand g1524 (n_1441, n_545, A[13]);
  nand g1525 (n_1442, A[12], n_545);
  nand g1526 (n_558, n_1185, n_1441, n_1442);
  xor g1528 (n_549, n_1191, A[21]);
  nand g1531 (n_1446, A[16], A[21]);
  nand g1532 (n_560, n_1192, n_1234, n_1446);
  xor g1534 (n_550, n_1447, n_546);
  nand g1536 (n_1449, n_546, A[20]);
  nand g1538 (n_562, n_1157, n_1449, n_1450);
  xor g1539 (n_1451, n_547, n_548);
  xor g1540 (n_553, n_1451, n_549);
  nand g1541 (n_1452, n_547, n_548);
  nand g1542 (n_1453, n_549, n_548);
  nand g1543 (n_1454, n_547, n_549);
  nand g1544 (n_563, n_1452, n_1453, n_1454);
  xor g1545 (n_1455, n_550, n_551);
  xor g1546 (n_554, n_1455, n_552);
  nand g1547 (n_1456, n_550, n_551);
  nand g1548 (n_1457, n_552, n_551);
  nand g1549 (n_1458, n_550, n_552);
  nand g1550 (n_566, n_1456, n_1457, n_1458);
  xor g1551 (n_1459, n_553, n_554);
  xor g1552 (n_86, n_1459, n_555);
  nand g1553 (n_1460, n_553, n_554);
  nand g1554 (n_1461, n_555, n_554);
  nand g1555 (n_1462, n_553, n_555);
  nand g1556 (n_37, n_1460, n_1461, n_1462);
  nand g1564 (n_571, n_1464, n_1465, n_1362);
  xor g1565 (n_1467, A[17], A[21]);
  xor g1566 (n_561, n_1467, A[22]);
  nand g1569 (n_1470, A[17], A[22]);
  nand g1570 (n_573, n_1234, n_1072, n_1470);
  xor g1571 (n_1471, n_558, n_559);
  xor g1572 (n_564, n_1471, n_560);
  nand g1573 (n_1472, n_558, n_559);
  nand g1574 (n_1473, n_560, n_559);
  nand g1575 (n_1474, n_558, n_560);
  nand g1576 (n_575, n_1472, n_1473, n_1474);
  xor g1577 (n_1475, n_561, n_562);
  xor g1578 (n_565, n_1475, n_563);
  nand g1579 (n_1476, n_561, n_562);
  nand g1580 (n_1477, n_563, n_562);
  nand g1581 (n_1478, n_561, n_563);
  nand g1582 (n_577, n_1476, n_1477, n_1478);
  xor g1583 (n_1479, n_564, n_565);
  xor g1584 (n_85, n_1479, n_566);
  nand g1585 (n_1480, n_564, n_565);
  nand g1586 (n_1481, n_566, n_565);
  nand g1587 (n_1482, n_564, n_566);
  nand g1588 (n_36, n_1480, n_1481, n_1482);
  xor g1598 (n_572, n_1391, A[22]);
  nand g1600 (n_1489, A[22], A[18]);
  nand g1602 (n_581, n_954, n_1489, n_990);
  xor g1603 (n_1491, A[23], n_570);
  xor g1604 (n_574, n_1491, n_571);
  nand g1605 (n_1492, A[23], n_570);
  nand g1606 (n_1493, n_571, n_570);
  nand g1607 (n_1494, A[23], n_571);
  nand g1608 (n_584, n_1492, n_1493, n_1494);
  xor g1609 (n_1495, n_572, n_573);
  xor g1610 (n_576, n_1495, n_574);
  nand g1611 (n_1496, n_572, n_573);
  nand g1612 (n_1497, n_574, n_573);
  nand g1613 (n_1498, n_572, n_574);
  nand g1614 (n_586, n_1496, n_1497, n_1498);
  xor g1615 (n_1499, n_575, n_576);
  xor g1616 (n_84, n_1499, n_577);
  nand g1617 (n_1500, n_575, n_576);
  nand g1618 (n_1501, n_577, n_576);
  nand g1619 (n_1502, n_575, n_577);
  nand g1620 (n_35, n_1500, n_1501, n_1502);
  xor g1622 (n_580, n_1387, A[16]);
  nand g1624 (n_1505, A[16], A[14]);
  nand g1626 (n_587, n_945, n_1505, n_1418);
  xor g1627 (n_1507, A[19], n_579);
  nand g1629 (n_1508, A[19], n_579);
  nand g1632 (n_589, n_1508, n_1509, n_1421);
  xor g1634 (n_583, n_1423, n_580);
  nand g1636 (n_1513, n_580, A[23]);
  nand g1637 (n_1514, A[20], n_580);
  nand g1638 (n_590, n_1029, n_1513, n_1514);
  xor g1639 (n_1515, n_581, n_582);
  xor g1640 (n_585, n_1515, n_583);
  nand g1641 (n_1516, n_581, n_582);
  nand g1642 (n_1517, n_583, n_582);
  nand g1643 (n_1518, n_581, n_583);
  nand g1644 (n_593, n_1516, n_1517, n_1518);
  xor g1645 (n_1519, n_584, n_585);
  xor g1646 (n_83, n_1519, n_586);
  nand g1647 (n_1520, n_584, n_585);
  nand g1648 (n_1521, n_586, n_585);
  nand g1649 (n_1522, n_584, n_586);
  nand g1650 (n_34, n_1520, n_1521, n_1522);
  xor g1658 (n_591, n_1447, n_587);
  nand g1660 (n_1529, n_587, A[20]);
  nand g1662 (n_597, n_1157, n_1529, n_1530);
  xor g1663 (n_1531, n_549, n_589);
  xor g1664 (n_592, n_1531, n_590);
  nand g1665 (n_1532, n_549, n_589);
  nand g1666 (n_1533, n_590, n_589);
  nand g1667 (n_1534, n_549, n_590);
  nand g1668 (n_600, n_1532, n_1533, n_1534);
  xor g1669 (n_1535, n_591, n_592);
  xor g1670 (n_82, n_1535, n_593);
  nand g1671 (n_1536, n_591, n_592);
  nand g1672 (n_1537, n_593, n_592);
  nand g1673 (n_1538, n_591, n_593);
  nand g1674 (n_33, n_1536, n_1537, n_1538);
  xor g1684 (n_599, n_1543, n_597);
  nand g1686 (n_1545, n_597, n_560);
  nand g1688 (n_607, n_1544, n_1545, n_1546);
  xor g1689 (n_1547, n_561, n_599);
  xor g1690 (n_81, n_1547, n_600);
  nand g1691 (n_1548, n_561, n_599);
  nand g1692 (n_1549, n_600, n_599);
  nand g1693 (n_1550, n_561, n_600);
  nand g1694 (n_32, n_1548, n_1549, n_1550);
  xor g1697 (n_1551, A[18], A[22]);
  xor g1698 (n_605, n_1551, A[23]);
  nand g1701 (n_1554, A[18], A[23]);
  nand g1702 (n_610, n_1489, n_1272, n_1554);
  nand g1706 (n_1557, n_573, A[18]);
  nand g1708 (n_611, n_1556, n_1557, n_1558);
  xor g1709 (n_1559, n_605, n_606);
  xor g1710 (n_80, n_1559, n_607);
  nand g1711 (n_1560, n_605, n_606);
  nand g1712 (n_1561, n_607, n_606);
  nand g1713 (n_1562, n_605, n_607);
  nand g1714 (n_31, n_1560, n_1561, n_1562);
  xor g1716 (n_609, n_1563, A[20]);
  nand g1719 (n_1566, A[19], A[20]);
  nand g1720 (n_613, n_1421, n_1157, n_1566);
  xor g1721 (n_1567, A[23], A[19]);
  xor g1722 (n_612, n_1567, n_609);
  nand g1723 (n_1568, A[23], A[19]);
  nand g1724 (n_1569, n_609, A[19]);
  nand g1725 (n_1570, A[23], n_609);
  nand g1726 (n_615, n_1568, n_1569, n_1570);
  xor g1727 (n_1571, n_610, n_611);
  xor g1728 (n_79, n_1571, n_612);
  nand g1729 (n_1572, n_610, n_611);
  nand g1730 (n_1573, n_612, n_611);
  nand g1731 (n_1574, n_610, n_612);
  nand g1732 (n_30, n_1572, n_1573, n_1574);
  xor g1739 (n_1579, n_613, n_425);
  xor g1740 (n_78, n_1579, n_615);
  nand g1741 (n_1580, n_613, n_425);
  nand g1742 (n_1581, n_615, n_425);
  nand g1743 (n_1582, n_613, n_615);
  nand g1744 (n_77, n_1580, n_1581, n_1582);
  nand g1751 (n_1586, A[22], n_443);
  nand g1752 (n_28, n_1584, n_1585, n_1586);
  nand g1760 (n_27, n_1588, n_1589, n_1030);
  xor g1762 (n_75, n_1591, A[22]);
  nand g1766 (n_74, n_1592, n_1272, n_1594);
  nor g11 (n_1610, A[0], A[2]);
  nand g12 (n_1605, A[0], A[2]);
  nor g13 (n_1606, n_68, A[3]);
  nand g14 (n_1607, n_68, A[3]);
  nor g15 (n_1616, A[4], n_117);
  nand g16 (n_1611, A[4], n_117);
  nor g17 (n_1612, A[5], n_116);
  nand g18 (n_1613, A[5], n_116);
  nor g19 (n_1622, n_67, n_115);
  nand g20 (n_1617, n_67, n_115);
  nor g21 (n_1618, n_66, n_114);
  nand g22 (n_1619, n_66, n_114);
  nor g23 (n_1628, n_65, n_113);
  nand g24 (n_1623, n_65, n_113);
  nor g25 (n_1624, n_64, n_112);
  nand g26 (n_1625, n_64, n_112);
  nor g27 (n_1634, n_63, n_111);
  nand g28 (n_1629, n_63, n_111);
  nor g29 (n_1630, n_62, n_110);
  nand g30 (n_1631, n_62, n_110);
  nor g31 (n_1640, n_61, n_109);
  nand g32 (n_1635, n_61, n_109);
  nor g33 (n_1636, n_60, n_108);
  nand g34 (n_1637, n_60, n_108);
  nor g35 (n_1646, n_59, n_107);
  nand g36 (n_1641, n_59, n_107);
  nor g37 (n_1642, n_58, n_106);
  nand g38 (n_1643, n_58, n_106);
  nor g39 (n_1652, n_57, n_105);
  nand g40 (n_1647, n_57, n_105);
  nor g41 (n_1648, n_56, n_104);
  nand g42 (n_1649, n_56, n_104);
  nor g43 (n_1658, n_55, n_103);
  nand g44 (n_1653, n_55, n_103);
  nor g45 (n_1654, n_54, n_102);
  nand g46 (n_1655, n_54, n_102);
  nor g47 (n_1664, n_53, n_101);
  nand g48 (n_1659, n_53, n_101);
  nor g49 (n_1660, n_52, n_100);
  nand g50 (n_1661, n_52, n_100);
  nor g51 (n_1670, n_51, n_99);
  nand g52 (n_1665, n_51, n_99);
  nor g53 (n_1666, n_50, n_98);
  nand g54 (n_1667, n_50, n_98);
  nor g55 (n_1676, n_49, n_97);
  nand g56 (n_1671, n_49, n_97);
  nor g57 (n_1672, n_48, n_96);
  nand g58 (n_1673, n_48, n_96);
  nor g59 (n_1682, n_47, n_95);
  nand g60 (n_1677, n_47, n_95);
  nor g61 (n_1678, n_46, n_94);
  nand g62 (n_1679, n_46, n_94);
  nor g63 (n_1688, n_45, n_93);
  nand g64 (n_1683, n_45, n_93);
  nor g65 (n_1684, n_44, n_92);
  nand g66 (n_1685, n_44, n_92);
  nor g67 (n_1694, n_43, n_91);
  nand g68 (n_1689, n_43, n_91);
  nor g69 (n_1690, n_42, n_90);
  nand g70 (n_1691, n_42, n_90);
  nor g71 (n_1700, n_41, n_89);
  nand g72 (n_1695, n_41, n_89);
  nor g73 (n_1696, n_40, n_88);
  nand g74 (n_1697, n_40, n_88);
  nor g75 (n_1706, n_39, n_87);
  nand g76 (n_1701, n_39, n_87);
  nor g77 (n_1702, n_38, n_86);
  nand g78 (n_1703, n_38, n_86);
  nor g79 (n_1712, n_37, n_85);
  nand g80 (n_1707, n_37, n_85);
  nor g81 (n_1708, n_36, n_84);
  nand g82 (n_1709, n_36, n_84);
  nor g83 (n_1718, n_35, n_83);
  nand g84 (n_1713, n_35, n_83);
  nor g85 (n_1714, n_34, n_82);
  nand g86 (n_1715, n_34, n_82);
  nor g87 (n_1724, n_33, n_81);
  nand g88 (n_1719, n_33, n_81);
  nor g89 (n_1720, n_32, n_80);
  nand g90 (n_1721, n_32, n_80);
  nor g91 (n_1730, n_31, n_79);
  nand g92 (n_1725, n_31, n_79);
  nor g93 (n_1726, n_30, n_78);
  nand g94 (n_1727, n_30, n_78);
  nor g95 (n_1736, n_29, n_77);
  nand g96 (n_1731, n_29, n_77);
  nor g97 (n_1732, n_28, n_76);
  nand g98 (n_1733, n_28, n_76);
  nor g99 (n_1740, n_27, n_75);
  nand g100 (n_1737, n_27, n_75);
  nor g106 (n_1608, n_1605, n_1606);
  nor g110 (n_1614, n_1611, n_1612);
  nor g113 (n_1750, n_1616, n_1612);
  nor g114 (n_1620, n_1617, n_1618);
  nor g117 (n_1752, n_1622, n_1618);
  nor g118 (n_1626, n_1623, n_1624);
  nor g121 (n_1760, n_1628, n_1624);
  nor g122 (n_1632, n_1629, n_1630);
  nor g125 (n_1762, n_1634, n_1630);
  nor g126 (n_1638, n_1635, n_1636);
  nor g129 (n_1770, n_1640, n_1636);
  nor g130 (n_1644, n_1641, n_1642);
  nor g133 (n_1772, n_1646, n_1642);
  nor g134 (n_1650, n_1647, n_1648);
  nor g137 (n_1780, n_1652, n_1648);
  nor g138 (n_1656, n_1653, n_1654);
  nor g141 (n_1782, n_1658, n_1654);
  nor g142 (n_1662, n_1659, n_1660);
  nor g145 (n_1790, n_1664, n_1660);
  nor g146 (n_1668, n_1665, n_1666);
  nor g149 (n_1792, n_1670, n_1666);
  nor g150 (n_1674, n_1671, n_1672);
  nor g153 (n_1800, n_1676, n_1672);
  nor g154 (n_1680, n_1677, n_1678);
  nor g157 (n_1802, n_1682, n_1678);
  nor g158 (n_1686, n_1683, n_1684);
  nor g161 (n_1810, n_1688, n_1684);
  nor g162 (n_1692, n_1689, n_1690);
  nor g165 (n_1812, n_1694, n_1690);
  nor g166 (n_1698, n_1695, n_1696);
  nor g169 (n_1820, n_1700, n_1696);
  nor g170 (n_1704, n_1701, n_1702);
  nor g173 (n_1822, n_1706, n_1702);
  nor g174 (n_1710, n_1707, n_1708);
  nor g177 (n_1830, n_1712, n_1708);
  nor g178 (n_1716, n_1713, n_1714);
  nor g181 (n_1832, n_1718, n_1714);
  nor g182 (n_1722, n_1719, n_1720);
  nor g185 (n_1840, n_1724, n_1720);
  nor g186 (n_1728, n_1725, n_1726);
  nor g189 (n_1842, n_1730, n_1726);
  nor g190 (n_1734, n_1731, n_1732);
  nor g193 (n_1850, n_1736, n_1732);
  nor g203 (n_1748, n_1622, n_1747);
  nand g212 (n_1860, n_1750, n_1752);
  nor g213 (n_1758, n_1634, n_1757);
  nand g222 (n_1867, n_1760, n_1762);
  nor g223 (n_1768, n_1646, n_1767);
  nand g232 (n_1875, n_1770, n_1772);
  nor g233 (n_1778, n_1658, n_1777);
  nand g242 (n_1882, n_1780, n_1782);
  nor g243 (n_1788, n_1670, n_1787);
  nand g252 (n_1890, n_1790, n_1792);
  nor g253 (n_1798, n_1682, n_1797);
  nand g262 (n_1897, n_1800, n_1802);
  nor g263 (n_1808, n_1694, n_1807);
  nand g1776 (n_1905, n_1810, n_1812);
  nor g1777 (n_1818, n_1706, n_1817);
  nand g1786 (n_1912, n_1820, n_1822);
  nor g1787 (n_1828, n_1718, n_1827);
  nand g1796 (n_1920, n_1830, n_1832);
  nor g1797 (n_1838, n_1730, n_1837);
  nand g1806 (n_1927, n_1840, n_1842);
  nor g1807 (n_1848, n_1740, n_1847);
  nand g1814 (n_2131, n_1611, n_1854);
  nand g1816 (n_2133, n_1747, n_1855);
  nand g1819 (n_2136, n_1858, n_1859);
  nand g1822 (n_1935, n_1862, n_1863);
  nor g1823 (n_1865, n_1640, n_1864);
  nor g1826 (n_1945, n_1640, n_1867);
  nor g1832 (n_1873, n_1871, n_1864);
  nor g1835 (n_1951, n_1867, n_1871);
  nor g1836 (n_1877, n_1875, n_1864);
  nor g1839 (n_1954, n_1867, n_1875);
  nor g1840 (n_1880, n_1664, n_1879);
  nor g1843 (n_2034, n_1664, n_1882);
  nor g1849 (n_1888, n_1886, n_1879);
  nor g1852 (n_2040, n_1882, n_1886);
  nor g1853 (n_1892, n_1890, n_1879);
  nor g1856 (n_1960, n_1882, n_1890);
  nor g1857 (n_1895, n_1688, n_1894);
  nor g1860 (n_1973, n_1688, n_1897);
  nor g1866 (n_1903, n_1901, n_1894);
  nor g1869 (n_1983, n_1897, n_1901);
  nor g1870 (n_1907, n_1905, n_1894);
  nor g1873 (n_1988, n_1897, n_1905);
  nor g1874 (n_1910, n_1712, n_1909);
  nor g1877 (n_2086, n_1712, n_1912);
  nor g1883 (n_1918, n_1916, n_1909);
  nor g1886 (n_2092, n_1912, n_1916);
  nor g1887 (n_1922, n_1920, n_1909);
  nor g1890 (n_1996, n_1912, n_1920);
  nor g1891 (n_1925, n_1736, n_1924);
  nor g1894 (n_2009, n_1736, n_1927);
  nor g1900 (n_1933, n_1931, n_1924);
  nor g1903 (n_2019, n_1927, n_1931);
  nand g1906 (n_2140, n_1623, n_1937);
  nand g1907 (n_1938, n_1760, n_1935);
  nand g1908 (n_2142, n_1757, n_1938);
  nand g1911 (n_2145, n_1941, n_1942);
  nand g1914 (n_2148, n_1864, n_1944);
  nand g1915 (n_1947, n_1945, n_1935);
  nand g1916 (n_2151, n_1946, n_1947);
  nand g1917 (n_1950, n_1948, n_1935);
  nand g1918 (n_2153, n_1949, n_1950);
  nand g1919 (n_1953, n_1951, n_1935);
  nand g1920 (n_2156, n_1952, n_1953);
  nand g1921 (n_1956, n_1954, n_1935);
  nand g1922 (n_2024, n_1955, n_1956);
  nor g1923 (n_1958, n_1676, n_1957);
  nand g1932 (n_2048, n_1800, n_1960);
  nor g1933 (n_1967, n_1965, n_1957);
  nor g1938 (n_1970, n_1897, n_1957);
  nand g1947 (n_2060, n_1960, n_1973);
  nand g1952 (n_2064, n_1960, n_1978);
  nand g1957 (n_2068, n_1960, n_1983);
  nand g1962 (n_2072, n_1960, n_1988);
  nor g1963 (n_1994, n_1724, n_1993);
  nand g1972 (n_2100, n_1840, n_1996);
  nor g1973 (n_2003, n_2001, n_1993);
  nor g1978 (n_2006, n_1927, n_1993);
  nand g1987 (n_2112, n_1996, n_2009);
  nand g1992 (n_2116, n_1996, n_2014);
  nand g1997 (n_2120, n_1996, n_2019);
  nand g2000 (n_2160, n_1647, n_2026);
  nand g2001 (n_2027, n_1780, n_2024);
  nand g2002 (n_2162, n_1777, n_2027);
  nand g2005 (n_2165, n_2030, n_2031);
  nand g2008 (n_2168, n_1879, n_2033);
  nand g2009 (n_2036, n_2034, n_2024);
  nand g2010 (n_2171, n_2035, n_2036);
  nand g2011 (n_2039, n_2037, n_2024);
  nand g2012 (n_2173, n_2038, n_2039);
  nand g2013 (n_2042, n_2040, n_2024);
  nand g2014 (n_2176, n_2041, n_2042);
  nand g2015 (n_2043, n_1960, n_2024);
  nand g2016 (n_2178, n_1957, n_2043);
  nand g2019 (n_2181, n_2046, n_2047);
  nand g2022 (n_2183, n_2050, n_2051);
  nand g2025 (n_2186, n_2054, n_2055);
  nand g2028 (n_2189, n_2058, n_2059);
  nand g2031 (n_2192, n_2062, n_2063);
  nand g2034 (n_2194, n_2066, n_2067);
  nand g2037 (n_2197, n_2070, n_2071);
  nand g2040 (n_2076, n_2074, n_2075);
  nand g2043 (n_2201, n_1695, n_2078);
  nand g2044 (n_2079, n_1820, n_2076);
  nand g2045 (n_2203, n_1817, n_2079);
  nand g2048 (n_2206, n_2082, n_2083);
  nand g2051 (n_2209, n_1909, n_2085);
  nand g2052 (n_2088, n_2086, n_2076);
  nand g2053 (n_2212, n_2087, n_2088);
  nand g2054 (n_2091, n_2089, n_2076);
  nand g2055 (n_2214, n_2090, n_2091);
  nand g2056 (n_2094, n_2092, n_2076);
  nand g2057 (n_2217, n_2093, n_2094);
  nand g2058 (n_2095, n_1996, n_2076);
  nand g2059 (n_2219, n_1993, n_2095);
  nand g2062 (n_2222, n_2098, n_2099);
  nand g2065 (n_2224, n_2102, n_2103);
  nand g2068 (n_2227, n_2106, n_2107);
  nand g2071 (n_2230, n_2110, n_2111);
  nand g2074 (n_2233, n_2114, n_2115);
  nand g2077 (n_2235, n_2118, n_2119);
  nand g2080 (n_2238, n_2122, n_2123);
  xnor g2092 (Z[5], n_2131, n_2132);
  xnor g2094 (Z[6], n_2133, n_2134);
  xnor g2097 (Z[7], n_2136, n_2137);
  xnor g2099 (Z[8], n_1935, n_2138);
  xnor g2102 (Z[9], n_2140, n_2141);
  xnor g2104 (Z[10], n_2142, n_2143);
  xnor g2107 (Z[11], n_2145, n_2146);
  xnor g2110 (Z[12], n_2148, n_2149);
  xnor g2113 (Z[13], n_2151, n_2152);
  xnor g2115 (Z[14], n_2153, n_2154);
  xnor g2118 (Z[15], n_2156, n_2157);
  xnor g2120 (Z[16], n_2024, n_2158);
  xnor g2123 (Z[17], n_2160, n_2161);
  xnor g2125 (Z[18], n_2162, n_2163);
  xnor g2128 (Z[19], n_2165, n_2166);
  xnor g2131 (Z[20], n_2168, n_2169);
  xnor g2134 (Z[21], n_2171, n_2172);
  xnor g2136 (Z[22], n_2173, n_2174);
  xnor g2139 (Z[23], n_2176, n_2177);
  xnor g2141 (Z[24], n_2178, n_2179);
  xnor g2144 (Z[25], n_2181, n_2182);
  xnor g2146 (Z[26], n_2183, n_2184);
  xnor g2149 (Z[27], n_2186, n_2187);
  xnor g2152 (Z[28], n_2189, n_2190);
  xnor g2155 (Z[29], n_2192, n_2193);
  xnor g2157 (Z[30], n_2194, n_2195);
  xnor g2160 (Z[31], n_2197, n_2198);
  xnor g2162 (Z[32], n_2076, n_2199);
  xnor g2165 (Z[33], n_2201, n_2202);
  xnor g2167 (Z[34], n_2203, n_2204);
  xnor g2170 (Z[35], n_2206, n_2207);
  xnor g2173 (Z[36], n_2209, n_2210);
  xnor g2176 (Z[37], n_2212, n_2213);
  xnor g2178 (Z[38], n_2214, n_2215);
  xnor g2181 (Z[39], n_2217, n_2218);
  xnor g2183 (Z[40], n_2219, n_2220);
  xnor g2186 (Z[41], n_2222, n_2223);
  xnor g2188 (Z[42], n_2224, n_2225);
  xnor g2191 (Z[43], n_2227, n_2228);
  xnor g2194 (Z[44], n_2230, n_2231);
  xnor g2197 (Z[45], n_2233, n_2234);
  xnor g2199 (Z[46], n_2235, n_2236);
  xnor g2202 (Z[47], n_2238, n_2239);
  or g2215 (n_1045, A[1], wc);
  not gc (wc, n_171);
  or g2216 (n_1046, A[1], wc0);
  not gc0 (wc0, A[2]);
  or g2217 (n_1070, wc1, A[24]);
  not gc1 (wc1, A[18]);
  or g2218 (n_1089, A[2], wc2);
  not gc2 (wc2, A[3]);
  or g2219 (n_1090, wc3, A[2]);
  not gc3 (wc3, A[1]);
  or g2220 (n_1157, wc4, A[24]);
  not gc4 (wc4, A[20]);
  xnor g2221 (n_1195, A[24], A[21]);
  or g2222 (n_1196, wc5, A[24]);
  not gc5 (wc5, A[21]);
  xnor g2223 (n_1215, A[6], A[5]);
  or g2224 (n_1216, A[5], wc6);
  not gc6 (wc6, A[6]);
  or g2225 (n_1253, A[6], wc7);
  not gc7 (wc7, A[7]);
  or g2226 (n_1254, wc8, A[6]);
  not gc8 (wc8, A[5]);
  or g2228 (n_1356, wc9, A[10]);
  not gc9 (wc9, A[9]);
  or g2229 (n_1357, A[10], wc10);
  not gc10 (wc10, A[14]);
  or g2231 (n_1385, wc11, A[11]);
  not gc11 (wc11, A[10]);
  or g2232 (n_1421, wc12, A[24]);
  not gc12 (wc12, A[19]);
  xnor g2233 (n_1447, A[24], A[20]);
  or g2235 (n_1464, wc13, A[14]);
  not gc13 (wc13, A[13]);
  or g2236 (n_1465, A[14], wc14);
  not gc14 (wc14, A[18]);
  or g2237 (n_1486, A[14], wc15);
  not gc15 (wc15, A[15]);
  or g2239 (n_1556, wc16, A[19]);
  not gc16 (wc16, A[18]);
  xnor g2240 (n_1563, A[24], A[19]);
  or g2242 (n_1584, A[21], wc17);
  not gc17 (wc17, A[22]);
  or g2244 (n_1588, A[22], wc18);
  not gc18 (wc18, A[23]);
  or g2245 (n_1589, wc19, A[22]);
  not gc19 (wc19, A[21]);
  xnor g2246 (n_1591, A[24], A[23]);
  or g2247 (n_1592, wc20, A[24]);
  not gc20 (wc20, A[23]);
  or g2248 (n_1594, wc21, A[24]);
  not gc21 (wc21, A[22]);
  xnor g2249 (n_350, n_1043, A[1]);
  xnor g2250 (n_373, n_1087, A[2]);
  xnor g2251 (n_454, n_1251, A[6]);
  xnor g2252 (n_505, n_1219, A[14]);
  or g2253 (n_533, A[10], wc22);
  not gc22 (wc22, n_1385);
  or g2254 (n_545, A[11], wc23);
  not gc23 (wc23, n_746);
  or g2255 (n_1422, A[24], wc24);
  not gc24 (wc24, n_534);
  xnor g2256 (n_559, n_1223, A[18]);
  xnor g2257 (n_570, n_1387, A[14]);
  nand g2258 (n_579, n_945, n_1486);
  xnor g2259 (n_1543, n_560, A[18]);
  or g2260 (n_1544, A[18], wc25);
  not gc25 (wc25, n_560);
  xnor g2261 (n_606, n_1391, n_573);
  or g2262 (n_1558, A[19], wc26);
  not gc26 (wc26, n_573);
  xnor g2263 (n_76, n_1271, A[21]);
  or g2265 (n_2125, wc27, n_1610);
  not gc27 (wc27, n_1605);
  xnor g2266 (n_525, n_1391, A[11]);
  or g2267 (n_1393, A[11], wc28);
  not gc28 (wc28, A[18]);
  or g2268 (n_1394, A[11], wc29);
  not gc29 (wc29, A[19]);
  xnor g2269 (n_538, n_1419, A[24]);
  or g2270 (n_1509, A[24], wc30);
  not gc30 (wc30, n_579);
  or g2271 (n_1530, A[24], wc31);
  not gc31 (wc31, n_587);
  xnor g2272 (n_29, n_1071, n_443);
  or g2273 (n_1585, A[21], wc32);
  not gc32 (wc32, n_443);
  and g2274 (n_1745, wc33, n_1607);
  not gc33 (wc33, n_1608);
  or g2275 (n_2128, wc34, n_1606);
  not gc34 (wc34, n_1607);
  xnor g2276 (n_582, n_1507, A[24]);
  and g2277 (n_1738, wc35, n_74);
  not gc35 (wc35, A[24]);
  or g2278 (n_1739, wc36, n_74);
  not gc36 (wc36, A[24]);
  not g2279 (Z[2], n_2125);
  or g2280 (n_1217, A[5], wc37);
  not gc37 (wc37, n_434);
  or g2281 (n_1450, A[24], wc38);
  not gc38 (wc38, n_546);
  or g2282 (n_1546, A[18], wc39);
  not gc39 (wc39, n_597);
  or g2285 (n_2129, wc40, n_1616);
  not gc40 (wc40, n_1611);
  or g2286 (n_2236, wc41, n_1740);
  not gc41 (wc41, n_1737);
  or g2287 (n_1337, A[24], wc42);
  not gc42 (wc42, n_491);
  and g2288 (n_1747, wc43, n_1613);
  not gc43 (wc43, n_1614);
  or g2289 (n_1854, n_1616, n_1745);
  or g2290 (n_1855, n_1745, wc44);
  not gc44 (wc44, n_1750);
  xor g2291 (Z[3], n_1605, n_2128);
  xor g2292 (Z[4], n_1745, n_2129);
  or g2293 (n_2132, wc45, n_1612);
  not gc45 (wc45, n_1613);
  or g2294 (n_2239, wc46, n_1738);
  not gc46 (wc46, n_1739);
  xnor g2295 (n_1335, n_490, A[24]);
  or g2296 (n_1336, A[24], wc47);
  not gc47 (wc47, n_490);
  and g2297 (n_1754, wc48, n_1619);
  not gc48 (wc48, n_1620);
  or g2298 (n_1856, wc49, n_1622);
  not gc49 (wc49, n_1750);
  or g2299 (n_2134, wc50, n_1622);
  not gc50 (wc50, n_1617);
  or g2300 (n_2137, wc51, n_1618);
  not gc51 (wc51, n_1619);
  or g2301 (n_2234, wc52, n_1732);
  not gc52 (wc52, n_1733);
  and g2302 (n_1858, wc53, n_1617);
  not gc53 (wc53, n_1748);
  and g2303 (n_1755, wc54, n_1752);
  not gc54 (wc54, n_1747);
  or g2304 (n_2138, wc55, n_1628);
  not gc55 (wc55, n_1623);
  or g2305 (n_2228, wc56, n_1726);
  not gc56 (wc56, n_1727);
  or g2306 (n_1069, A[24], wc57);
  not gc57 (wc57, n_358);
  xnor g2307 (n_1155, n_401, A[24]);
  or g2308 (n_1156, A[24], wc58);
  not gc58 (wc58, n_401);
  xnor g2309 (n_1303, n_475, A[24]);
  or g2310 (n_1304, A[24], wc59);
  not gc59 (wc59, n_475);
  and g2311 (n_1757, wc60, n_1625);
  not gc60 (wc60, n_1626);
  and g2312 (n_1847, wc61, n_1733);
  not gc61 (wc61, n_1734);
  and g2313 (n_1862, wc62, n_1754);
  not gc62 (wc62, n_1755);
  or g2314 (n_1931, wc63, n_1740);
  not gc63 (wc63, n_1850);
  or g2315 (n_1859, n_1745, n_1856);
  or g2316 (n_1863, n_1860, n_1745);
  or g2317 (n_2141, wc64, n_1624);
  not gc64 (wc64, n_1625);
  or g2318 (n_2231, wc65, n_1736);
  not gc65 (wc65, n_1731);
  xnor g2319 (n_364, n_1067, A[24]);
  or g2320 (n_1939, wc66, n_1634);
  not gc66 (wc66, n_1760);
  or g2321 (n_2143, wc67, n_1634);
  not gc67 (wc67, n_1629);
  and g2322 (n_1837, wc68, n_1721);
  not gc68 (wc68, n_1722);
  and g2323 (n_1844, wc69, n_1727);
  not gc69 (wc69, n_1728);
  and g2324 (n_1941, wc70, n_1629);
  not gc70 (wc70, n_1758);
  or g2325 (n_2001, wc71, n_1730);
  not gc71 (wc71, n_1840);
  and g2326 (n_1932, wc72, n_1737);
  not gc72 (wc72, n_1848);
  or g2327 (n_1937, wc73, n_1628);
  not gc73 (wc73, n_1935);
  or g2328 (n_2152, wc74, n_1636);
  not gc74 (wc74, n_1637);
  or g2329 (n_2218, wc75, n_1714);
  not gc75 (wc75, n_1715);
  or g2330 (n_2220, wc76, n_1724);
  not gc76 (wc76, n_1719);
  or g2331 (n_2223, wc77, n_1720);
  not gc77 (wc77, n_1721);
  or g2332 (n_2225, wc78, n_1730);
  not gc78 (wc78, n_1725);
  and g2333 (n_1764, wc79, n_1631);
  not gc79 (wc79, n_1632);
  and g2334 (n_1767, wc80, n_1637);
  not gc80 (wc80, n_1638);
  and g2335 (n_1845, wc81, n_1842);
  not gc81 (wc81, n_1837);
  and g2336 (n_2014, wc82, n_1850);
  not gc82 (wc82, n_1927);
  or g2337 (n_1942, n_1939, wc83);
  not gc83 (wc83, n_1935);
  or g2338 (n_2146, wc84, n_1630);
  not gc84 (wc84, n_1631);
  or g2339 (n_2149, wc85, n_1640);
  not gc85 (wc85, n_1635);
  and g2340 (n_1827, wc86, n_1709);
  not gc86 (wc86, n_1710);
  and g2341 (n_1834, wc87, n_1715);
  not gc87 (wc87, n_1716);
  and g2342 (n_1765, wc88, n_1762);
  not gc88 (wc88, n_1757);
  or g2343 (n_1871, wc89, n_1646);
  not gc89 (wc89, n_1770);
  or g2344 (n_1916, wc90, n_1718);
  not gc90 (wc90, n_1830);
  and g2345 (n_2002, wc91, n_1725);
  not gc91 (wc91, n_1838);
  and g2346 (n_1924, wc92, n_1844);
  not gc92 (wc92, n_1845);
  and g2347 (n_1948, wc93, n_1770);
  not gc93 (wc93, n_1867);
  or g2348 (n_2154, wc94, n_1646);
  not gc94 (wc94, n_1641);
  or g2349 (n_2210, wc95, n_1712);
  not gc95 (wc95, n_1707);
  or g2350 (n_2213, wc96, n_1708);
  not gc96 (wc96, n_1709);
  or g2351 (n_2215, wc97, n_1718);
  not gc97 (wc97, n_1713);
  and g2352 (n_1774, wc98, n_1643);
  not gc98 (wc98, n_1644);
  and g2353 (n_1864, wc99, n_1764);
  not gc99 (wc99, n_1765);
  and g2354 (n_1872, wc100, n_1641);
  not gc100 (wc100, n_1768);
  and g2355 (n_1835, wc101, n_1832);
  not gc101 (wc101, n_1827);
  and g2356 (n_1929, wc102, n_1850);
  not gc102 (wc102, n_1924);
  or g2357 (n_1944, wc103, n_1867);
  not gc103 (wc103, n_1935);
  or g2358 (n_2157, wc104, n_1642);
  not gc104 (wc104, n_1643);
  and g2359 (n_1777, wc105, n_1649);
  not gc105 (wc105, n_1650);
  and g2360 (n_1775, wc106, n_1772);
  not gc106 (wc106, n_1767);
  and g2361 (n_1917, wc107, n_1713);
  not gc107 (wc107, n_1828);
  and g2362 (n_1921, wc108, n_1834);
  not gc108 (wc108, n_1835);
  and g2363 (n_1869, wc109, n_1770);
  not gc109 (wc109, n_1864);
  and g2364 (n_2011, wc110, n_1731);
  not gc110 (wc110, n_1925);
  and g2365 (n_2016, wc111, n_1847);
  not gc111 (wc111, n_1929);
  and g2366 (n_2021, n_1932, wc112);
  not gc112 (wc112, n_1933);
  or g2367 (n_2158, wc113, n_1652);
  not gc113 (wc113, n_1647);
  or g2368 (n_2161, wc114, n_1648);
  not gc114 (wc114, n_1649);
  and g2369 (n_1876, wc115, n_1774);
  not gc115 (wc115, n_1775);
  and g2370 (n_1946, wc116, n_1635);
  not gc116 (wc116, n_1865);
  and g2371 (n_1949, wc117, n_1767);
  not gc117 (wc117, n_1869);
  and g2372 (n_1952, n_1872, wc118);
  not gc118 (wc118, n_1873);
  or g2373 (n_2169, wc119, n_1664);
  not gc119 (wc119, n_1659);
  and g2374 (n_1784, wc120, n_1655);
  not gc120 (wc120, n_1656);
  and g2375 (n_1787, wc121, n_1661);
  not gc121 (wc121, n_1662);
  and g2376 (n_1794, wc122, n_1667);
  not gc122 (wc122, n_1668);
  and g2377 (n_1824, wc123, n_1703);
  not gc123 (wc123, n_1704);
  and g2378 (n_2030, wc124, n_1653);
  not gc124 (wc124, n_1778);
  or g2379 (n_2028, wc125, n_1658);
  not gc125 (wc125, n_1780);
  or g2380 (n_1886, wc126, n_1670);
  not gc126 (wc126, n_1790);
  or g2381 (n_2163, wc127, n_1658);
  not gc127 (wc127, n_1653);
  or g2382 (n_2166, wc128, n_1654);
  not gc128 (wc128, n_1655);
  or g2383 (n_2172, wc129, n_1660);
  not gc129 (wc129, n_1661);
  or g2384 (n_2174, wc130, n_1670);
  not gc130 (wc130, n_1665);
  or g2385 (n_2177, wc131, n_1666);
  not gc131 (wc131, n_1667);
  or g2386 (n_2179, wc132, n_1676);
  not gc132 (wc132, n_1671);
  or g2387 (n_2204, wc133, n_1706);
  not gc133 (wc133, n_1701);
  or g2388 (n_2207, wc134, n_1702);
  not gc134 (wc134, n_1703);
  and g2389 (n_1785, wc135, n_1782);
  not gc135 (wc135, n_1777);
  and g2390 (n_1795, wc136, n_1792);
  not gc136 (wc136, n_1787);
  and g2391 (n_1955, n_1876, wc137);
  not gc137 (wc137, n_1877);
  and g2392 (n_2037, wc138, n_1790);
  not gc138 (wc138, n_1882);
  and g2393 (n_1797, wc139, n_1673);
  not gc139 (wc139, n_1674);
  and g2394 (n_1804, wc140, n_1679);
  not gc140 (wc140, n_1680);
  and g2395 (n_1807, wc141, n_1685);
  not gc141 (wc141, n_1686);
  and g2396 (n_1814, wc142, n_1691);
  not gc142 (wc142, n_1692);
  and g2397 (n_1817, wc143, n_1697);
  not gc143 (wc143, n_1698);
  and g2398 (n_1879, wc144, n_1784);
  not gc144 (wc144, n_1785);
  and g2399 (n_1887, wc145, n_1665);
  not gc145 (wc145, n_1788);
  and g2400 (n_1891, wc146, n_1794);
  not gc146 (wc146, n_1795);
  or g2401 (n_1965, wc147, n_1682);
  not gc147 (wc147, n_1800);
  or g2402 (n_1901, wc148, n_1694);
  not gc148 (wc148, n_1810);
  or g2403 (n_2080, wc149, n_1706);
  not gc149 (wc149, n_1820);
  or g2404 (n_2044, wc150, n_1676);
  not gc150 (wc150, n_1960);
  or g2405 (n_2182, wc151, n_1672);
  not gc151 (wc151, n_1673);
  or g2406 (n_2184, wc152, n_1682);
  not gc152 (wc152, n_1677);
  or g2407 (n_2187, wc153, n_1678);
  not gc153 (wc153, n_1679);
  or g2408 (n_2190, wc154, n_1688);
  not gc154 (wc154, n_1683);
  or g2409 (n_2193, wc155, n_1684);
  not gc155 (wc155, n_1685);
  or g2410 (n_2195, wc156, n_1694);
  not gc156 (wc156, n_1689);
  or g2411 (n_2198, wc157, n_1690);
  not gc157 (wc157, n_1691);
  or g2412 (n_2199, wc158, n_1700);
  not gc158 (wc158, n_1695);
  or g2413 (n_2202, wc159, n_1696);
  not gc159 (wc159, n_1697);
  and g2414 (n_1805, wc160, n_1802);
  not gc160 (wc160, n_1797);
  and g2415 (n_1815, wc161, n_1812);
  not gc161 (wc161, n_1807);
  and g2416 (n_1825, wc162, n_1822);
  not gc162 (wc162, n_1817);
  and g2417 (n_1884, wc163, n_1790);
  not gc163 (wc163, n_1879);
  and g2418 (n_1978, wc164, n_1810);
  not gc164 (wc164, n_1897);
  and g2419 (n_2089, wc165, n_1830);
  not gc165 (wc165, n_1912);
  or g2420 (n_2026, wc166, n_1652);
  not gc166 (wc166, n_2024);
  or g2421 (n_2031, n_2028, wc167);
  not gc167 (wc167, n_2024);
  or g2422 (n_2033, wc168, n_1882);
  not gc168 (wc168, n_2024);
  and g2423 (n_1966, wc169, n_1677);
  not gc169 (wc169, n_1798);
  and g2424 (n_1894, wc170, n_1804);
  not gc170 (wc170, n_1805);
  and g2425 (n_1902, wc171, n_1689);
  not gc171 (wc171, n_1808);
  and g2426 (n_1906, wc172, n_1814);
  not gc172 (wc172, n_1815);
  and g2427 (n_2082, wc173, n_1701);
  not gc173 (wc173, n_1818);
  and g2428 (n_1909, wc174, n_1824);
  not gc174 (wc174, n_1825);
  and g2429 (n_2035, wc175, n_1659);
  not gc175 (wc175, n_1880);
  and g2430 (n_2038, wc176, n_1787);
  not gc176 (wc176, n_1884);
  and g2431 (n_2041, n_1887, wc177);
  not gc177 (wc177, n_1888);
  and g2432 (n_1957, n_1891, wc178);
  not gc178 (wc178, n_1892);
  or g2433 (n_2052, n_1965, wc179);
  not gc179 (wc179, n_1960);
  or g2434 (n_2056, wc180, n_1897);
  not gc180 (wc180, n_1960);
  or g2435 (n_2096, wc181, n_1724);
  not gc181 (wc181, n_1996);
  or g2436 (n_2104, n_2001, wc182);
  not gc182 (wc182, n_1996);
  or g2437 (n_2108, wc183, n_1927);
  not gc183 (wc183, n_1996);
  or g2438 (n_2047, n_2044, wc184);
  not gc184 (wc184, n_2024);
  or g2439 (n_2051, n_2048, wc185);
  not gc185 (wc185, n_2024);
  and g2440 (n_1899, wc186, n_1810);
  not gc186 (wc186, n_1894);
  and g2441 (n_1914, wc187, n_1830);
  not gc187 (wc187, n_1909);
  and g2442 (n_1963, wc188, n_1800);
  not gc188 (wc188, n_1957);
  and g2443 (n_1976, wc189, n_1973);
  not gc189 (wc189, n_1957);
  and g2444 (n_1981, wc190, n_1978);
  not gc190 (wc190, n_1957);
  and g2445 (n_1986, wc191, n_1983);
  not gc191 (wc191, n_1957);
  and g2446 (n_1991, wc192, n_1988);
  not gc192 (wc192, n_1957);
  and g2447 (n_1975, wc193, n_1683);
  not gc193 (wc193, n_1895);
  and g2448 (n_1980, wc194, n_1807);
  not gc194 (wc194, n_1899);
  and g2449 (n_1985, n_1902, wc195);
  not gc195 (wc195, n_1903);
  and g2450 (n_1990, n_1906, wc196);
  not gc196 (wc196, n_1907);
  and g2451 (n_2087, wc197, n_1707);
  not gc197 (wc197, n_1910);
  and g2452 (n_2090, wc198, n_1827);
  not gc198 (wc198, n_1914);
  and g2453 (n_2093, n_1917, wc199);
  not gc199 (wc199, n_1918);
  and g2454 (n_1993, n_1921, wc200);
  not gc200 (wc200, n_1922);
  and g2455 (n_2046, wc201, n_1671);
  not gc201 (wc201, n_1958);
  and g2456 (n_2050, wc202, n_1797);
  not gc202 (wc202, n_1963);
  and g2457 (n_2054, n_1966, wc203);
  not gc203 (wc203, n_1967);
  and g2458 (n_2058, n_1894, wc204);
  not gc204 (wc204, n_1970);
  or g2459 (n_2055, n_2052, wc205);
  not gc205 (wc205, n_2024);
  or g2460 (n_2059, n_2056, wc206);
  not gc206 (wc206, n_2024);
  or g2461 (n_2063, n_2060, wc207);
  not gc207 (wc207, n_2024);
  or g2462 (n_2067, n_2064, wc208);
  not gc208 (wc208, n_2024);
  or g2463 (n_2071, n_2068, wc209);
  not gc209 (wc209, n_2024);
  or g2464 (n_2075, n_2072, wc210);
  not gc210 (wc210, n_2024);
  and g2465 (n_1999, wc211, n_1840);
  not gc211 (wc211, n_1993);
  and g2466 (n_2012, wc212, n_2009);
  not gc212 (wc212, n_1993);
  and g2467 (n_2017, wc213, n_2014);
  not gc213 (wc213, n_1993);
  and g2468 (n_2022, wc214, n_2019);
  not gc214 (wc214, n_1993);
  and g2469 (n_2062, n_1975, wc215);
  not gc215 (wc215, n_1976);
  and g2470 (n_2066, n_1980, wc216);
  not gc216 (wc216, n_1981);
  and g2471 (n_2070, n_1985, wc217);
  not gc217 (wc217, n_1986);
  and g2472 (n_2074, n_1990, wc218);
  not gc218 (wc218, n_1991);
  and g2473 (n_2098, wc219, n_1719);
  not gc219 (wc219, n_1994);
  and g2474 (n_2102, wc220, n_1837);
  not gc220 (wc220, n_1999);
  and g2475 (n_2106, n_2002, wc221);
  not gc221 (wc221, n_2003);
  and g2476 (n_2110, n_1924, wc222);
  not gc222 (wc222, n_2006);
  and g2477 (n_2114, wc223, n_2011);
  not gc223 (wc223, n_2012);
  and g2478 (n_2118, wc224, n_2016);
  not gc224 (wc224, n_2017);
  and g2479 (n_2122, wc225, n_2021);
  not gc225 (wc225, n_2022);
  or g2480 (n_2078, wc226, n_1700);
  not gc226 (wc226, n_2076);
  or g2481 (n_2083, n_2080, wc227);
  not gc227 (wc227, n_2076);
  or g2482 (n_2085, wc228, n_1912);
  not gc228 (wc228, n_2076);
  or g2483 (n_2099, n_2096, wc229);
  not gc229 (wc229, n_2076);
  or g2484 (n_2103, wc230, n_2100);
  not gc230 (wc230, n_2076);
  or g2485 (n_2107, n_2104, wc231);
  not gc231 (wc231, n_2076);
  or g2486 (n_2111, n_2108, wc232);
  not gc232 (wc232, n_2076);
  or g2487 (n_2115, wc233, n_2112);
  not gc233 (wc233, n_2076);
  or g2488 (n_2119, wc234, n_2116);
  not gc234 (wc234, n_2076);
  or g2489 (n_2123, wc235, n_2120);
  not gc235 (wc235, n_2076);
endmodule

module mult_signed_const_5753_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_5753_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_6020_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_74, n_75, n_76, n_77;
  wire n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85;
  wire n_86, n_87, n_88, n_89, n_90, n_91, n_92, n_93;
  wire n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101;
  wire n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109;
  wire n_110, n_111, n_112, n_113, n_114, n_115, n_116, n_117;
  wire n_118, n_119, n_171, n_172, n_173, n_174, n_176, n_179;
  wire n_180, n_181, n_184, n_185, n_189, n_190, n_195, n_196;
  wire n_197, n_201, n_202, n_203, n_204, n_205, n_208, n_210;
  wire n_211, n_212, n_213, n_218, n_219, n_220, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_232, n_234, n_235, n_236;
  wire n_237, n_238, n_239, n_240, n_243, n_244, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_258, n_259, n_261;
  wire n_262, n_263, n_271, n_272, n_273, n_274, n_275, n_276;
  wire n_277, n_278, n_284, n_285, n_286, n_287, n_288, n_289;
  wire n_290, n_291, n_292, n_293, n_294, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_315, n_316, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_327, n_333, n_335;
  wire n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_346, n_350, n_352, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_372, n_373, n_374, n_375, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_393, n_394, n_395;
  wire n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403;
  wire n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411;
  wire n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419;
  wire n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_431, n_434, n_435, n_436, n_437;
  wire n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445;
  wire n_446, n_447, n_448, n_449, n_450, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_488, n_489, n_490, n_491;
  wire n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499;
  wire n_500, n_501, n_504, n_505, n_506, n_507, n_508, n_509;
  wire n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_533, n_534, n_535, n_536, n_537;
  wire n_538, n_539, n_540, n_541, n_542, n_543, n_544, n_545;
  wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
  wire n_554, n_555, n_558, n_559, n_560, n_561, n_562, n_563;
  wire n_564, n_565, n_566, n_570, n_571, n_572, n_573, n_574;
  wire n_575, n_576, n_577, n_579, n_580, n_582, n_583, n_584;
  wire n_585, n_586, n_587, n_589, n_590, n_591, n_592, n_593;
  wire n_596, n_597, n_599, n_600, n_605, n_606, n_607, n_610;
  wire n_611, n_612, n_614, n_615, n_618, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_642, n_643, n_647, n_648, n_649, n_650, n_651, n_652;
  wire n_653, n_654, n_659, n_660, n_661, n_662, n_663, n_664;
  wire n_665, n_666, n_671, n_672, n_673, n_674, n_675, n_676;
  wire n_677, n_678, n_685, n_686, n_687, n_688, n_689, n_690;
  wire n_691, n_692, n_693, n_694, n_699, n_700, n_701, n_702;
  wire n_703, n_704, n_705, n_706, n_707, n_708, n_709, n_710;
  wire n_711, n_712, n_713, n_714, n_723, n_724, n_725, n_726;
  wire n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734;
  wire n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748;
  wire n_749, n_750, n_751, n_752, n_753, n_754, n_765, n_766;
  wire n_767, n_768, n_769, n_770, n_771, n_772, n_773, n_774;
  wire n_775, n_776, n_777, n_778, n_786, n_787, n_791, n_792;
  wire n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800;
  wire n_801, n_802, n_803, n_804, n_805, n_806, n_811, n_817;
  wire n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825;
  wire n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833;
  wire n_834, n_847, n_848, n_849, n_850, n_851, n_852, n_853;
  wire n_854, n_855, n_856, n_857, n_858, n_859, n_860, n_861;
  wire n_862, n_873, n_874, n_875, n_876, n_877, n_878, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_894, n_903, n_904, n_906;
  wire n_907, n_908, n_909, n_911, n_912, n_913, n_914, n_915;
  wire n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923;
  wire n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_941;
  wire n_942, n_943, n_944, n_946, n_947, n_948, n_949, n_950;
  wire n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958;
  wire n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966;
  wire n_973, n_974, n_975, n_976, n_979, n_981, n_982, n_983;
  wire n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991;
  wire n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999;
  wire n_1000, n_1001, n_1002, n_1015, n_1017, n_1018, n_1019, n_1020;
  wire n_1021, n_1022, n_1023, n_1025, n_1026, n_1027, n_1028, n_1029;
  wire n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037;
  wire n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1045, n_1046;
  wire n_1047, n_1048, n_1050, n_1055, n_1056, n_1057, n_1059, n_1060;
  wire n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068;
  wire n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
  wire n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084;
  wire n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092;
  wire n_1093, n_1094, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103;
  wire n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111;
  wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119;
  wire n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127;
  wire n_1128, n_1129, n_1130, n_1133, n_1134, n_1135, n_1136, n_1137;
  wire n_1138, n_1139, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147;
  wire n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155;
  wire n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164;
  wire n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172;
  wire n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180;
  wire n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188;
  wire n_1189, n_1190, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198;
  wire n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206;
  wire n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214;
  wire n_1215, n_1216, n_1217, n_1219, n_1220, n_1221, n_1223, n_1224;
  wire n_1225, n_1226, n_1227, n_1228, n_1229, n_1231, n_1232, n_1234;
  wire n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242;
  wire n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250;
  wire n_1253, n_1255, n_1256, n_1257, n_1259, n_1260, n_1261, n_1262;
  wire n_1263, n_1264, n_1265, n_1267, n_1268, n_1270, n_1271, n_1272;
  wire n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280;
  wire n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1291, n_1292;
  wire n_1294, n_1295, n_1296, n_1297, n_1302, n_1303, n_1304, n_1305;
  wire n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313;
  wire n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321;
  wire n_1322, n_1326, n_1327, n_1329, n_1330, n_1331, n_1332, n_1333;
  wire n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342;
  wire n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350;
  wire n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1359, n_1360;
  wire n_1362, n_1363, n_1364, n_1366, n_1367, n_1368, n_1369, n_1370;
  wire n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378;
  wire n_1379, n_1380, n_1381, n_1382, n_1383, n_1387, n_1388, n_1389;
  wire n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1397, n_1398;
  wire n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406;
  wire n_1407, n_1408, n_1409, n_1410, n_1418, n_1422, n_1423, n_1424;
  wire n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432;
  wire n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1443, n_1447;
  wire n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455;
  wire n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463;
  wire n_1464, n_1465, n_1466, n_1467, n_1468, n_1470, n_1471, n_1472;
  wire n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480;
  wire n_1481, n_1482, n_1486, n_1487, n_1489, n_1490, n_1491, n_1492;
  wire n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500;
  wire n_1501, n_1502, n_1505, n_1511, n_1512, n_1513, n_1514, n_1515;
  wire n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1526;
  wire n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536;
  wire n_1537, n_1538, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548;
  wire n_1549, n_1550, n_1551, n_1554, n_1556, n_1557, n_1558, n_1559;
  wire n_1560, n_1561, n_1562, n_1567, n_1569, n_1570, n_1571, n_1572;
  wire n_1573, n_1574, n_1575, n_1578, n_1579, n_1580, n_1581, n_1582;
  wire n_1583, n_1584, n_1585, n_1586, n_1588, n_1589, n_1590, n_1591;
  wire n_1592, n_1594, n_1605, n_1606, n_1607, n_1608, n_1610, n_1611;
  wire n_1612, n_1613, n_1614, n_1616, n_1617, n_1618, n_1619, n_1620;
  wire n_1622, n_1623, n_1624, n_1625, n_1626, n_1628, n_1629, n_1630;
  wire n_1631, n_1632, n_1634, n_1635, n_1636, n_1637, n_1638, n_1640;
  wire n_1641, n_1642, n_1643, n_1644, n_1646, n_1647, n_1648, n_1649;
  wire n_1650, n_1652, n_1653, n_1654, n_1655, n_1656, n_1658, n_1659;
  wire n_1660, n_1661, n_1662, n_1664, n_1665, n_1666, n_1667, n_1668;
  wire n_1670, n_1671, n_1672, n_1673, n_1674, n_1676, n_1677, n_1678;
  wire n_1679, n_1680, n_1682, n_1683, n_1684, n_1685, n_1686, n_1688;
  wire n_1689, n_1690, n_1691, n_1692, n_1694, n_1695, n_1696, n_1697;
  wire n_1698, n_1700, n_1701, n_1702, n_1703, n_1704, n_1706, n_1707;
  wire n_1708, n_1709, n_1710, n_1712, n_1713, n_1714, n_1715, n_1716;
  wire n_1718, n_1719, n_1720, n_1721, n_1722, n_1724, n_1725, n_1726;
  wire n_1727, n_1728, n_1730, n_1731, n_1732, n_1733, n_1734, n_1736;
  wire n_1737, n_1738, n_1739, n_1740, n_1745, n_1747, n_1748, n_1750;
  wire n_1752, n_1754, n_1755, n_1757, n_1758, n_1760, n_1762, n_1764;
  wire n_1765, n_1767, n_1768, n_1770, n_1772, n_1774, n_1775, n_1777;
  wire n_1778, n_1780, n_1782, n_1784, n_1785, n_1787, n_1788, n_1790;
  wire n_1792, n_1794, n_1795, n_1797, n_1798, n_1800, n_1802, n_1804;
  wire n_1805, n_1807, n_1808, n_1810, n_1812, n_1814, n_1815, n_1817;
  wire n_1818, n_1820, n_1822, n_1824, n_1825, n_1827, n_1828, n_1830;
  wire n_1832, n_1834, n_1835, n_1837, n_1838, n_1840, n_1842, n_1844;
  wire n_1845, n_1847, n_1848, n_1850, n_1854, n_1855, n_1856, n_1858;
  wire n_1859, n_1860, n_1862, n_1863, n_1864, n_1865, n_1867, n_1869;
  wire n_1871, n_1872, n_1873, n_1875, n_1876, n_1877, n_1879, n_1880;
  wire n_1882, n_1884, n_1886, n_1887, n_1888, n_1890, n_1891, n_1892;
  wire n_1894, n_1895, n_1897, n_1899, n_1901, n_1902, n_1903, n_1905;
  wire n_1906, n_1907, n_1909, n_1910, n_1912, n_1914, n_1916, n_1917;
  wire n_1918, n_1920, n_1921, n_1922, n_1924, n_1925, n_1927, n_1929;
  wire n_1931, n_1932, n_1933, n_1935, n_1937, n_1938, n_1939, n_1941;
  wire n_1942, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950;
  wire n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958;
  wire n_1960, n_1963, n_1965, n_1966, n_1967, n_1970, n_1973, n_1975;
  wire n_1976, n_1978, n_1980, n_1981, n_1983, n_1985, n_1986, n_1988;
  wire n_1990, n_1991, n_1993, n_1994, n_1996, n_1999, n_2001, n_2002;
  wire n_2003, n_2006, n_2009, n_2011, n_2012, n_2014, n_2016, n_2017;
  wire n_2019, n_2021, n_2022, n_2024, n_2026, n_2027, n_2028, n_2030;
  wire n_2031, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039;
  wire n_2040, n_2041, n_2042, n_2043, n_2044, n_2046, n_2047, n_2048;
  wire n_2050, n_2051, n_2052, n_2054, n_2055, n_2056, n_2058, n_2059;
  wire n_2060, n_2062, n_2063, n_2064, n_2066, n_2067, n_2068, n_2070;
  wire n_2071, n_2072, n_2074, n_2075, n_2076, n_2078, n_2079, n_2080;
  wire n_2082, n_2083, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090;
  wire n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2098, n_2099;
  wire n_2100, n_2102, n_2103, n_2104, n_2106, n_2107, n_2108, n_2110;
  wire n_2111, n_2112, n_2114, n_2115, n_2116, n_2118, n_2119, n_2120;
  wire n_2122, n_2123, n_2125, n_2128, n_2129, n_2131, n_2132, n_2133;
  wire n_2134, n_2136, n_2137, n_2138, n_2140, n_2141, n_2142, n_2143;
  wire n_2145, n_2146, n_2148, n_2149, n_2151, n_2152, n_2153, n_2154;
  wire n_2156, n_2157, n_2158, n_2160, n_2161, n_2162, n_2163, n_2165;
  wire n_2166, n_2168, n_2169, n_2171, n_2172, n_2173, n_2174, n_2176;
  wire n_2177, n_2178, n_2179, n_2181, n_2182, n_2183, n_2184, n_2186;
  wire n_2187, n_2189, n_2190, n_2192, n_2193, n_2194, n_2195, n_2197;
  wire n_2198, n_2199, n_2201, n_2202, n_2203, n_2204, n_2206, n_2207;
  wire n_2209, n_2210, n_2212, n_2213, n_2214, n_2215, n_2217, n_2218;
  wire n_2219, n_2220, n_2222, n_2223, n_2224, n_2225, n_2227, n_2228;
  wire n_2230, n_2231, n_2233, n_2234, n_2235, n_2236, n_2238, n_2239;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_69, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_623, A[1], n_171);
  xor g270 (n_117, n_623, A[2]);
  nand g3 (n_624, A[1], n_171);
  nand g271 (n_625, A[2], n_171);
  nand g272 (n_626, A[1], A[2]);
  nand g273 (n_172, n_624, n_625, n_626);
  xor g274 (n_627, A[2], A[3]);
  xor g275 (n_116, n_627, n_172);
  nand g276 (n_628, A[2], A[3]);
  nand g4 (n_629, n_172, A[3]);
  nand g277 (n_630, A[2], n_172);
  nand g278 (n_174, n_628, n_629, n_630);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_176, A[0], A[3]);
  xor g281 (n_631, A[4], n_173);
  xor g282 (n_115, n_631, n_174);
  nand g283 (n_632, A[4], n_173);
  nand g284 (n_633, n_174, n_173);
  nand g5 (n_634, A[4], n_174);
  nand g6 (n_66, n_632, n_633, n_634);
  xor g287 (n_635, n_69, A[4]);
  xor g288 (n_71, n_635, n_176);
  nand g289 (n_636, n_69, A[4]);
  nand g290 (n_637, n_176, A[4]);
  nand g291 (n_638, n_69, n_176);
  nand g292 (n_180, n_636, n_637, n_638);
  xor g293 (n_639, A[5], n_71);
  xor g294 (n_114, n_639, A[7]);
  nand g295 (n_640, A[5], n_71);
  nand g296 (n_641, A[7], n_71);
  nand g297 (n_642, A[5], A[7]);
  nand g298 (n_181, n_640, n_641, n_642);
  xor g299 (n_643, A[1], A[2]);
  xor g300 (n_179, n_643, n_171);
  xor g305 (n_647, n_179, A[5]);
  xor g306 (n_65, n_647, A[6]);
  nand g307 (n_648, n_179, A[5]);
  nand g308 (n_649, A[6], A[5]);
  nand g309 (n_650, n_179, A[6]);
  nand g310 (n_184, n_648, n_649, n_650);
  xor g311 (n_651, n_180, A[8]);
  xor g312 (n_113, n_651, n_181);
  nand g313 (n_652, n_180, A[8]);
  nand g314 (n_653, n_181, A[8]);
  nand g315 (n_654, n_180, n_181);
  nand g316 (n_64, n_652, n_653, n_654);
  xor g323 (n_659, n_116, A[6]);
  xor g324 (n_185, n_659, A[7]);
  nand g325 (n_660, n_116, A[6]);
  nand g326 (n_661, A[7], A[6]);
  nand g327 (n_662, n_116, A[7]);
  nand g328 (n_189, n_660, n_661, n_662);
  xor g329 (n_663, A[9], n_184);
  xor g330 (n_112, n_663, n_185);
  nand g331 (n_664, A[9], n_184);
  nand g332 (n_665, n_185, n_184);
  nand g333 (n_666, A[9], n_185);
  nand g334 (n_63, n_664, n_665, n_666);
  xor g343 (n_671, A[7], A[8]);
  xor g344 (n_190, n_671, A[10]);
  nand g345 (n_672, A[7], A[8]);
  nand g346 (n_673, A[10], A[8]);
  nand g347 (n_674, A[7], A[10]);
  nand g348 (n_196, n_672, n_673, n_674);
  xor g349 (n_675, n_115, n_189);
  xor g350 (n_111, n_675, n_190);
  nand g351 (n_676, n_115, n_189);
  nand g352 (n_677, n_190, n_189);
  nand g353 (n_678, n_115, n_190);
  nand g354 (n_62, n_676, n_677, n_678);
  xor g364 (n_195, n_639, A[8]);
  nand g366 (n_685, A[8], n_71);
  nand g367 (n_686, A[5], A[8]);
  nand g368 (n_202, n_640, n_685, n_686);
  xor g369 (n_687, n_66, A[9]);
  xor g370 (n_197, n_687, A[11]);
  nand g371 (n_688, n_66, A[9]);
  nand g372 (n_689, A[11], A[9]);
  nand g373 (n_690, n_66, A[11]);
  nand g374 (n_203, n_688, n_689, n_690);
  xor g375 (n_691, n_195, n_196);
  xor g376 (n_110, n_691, n_197);
  nand g377 (n_692, n_195, n_196);
  nand g378 (n_693, n_197, n_196);
  nand g379 (n_694, n_195, n_197);
  nand g380 (n_61, n_692, n_693, n_694);
  xor g387 (n_699, n_117, A[5]);
  xor g388 (n_201, n_699, n_180);
  nand g389 (n_700, n_117, A[5]);
  nand g390 (n_701, n_180, A[5]);
  nand g391 (n_702, n_117, n_180);
  nand g392 (n_208, n_700, n_701, n_702);
  xor g393 (n_703, A[6], A[10]);
  xor g394 (n_204, n_703, A[9]);
  nand g395 (n_704, A[6], A[10]);
  nand g396 (n_705, A[9], A[10]);
  nand g397 (n_706, A[6], A[9]);
  nand g398 (n_210, n_704, n_705, n_706);
  xor g399 (n_707, n_201, A[12]);
  xor g400 (n_205, n_707, n_202);
  nand g401 (n_708, n_201, A[12]);
  nand g402 (n_709, n_202, A[12]);
  nand g403 (n_710, n_201, n_202);
  nand g404 (n_212, n_708, n_709, n_710);
  xor g405 (n_711, n_203, n_204);
  xor g406 (n_109, n_711, n_205);
  nand g407 (n_712, n_203, n_204);
  nand g408 (n_713, n_205, n_204);
  nand g409 (n_714, n_203, n_205);
  nand g410 (n_60, n_712, n_713, n_714);
  xor g423 (n_723, A[11], A[10]);
  xor g424 (n_211, n_723, A[13]);
  nand g425 (n_724, A[11], A[10]);
  nand g426 (n_725, A[13], A[10]);
  nand g427 (n_726, A[11], A[13]);
  nand g428 (n_219, n_724, n_725, n_726);
  xor g429 (n_727, n_208, n_185);
  xor g430 (n_213, n_727, n_210);
  nand g431 (n_728, n_208, n_185);
  nand g432 (n_729, n_210, n_185);
  nand g433 (n_730, n_208, n_210);
  nand g434 (n_67, n_728, n_729, n_730);
  xor g435 (n_731, n_211, n_212);
  xor g436 (n_108, n_731, n_213);
  nand g437 (n_732, n_211, n_212);
  nand g438 (n_733, n_213, n_212);
  nand g439 (n_734, n_211, n_213);
  nand g440 (n_59, n_732, n_733, n_734);
  xor g450 (n_218, n_671, n_115);
  nand g452 (n_741, n_115, A[8]);
  nand g453 (n_742, A[7], n_115);
  nand g454 (n_223, n_672, n_741, n_742);
  xor g455 (n_743, A[11], A[12]);
  xor g456 (n_220, n_743, n_189);
  nand g457 (n_744, A[11], A[12]);
  nand g458 (n_745, n_189, A[12]);
  nand g459 (n_746, A[11], n_189);
  nand g460 (n_224, n_744, n_745, n_746);
  xor g461 (n_747, A[14], n_218);
  xor g462 (n_68, n_747, n_219);
  nand g463 (n_748, A[14], n_218);
  nand g464 (n_749, n_219, n_218);
  nand g465 (n_750, A[14], n_219);
  nand g466 (n_227, n_748, n_749, n_750);
  xor g467 (n_751, n_220, n_67);
  xor g468 (n_107, n_751, n_68);
  nand g469 (n_752, n_220, n_67);
  nand g470 (n_753, n_68, n_67);
  nand g471 (n_754, n_220, n_68);
  nand g472 (n_58, n_752, n_753, n_754);
  xor g488 (n_225, n_687, A[13]);
  nand g490 (n_765, A[13], n_66);
  nand g491 (n_766, A[9], A[13]);
  nand g492 (n_234, n_688, n_765, n_766);
  xor g493 (n_767, A[12], A[15]);
  xor g494 (n_226, n_767, n_195);
  nand g495 (n_768, A[12], A[15]);
  nand g496 (n_769, n_195, A[15]);
  nand g497 (n_770, A[12], n_195);
  nand g498 (n_237, n_768, n_769, n_770);
  xor g499 (n_771, n_223, n_224);
  xor g500 (n_228, n_771, n_225);
  nand g501 (n_772, n_223, n_224);
  nand g502 (n_773, n_225, n_224);
  nand g503 (n_774, n_223, n_225);
  nand g504 (n_239, n_772, n_773, n_774);
  xor g505 (n_775, n_226, n_227);
  xor g506 (n_106, n_775, n_228);
  nand g507 (n_776, n_226, n_227);
  nand g508 (n_777, n_228, n_227);
  nand g509 (n_778, n_226, n_228);
  nand g510 (n_57, n_776, n_777, n_778);
  xor g518 (n_232, n_647, n_180);
  nand g521 (n_786, n_179, n_180);
  nand g522 (n_243, n_648, n_701, n_786);
  xor g523 (n_787, A[6], A[9]);
  xor g524 (n_235, n_787, A[10]);
  xor g529 (n_791, n_232, A[14]);
  xor g530 (n_236, n_791, A[13]);
  nand g531 (n_792, n_232, A[14]);
  nand g532 (n_793, A[13], A[14]);
  nand g533 (n_794, n_232, A[13]);
  nand g534 (n_247, n_792, n_793, n_794);
  xor g535 (n_795, n_202, A[16]);
  xor g536 (n_238, n_795, n_234);
  nand g537 (n_796, n_202, A[16]);
  nand g538 (n_797, n_234, A[16]);
  nand g539 (n_798, n_202, n_234);
  nand g540 (n_249, n_796, n_797, n_798);
  xor g541 (n_799, n_235, n_236);
  xor g542 (n_240, n_799, n_237);
  nand g543 (n_800, n_235, n_236);
  nand g544 (n_801, n_237, n_236);
  nand g545 (n_802, n_235, n_237);
  nand g546 (n_250, n_800, n_801, n_802);
  xor g547 (n_803, n_238, n_239);
  xor g548 (n_105, n_803, n_240);
  nand g549 (n_804, n_238, n_239);
  nand g550 (n_805, n_240, n_239);
  nand g551 (n_806, n_238, n_240);
  nand g552 (n_56, n_804, n_805, n_806);
  xor g559 (n_811, n_116, A[7]);
  xor g560 (n_244, n_811, A[6]);
  xor g566 (n_246, n_723, A[14]);
  nand g568 (n_817, A[14], A[11]);
  nand g569 (n_818, A[10], A[14]);
  nand g570 (n_258, n_724, n_817, n_818);
  xor g571 (n_819, n_243, n_244);
  xor g572 (n_248, n_819, A[15]);
  nand g573 (n_820, n_243, n_244);
  nand g574 (n_821, A[15], n_244);
  nand g575 (n_822, n_243, A[15]);
  nand g576 (n_259, n_820, n_821, n_822);
  xor g577 (n_823, n_210, A[17]);
  xor g578 (n_251, n_823, n_246);
  nand g579 (n_824, n_210, A[17]);
  nand g580 (n_825, n_246, A[17]);
  nand g581 (n_826, n_210, n_246);
  nand g582 (n_262, n_824, n_825, n_826);
  xor g583 (n_827, n_247, n_248);
  xor g584 (n_252, n_827, n_249);
  nand g585 (n_828, n_247, n_248);
  nand g586 (n_829, n_249, n_248);
  nand g587 (n_830, n_247, n_249);
  nand g588 (n_119, n_828, n_829, n_830);
  xor g589 (n_831, n_250, n_251);
  xor g590 (n_104, n_831, n_252);
  nand g591 (n_832, n_250, n_251);
  nand g592 (n_833, n_252, n_251);
  nand g593 (n_834, n_250, n_252);
  nand g594 (n_55, n_832, n_833, n_834);
  xor g615 (n_847, A[15], n_218);
  xor g616 (n_261, n_847, A[16]);
  nand g617 (n_848, A[15], n_218);
  nand g618 (n_849, A[16], n_218);
  nand g619 (n_850, A[15], A[16]);
  nand g620 (n_272, n_848, n_849, n_850);
  xor g621 (n_851, A[18], n_258);
  xor g622 (n_118, n_851, n_259);
  nand g623 (n_852, A[18], n_258);
  nand g624 (n_853, n_259, n_258);
  nand g625 (n_854, A[18], n_259);
  nand g626 (n_274, n_852, n_853, n_854);
  xor g627 (n_855, n_220, n_261);
  xor g628 (n_263, n_855, n_262);
  nand g629 (n_856, n_220, n_261);
  nand g630 (n_857, n_262, n_261);
  nand g631 (n_858, n_220, n_262);
  nand g632 (n_277, n_856, n_857, n_858);
  xor g633 (n_859, n_118, n_119);
  xor g634 (n_103, n_859, n_263);
  nand g635 (n_860, n_118, n_119);
  nand g636 (n_861, n_263, n_119);
  nand g637 (n_862, n_118, n_263);
  nand g638 (n_54, n_860, n_861, n_862);
  xor g654 (n_271, n_687, A[12]);
  nand g656 (n_873, A[12], n_66);
  nand g657 (n_874, A[9], A[12]);
  nand g658 (n_285, n_688, n_873, n_874);
  xor g659 (n_875, A[13], n_195);
  xor g660 (n_273, n_875, A[16]);
  nand g661 (n_876, A[13], n_195);
  nand g662 (n_877, A[16], n_195);
  nand g663 (n_878, A[13], A[16]);
  nand g664 (n_287, n_876, n_877, n_878);
  xor g666 (n_275, n_771, A[17]);
  nand g668 (n_881, A[17], n_224);
  nand g669 (n_882, n_223, A[17]);
  nand g670 (n_288, n_772, n_881, n_882);
  xor g671 (n_883, n_271, A[19]);
  xor g672 (n_276, n_883, n_272);
  nand g673 (n_884, n_271, A[19]);
  nand g674 (n_885, n_272, A[19]);
  nand g675 (n_886, n_271, n_272);
  nand g676 (n_291, n_884, n_885, n_886);
  xor g677 (n_887, n_273, n_274);
  xor g678 (n_278, n_887, n_275);
  nand g679 (n_888, n_273, n_274);
  nand g680 (n_889, n_275, n_274);
  nand g681 (n_890, n_273, n_275);
  nand g682 (n_293, n_888, n_889, n_890);
  xor g683 (n_891, n_276, n_277);
  xor g684 (n_102, n_891, n_278);
  nand g685 (n_892, n_276, n_277);
  nand g686 (n_893, n_278, n_277);
  nand g687 (n_894, n_276, n_278);
  nand g688 (n_53, n_892, n_893, n_894);
  xor g701 (n_903, n_180, A[10]);
  xor g702 (n_284, n_903, A[9]);
  nand g703 (n_904, n_180, A[10]);
  nand g705 (n_906, n_180, A[9]);
  nand g706 (n_299, n_904, n_705, n_906);
  xor g707 (n_907, A[13], n_65);
  xor g708 (n_286, n_907, A[14]);
  nand g709 (n_908, A[13], n_65);
  nand g710 (n_909, A[14], n_65);
  nand g712 (n_301, n_908, n_909, n_793);
  xor g713 (n_911, n_202, n_284);
  xor g714 (n_290, n_911, n_285);
  nand g715 (n_912, n_202, n_284);
  nand g716 (n_913, n_285, n_284);
  nand g717 (n_914, n_202, n_285);
  nand g718 (n_304, n_912, n_913, n_914);
  xor g719 (n_915, A[18], A[20]);
  xor g720 (n_289, n_915, A[17]);
  nand g721 (n_916, A[18], A[20]);
  nand g722 (n_917, A[17], A[20]);
  nand g723 (n_918, A[18], A[17]);
  nand g724 (n_303, n_916, n_917, n_918);
  xor g725 (n_919, n_286, n_287);
  xor g726 (n_292, n_919, n_288);
  nand g727 (n_920, n_286, n_287);
  nand g728 (n_921, n_288, n_287);
  nand g729 (n_922, n_286, n_288);
  nand g730 (n_307, n_920, n_921, n_922);
  xor g731 (n_923, n_289, n_290);
  xor g732 (n_294, n_923, n_291);
  nand g733 (n_924, n_289, n_290);
  nand g734 (n_925, n_291, n_290);
  nand g735 (n_926, n_289, n_291);
  nand g736 (n_309, n_924, n_925, n_926);
  xor g737 (n_927, n_292, n_293);
  xor g738 (n_101, n_927, n_294);
  nand g739 (n_928, n_292, n_293);
  nand g740 (n_929, n_294, n_293);
  nand g741 (n_930, n_292, n_294);
  nand g742 (n_52, n_928, n_929, n_930);
  xor g756 (n_300, n_723, n_184);
  nand g758 (n_941, n_184, A[10]);
  nand g759 (n_942, A[11], n_184);
  nand g760 (n_316, n_724, n_941, n_942);
  xor g761 (n_943, A[14], A[15]);
  xor g762 (n_302, n_943, n_244);
  nand g763 (n_944, A[14], A[15]);
  nand g765 (n_946, A[14], n_244);
  nand g766 (n_318, n_944, n_821, n_946);
  xor g767 (n_947, n_299, n_300);
  xor g768 (n_306, n_947, A[19]);
  nand g769 (n_948, n_299, n_300);
  nand g770 (n_949, A[19], n_300);
  nand g771 (n_950, n_299, A[19]);
  nand g772 (n_319, n_948, n_949, n_950);
  xor g773 (n_951, A[18], n_301);
  xor g774 (n_305, n_951, A[21]);
  nand g775 (n_952, A[18], n_301);
  nand g776 (n_953, A[21], n_301);
  nand g777 (n_954, A[18], A[21]);
  nand g778 (n_322, n_952, n_953, n_954);
  xor g779 (n_955, n_302, n_303);
  xor g780 (n_308, n_955, n_304);
  nand g781 (n_956, n_302, n_303);
  nand g782 (n_957, n_304, n_303);
  nand g783 (n_958, n_302, n_304);
  nand g784 (n_324, n_956, n_957, n_958);
  xor g785 (n_959, n_305, n_306);
  xor g786 (n_310, n_959, n_307);
  nand g787 (n_960, n_305, n_306);
  nand g788 (n_961, n_307, n_306);
  nand g789 (n_962, n_305, n_307);
  nand g790 (n_327, n_960, n_961, n_962);
  xor g791 (n_963, n_308, n_309);
  xor g792 (n_100, n_963, n_310);
  nand g793 (n_964, n_308, n_309);
  nand g794 (n_965, n_310, n_309);
  nand g795 (n_966, n_308, n_310);
  nand g796 (n_51, n_964, n_965, n_966);
  xor g806 (n_315, n_671, A[11]);
  nand g808 (n_973, A[11], A[8]);
  nand g809 (n_974, A[7], A[11]);
  nand g810 (n_333, n_672, n_973, n_974);
  xor g811 (n_975, n_115, A[12]);
  xor g812 (n_317, n_975, n_189);
  nand g813 (n_976, n_115, A[12]);
  nand g816 (n_335, n_976, n_745, n_676);
  xor g817 (n_979, A[15], A[16]);
  xor g818 (n_320, n_979, n_315);
  nand g820 (n_981, n_315, A[16]);
  nand g821 (n_982, A[15], n_315);
  nand g822 (n_337, n_850, n_981, n_982);
  xor g823 (n_983, A[20], A[19]);
  xor g824 (n_321, n_983, n_316);
  nand g825 (n_984, A[20], A[19]);
  nand g826 (n_985, n_316, A[19]);
  nand g827 (n_986, A[20], n_316);
  nand g828 (n_338, n_984, n_985, n_986);
  xor g829 (n_987, n_317, n_318);
  xor g830 (n_323, n_987, A[22]);
  nand g831 (n_988, n_317, n_318);
  nand g832 (n_989, A[22], n_318);
  nand g833 (n_990, n_317, A[22]);
  nand g834 (n_340, n_988, n_989, n_990);
  xor g835 (n_991, n_319, n_320);
  xor g836 (n_325, n_991, n_321);
  nand g837 (n_992, n_319, n_320);
  nand g838 (n_993, n_321, n_320);
  nand g839 (n_994, n_319, n_321);
  nand g840 (n_343, n_992, n_993, n_994);
  xor g841 (n_995, n_322, n_323);
  xor g842 (n_326, n_995, n_324);
  nand g843 (n_996, n_322, n_323);
  nand g844 (n_997, n_324, n_323);
  nand g845 (n_998, n_322, n_324);
  nand g846 (n_345, n_996, n_997, n_998);
  xor g847 (n_999, n_325, n_326);
  xor g848 (n_99, n_999, n_327);
  nand g849 (n_1000, n_325, n_326);
  nand g850 (n_1001, n_327, n_326);
  nand g851 (n_1002, n_325, n_327);
  nand g852 (n_50, n_1000, n_1001, n_1002);
  xor g873 (n_1015, A[12], n_195);
  xor g874 (n_336, n_1015, n_333);
  nand g876 (n_1017, n_333, n_195);
  nand g877 (n_1018, A[12], n_333);
  nand g878 (n_357, n_770, n_1017, n_1018);
  xor g879 (n_1019, A[16], n_225);
  xor g880 (n_341, n_1019, n_335);
  nand g881 (n_1020, A[16], n_225);
  nand g882 (n_1021, n_335, n_225);
  nand g883 (n_1022, A[16], n_335);
  nand g884 (n_358, n_1020, n_1021, n_1022);
  xor g885 (n_1023, A[17], A[20]);
  xor g886 (n_339, n_1023, A[23]);
  nand g888 (n_1025, A[23], A[20]);
  nand g889 (n_1026, A[17], A[23]);
  nand g890 (n_360, n_917, n_1025, n_1026);
  xor g891 (n_1027, A[21], n_336);
  xor g892 (n_342, n_1027, n_337);
  nand g893 (n_1028, A[21], n_336);
  nand g894 (n_1029, n_337, n_336);
  nand g895 (n_1030, A[21], n_337);
  nand g896 (n_362, n_1028, n_1029, n_1030);
  xor g897 (n_1031, n_338, n_339);
  xor g898 (n_344, n_1031, n_340);
  nand g899 (n_1032, n_338, n_339);
  nand g900 (n_1033, n_340, n_339);
  nand g901 (n_1034, n_338, n_340);
  nand g902 (n_365, n_1032, n_1033, n_1034);
  xor g903 (n_1035, n_341, n_342);
  xor g904 (n_346, n_1035, n_343);
  nand g905 (n_1036, n_341, n_342);
  nand g906 (n_1037, n_343, n_342);
  nand g907 (n_1038, n_341, n_343);
  nand g908 (n_367, n_1036, n_1037, n_1038);
  xor g909 (n_1039, n_344, n_345);
  xor g910 (n_98, n_1039, n_346);
  nand g911 (n_1040, n_344, n_345);
  nand g912 (n_1041, n_346, n_345);
  nand g913 (n_1042, n_344, n_346);
  nand g914 (n_49, n_1040, n_1041, n_1042);
  xor g917 (n_1043, A[2], n_171);
  nand g922 (n_372, n_625, n_1045, n_1046);
  xor g923 (n_1047, n_350, A[5]);
  xor g924 (n_352, n_1047, n_180);
  nand g925 (n_1048, n_350, A[5]);
  nand g927 (n_1050, n_350, n_180);
  nand g928 (n_374, n_1048, n_701, n_1050);
  xor g935 (n_1055, A[14], n_352);
  xor g936 (n_356, n_1055, A[13]);
  nand g937 (n_1056, A[14], n_352);
  nand g938 (n_1057, A[13], n_352);
  nand g940 (n_378, n_1056, n_1057, n_793);
  xor g941 (n_1059, n_202, n_235);
  xor g942 (n_359, n_1059, A[18]);
  nand g943 (n_1060, n_202, n_235);
  nand g944 (n_1061, A[18], n_235);
  nand g945 (n_1062, n_202, A[18]);
  nand g946 (n_381, n_1060, n_1061, n_1062);
  xor g947 (n_1063, n_234, A[17]);
  nand g949 (n_1064, n_234, A[17]);
  nand g952 (n_382, n_1064, n_1065, n_1066);
  xor g953 (n_1067, n_356, A[22]);
  xor g954 (n_363, n_1067, A[21]);
  nand g955 (n_1068, n_356, A[22]);
  nand g956 (n_1069, A[21], A[22]);
  nand g957 (n_1070, n_356, A[21]);
  nand g958 (n_384, n_1068, n_1069, n_1070);
  xor g959 (n_1071, n_357, n_358);
  xor g960 (n_364, n_1071, n_359);
  nand g961 (n_1072, n_357, n_358);
  nand g962 (n_1073, n_359, n_358);
  nand g963 (n_1074, n_357, n_359);
  nand g964 (n_386, n_1072, n_1073, n_1074);
  xor g965 (n_1075, n_360, n_361);
  xor g966 (n_366, n_1075, n_362);
  nand g967 (n_1076, n_360, n_361);
  nand g968 (n_1077, n_362, n_361);
  nand g969 (n_1078, n_360, n_362);
  nand g970 (n_388, n_1076, n_1077, n_1078);
  xor g971 (n_1079, n_363, n_364);
  xor g972 (n_368, n_1079, n_365);
  nand g973 (n_1080, n_363, n_364);
  nand g974 (n_1081, n_365, n_364);
  nand g975 (n_1082, n_363, n_365);
  nand g976 (n_390, n_1080, n_1081, n_1082);
  xor g977 (n_1083, n_366, n_367);
  xor g978 (n_97, n_1083, n_368);
  nand g979 (n_1084, n_366, n_367);
  nand g980 (n_1085, n_368, n_367);
  nand g981 (n_1086, n_366, n_368);
  nand g982 (n_48, n_1084, n_1085, n_1086);
  xor g985 (n_1087, A[1], A[3]);
  nand g987 (n_1088, A[1], A[3]);
  nand g990 (n_393, n_1088, n_1089, n_1090);
  xor g991 (n_1091, n_372, n_373);
  xor g992 (n_375, n_1091, A[7]);
  nand g993 (n_1092, n_372, n_373);
  nand g994 (n_1093, A[7], n_373);
  nand g995 (n_1094, n_372, A[7]);
  nand g996 (n_396, n_1092, n_1093, n_1094);
  xor g998 (n_377, n_703, A[11]);
  nand g1001 (n_1098, A[6], A[11]);
  nand g1002 (n_397, n_704, n_724, n_1098);
  xor g1003 (n_1099, n_374, n_375);
  xor g1004 (n_379, n_1099, A[14]);
  nand g1005 (n_1100, n_374, n_375);
  nand g1006 (n_1101, A[14], n_375);
  nand g1007 (n_1102, n_374, A[14]);
  nand g1008 (n_398, n_1100, n_1101, n_1102);
  xor g1009 (n_1103, A[15], n_210);
  xor g1010 (n_380, n_1103, n_377);
  nand g1011 (n_1104, A[15], n_210);
  nand g1012 (n_1105, n_377, n_210);
  nand g1013 (n_1106, A[15], n_377);
  nand g1014 (n_401, n_1104, n_1105, n_1106);
  xor g1015 (n_1107, A[19], n_378);
  xor g1016 (n_383, n_1107, A[18]);
  nand g1017 (n_1108, A[19], n_378);
  nand g1018 (n_1109, A[18], n_378);
  nand g1019 (n_1110, A[19], A[18]);
  nand g1020 (n_402, n_1108, n_1109, n_1110);
  xor g1021 (n_1111, A[22], n_379);
  xor g1022 (n_385, n_1111, A[23]);
  nand g1023 (n_1112, A[22], n_379);
  nand g1024 (n_1113, A[23], n_379);
  nand g1025 (n_1114, A[22], A[23]);
  nand g1026 (n_404, n_1112, n_1113, n_1114);
  xor g1027 (n_1115, n_380, n_381);
  xor g1028 (n_387, n_1115, n_382);
  nand g1029 (n_1116, n_380, n_381);
  nand g1030 (n_1117, n_382, n_381);
  nand g1031 (n_1118, n_380, n_382);
  nand g1032 (n_407, n_1116, n_1117, n_1118);
  xor g1033 (n_1119, n_383, n_384);
  xor g1034 (n_389, n_1119, n_385);
  nand g1035 (n_1120, n_383, n_384);
  nand g1036 (n_1121, n_385, n_384);
  nand g1037 (n_1122, n_383, n_385);
  nand g1038 (n_409, n_1120, n_1121, n_1122);
  xor g1039 (n_1123, n_386, n_387);
  xor g1040 (n_391, n_1123, n_388);
  nand g1041 (n_1124, n_386, n_387);
  nand g1042 (n_1125, n_388, n_387);
  nand g1043 (n_1126, n_386, n_388);
  nand g1044 (n_412, n_1124, n_1125, n_1126);
  xor g1045 (n_1127, n_389, n_390);
  xor g1046 (n_96, n_1127, n_391);
  nand g1047 (n_1128, n_389, n_390);
  nand g1048 (n_1129, n_391, n_390);
  nand g1049 (n_1130, n_389, n_391);
  nand g1050 (n_47, n_1128, n_1129, n_1130);
  xor g1052 (n_394, n_627, A[4]);
  nand g1054 (n_1133, A[4], A[2]);
  nand g1055 (n_1134, A[3], A[4]);
  nand g1056 (n_413, n_628, n_1133, n_1134);
  xor g1057 (n_1135, n_393, n_394);
  xor g1058 (n_395, n_1135, A[7]);
  nand g1059 (n_1136, n_393, n_394);
  nand g1060 (n_1137, A[7], n_394);
  nand g1061 (n_1138, n_393, A[7]);
  nand g1062 (n_415, n_1136, n_1137, n_1138);
  xor g1063 (n_1139, A[8], A[11]);
  xor g1064 (n_399, n_1139, A[12]);
  nand g1067 (n_1142, A[8], A[12]);
  nand g1068 (n_417, n_973, n_744, n_1142);
  xor g1069 (n_1143, n_395, n_396);
  xor g1070 (n_400, n_1143, A[15]);
  nand g1071 (n_1144, n_395, n_396);
  nand g1072 (n_1145, A[15], n_396);
  nand g1073 (n_1146, n_395, A[15]);
  nand g1074 (n_419, n_1144, n_1145, n_1146);
  xor g1075 (n_1147, n_397, A[16]);
  xor g1076 (n_403, n_1147, n_398);
  nand g1077 (n_1148, n_397, A[16]);
  nand g1078 (n_1149, n_398, A[16]);
  nand g1079 (n_1150, n_397, n_398);
  nand g1080 (n_420, n_1148, n_1149, n_1150);
  xor g1082 (n_405, n_1151, n_399);
  nand g1084 (n_1153, n_399, A[19]);
  nand g1086 (n_421, n_1152, n_1153, n_1154);
  xor g1087 (n_1155, A[20], A[23]);
  xor g1088 (n_406, n_1155, n_400);
  nand g1090 (n_1157, n_400, A[23]);
  nand g1091 (n_1158, A[20], n_400);
  nand g1092 (n_422, n_1025, n_1157, n_1158);
  xor g1093 (n_1159, n_401, n_402);
  xor g1094 (n_408, n_1159, n_403);
  nand g1095 (n_1160, n_401, n_402);
  nand g1096 (n_1161, n_403, n_402);
  nand g1097 (n_1162, n_401, n_403);
  nand g1098 (n_426, n_1160, n_1161, n_1162);
  xor g1099 (n_1163, n_404, n_405);
  xor g1100 (n_410, n_1163, n_406);
  nand g1101 (n_1164, n_404, n_405);
  nand g1102 (n_1165, n_406, n_405);
  nand g1103 (n_1166, n_404, n_406);
  nand g1104 (n_429, n_1164, n_1165, n_1166);
  xor g1105 (n_1167, n_407, n_408);
  xor g1106 (n_411, n_1167, n_409);
  nand g1107 (n_1168, n_407, n_408);
  nand g1108 (n_1169, n_409, n_408);
  nand g1109 (n_1170, n_407, n_409);
  nand g1110 (n_431, n_1168, n_1169, n_1170);
  xor g1111 (n_1171, n_410, n_411);
  xor g1112 (n_95, n_1171, n_412);
  nand g1113 (n_1172, n_410, n_411);
  nand g1114 (n_1173, n_412, n_411);
  nand g1115 (n_1174, n_410, n_412);
  nand g1116 (n_46, n_1172, n_1173, n_1174);
  xor g1117 (n_1175, A[4], A[5]);
  xor g1118 (n_414, n_1175, n_413);
  nand g1119 (n_1176, A[4], A[5]);
  nand g1120 (n_1177, n_413, A[5]);
  nand g1121 (n_1178, A[4], n_413);
  nand g1122 (n_434, n_1176, n_1177, n_1178);
  xor g1123 (n_1179, A[8], A[9]);
  xor g1124 (n_416, n_1179, n_414);
  nand g1125 (n_1180, A[8], A[9]);
  nand g1126 (n_1181, n_414, A[9]);
  nand g1127 (n_1182, A[8], n_414);
  nand g1128 (n_436, n_1180, n_1181, n_1182);
  xor g1129 (n_1183, A[13], A[12]);
  xor g1130 (n_418, n_1183, n_415);
  nand g1131 (n_1184, A[13], A[12]);
  nand g1132 (n_1185, n_415, A[12]);
  nand g1133 (n_1186, A[13], n_415);
  nand g1134 (n_438, n_1184, n_1185, n_1186);
  xor g1136 (n_424, n_1187, n_416);
  nand g1139 (n_1190, A[16], n_416);
  nand g1140 (n_441, n_1188, n_1189, n_1190);
  xor g1142 (n_423, n_1023, n_417);
  nand g1144 (n_1193, n_417, A[20]);
  nand g1145 (n_1194, A[17], n_417);
  nand g1146 (n_439, n_917, n_1193, n_1194);
  xor g1147 (n_1195, n_418, A[21]);
  xor g1148 (n_425, n_1195, n_419);
  nand g1149 (n_1196, n_418, A[21]);
  nand g1150 (n_1197, n_419, A[21]);
  nand g1151 (n_1198, n_418, n_419);
  nand g1152 (n_442, n_1196, n_1197, n_1198);
  xor g1153 (n_1199, n_420, n_421);
  xor g1154 (n_427, n_1199, n_422);
  nand g1155 (n_1200, n_420, n_421);
  nand g1156 (n_1201, n_422, n_421);
  nand g1157 (n_1202, n_420, n_422);
  nand g1158 (n_445, n_1200, n_1201, n_1202);
  xor g1159 (n_1203, n_423, n_424);
  xor g1160 (n_428, n_1203, n_425);
  nand g1161 (n_1204, n_423, n_424);
  nand g1162 (n_1205, n_425, n_424);
  nand g1163 (n_1206, n_423, n_425);
  nand g1164 (n_447, n_1204, n_1205, n_1206);
  xor g1165 (n_1207, n_426, n_427);
  xor g1166 (n_430, n_1207, n_428);
  nand g1167 (n_1208, n_426, n_427);
  nand g1168 (n_1209, n_428, n_427);
  nand g1169 (n_1210, n_426, n_428);
  nand g1170 (n_450, n_1208, n_1209, n_1210);
  xor g1171 (n_1211, n_429, n_430);
  xor g1172 (n_94, n_1211, n_431);
  nand g1173 (n_1212, n_429, n_430);
  nand g1174 (n_1213, n_431, n_430);
  nand g1175 (n_1214, n_429, n_431);
  nand g1176 (n_45, n_1212, n_1213, n_1214);
  xor g1180 (n_435, n_1215, A[9]);
  nand g1184 (n_455, n_1216, n_1217, n_706);
  xor g1185 (n_1219, A[10], n_434);
  xor g1186 (n_437, n_1219, A[14]);
  nand g1187 (n_1220, A[10], n_434);
  nand g1188 (n_1221, A[14], n_434);
  nand g1190 (n_457, n_1220, n_1221, n_818);
  xor g1191 (n_1223, A[13], n_435);
  xor g1192 (n_440, n_1223, n_436);
  nand g1193 (n_1224, A[13], n_435);
  nand g1194 (n_1225, n_436, n_435);
  nand g1195 (n_1226, A[13], n_436);
  nand g1196 (n_458, n_1224, n_1225, n_1226);
  xor g1197 (n_1227, A[18], n_437);
  xor g1198 (n_443, n_1227, A[17]);
  nand g1199 (n_1228, A[18], n_437);
  nand g1200 (n_1229, A[17], n_437);
  nand g1202 (n_460, n_1228, n_1229, n_918);
  xor g1203 (n_1231, n_438, A[21]);
  xor g1204 (n_444, n_1231, A[22]);
  nand g1205 (n_1232, n_438, A[21]);
  nand g1207 (n_1234, n_438, A[22]);
  nand g1208 (n_462, n_1232, n_1069, n_1234);
  xor g1209 (n_1235, n_439, n_440);
  xor g1210 (n_446, n_1235, n_441);
  nand g1211 (n_1236, n_439, n_440);
  nand g1212 (n_1237, n_441, n_440);
  nand g1213 (n_1238, n_439, n_441);
  nand g1214 (n_464, n_1236, n_1237, n_1238);
  xor g1215 (n_1239, n_442, n_443);
  xor g1216 (n_448, n_1239, n_444);
  nand g1217 (n_1240, n_442, n_443);
  nand g1218 (n_1241, n_444, n_443);
  nand g1219 (n_1242, n_442, n_444);
  nand g1220 (n_466, n_1240, n_1241, n_1242);
  xor g1221 (n_1243, n_445, n_446);
  xor g1222 (n_449, n_1243, n_447);
  nand g1223 (n_1244, n_445, n_446);
  nand g1224 (n_1245, n_447, n_446);
  nand g1225 (n_1246, n_445, n_447);
  nand g1226 (n_469, n_1244, n_1245, n_1246);
  xor g1227 (n_1247, n_448, n_449);
  xor g1228 (n_93, n_1247, n_450);
  nand g1229 (n_1248, n_448, n_449);
  nand g1230 (n_1249, n_450, n_449);
  nand g1231 (n_1250, n_448, n_450);
  nand g1232 (n_44, n_1248, n_1249, n_1250);
  nand g1238 (n_1253, A[10], A[5]);
  nand g1240 (n_472, n_649, n_1253, n_704);
  xor g1242 (n_456, n_1255, A[14]);
  nand g1246 (n_473, n_1256, n_1257, n_817);
  xor g1247 (n_1259, A[15], n_454);
  xor g1248 (n_459, n_1259, n_455);
  nand g1249 (n_1260, A[15], n_454);
  nand g1250 (n_1261, n_455, n_454);
  nand g1251 (n_1262, A[15], n_455);
  nand g1252 (n_475, n_1260, n_1261, n_1262);
  xor g1253 (n_1263, A[19], n_456);
  xor g1254 (n_461, n_1263, A[18]);
  nand g1255 (n_1264, A[19], n_456);
  nand g1256 (n_1265, A[18], n_456);
  nand g1258 (n_477, n_1264, n_1265, n_1110);
  xor g1259 (n_1267, n_457, A[22]);
  xor g1260 (n_463, n_1267, A[23]);
  nand g1261 (n_1268, n_457, A[22]);
  nand g1263 (n_1270, n_457, A[23]);
  nand g1264 (n_479, n_1268, n_1114, n_1270);
  xor g1265 (n_1271, n_458, n_459);
  xor g1266 (n_465, n_1271, n_460);
  nand g1267 (n_1272, n_458, n_459);
  nand g1268 (n_1273, n_460, n_459);
  nand g1269 (n_1274, n_458, n_460);
  nand g1270 (n_481, n_1272, n_1273, n_1274);
  xor g1271 (n_1275, n_461, n_462);
  xor g1272 (n_467, n_1275, n_463);
  nand g1273 (n_1276, n_461, n_462);
  nand g1274 (n_1277, n_463, n_462);
  nand g1275 (n_1278, n_461, n_463);
  nand g1276 (n_483, n_1276, n_1277, n_1278);
  xor g1277 (n_1279, n_464, n_465);
  xor g1278 (n_468, n_1279, n_466);
  nand g1279 (n_1280, n_464, n_465);
  nand g1280 (n_1281, n_466, n_465);
  nand g1281 (n_1282, n_464, n_466);
  nand g1282 (n_486, n_1280, n_1281, n_1282);
  xor g1283 (n_1283, n_467, n_468);
  xor g1284 (n_92, n_1283, n_469);
  nand g1285 (n_1284, n_467, n_468);
  nand g1286 (n_1285, n_469, n_468);
  nand g1287 (n_1286, n_467, n_469);
  nand g1288 (n_43, n_1284, n_1285, n_1286);
  xor g1295 (n_1291, A[7], A[12]);
  xor g1296 (n_474, n_1291, A[15]);
  nand g1297 (n_1292, A[7], A[12]);
  nand g1299 (n_1294, A[7], A[15]);
  nand g1300 (n_489, n_1292, n_768, n_1294);
  xor g1301 (n_1295, n_315, n_472);
  xor g1302 (n_476, n_1295, A[16]);
  nand g1303 (n_1296, n_315, n_472);
  nand g1304 (n_1297, A[16], n_472);
  nand g1306 (n_490, n_1296, n_1297, n_981);
  xor g1308 (n_478, n_1151, A[20]);
  nand g1312 (n_491, n_1152, n_984, n_1302);
  xor g1313 (n_1303, n_473, A[23]);
  xor g1314 (n_480, n_1303, n_474);
  nand g1315 (n_1304, n_473, A[23]);
  nand g1316 (n_1305, n_474, A[23]);
  nand g1317 (n_1306, n_473, n_474);
  nand g1318 (n_493, n_1304, n_1305, n_1306);
  xor g1319 (n_1307, n_475, n_476);
  xor g1320 (n_482, n_1307, n_477);
  nand g1321 (n_1308, n_475, n_476);
  nand g1322 (n_1309, n_477, n_476);
  nand g1323 (n_1310, n_475, n_477);
  nand g1324 (n_496, n_1308, n_1309, n_1310);
  xor g1325 (n_1311, n_478, n_479);
  xor g1326 (n_484, n_1311, n_480);
  nand g1327 (n_1312, n_478, n_479);
  nand g1328 (n_1313, n_480, n_479);
  nand g1329 (n_1314, n_478, n_480);
  nand g1330 (n_498, n_1312, n_1313, n_1314);
  xor g1331 (n_1315, n_481, n_482);
  xor g1332 (n_485, n_1315, n_483);
  nand g1333 (n_1316, n_481, n_482);
  nand g1334 (n_1317, n_483, n_482);
  nand g1335 (n_1318, n_481, n_483);
  nand g1336 (n_501, n_1316, n_1317, n_1318);
  xor g1337 (n_1319, n_484, n_485);
  xor g1338 (n_91, n_1319, n_486);
  nand g1339 (n_1320, n_484, n_485);
  nand g1340 (n_1321, n_486, n_485);
  nand g1341 (n_1322, n_484, n_486);
  nand g1342 (n_42, n_1320, n_1321, n_1322);
  xor g1344 (n_488, n_1179, A[13]);
  nand g1347 (n_1326, A[8], A[13]);
  nand g1348 (n_504, n_1180, n_766, n_1326);
  xor g1349 (n_1327, A[12], n_333);
  xor g1350 (n_492, n_1327, A[16]);
  nand g1352 (n_1329, A[16], n_333);
  nand g1353 (n_1330, A[12], A[16]);
  nand g1354 (n_506, n_1018, n_1329, n_1330);
  xor g1356 (n_494, n_1331, A[17]);
  nand g1358 (n_1333, A[17], n_488);
  nand g1360 (n_507, n_1332, n_1333, n_1065);
  xor g1361 (n_1335, A[20], A[21]);
  xor g1362 (n_495, n_1335, n_489);
  nand g1363 (n_1336, A[20], A[21]);
  nand g1364 (n_1337, n_489, A[21]);
  nand g1365 (n_1338, A[20], n_489);
  nand g1366 (n_509, n_1336, n_1337, n_1338);
  xor g1367 (n_1339, n_490, n_491);
  xor g1368 (n_497, n_1339, n_492);
  nand g1369 (n_1340, n_490, n_491);
  nand g1370 (n_1341, n_492, n_491);
  nand g1371 (n_1342, n_490, n_492);
  nand g1372 (n_512, n_1340, n_1341, n_1342);
  xor g1373 (n_1343, n_493, n_494);
  xor g1374 (n_499, n_1343, n_495);
  nand g1375 (n_1344, n_493, n_494);
  nand g1376 (n_1345, n_495, n_494);
  nand g1377 (n_1346, n_493, n_495);
  nand g1378 (n_513, n_1344, n_1345, n_1346);
  xor g1379 (n_1347, n_496, n_497);
  xor g1380 (n_500, n_1347, n_498);
  nand g1381 (n_1348, n_496, n_497);
  nand g1382 (n_1349, n_498, n_497);
  nand g1383 (n_1350, n_496, n_498);
  nand g1384 (n_516, n_1348, n_1349, n_1350);
  xor g1385 (n_1351, n_499, n_500);
  xor g1386 (n_90, n_1351, n_501);
  nand g1387 (n_1352, n_499, n_500);
  nand g1388 (n_1353, n_501, n_500);
  nand g1389 (n_1354, n_499, n_501);
  nand g1390 (n_41, n_1352, n_1353, n_1354);
  xor g1393 (n_1355, A[9], A[14]);
  xor g1394 (n_505, n_1355, A[13]);
  nand g1395 (n_1356, A[9], A[14]);
  nand g1398 (n_520, n_1356, n_793, n_766);
  xor g1400 (n_508, n_1359, A[17]);
  nand g1404 (n_523, n_1360, n_918, n_1362);
  xor g1405 (n_1363, n_504, A[21]);
  xor g1406 (n_510, n_1363, A[22]);
  nand g1407 (n_1364, n_504, A[21]);
  nand g1409 (n_1366, n_504, A[22]);
  nand g1410 (n_525, n_1364, n_1069, n_1366);
  xor g1411 (n_1367, n_505, n_506);
  xor g1412 (n_511, n_1367, n_507);
  nand g1413 (n_1368, n_505, n_506);
  nand g1414 (n_1369, n_507, n_506);
  nand g1415 (n_1370, n_505, n_507);
  nand g1416 (n_526, n_1368, n_1369, n_1370);
  xor g1417 (n_1371, n_508, n_509);
  xor g1418 (n_514, n_1371, n_510);
  nand g1419 (n_1372, n_508, n_509);
  nand g1420 (n_1373, n_510, n_509);
  nand g1421 (n_1374, n_508, n_510);
  nand g1422 (n_529, n_1372, n_1373, n_1374);
  xor g1423 (n_1375, n_511, n_512);
  xor g1424 (n_515, n_1375, n_513);
  nand g1425 (n_1376, n_511, n_512);
  nand g1426 (n_1377, n_513, n_512);
  nand g1427 (n_1378, n_511, n_513);
  nand g1428 (n_531, n_1376, n_1377, n_1378);
  xor g1429 (n_1379, n_514, n_515);
  xor g1430 (n_89, n_1379, n_516);
  nand g1431 (n_1380, n_514, n_515);
  nand g1432 (n_1381, n_516, n_515);
  nand g1433 (n_1382, n_514, n_516);
  nand g1434 (n_40, n_1380, n_1381, n_1382);
  xor g1437 (n_1383, A[10], A[14]);
  xor g1438 (n_521, n_1383, A[10]);
  xor g1444 (n_522, n_1387, A[19]);
  nand g1446 (n_1389, A[19], A[15]);
  nand g1448 (n_535, n_1388, n_1389, n_1390);
  xor g1449 (n_1391, A[18], n_520);
  xor g1450 (n_524, n_1391, n_521);
  nand g1451 (n_1392, A[18], n_520);
  nand g1452 (n_1393, n_521, n_520);
  nand g1453 (n_1394, A[18], n_521);
  nand g1454 (n_538, n_1392, n_1393, n_1394);
  xor g1455 (n_1395, A[23], A[22]);
  xor g1456 (n_527, n_1395, n_522);
  nand g1458 (n_1397, n_522, A[22]);
  nand g1459 (n_1398, A[23], n_522);
  nand g1460 (n_540, n_1114, n_1397, n_1398);
  xor g1461 (n_1399, n_523, n_524);
  xor g1462 (n_528, n_1399, n_525);
  nand g1463 (n_1400, n_523, n_524);
  nand g1464 (n_1401, n_525, n_524);
  nand g1465 (n_1402, n_523, n_525);
  nand g1466 (n_541, n_1400, n_1401, n_1402);
  xor g1467 (n_1403, n_526, n_527);
  xor g1468 (n_530, n_1403, n_528);
  nand g1469 (n_1404, n_526, n_527);
  nand g1470 (n_1405, n_528, n_527);
  nand g1471 (n_1406, n_526, n_528);
  nand g1472 (n_544, n_1404, n_1405, n_1406);
  xor g1473 (n_1407, n_529, n_530);
  xor g1474 (n_88, n_1407, n_531);
  nand g1475 (n_1408, n_529, n_530);
  nand g1476 (n_1409, n_531, n_530);
  nand g1477 (n_1410, n_529, n_531);
  nand g1478 (n_39, n_1408, n_1409, n_1410);
  xor g1480 (n_534, n_743, A[11]);
  nand g1490 (n_547, n_850, n_1188, n_1418);
  xor g1492 (n_537, n_983, A[23]);
  nand g1495 (n_1422, A[19], A[23]);
  nand g1496 (n_549, n_984, n_1025, n_1422);
  xor g1497 (n_1423, n_533, n_534);
  xor g1498 (n_539, n_1423, n_535);
  nand g1499 (n_1424, n_533, n_534);
  nand g1500 (n_1425, n_535, n_534);
  nand g1501 (n_1426, n_533, n_535);
  nand g1502 (n_551, n_1424, n_1425, n_1426);
  xor g1503 (n_1427, n_536, n_537);
  xor g1504 (n_542, n_1427, n_538);
  nand g1505 (n_1428, n_536, n_537);
  nand g1506 (n_1429, n_538, n_537);
  nand g1507 (n_1430, n_536, n_538);
  nand g1508 (n_552, n_1428, n_1429, n_1430);
  xor g1509 (n_1431, n_539, n_540);
  xor g1510 (n_543, n_1431, n_541);
  nand g1511 (n_1432, n_539, n_540);
  nand g1512 (n_1433, n_541, n_540);
  nand g1513 (n_1434, n_539, n_541);
  nand g1514 (n_555, n_1432, n_1433, n_1434);
  xor g1515 (n_1435, n_542, n_543);
  xor g1516 (n_87, n_1435, n_544);
  nand g1517 (n_1436, n_542, n_543);
  nand g1518 (n_1437, n_544, n_543);
  nand g1519 (n_1438, n_542, n_544);
  nand g1520 (n_38, n_1436, n_1437, n_1438);
  xor g1522 (n_546, n_1183, A[16]);
  nand g1526 (n_558, n_1184, n_1330, n_878);
  xor g1528 (n_548, n_1443, A[20]);
  nand g1532 (n_559, n_1065, n_917, n_1302);
  xor g1533 (n_1447, A[21], n_545);
  xor g1534 (n_550, n_1447, n_546);
  nand g1535 (n_1448, A[21], n_545);
  nand g1536 (n_1449, n_546, n_545);
  nand g1537 (n_1450, A[21], n_546);
  nand g1538 (n_562, n_1448, n_1449, n_1450);
  xor g1539 (n_1451, n_547, n_548);
  xor g1540 (n_553, n_1451, n_549);
  nand g1541 (n_1452, n_547, n_548);
  nand g1542 (n_1453, n_549, n_548);
  nand g1543 (n_1454, n_547, n_549);
  nand g1544 (n_563, n_1452, n_1453, n_1454);
  xor g1545 (n_1455, n_550, n_551);
  xor g1546 (n_554, n_1455, n_552);
  nand g1547 (n_1456, n_550, n_551);
  nand g1548 (n_1457, n_552, n_551);
  nand g1549 (n_1458, n_550, n_552);
  nand g1550 (n_566, n_1456, n_1457, n_1458);
  xor g1551 (n_1459, n_553, n_554);
  xor g1552 (n_86, n_1459, n_555);
  nand g1553 (n_1460, n_553, n_554);
  nand g1554 (n_1461, n_555, n_554);
  nand g1555 (n_1462, n_553, n_555);
  nand g1556 (n_37, n_1460, n_1461, n_1462);
  xor g1560 (n_560, n_1463, A[18]);
  nand g1563 (n_1466, A[13], A[18]);
  nand g1564 (n_570, n_1464, n_1465, n_1466);
  xor g1565 (n_1467, A[17], A[21]);
  xor g1566 (n_561, n_1467, A[22]);
  nand g1567 (n_1468, A[17], A[21]);
  nand g1569 (n_1470, A[17], A[22]);
  nand g1570 (n_572, n_1468, n_1069, n_1470);
  xor g1571 (n_1471, n_558, n_559);
  xor g1572 (n_564, n_1471, n_560);
  nand g1573 (n_1472, n_558, n_559);
  nand g1574 (n_1473, n_560, n_559);
  nand g1575 (n_1474, n_558, n_560);
  nand g1576 (n_574, n_1472, n_1473, n_1474);
  xor g1577 (n_1475, n_561, n_562);
  xor g1578 (n_565, n_1475, n_563);
  nand g1579 (n_1476, n_561, n_562);
  nand g1580 (n_1477, n_563, n_562);
  nand g1581 (n_1478, n_561, n_563);
  nand g1582 (n_577, n_1476, n_1477, n_1478);
  xor g1583 (n_1479, n_564, n_565);
  xor g1584 (n_85, n_1479, n_566);
  nand g1585 (n_1480, n_564, n_565);
  nand g1586 (n_1481, n_566, n_565);
  nand g1587 (n_1482, n_564, n_566);
  nand g1588 (n_36, n_1480, n_1481, n_1482);
  xor g1597 (n_1487, A[19], A[18]);
  xor g1598 (n_573, n_1487, A[22]);
  nand g1600 (n_1489, A[22], A[18]);
  nand g1601 (n_1490, A[19], A[22]);
  nand g1602 (n_582, n_1110, n_1489, n_1490);
  xor g1603 (n_1491, A[23], n_570);
  xor g1604 (n_575, n_1491, n_571);
  nand g1605 (n_1492, A[23], n_570);
  nand g1606 (n_1493, n_571, n_570);
  nand g1607 (n_1494, A[23], n_571);
  nand g1608 (n_583, n_1492, n_1493, n_1494);
  xor g1609 (n_1495, n_572, n_573);
  xor g1610 (n_576, n_1495, n_574);
  nand g1611 (n_1496, n_572, n_573);
  nand g1612 (n_1497, n_574, n_573);
  nand g1613 (n_1498, n_572, n_574);
  nand g1614 (n_586, n_1496, n_1497, n_1498);
  xor g1615 (n_1499, n_575, n_576);
  xor g1616 (n_84, n_1499, n_577);
  nand g1617 (n_1500, n_575, n_576);
  nand g1618 (n_1501, n_577, n_576);
  nand g1619 (n_1502, n_575, n_577);
  nand g1620 (n_35, n_1500, n_1501, n_1502);
  xor g1622 (n_580, n_979, A[14]);
  nand g1624 (n_1505, A[14], A[16]);
  nand g1626 (n_587, n_850, n_1505, n_944);
  xor g1633 (n_1511, A[23], n_579);
  xor g1634 (n_584, n_1511, n_580);
  nand g1635 (n_1512, A[23], n_579);
  nand g1636 (n_1513, n_580, n_579);
  nand g1637 (n_1514, A[23], n_580);
  nand g1638 (n_591, n_1512, n_1513, n_1514);
  xor g1639 (n_1515, n_478, n_582);
  xor g1640 (n_585, n_1515, n_583);
  nand g1641 (n_1516, n_478, n_582);
  nand g1642 (n_1517, n_583, n_582);
  nand g1643 (n_1518, n_478, n_583);
  nand g1644 (n_593, n_1516, n_1517, n_1518);
  xor g1645 (n_1519, n_584, n_585);
  xor g1646 (n_83, n_1519, n_586);
  nand g1647 (n_1520, n_584, n_585);
  nand g1648 (n_1521, n_586, n_585);
  nand g1649 (n_1522, n_584, n_586);
  nand g1650 (n_34, n_1520, n_1521, n_1522);
  xor g1652 (n_589, n_1187, A[17]);
  nand g1655 (n_1526, A[16], A[17]);
  nand g1656 (n_596, n_1188, n_1065, n_1526);
  xor g1658 (n_590, n_1335, n_587);
  nand g1660 (n_1529, n_587, A[21]);
  nand g1661 (n_1530, A[20], n_587);
  nand g1662 (n_597, n_1336, n_1529, n_1530);
  xor g1663 (n_1531, n_491, n_589);
  xor g1664 (n_592, n_1531, n_590);
  nand g1665 (n_1532, n_491, n_589);
  nand g1666 (n_1533, n_590, n_589);
  nand g1667 (n_1534, n_491, n_590);
  nand g1668 (n_600, n_1532, n_1533, n_1534);
  xor g1669 (n_1535, n_591, n_592);
  xor g1670 (n_82, n_1535, n_593);
  nand g1671 (n_1536, n_591, n_592);
  nand g1672 (n_1537, n_593, n_592);
  nand g1673 (n_1538, n_591, n_593);
  nand g1674 (n_33, n_1536, n_1537, n_1538);
  xor g1684 (n_599, n_1543, n_597);
  nand g1686 (n_1545, n_597, n_596);
  nand g1688 (n_607, n_1544, n_1545, n_1546);
  xor g1689 (n_1547, n_561, n_599);
  xor g1690 (n_81, n_1547, n_600);
  nand g1691 (n_1548, n_561, n_599);
  nand g1692 (n_1549, n_600, n_599);
  nand g1693 (n_1550, n_561, n_600);
  nand g1694 (n_32, n_1548, n_1549, n_1550);
  xor g1697 (n_1551, A[18], A[22]);
  xor g1698 (n_605, n_1551, A[23]);
  nand g1701 (n_1554, A[18], A[23]);
  nand g1702 (n_610, n_1489, n_1114, n_1554);
  nand g1706 (n_1557, n_572, A[18]);
  nand g1708 (n_612, n_1556, n_1557, n_1558);
  xor g1709 (n_1559, n_605, n_606);
  xor g1710 (n_80, n_1559, n_607);
  nand g1711 (n_1560, n_605, n_606);
  nand g1712 (n_1561, n_607, n_606);
  nand g1713 (n_1562, n_605, n_607);
  nand g1714 (n_31, n_1560, n_1561, n_1562);
  xor g1721 (n_1567, A[23], A[19]);
  xor g1722 (n_611, n_1567, n_478);
  nand g1724 (n_1569, n_478, A[19]);
  nand g1725 (n_1570, A[23], n_478);
  nand g1726 (n_615, n_1422, n_1569, n_1570);
  xor g1727 (n_1571, n_610, n_611);
  xor g1728 (n_79, n_1571, n_612);
  nand g1729 (n_1572, n_610, n_611);
  nand g1730 (n_1573, n_612, n_611);
  nand g1731 (n_1574, n_610, n_612);
  nand g1732 (n_30, n_1572, n_1573, n_1574);
  xor g1734 (n_614, n_1575, A[21]);
  nand g1738 (n_618, n_1302, n_1336, n_1578);
  xor g1739 (n_1579, n_491, n_614);
  xor g1740 (n_78, n_1579, n_615);
  nand g1741 (n_1580, n_491, n_614);
  nand g1742 (n_1581, n_615, n_614);
  nand g1743 (n_1582, n_491, n_615);
  nand g1744 (n_77, n_1580, n_1581, n_1582);
  xor g1748 (n_29, n_1583, n_618);
  nand g1751 (n_1586, A[22], n_618);
  nand g1752 (n_28, n_1584, n_1585, n_1586);
  nand g1759 (n_1590, A[23], A[21]);
  nand g1760 (n_27, n_1588, n_1589, n_1590);
  xor g1762 (n_75, n_1591, A[22]);
  nand g1766 (n_74, n_1592, n_1114, n_1594);
  nor g11 (n_1610, A[0], A[2]);
  nand g12 (n_1605, A[0], A[2]);
  nor g13 (n_1606, n_69, A[3]);
  nand g14 (n_1607, n_69, A[3]);
  nor g15 (n_1616, A[4], n_117);
  nand g16 (n_1611, A[4], n_117);
  nor g17 (n_1612, A[5], n_116);
  nand g18 (n_1613, A[5], n_116);
  nor g19 (n_1622, A[6], n_115);
  nand g20 (n_1617, A[6], n_115);
  nor g21 (n_1618, n_66, n_114);
  nand g22 (n_1619, n_66, n_114);
  nor g23 (n_1628, n_65, n_113);
  nand g24 (n_1623, n_65, n_113);
  nor g25 (n_1624, n_64, n_112);
  nand g26 (n_1625, n_64, n_112);
  nor g27 (n_1634, n_63, n_111);
  nand g28 (n_1629, n_63, n_111);
  nor g29 (n_1630, n_62, n_110);
  nand g30 (n_1631, n_62, n_110);
  nor g31 (n_1640, n_61, n_109);
  nand g32 (n_1635, n_61, n_109);
  nor g33 (n_1636, n_60, n_108);
  nand g34 (n_1637, n_60, n_108);
  nor g35 (n_1646, n_59, n_107);
  nand g36 (n_1641, n_59, n_107);
  nor g37 (n_1642, n_58, n_106);
  nand g38 (n_1643, n_58, n_106);
  nor g39 (n_1652, n_57, n_105);
  nand g40 (n_1647, n_57, n_105);
  nor g41 (n_1648, n_56, n_104);
  nand g42 (n_1649, n_56, n_104);
  nor g43 (n_1658, n_55, n_103);
  nand g44 (n_1653, n_55, n_103);
  nor g45 (n_1654, n_54, n_102);
  nand g46 (n_1655, n_54, n_102);
  nor g47 (n_1664, n_53, n_101);
  nand g48 (n_1659, n_53, n_101);
  nor g49 (n_1660, n_52, n_100);
  nand g50 (n_1661, n_52, n_100);
  nor g51 (n_1670, n_51, n_99);
  nand g52 (n_1665, n_51, n_99);
  nor g53 (n_1666, n_50, n_98);
  nand g54 (n_1667, n_50, n_98);
  nor g55 (n_1676, n_49, n_97);
  nand g56 (n_1671, n_49, n_97);
  nor g57 (n_1672, n_48, n_96);
  nand g58 (n_1673, n_48, n_96);
  nor g59 (n_1682, n_47, n_95);
  nand g60 (n_1677, n_47, n_95);
  nor g61 (n_1678, n_46, n_94);
  nand g62 (n_1679, n_46, n_94);
  nor g63 (n_1688, n_45, n_93);
  nand g64 (n_1683, n_45, n_93);
  nor g65 (n_1684, n_44, n_92);
  nand g66 (n_1685, n_44, n_92);
  nor g67 (n_1694, n_43, n_91);
  nand g68 (n_1689, n_43, n_91);
  nor g69 (n_1690, n_42, n_90);
  nand g70 (n_1691, n_42, n_90);
  nor g71 (n_1700, n_41, n_89);
  nand g72 (n_1695, n_41, n_89);
  nor g73 (n_1696, n_40, n_88);
  nand g74 (n_1697, n_40, n_88);
  nor g75 (n_1706, n_39, n_87);
  nand g76 (n_1701, n_39, n_87);
  nor g77 (n_1702, n_38, n_86);
  nand g78 (n_1703, n_38, n_86);
  nor g79 (n_1712, n_37, n_85);
  nand g80 (n_1707, n_37, n_85);
  nor g81 (n_1708, n_36, n_84);
  nand g82 (n_1709, n_36, n_84);
  nor g83 (n_1718, n_35, n_83);
  nand g84 (n_1713, n_35, n_83);
  nor g85 (n_1714, n_34, n_82);
  nand g86 (n_1715, n_34, n_82);
  nor g87 (n_1724, n_33, n_81);
  nand g88 (n_1719, n_33, n_81);
  nor g89 (n_1720, n_32, n_80);
  nand g90 (n_1721, n_32, n_80);
  nor g91 (n_1730, n_31, n_79);
  nand g92 (n_1725, n_31, n_79);
  nor g93 (n_1726, n_30, n_78);
  nand g94 (n_1727, n_30, n_78);
  nor g95 (n_1736, n_29, n_77);
  nand g96 (n_1731, n_29, n_77);
  nor g97 (n_1732, n_28, n_76);
  nand g98 (n_1733, n_28, n_76);
  nor g99 (n_1740, n_27, n_75);
  nand g100 (n_1737, n_27, n_75);
  nor g106 (n_1608, n_1605, n_1606);
  nor g110 (n_1614, n_1611, n_1612);
  nor g113 (n_1750, n_1616, n_1612);
  nor g114 (n_1620, n_1617, n_1618);
  nor g117 (n_1752, n_1622, n_1618);
  nor g118 (n_1626, n_1623, n_1624);
  nor g121 (n_1760, n_1628, n_1624);
  nor g122 (n_1632, n_1629, n_1630);
  nor g125 (n_1762, n_1634, n_1630);
  nor g126 (n_1638, n_1635, n_1636);
  nor g129 (n_1770, n_1640, n_1636);
  nor g130 (n_1644, n_1641, n_1642);
  nor g133 (n_1772, n_1646, n_1642);
  nor g134 (n_1650, n_1647, n_1648);
  nor g137 (n_1780, n_1652, n_1648);
  nor g138 (n_1656, n_1653, n_1654);
  nor g141 (n_1782, n_1658, n_1654);
  nor g142 (n_1662, n_1659, n_1660);
  nor g145 (n_1790, n_1664, n_1660);
  nor g146 (n_1668, n_1665, n_1666);
  nor g149 (n_1792, n_1670, n_1666);
  nor g150 (n_1674, n_1671, n_1672);
  nor g153 (n_1800, n_1676, n_1672);
  nor g154 (n_1680, n_1677, n_1678);
  nor g157 (n_1802, n_1682, n_1678);
  nor g158 (n_1686, n_1683, n_1684);
  nor g161 (n_1810, n_1688, n_1684);
  nor g162 (n_1692, n_1689, n_1690);
  nor g165 (n_1812, n_1694, n_1690);
  nor g166 (n_1698, n_1695, n_1696);
  nor g169 (n_1820, n_1700, n_1696);
  nor g170 (n_1704, n_1701, n_1702);
  nor g173 (n_1822, n_1706, n_1702);
  nor g174 (n_1710, n_1707, n_1708);
  nor g177 (n_1830, n_1712, n_1708);
  nor g178 (n_1716, n_1713, n_1714);
  nor g181 (n_1832, n_1718, n_1714);
  nor g182 (n_1722, n_1719, n_1720);
  nor g185 (n_1840, n_1724, n_1720);
  nor g186 (n_1728, n_1725, n_1726);
  nor g189 (n_1842, n_1730, n_1726);
  nor g190 (n_1734, n_1731, n_1732);
  nor g193 (n_1850, n_1736, n_1732);
  nor g203 (n_1748, n_1622, n_1747);
  nand g212 (n_1860, n_1750, n_1752);
  nor g213 (n_1758, n_1634, n_1757);
  nand g222 (n_1867, n_1760, n_1762);
  nor g223 (n_1768, n_1646, n_1767);
  nand g232 (n_1875, n_1770, n_1772);
  nor g233 (n_1778, n_1658, n_1777);
  nand g242 (n_1882, n_1780, n_1782);
  nor g243 (n_1788, n_1670, n_1787);
  nand g252 (n_1890, n_1790, n_1792);
  nor g253 (n_1798, n_1682, n_1797);
  nand g262 (n_1897, n_1800, n_1802);
  nor g263 (n_1808, n_1694, n_1807);
  nand g1776 (n_1905, n_1810, n_1812);
  nor g1777 (n_1818, n_1706, n_1817);
  nand g1786 (n_1912, n_1820, n_1822);
  nor g1787 (n_1828, n_1718, n_1827);
  nand g1796 (n_1920, n_1830, n_1832);
  nor g1797 (n_1838, n_1730, n_1837);
  nand g1806 (n_1927, n_1840, n_1842);
  nor g1807 (n_1848, n_1740, n_1847);
  nand g1814 (n_2131, n_1611, n_1854);
  nand g1816 (n_2133, n_1747, n_1855);
  nand g1819 (n_2136, n_1858, n_1859);
  nand g1822 (n_1935, n_1862, n_1863);
  nor g1823 (n_1865, n_1640, n_1864);
  nor g1826 (n_1945, n_1640, n_1867);
  nor g1832 (n_1873, n_1871, n_1864);
  nor g1835 (n_1951, n_1867, n_1871);
  nor g1836 (n_1877, n_1875, n_1864);
  nor g1839 (n_1954, n_1867, n_1875);
  nor g1840 (n_1880, n_1664, n_1879);
  nor g1843 (n_2034, n_1664, n_1882);
  nor g1849 (n_1888, n_1886, n_1879);
  nor g1852 (n_2040, n_1882, n_1886);
  nor g1853 (n_1892, n_1890, n_1879);
  nor g1856 (n_1960, n_1882, n_1890);
  nor g1857 (n_1895, n_1688, n_1894);
  nor g1860 (n_1973, n_1688, n_1897);
  nor g1866 (n_1903, n_1901, n_1894);
  nor g1869 (n_1983, n_1897, n_1901);
  nor g1870 (n_1907, n_1905, n_1894);
  nor g1873 (n_1988, n_1897, n_1905);
  nor g1874 (n_1910, n_1712, n_1909);
  nor g1877 (n_2086, n_1712, n_1912);
  nor g1883 (n_1918, n_1916, n_1909);
  nor g1886 (n_2092, n_1912, n_1916);
  nor g1887 (n_1922, n_1920, n_1909);
  nor g1890 (n_1996, n_1912, n_1920);
  nor g1891 (n_1925, n_1736, n_1924);
  nor g1894 (n_2009, n_1736, n_1927);
  nor g1900 (n_1933, n_1931, n_1924);
  nor g1903 (n_2019, n_1927, n_1931);
  nand g1906 (n_2140, n_1623, n_1937);
  nand g1907 (n_1938, n_1760, n_1935);
  nand g1908 (n_2142, n_1757, n_1938);
  nand g1911 (n_2145, n_1941, n_1942);
  nand g1914 (n_2148, n_1864, n_1944);
  nand g1915 (n_1947, n_1945, n_1935);
  nand g1916 (n_2151, n_1946, n_1947);
  nand g1917 (n_1950, n_1948, n_1935);
  nand g1918 (n_2153, n_1949, n_1950);
  nand g1919 (n_1953, n_1951, n_1935);
  nand g1920 (n_2156, n_1952, n_1953);
  nand g1921 (n_1956, n_1954, n_1935);
  nand g1922 (n_2024, n_1955, n_1956);
  nor g1923 (n_1958, n_1676, n_1957);
  nand g1932 (n_2048, n_1800, n_1960);
  nor g1933 (n_1967, n_1965, n_1957);
  nor g1938 (n_1970, n_1897, n_1957);
  nand g1947 (n_2060, n_1960, n_1973);
  nand g1952 (n_2064, n_1960, n_1978);
  nand g1957 (n_2068, n_1960, n_1983);
  nand g1962 (n_2072, n_1960, n_1988);
  nor g1963 (n_1994, n_1724, n_1993);
  nand g1972 (n_2100, n_1840, n_1996);
  nor g1973 (n_2003, n_2001, n_1993);
  nor g1978 (n_2006, n_1927, n_1993);
  nand g1987 (n_2112, n_1996, n_2009);
  nand g1992 (n_2116, n_1996, n_2014);
  nand g1997 (n_2120, n_1996, n_2019);
  nand g2000 (n_2160, n_1647, n_2026);
  nand g2001 (n_2027, n_1780, n_2024);
  nand g2002 (n_2162, n_1777, n_2027);
  nand g2005 (n_2165, n_2030, n_2031);
  nand g2008 (n_2168, n_1879, n_2033);
  nand g2009 (n_2036, n_2034, n_2024);
  nand g2010 (n_2171, n_2035, n_2036);
  nand g2011 (n_2039, n_2037, n_2024);
  nand g2012 (n_2173, n_2038, n_2039);
  nand g2013 (n_2042, n_2040, n_2024);
  nand g2014 (n_2176, n_2041, n_2042);
  nand g2015 (n_2043, n_1960, n_2024);
  nand g2016 (n_2178, n_1957, n_2043);
  nand g2019 (n_2181, n_2046, n_2047);
  nand g2022 (n_2183, n_2050, n_2051);
  nand g2025 (n_2186, n_2054, n_2055);
  nand g2028 (n_2189, n_2058, n_2059);
  nand g2031 (n_2192, n_2062, n_2063);
  nand g2034 (n_2194, n_2066, n_2067);
  nand g2037 (n_2197, n_2070, n_2071);
  nand g2040 (n_2076, n_2074, n_2075);
  nand g2043 (n_2201, n_1695, n_2078);
  nand g2044 (n_2079, n_1820, n_2076);
  nand g2045 (n_2203, n_1817, n_2079);
  nand g2048 (n_2206, n_2082, n_2083);
  nand g2051 (n_2209, n_1909, n_2085);
  nand g2052 (n_2088, n_2086, n_2076);
  nand g2053 (n_2212, n_2087, n_2088);
  nand g2054 (n_2091, n_2089, n_2076);
  nand g2055 (n_2214, n_2090, n_2091);
  nand g2056 (n_2094, n_2092, n_2076);
  nand g2057 (n_2217, n_2093, n_2094);
  nand g2058 (n_2095, n_1996, n_2076);
  nand g2059 (n_2219, n_1993, n_2095);
  nand g2062 (n_2222, n_2098, n_2099);
  nand g2065 (n_2224, n_2102, n_2103);
  nand g2068 (n_2227, n_2106, n_2107);
  nand g2071 (n_2230, n_2110, n_2111);
  nand g2074 (n_2233, n_2114, n_2115);
  nand g2077 (n_2235, n_2118, n_2119);
  nand g2080 (n_2238, n_2122, n_2123);
  xnor g2092 (Z[5], n_2131, n_2132);
  xnor g2094 (Z[6], n_2133, n_2134);
  xnor g2097 (Z[7], n_2136, n_2137);
  xnor g2099 (Z[8], n_1935, n_2138);
  xnor g2102 (Z[9], n_2140, n_2141);
  xnor g2104 (Z[10], n_2142, n_2143);
  xnor g2107 (Z[11], n_2145, n_2146);
  xnor g2110 (Z[12], n_2148, n_2149);
  xnor g2113 (Z[13], n_2151, n_2152);
  xnor g2115 (Z[14], n_2153, n_2154);
  xnor g2118 (Z[15], n_2156, n_2157);
  xnor g2120 (Z[16], n_2024, n_2158);
  xnor g2123 (Z[17], n_2160, n_2161);
  xnor g2125 (Z[18], n_2162, n_2163);
  xnor g2128 (Z[19], n_2165, n_2166);
  xnor g2131 (Z[20], n_2168, n_2169);
  xnor g2134 (Z[21], n_2171, n_2172);
  xnor g2136 (Z[22], n_2173, n_2174);
  xnor g2139 (Z[23], n_2176, n_2177);
  xnor g2141 (Z[24], n_2178, n_2179);
  xnor g2144 (Z[25], n_2181, n_2182);
  xnor g2146 (Z[26], n_2183, n_2184);
  xnor g2149 (Z[27], n_2186, n_2187);
  xnor g2152 (Z[28], n_2189, n_2190);
  xnor g2155 (Z[29], n_2192, n_2193);
  xnor g2157 (Z[30], n_2194, n_2195);
  xnor g2160 (Z[31], n_2197, n_2198);
  xnor g2162 (Z[32], n_2076, n_2199);
  xnor g2165 (Z[33], n_2201, n_2202);
  xnor g2167 (Z[34], n_2203, n_2204);
  xnor g2170 (Z[35], n_2206, n_2207);
  xnor g2173 (Z[36], n_2209, n_2210);
  xnor g2176 (Z[37], n_2212, n_2213);
  xnor g2178 (Z[38], n_2214, n_2215);
  xnor g2181 (Z[39], n_2217, n_2218);
  xnor g2183 (Z[40], n_2219, n_2220);
  xnor g2186 (Z[41], n_2222, n_2223);
  xnor g2188 (Z[42], n_2224, n_2225);
  xnor g2191 (Z[43], n_2227, n_2228);
  xnor g2194 (Z[44], n_2230, n_2231);
  xnor g2197 (Z[45], n_2233, n_2234);
  xnor g2199 (Z[46], n_2235, n_2236);
  xnor g2202 (Z[47], n_2238, n_2239);
  or g2215 (n_1045, A[1], wc);
  not gc (wc, n_171);
  or g2216 (n_1046, A[1], wc0);
  not gc0 (wc0, A[2]);
  or g2217 (n_1065, wc1, A[24]);
  not gc1 (wc1, A[17]);
  or g2218 (n_1089, A[2], wc2);
  not gc2 (wc2, A[3]);
  or g2219 (n_1090, wc3, A[2]);
  not gc3 (wc3, A[1]);
  xnor g2220 (n_1151, A[24], A[19]);
  or g2221 (n_1152, wc4, A[24]);
  not gc4 (wc4, A[19]);
  xnor g2222 (n_1187, A[24], A[16]);
  or g2223 (n_1188, wc5, A[24]);
  not gc5 (wc5, A[16]);
  xnor g2224 (n_1215, A[6], A[5]);
  or g2225 (n_1216, A[5], wc6);
  not gc6 (wc6, A[6]);
  or g2226 (n_1217, A[5], wc7);
  not gc7 (wc7, A[9]);
  xnor g2228 (n_1255, A[11], A[7]);
  or g2229 (n_1256, A[7], wc8);
  not gc8 (wc8, A[11]);
  or g2230 (n_1257, A[7], wc9);
  not gc9 (wc9, A[14]);
  or g2231 (n_1302, wc10, A[24]);
  not gc10 (wc10, A[20]);
  xnor g2232 (n_1359, A[18], A[10]);
  or g2233 (n_1360, A[10], wc11);
  not gc11 (wc11, A[18]);
  or g2234 (n_1362, A[10], wc12);
  not gc12 (wc12, A[17]);
  xnor g2236 (n_1387, A[15], A[11]);
  or g2237 (n_1388, A[11], wc13);
  not gc13 (wc13, A[15]);
  or g2238 (n_1390, A[11], wc14);
  not gc14 (wc14, A[19]);
  xnor g2240 (n_536, n_979, A[24]);
  or g2241 (n_1418, wc15, A[24]);
  not gc15 (wc15, A[15]);
  xnor g2242 (n_1443, A[24], A[17]);
  xnor g2243 (n_1463, A[14], A[13]);
  or g2244 (n_1464, wc16, A[14]);
  not gc16 (wc16, A[13]);
  or g2245 (n_1465, A[14], wc17);
  not gc17 (wc17, A[18]);
  or g2246 (n_1486, A[14], wc18);
  not gc18 (wc18, A[15]);
  or g2248 (n_1556, wc19, A[19]);
  not gc19 (wc19, A[18]);
  xnor g2249 (n_1575, A[24], A[20]);
  or g2250 (n_1578, wc20, A[24]);
  not gc20 (wc20, A[21]);
  xnor g2251 (n_1583, A[22], A[21]);
  or g2252 (n_1584, A[21], wc21);
  not gc21 (wc21, A[22]);
  or g2254 (n_1588, A[22], wc22);
  not gc22 (wc22, A[23]);
  or g2255 (n_1589, wc23, A[22]);
  not gc23 (wc23, A[21]);
  xnor g2256 (n_1591, A[24], A[23]);
  or g2257 (n_1592, wc24, A[24]);
  not gc24 (wc24, A[23]);
  or g2258 (n_1594, wc25, A[24]);
  not gc25 (wc25, A[22]);
  xnor g2259 (n_350, n_1043, A[1]);
  xnor g2260 (n_373, n_1087, A[2]);
  or g2261 (n_1154, A[24], wc26);
  not gc26 (wc26, n_399);
  xnor g2262 (n_454, n_1215, A[10]);
  xnor g2263 (n_1331, n_488, A[24]);
  or g2264 (n_1332, A[24], wc27);
  not gc27 (wc27, n_488);
  or g2265 (n_533, A[10], wc28);
  not gc28 (wc28, n_818);
  or g2266 (n_545, A[11], wc29);
  not gc29 (wc29, n_744);
  xnor g2267 (n_571, n_943, A[14]);
  nand g2268 (n_579, n_944, n_1486);
  xnor g2269 (n_606, n_572, n_1487);
  or g2270 (n_1558, A[19], wc30);
  not gc30 (wc30, n_572);
  xnor g2271 (n_76, n_1395, A[21]);
  or g2273 (n_2125, wc31, n_1610);
  not gc31 (wc31, n_1605);
  xnor g2274 (n_1543, n_596, A[18]);
  or g2275 (n_1544, A[18], wc32);
  not gc32 (wc32, n_596);
  or g2276 (n_1585, A[21], wc33);
  not gc33 (wc33, n_618);
  and g2277 (n_1745, wc34, n_1607);
  not gc34 (wc34, n_1608);
  or g2278 (n_2128, wc35, n_1606);
  not gc35 (wc35, n_1607);
  and g2279 (n_1738, wc36, n_74);
  not gc36 (wc36, A[24]);
  or g2280 (n_1739, wc37, n_74);
  not gc37 (wc37, A[24]);
  not g2281 (Z[2], n_2125);
  or g2282 (n_1189, A[24], wc38);
  not gc38 (wc38, n_416);
  or g2283 (n_1546, A[18], wc39);
  not gc39 (wc39, n_597);
  or g2286 (n_2129, wc40, n_1616);
  not gc40 (wc40, n_1611);
  or g2287 (n_2236, wc41, n_1740);
  not gc41 (wc41, n_1737);
  and g2288 (n_1747, wc42, n_1613);
  not gc42 (wc42, n_1614);
  or g2289 (n_1854, n_1616, n_1745);
  or g2290 (n_1855, n_1745, wc43);
  not gc43 (wc43, n_1750);
  xor g2291 (Z[3], n_1605, n_2128);
  xor g2292 (Z[4], n_1745, n_2129);
  or g2293 (n_2132, wc44, n_1612);
  not gc44 (wc44, n_1613);
  or g2294 (n_2239, wc45, n_1738);
  not gc45 (wc45, n_1739);
  or g2295 (n_2234, wc46, n_1732);
  not gc46 (wc46, n_1733);
  and g2296 (n_1858, wc47, n_1617);
  not gc47 (wc47, n_1748);
  or g2297 (n_1856, wc48, n_1622);
  not gc48 (wc48, n_1750);
  or g2298 (n_2134, wc49, n_1622);
  not gc49 (wc49, n_1617);
  or g2299 (n_2138, wc50, n_1628);
  not gc50 (wc50, n_1623);
  or g2300 (n_2228, wc51, n_1726);
  not gc51 (wc51, n_1727);
  or g2301 (n_1066, A[24], wc52);
  not gc52 (wc52, n_234);
  and g2302 (n_1754, wc53, n_1619);
  not gc53 (wc53, n_1620);
  and g2303 (n_1757, wc54, n_1625);
  not gc54 (wc54, n_1626);
  and g2304 (n_1847, wc55, n_1733);
  not gc55 (wc55, n_1734);
  or g2305 (n_1931, wc56, n_1740);
  not gc56 (wc56, n_1850);
  or g2306 (n_2137, wc57, n_1618);
  not gc57 (wc57, n_1619);
  or g2307 (n_2141, wc58, n_1624);
  not gc58 (wc58, n_1625);
  or g2308 (n_2231, wc59, n_1736);
  not gc59 (wc59, n_1731);
  xnor g2309 (n_361, n_1063, A[24]);
  and g2310 (n_1755, wc60, n_1752);
  not gc60 (wc60, n_1747);
  or g2311 (n_1939, wc61, n_1634);
  not gc61 (wc61, n_1760);
  or g2312 (n_1859, n_1745, n_1856);
  or g2313 (n_2143, wc62, n_1634);
  not gc62 (wc62, n_1629);
  or g2314 (n_2223, wc63, n_1720);
  not gc63 (wc63, n_1721);
  and g2315 (n_1834, wc64, n_1715);
  not gc64 (wc64, n_1716);
  and g2316 (n_1837, wc65, n_1721);
  not gc65 (wc65, n_1722);
  and g2317 (n_1844, wc66, n_1727);
  not gc66 (wc66, n_1728);
  and g2318 (n_1862, wc67, n_1754);
  not gc67 (wc67, n_1755);
  and g2319 (n_1941, wc68, n_1629);
  not gc68 (wc68, n_1758);
  or g2320 (n_2001, wc69, n_1730);
  not gc69 (wc69, n_1840);
  and g2321 (n_1932, wc70, n_1737);
  not gc70 (wc70, n_1848);
  or g2322 (n_1863, n_1860, n_1745);
  or g2323 (n_2215, wc71, n_1718);
  not gc71 (wc71, n_1713);
  or g2324 (n_2218, wc72, n_1714);
  not gc72 (wc72, n_1715);
  or g2325 (n_2220, wc73, n_1724);
  not gc73 (wc73, n_1719);
  or g2326 (n_2225, wc74, n_1730);
  not gc74 (wc74, n_1725);
  and g2327 (n_1764, wc75, n_1631);
  not gc75 (wc75, n_1632);
  and g2328 (n_1827, wc76, n_1709);
  not gc76 (wc76, n_1710);
  or g2329 (n_1916, wc77, n_1718);
  not gc77 (wc77, n_1830);
  and g2330 (n_1845, wc78, n_1842);
  not gc78 (wc78, n_1837);
  and g2331 (n_2014, wc79, n_1850);
  not gc79 (wc79, n_1927);
  or g2332 (n_2146, wc80, n_1630);
  not gc80 (wc80, n_1631);
  or g2333 (n_2154, wc81, n_1646);
  not gc81 (wc81, n_1641);
  or g2334 (n_2207, wc82, n_1702);
  not gc82 (wc82, n_1703);
  or g2335 (n_2210, wc83, n_1712);
  not gc83 (wc83, n_1707);
  or g2336 (n_2213, wc84, n_1708);
  not gc84 (wc84, n_1709);
  and g2337 (n_1767, wc85, n_1637);
  not gc85 (wc85, n_1638);
  and g2338 (n_1774, wc86, n_1643);
  not gc86 (wc86, n_1644);
  and g2339 (n_1824, wc87, n_1703);
  not gc87 (wc87, n_1704);
  and g2340 (n_1765, wc88, n_1762);
  not gc88 (wc88, n_1757);
  or g2341 (n_1871, wc89, n_1646);
  not gc89 (wc89, n_1770);
  and g2342 (n_1835, wc90, n_1832);
  not gc90 (wc90, n_1827);
  and g2343 (n_2002, wc91, n_1725);
  not gc91 (wc91, n_1838);
  and g2344 (n_1924, wc92, n_1844);
  not gc92 (wc92, n_1845);
  or g2345 (n_1937, wc93, n_1628);
  not gc93 (wc93, n_1935);
  or g2346 (n_1942, n_1939, wc94);
  not gc94 (wc94, n_1935);
  or g2347 (n_2149, wc95, n_1640);
  not gc95 (wc95, n_1635);
  or g2348 (n_2152, wc96, n_1636);
  not gc96 (wc96, n_1637);
  or g2349 (n_2157, wc97, n_1642);
  not gc97 (wc97, n_1643);
  or g2350 (n_2204, wc98, n_1706);
  not gc98 (wc98, n_1701);
  and g2351 (n_1864, wc99, n_1764);
  not gc99 (wc99, n_1765);
  and g2352 (n_1775, wc100, n_1772);
  not gc100 (wc100, n_1767);
  and g2353 (n_1917, wc101, n_1713);
  not gc101 (wc101, n_1828);
  and g2354 (n_1921, wc102, n_1834);
  not gc102 (wc102, n_1835);
  and g2355 (n_1948, wc103, n_1770);
  not gc103 (wc103, n_1867);
  and g2356 (n_1929, wc104, n_1850);
  not gc104 (wc104, n_1924);
  or g2357 (n_1944, wc105, n_1867);
  not gc105 (wc105, n_1935);
  and g2358 (n_1777, wc106, n_1649);
  not gc106 (wc106, n_1650);
  and g2359 (n_1872, wc107, n_1641);
  not gc107 (wc107, n_1768);
  and g2360 (n_1876, wc108, n_1774);
  not gc108 (wc108, n_1775);
  and g2361 (n_1869, wc109, n_1770);
  not gc109 (wc109, n_1864);
  and g2362 (n_2011, wc110, n_1731);
  not gc110 (wc110, n_1925);
  and g2363 (n_2016, wc111, n_1847);
  not gc111 (wc111, n_1929);
  and g2364 (n_2021, n_1932, wc112);
  not gc112 (wc112, n_1933);
  or g2365 (n_2158, wc113, n_1652);
  not gc113 (wc113, n_1647);
  or g2366 (n_2161, wc114, n_1648);
  not gc114 (wc114, n_1649);
  and g2367 (n_1946, wc115, n_1635);
  not gc115 (wc115, n_1865);
  and g2368 (n_1949, wc116, n_1767);
  not gc116 (wc116, n_1869);
  or g2369 (n_2169, wc117, n_1664);
  not gc117 (wc117, n_1659);
  and g2370 (n_1784, wc118, n_1655);
  not gc118 (wc118, n_1656);
  and g2371 (n_1787, wc119, n_1661);
  not gc119 (wc119, n_1662);
  and g2372 (n_1814, wc120, n_1691);
  not gc120 (wc120, n_1692);
  and g2373 (n_1817, wc121, n_1697);
  not gc121 (wc121, n_1698);
  and g2374 (n_2030, wc122, n_1653);
  not gc122 (wc122, n_1778);
  or g2375 (n_2028, wc123, n_1658);
  not gc123 (wc123, n_1780);
  or g2376 (n_2080, wc124, n_1706);
  not gc124 (wc124, n_1820);
  and g2377 (n_1952, n_1872, wc125);
  not gc125 (wc125, n_1873);
  and g2378 (n_1955, n_1876, wc126);
  not gc126 (wc126, n_1877);
  or g2379 (n_2163, wc127, n_1658);
  not gc127 (wc127, n_1653);
  or g2380 (n_2166, wc128, n_1654);
  not gc128 (wc128, n_1655);
  or g2381 (n_2172, wc129, n_1660);
  not gc129 (wc129, n_1661);
  or g2382 (n_2193, wc130, n_1684);
  not gc130 (wc130, n_1685);
  or g2383 (n_2195, wc131, n_1694);
  not gc131 (wc131, n_1689);
  or g2384 (n_2198, wc132, n_1690);
  not gc132 (wc132, n_1691);
  or g2385 (n_2199, wc133, n_1700);
  not gc133 (wc133, n_1695);
  or g2386 (n_2202, wc134, n_1696);
  not gc134 (wc134, n_1697);
  and g2387 (n_1785, wc135, n_1782);
  not gc135 (wc135, n_1777);
  or g2388 (n_1886, wc136, n_1670);
  not gc136 (wc136, n_1790);
  and g2389 (n_1825, wc137, n_1822);
  not gc137 (wc137, n_1817);
  and g2390 (n_2037, wc138, n_1790);
  not gc138 (wc138, n_1882);
  and g2391 (n_2089, wc139, n_1830);
  not gc139 (wc139, n_1912);
  or g2392 (n_2174, wc140, n_1670);
  not gc140 (wc140, n_1665);
  and g2393 (n_1794, wc141, n_1667);
  not gc141 (wc141, n_1668);
  and g2394 (n_1797, wc142, n_1673);
  not gc142 (wc142, n_1674);
  and g2395 (n_1804, wc143, n_1679);
  not gc143 (wc143, n_1680);
  and g2396 (n_1807, wc144, n_1685);
  not gc144 (wc144, n_1686);
  and g2397 (n_1879, wc145, n_1784);
  not gc145 (wc145, n_1785);
  and g2398 (n_1887, wc146, n_1665);
  not gc146 (wc146, n_1788);
  or g2399 (n_1965, wc147, n_1682);
  not gc147 (wc147, n_1800);
  or g2400 (n_1901, wc148, n_1694);
  not gc148 (wc148, n_1810);
  and g2401 (n_2082, wc149, n_1701);
  not gc149 (wc149, n_1818);
  and g2402 (n_1909, wc150, n_1824);
  not gc150 (wc150, n_1825);
  or g2403 (n_2096, wc151, n_1724);
  not gc151 (wc151, n_1996);
  or g2404 (n_2104, n_2001, wc152);
  not gc152 (wc152, n_1996);
  or g2405 (n_2108, wc153, n_1927);
  not gc153 (wc153, n_1996);
  or g2406 (n_2026, wc154, n_1652);
  not gc154 (wc154, n_2024);
  or g2407 (n_2031, n_2028, wc155);
  not gc155 (wc155, n_2024);
  or g2408 (n_2033, wc156, n_1882);
  not gc156 (wc156, n_2024);
  or g2409 (n_2177, wc157, n_1666);
  not gc157 (wc157, n_1667);
  or g2410 (n_2179, wc158, n_1676);
  not gc158 (wc158, n_1671);
  or g2411 (n_2182, wc159, n_1672);
  not gc159 (wc159, n_1673);
  or g2412 (n_2184, wc160, n_1682);
  not gc160 (wc160, n_1677);
  or g2413 (n_2187, wc161, n_1678);
  not gc161 (wc161, n_1679);
  or g2414 (n_2190, wc162, n_1688);
  not gc162 (wc162, n_1683);
  and g2415 (n_1795, wc163, n_1792);
  not gc163 (wc163, n_1787);
  and g2416 (n_1805, wc164, n_1802);
  not gc164 (wc164, n_1797);
  and g2417 (n_1815, wc165, n_1812);
  not gc165 (wc165, n_1807);
  and g2418 (n_1884, wc166, n_1790);
  not gc166 (wc166, n_1879);
  and g2419 (n_1978, wc167, n_1810);
  not gc167 (wc167, n_1897);
  and g2420 (n_1914, wc168, n_1830);
  not gc168 (wc168, n_1909);
  and g2421 (n_1891, wc169, n_1794);
  not gc169 (wc169, n_1795);
  and g2422 (n_1966, wc170, n_1677);
  not gc170 (wc170, n_1798);
  and g2423 (n_1894, wc171, n_1804);
  not gc171 (wc171, n_1805);
  and g2424 (n_1902, wc172, n_1689);
  not gc172 (wc172, n_1808);
  and g2425 (n_1906, wc173, n_1814);
  not gc173 (wc173, n_1815);
  and g2426 (n_2035, wc174, n_1659);
  not gc174 (wc174, n_1880);
  and g2427 (n_2038, wc175, n_1787);
  not gc175 (wc175, n_1884);
  and g2428 (n_2041, n_1887, wc176);
  not gc176 (wc176, n_1888);
  and g2429 (n_2087, wc177, n_1707);
  not gc177 (wc177, n_1910);
  and g2430 (n_2090, wc178, n_1827);
  not gc178 (wc178, n_1914);
  and g2431 (n_2093, n_1917, wc179);
  not gc179 (wc179, n_1918);
  and g2432 (n_1993, n_1921, wc180);
  not gc180 (wc180, n_1922);
  or g2433 (n_2044, wc181, n_1676);
  not gc181 (wc181, n_1960);
  or g2434 (n_2052, n_1965, wc182);
  not gc182 (wc182, n_1960);
  or g2435 (n_2056, wc183, n_1897);
  not gc183 (wc183, n_1960);
  and g2436 (n_1899, wc184, n_1810);
  not gc184 (wc184, n_1894);
  and g2437 (n_1999, wc185, n_1840);
  not gc185 (wc185, n_1993);
  and g2438 (n_2012, wc186, n_2009);
  not gc186 (wc186, n_1993);
  and g2439 (n_2017, wc187, n_2014);
  not gc187 (wc187, n_1993);
  and g2440 (n_2022, wc188, n_2019);
  not gc188 (wc188, n_1993);
  and g2441 (n_1957, n_1891, wc189);
  not gc189 (wc189, n_1892);
  and g2442 (n_1975, wc190, n_1683);
  not gc190 (wc190, n_1895);
  and g2443 (n_1980, wc191, n_1807);
  not gc191 (wc191, n_1899);
  and g2444 (n_1985, n_1902, wc192);
  not gc192 (wc192, n_1903);
  and g2445 (n_1990, n_1906, wc193);
  not gc193 (wc193, n_1907);
  and g2446 (n_2098, wc194, n_1719);
  not gc194 (wc194, n_1994);
  and g2447 (n_2102, wc195, n_1837);
  not gc195 (wc195, n_1999);
  and g2448 (n_2106, n_2002, wc196);
  not gc196 (wc196, n_2003);
  and g2449 (n_2110, n_1924, wc197);
  not gc197 (wc197, n_2006);
  and g2450 (n_2114, wc198, n_2011);
  not gc198 (wc198, n_2012);
  and g2451 (n_2118, wc199, n_2016);
  not gc199 (wc199, n_2017);
  and g2452 (n_2122, wc200, n_2021);
  not gc200 (wc200, n_2022);
  or g2453 (n_2047, n_2044, wc201);
  not gc201 (wc201, n_2024);
  or g2454 (n_2051, n_2048, wc202);
  not gc202 (wc202, n_2024);
  or g2455 (n_2055, n_2052, wc203);
  not gc203 (wc203, n_2024);
  or g2456 (n_2059, n_2056, wc204);
  not gc204 (wc204, n_2024);
  or g2457 (n_2063, n_2060, wc205);
  not gc205 (wc205, n_2024);
  or g2458 (n_2067, n_2064, wc206);
  not gc206 (wc206, n_2024);
  or g2459 (n_2071, n_2068, wc207);
  not gc207 (wc207, n_2024);
  or g2460 (n_2075, n_2072, wc208);
  not gc208 (wc208, n_2024);
  and g2461 (n_1963, wc209, n_1800);
  not gc209 (wc209, n_1957);
  and g2462 (n_1976, wc210, n_1973);
  not gc210 (wc210, n_1957);
  and g2463 (n_1981, wc211, n_1978);
  not gc211 (wc211, n_1957);
  and g2464 (n_1986, wc212, n_1983);
  not gc212 (wc212, n_1957);
  and g2465 (n_1991, wc213, n_1988);
  not gc213 (wc213, n_1957);
  and g2466 (n_2046, wc214, n_1671);
  not gc214 (wc214, n_1958);
  and g2467 (n_2050, wc215, n_1797);
  not gc215 (wc215, n_1963);
  and g2468 (n_2054, n_1966, wc216);
  not gc216 (wc216, n_1967);
  and g2469 (n_2058, n_1894, wc217);
  not gc217 (wc217, n_1970);
  and g2470 (n_2062, wc218, n_1975);
  not gc218 (wc218, n_1976);
  and g2471 (n_2066, wc219, n_1980);
  not gc219 (wc219, n_1981);
  and g2472 (n_2070, wc220, n_1985);
  not gc220 (wc220, n_1986);
  and g2473 (n_2074, wc221, n_1990);
  not gc221 (wc221, n_1991);
  or g2474 (n_2078, wc222, n_1700);
  not gc222 (wc222, n_2076);
  or g2475 (n_2083, n_2080, wc223);
  not gc223 (wc223, n_2076);
  or g2476 (n_2085, wc224, n_1912);
  not gc224 (wc224, n_2076);
  or g2477 (n_2099, n_2096, wc225);
  not gc225 (wc225, n_2076);
  or g2478 (n_2103, wc226, n_2100);
  not gc226 (wc226, n_2076);
  or g2479 (n_2107, n_2104, wc227);
  not gc227 (wc227, n_2076);
  or g2480 (n_2111, n_2108, wc228);
  not gc228 (wc228, n_2076);
  or g2481 (n_2115, wc229, n_2112);
  not gc229 (wc229, n_2076);
  or g2482 (n_2119, wc230, n_2116);
  not gc230 (wc230, n_2076);
  or g2483 (n_2123, wc231, n_2120);
  not gc231 (wc231, n_2076);
endmodule

module mult_signed_const_6020_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_6020_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

