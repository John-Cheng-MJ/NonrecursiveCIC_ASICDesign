module add_signed_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [23:0] A, B;
  output [21:0] Z;
  wire [23:0] A, B;
  wire [21:0] Z;
  wire n_73, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123;
  wire n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131;
  wire n_132, n_133, n_134, n_135, n_136, n_137, n_138, n_139;
  wire n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147;
  wire n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155;
  wire n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163;
  wire n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171;
  wire n_172, n_173, n_174, n_175, n_176, n_180;
  nand g4 (n_73, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_77, A[1], B[1]);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_117, A[9], B[9]);
  nand g59 (n_118, A[9], n_116);
  nand g60 (n_119, B[9], n_116);
  nand g61 (n_121, n_117, n_118, n_119);
  xor g62 (n_120, A[9], B[9]);
  xor g63 (Z[9], n_116, n_120);
  nand g64 (n_122, A[10], B[10]);
  nand g65 (n_123, A[10], n_121);
  nand g66 (n_124, B[10], n_121);
  nand g67 (n_126, n_122, n_123, n_124);
  xor g68 (n_125, A[10], B[10]);
  xor g69 (Z[10], n_121, n_125);
  nand g70 (n_127, A[11], B[11]);
  nand g71 (n_128, A[11], n_126);
  nand g72 (n_129, B[11], n_126);
  nand g73 (n_131, n_127, n_128, n_129);
  xor g74 (n_130, A[11], B[11]);
  xor g75 (Z[11], n_126, n_130);
  nand g76 (n_132, A[12], B[12]);
  nand g77 (n_133, A[12], n_131);
  nand g78 (n_134, B[12], n_131);
  nand g79 (n_136, n_132, n_133, n_134);
  xor g80 (n_135, A[12], B[12]);
  xor g81 (Z[12], n_131, n_135);
  nand g82 (n_137, A[13], B[13]);
  nand g83 (n_138, A[13], n_136);
  nand g84 (n_139, B[13], n_136);
  nand g85 (n_141, n_137, n_138, n_139);
  xor g86 (n_140, A[13], B[13]);
  xor g87 (Z[13], n_136, n_140);
  nand g88 (n_142, A[14], B[14]);
  nand g89 (n_143, A[14], n_141);
  nand g90 (n_144, B[14], n_141);
  nand g91 (n_146, n_142, n_143, n_144);
  xor g92 (n_145, A[14], B[14]);
  xor g93 (Z[14], n_141, n_145);
  nand g94 (n_147, A[15], B[15]);
  nand g95 (n_148, A[15], n_146);
  nand g96 (n_149, B[15], n_146);
  nand g97 (n_151, n_147, n_148, n_149);
  xor g98 (n_150, A[15], B[15]);
  xor g99 (Z[15], n_146, n_150);
  nand g100 (n_152, A[16], B[16]);
  nand g101 (n_153, A[16], n_151);
  nand g102 (n_154, B[16], n_151);
  nand g103 (n_156, n_152, n_153, n_154);
  xor g104 (n_155, A[16], B[16]);
  xor g105 (Z[16], n_151, n_155);
  nand g106 (n_157, A[17], B[17]);
  nand g107 (n_158, A[17], n_156);
  nand g108 (n_159, B[17], n_156);
  nand g109 (n_161, n_157, n_158, n_159);
  xor g110 (n_160, A[17], B[17]);
  xor g111 (Z[17], n_156, n_160);
  nand g112 (n_162, A[18], B[18]);
  nand g113 (n_163, A[18], n_161);
  nand g114 (n_164, B[18], n_161);
  nand g115 (n_166, n_162, n_163, n_164);
  xor g116 (n_165, A[18], B[18]);
  xor g117 (Z[18], n_161, n_165);
  nand g118 (n_167, A[19], B[19]);
  nand g119 (n_168, A[19], n_166);
  nand g120 (n_169, B[19], n_166);
  nand g121 (n_171, n_167, n_168, n_169);
  xor g122 (n_170, A[19], B[19]);
  xor g123 (Z[19], n_166, n_170);
  nand g124 (n_172, A[20], B[20]);
  nand g125 (n_173, A[20], n_171);
  nand g126 (n_174, B[20], n_171);
  nand g127 (n_176, n_172, n_173, n_174);
  xor g128 (n_175, A[20], B[20]);
  xor g129 (Z[20], n_171, n_175);
  xor g135 (Z[21], n_176, n_180);
  xor g137 (n_180, A[21], B[21]);
  or g138 (n_78, wc, n_73);
  not gc (wc, A[1]);
  or g139 (n_79, wc0, n_73);
  not gc0 (wc0, B[1]);
  xnor g140 (Z[1], n_73, n_80);
endmodule

module add_signed_GENERIC(A, B, Z);
  input [23:0] A, B;
  output [21:0] Z;
  wire [23:0] A, B;
  wire [21:0] Z;
  add_signed_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3151_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  wire n_76, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_188;
  nand g4 (n_76, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_120, A[9], B[9]);
  nand g59 (n_121, A[9], n_119);
  nand g60 (n_122, B[9], n_119);
  nand g61 (n_124, n_120, n_121, n_122);
  xor g62 (n_123, A[9], B[9]);
  xor g63 (Z[9], n_119, n_123);
  nand g64 (n_125, A[10], B[10]);
  nand g65 (n_126, A[10], n_124);
  nand g66 (n_127, B[10], n_124);
  nand g67 (n_129, n_125, n_126, n_127);
  xor g68 (n_128, A[10], B[10]);
  xor g69 (Z[10], n_124, n_128);
  nand g70 (n_130, A[11], B[11]);
  nand g71 (n_131, A[11], n_129);
  nand g72 (n_132, B[11], n_129);
  nand g73 (n_134, n_130, n_131, n_132);
  xor g74 (n_133, A[11], B[11]);
  xor g75 (Z[11], n_129, n_133);
  nand g76 (n_135, A[12], B[12]);
  nand g77 (n_136, A[12], n_134);
  nand g78 (n_137, B[12], n_134);
  nand g79 (n_139, n_135, n_136, n_137);
  xor g80 (n_138, A[12], B[12]);
  xor g81 (Z[12], n_134, n_138);
  nand g82 (n_140, A[13], B[13]);
  nand g83 (n_141, A[13], n_139);
  nand g84 (n_142, B[13], n_139);
  nand g85 (n_144, n_140, n_141, n_142);
  xor g86 (n_143, A[13], B[13]);
  xor g87 (Z[13], n_139, n_143);
  nand g88 (n_145, A[14], B[14]);
  nand g89 (n_146, A[14], n_144);
  nand g90 (n_147, B[14], n_144);
  nand g91 (n_149, n_145, n_146, n_147);
  xor g92 (n_148, A[14], B[14]);
  xor g93 (Z[14], n_144, n_148);
  nand g94 (n_150, A[15], B[15]);
  nand g95 (n_151, A[15], n_149);
  nand g96 (n_152, B[15], n_149);
  nand g97 (n_154, n_150, n_151, n_152);
  xor g98 (n_153, A[15], B[15]);
  xor g99 (Z[15], n_149, n_153);
  nand g100 (n_155, A[16], B[16]);
  nand g101 (n_156, A[16], n_154);
  nand g102 (n_157, B[16], n_154);
  nand g103 (n_159, n_155, n_156, n_157);
  xor g104 (n_158, A[16], B[16]);
  xor g105 (Z[16], n_154, n_158);
  nand g106 (n_160, A[17], B[17]);
  nand g107 (n_161, A[17], n_159);
  nand g108 (n_162, B[17], n_159);
  nand g109 (n_164, n_160, n_161, n_162);
  xor g110 (n_163, A[17], B[17]);
  xor g111 (Z[17], n_159, n_163);
  nand g112 (n_165, A[18], B[18]);
  nand g113 (n_166, A[18], n_164);
  nand g114 (n_167, B[18], n_164);
  nand g115 (n_169, n_165, n_166, n_167);
  xor g116 (n_168, A[18], B[18]);
  xor g117 (Z[18], n_164, n_168);
  nand g118 (n_170, A[19], B[19]);
  nand g119 (n_171, A[19], n_169);
  nand g120 (n_172, B[19], n_169);
  nand g121 (n_174, n_170, n_171, n_172);
  xor g122 (n_173, A[19], B[19]);
  xor g123 (Z[19], n_169, n_173);
  nand g124 (n_175, A[20], B[20]);
  nand g125 (n_176, A[20], n_174);
  nand g126 (n_177, B[20], n_174);
  nand g127 (n_179, n_175, n_176, n_177);
  xor g128 (n_178, A[20], B[20]);
  xor g129 (Z[20], n_174, n_178);
  nand g130 (n_180, A[21], B[21]);
  nand g131 (n_181, A[21], n_179);
  nand g132 (n_182, B[21], n_179);
  nand g133 (n_184, n_180, n_181, n_182);
  xor g134 (n_183, A[21], B[21]);
  xor g135 (Z[21], n_179, n_183);
  xor g141 (Z[22], n_184, n_188);
  xor g143 (n_188, A[22], B[22]);
  or g144 (n_81, wc, n_76);
  not gc (wc, A[1]);
  or g145 (n_82, wc0, n_76);
  not gc0 (wc0, B[1]);
  xnor g146 (Z[1], n_76, n_83);
endmodule

module add_signed_3151_GENERIC(A, B, Z);
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  add_signed_3151_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3151_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  wire n_76, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_188;
  nand g4 (n_76, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_120, A[9], B[9]);
  nand g59 (n_121, A[9], n_119);
  nand g60 (n_122, B[9], n_119);
  nand g61 (n_124, n_120, n_121, n_122);
  xor g62 (n_123, A[9], B[9]);
  xor g63 (Z[9], n_119, n_123);
  nand g64 (n_125, A[10], B[10]);
  nand g65 (n_126, A[10], n_124);
  nand g66 (n_127, B[10], n_124);
  nand g67 (n_129, n_125, n_126, n_127);
  xor g68 (n_128, A[10], B[10]);
  xor g69 (Z[10], n_124, n_128);
  nand g70 (n_130, A[11], B[11]);
  nand g71 (n_131, A[11], n_129);
  nand g72 (n_132, B[11], n_129);
  nand g73 (n_134, n_130, n_131, n_132);
  xor g74 (n_133, A[11], B[11]);
  xor g75 (Z[11], n_129, n_133);
  nand g76 (n_135, A[12], B[12]);
  nand g77 (n_136, A[12], n_134);
  nand g78 (n_137, B[12], n_134);
  nand g79 (n_139, n_135, n_136, n_137);
  xor g80 (n_138, A[12], B[12]);
  xor g81 (Z[12], n_134, n_138);
  nand g82 (n_140, A[13], B[13]);
  nand g83 (n_141, A[13], n_139);
  nand g84 (n_142, B[13], n_139);
  nand g85 (n_144, n_140, n_141, n_142);
  xor g86 (n_143, A[13], B[13]);
  xor g87 (Z[13], n_139, n_143);
  nand g88 (n_145, A[14], B[14]);
  nand g89 (n_146, A[14], n_144);
  nand g90 (n_147, B[14], n_144);
  nand g91 (n_149, n_145, n_146, n_147);
  xor g92 (n_148, A[14], B[14]);
  xor g93 (Z[14], n_144, n_148);
  nand g94 (n_150, A[15], B[15]);
  nand g95 (n_151, A[15], n_149);
  nand g96 (n_152, B[15], n_149);
  nand g97 (n_154, n_150, n_151, n_152);
  xor g98 (n_153, A[15], B[15]);
  xor g99 (Z[15], n_149, n_153);
  nand g100 (n_155, A[16], B[16]);
  nand g101 (n_156, A[16], n_154);
  nand g102 (n_157, B[16], n_154);
  nand g103 (n_159, n_155, n_156, n_157);
  xor g104 (n_158, A[16], B[16]);
  xor g105 (Z[16], n_154, n_158);
  nand g106 (n_160, A[17], B[17]);
  nand g107 (n_161, A[17], n_159);
  nand g108 (n_162, B[17], n_159);
  nand g109 (n_164, n_160, n_161, n_162);
  xor g110 (n_163, A[17], B[17]);
  xor g111 (Z[17], n_159, n_163);
  nand g112 (n_165, A[18], B[18]);
  nand g113 (n_166, A[18], n_164);
  nand g114 (n_167, B[18], n_164);
  nand g115 (n_169, n_165, n_166, n_167);
  xor g116 (n_168, A[18], B[18]);
  xor g117 (Z[18], n_164, n_168);
  nand g118 (n_170, A[19], B[19]);
  nand g119 (n_171, A[19], n_169);
  nand g120 (n_172, B[19], n_169);
  nand g121 (n_174, n_170, n_171, n_172);
  xor g122 (n_173, A[19], B[19]);
  xor g123 (Z[19], n_169, n_173);
  nand g124 (n_175, A[20], B[20]);
  nand g125 (n_176, A[20], n_174);
  nand g126 (n_177, B[20], n_174);
  nand g127 (n_179, n_175, n_176, n_177);
  xor g128 (n_178, A[20], B[20]);
  xor g129 (Z[20], n_174, n_178);
  nand g130 (n_180, A[21], B[21]);
  nand g131 (n_181, A[21], n_179);
  nand g132 (n_182, B[21], n_179);
  nand g133 (n_184, n_180, n_181, n_182);
  xor g134 (n_183, A[21], B[21]);
  xor g135 (Z[21], n_179, n_183);
  xor g141 (Z[22], n_184, n_188);
  xor g143 (n_188, A[22], B[22]);
  or g144 (n_81, wc, n_76);
  not gc (wc, A[1]);
  or g145 (n_82, wc0, n_76);
  not gc0 (wc0, B[1]);
  xnor g146 (Z[1], n_76, n_83);
endmodule

module add_signed_3151_1_GENERIC(A, B, Z);
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  add_signed_3151_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3151_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  wire n_76, n_80, n_81, n_82, n_83, n_84, n_85, n_86;
  wire n_87, n_88, n_89, n_90, n_91, n_92, n_93, n_94;
  wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174;
  wire n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182;
  wire n_183, n_184, n_188;
  nand g4 (n_76, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_80, A[1], B[1]);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_120, A[9], B[9]);
  nand g59 (n_121, A[9], n_119);
  nand g60 (n_122, B[9], n_119);
  nand g61 (n_124, n_120, n_121, n_122);
  xor g62 (n_123, A[9], B[9]);
  xor g63 (Z[9], n_119, n_123);
  nand g64 (n_125, A[10], B[10]);
  nand g65 (n_126, A[10], n_124);
  nand g66 (n_127, B[10], n_124);
  nand g67 (n_129, n_125, n_126, n_127);
  xor g68 (n_128, A[10], B[10]);
  xor g69 (Z[10], n_124, n_128);
  nand g70 (n_130, A[11], B[11]);
  nand g71 (n_131, A[11], n_129);
  nand g72 (n_132, B[11], n_129);
  nand g73 (n_134, n_130, n_131, n_132);
  xor g74 (n_133, A[11], B[11]);
  xor g75 (Z[11], n_129, n_133);
  nand g76 (n_135, A[12], B[12]);
  nand g77 (n_136, A[12], n_134);
  nand g78 (n_137, B[12], n_134);
  nand g79 (n_139, n_135, n_136, n_137);
  xor g80 (n_138, A[12], B[12]);
  xor g81 (Z[12], n_134, n_138);
  nand g82 (n_140, A[13], B[13]);
  nand g83 (n_141, A[13], n_139);
  nand g84 (n_142, B[13], n_139);
  nand g85 (n_144, n_140, n_141, n_142);
  xor g86 (n_143, A[13], B[13]);
  xor g87 (Z[13], n_139, n_143);
  nand g88 (n_145, A[14], B[14]);
  nand g89 (n_146, A[14], n_144);
  nand g90 (n_147, B[14], n_144);
  nand g91 (n_149, n_145, n_146, n_147);
  xor g92 (n_148, A[14], B[14]);
  xor g93 (Z[14], n_144, n_148);
  nand g94 (n_150, A[15], B[15]);
  nand g95 (n_151, A[15], n_149);
  nand g96 (n_152, B[15], n_149);
  nand g97 (n_154, n_150, n_151, n_152);
  xor g98 (n_153, A[15], B[15]);
  xor g99 (Z[15], n_149, n_153);
  nand g100 (n_155, A[16], B[16]);
  nand g101 (n_156, A[16], n_154);
  nand g102 (n_157, B[16], n_154);
  nand g103 (n_159, n_155, n_156, n_157);
  xor g104 (n_158, A[16], B[16]);
  xor g105 (Z[16], n_154, n_158);
  nand g106 (n_160, A[17], B[17]);
  nand g107 (n_161, A[17], n_159);
  nand g108 (n_162, B[17], n_159);
  nand g109 (n_164, n_160, n_161, n_162);
  xor g110 (n_163, A[17], B[17]);
  xor g111 (Z[17], n_159, n_163);
  nand g112 (n_165, A[18], B[18]);
  nand g113 (n_166, A[18], n_164);
  nand g114 (n_167, B[18], n_164);
  nand g115 (n_169, n_165, n_166, n_167);
  xor g116 (n_168, A[18], B[18]);
  xor g117 (Z[18], n_164, n_168);
  nand g118 (n_170, A[19], B[19]);
  nand g119 (n_171, A[19], n_169);
  nand g120 (n_172, B[19], n_169);
  nand g121 (n_174, n_170, n_171, n_172);
  xor g122 (n_173, A[19], B[19]);
  xor g123 (Z[19], n_169, n_173);
  nand g124 (n_175, A[20], B[20]);
  nand g125 (n_176, A[20], n_174);
  nand g126 (n_177, B[20], n_174);
  nand g127 (n_179, n_175, n_176, n_177);
  xor g128 (n_178, A[20], B[20]);
  xor g129 (Z[20], n_174, n_178);
  nand g130 (n_180, A[21], B[21]);
  nand g131 (n_181, A[21], n_179);
  nand g132 (n_182, B[21], n_179);
  nand g133 (n_184, n_180, n_181, n_182);
  xor g134 (n_183, A[21], B[21]);
  xor g135 (Z[21], n_179, n_183);
  xor g141 (Z[22], n_184, n_188);
  xor g143 (n_188, A[22], B[22]);
  or g144 (n_81, wc, n_76);
  not gc (wc, A[1]);
  or g145 (n_82, wc0, n_76);
  not gc0 (wc0, B[1]);
  xnor g146 (Z[1], n_76, n_83);
endmodule

module add_signed_3151_2_GENERIC(A, B, Z);
  input [24:0] A, B;
  output [22:0] Z;
  wire [24:0] A, B;
  wire [22:0] Z;
  add_signed_3151_2_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3180_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  wire n_79, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_196;
  nand g4 (n_79, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_83, A[1], B[1]);
  nand g13 (n_87, n_83, n_84, n_85);
  xor g14 (n_86, A[1], B[1]);
  nand g16 (n_88, A[2], B[2]);
  nand g17 (n_89, A[2], n_87);
  nand g18 (n_90, B[2], n_87);
  nand g19 (n_92, n_88, n_89, n_90);
  xor g20 (n_91, A[2], B[2]);
  xor g21 (Z[2], n_87, n_91);
  nand g22 (n_93, A[3], B[3]);
  nand g23 (n_94, A[3], n_92);
  nand g24 (n_95, B[3], n_92);
  nand g25 (n_97, n_93, n_94, n_95);
  xor g26 (n_96, A[3], B[3]);
  xor g27 (Z[3], n_92, n_96);
  nand g28 (n_98, A[4], B[4]);
  nand g29 (n_99, A[4], n_97);
  nand g30 (n_100, B[4], n_97);
  nand g31 (n_102, n_98, n_99, n_100);
  xor g32 (n_101, A[4], B[4]);
  xor g33 (Z[4], n_97, n_101);
  nand g34 (n_103, A[5], B[5]);
  nand g35 (n_104, A[5], n_102);
  nand g36 (n_105, B[5], n_102);
  nand g37 (n_107, n_103, n_104, n_105);
  xor g38 (n_106, A[5], B[5]);
  xor g39 (Z[5], n_102, n_106);
  nand g40 (n_108, A[6], B[6]);
  nand g41 (n_109, A[6], n_107);
  nand g42 (n_110, B[6], n_107);
  nand g43 (n_112, n_108, n_109, n_110);
  xor g44 (n_111, A[6], B[6]);
  xor g45 (Z[6], n_107, n_111);
  nand g46 (n_113, A[7], B[7]);
  nand g47 (n_114, A[7], n_112);
  nand g48 (n_115, B[7], n_112);
  nand g49 (n_117, n_113, n_114, n_115);
  xor g50 (n_116, A[7], B[7]);
  xor g51 (Z[7], n_112, n_116);
  nand g52 (n_118, A[8], B[8]);
  nand g53 (n_119, A[8], n_117);
  nand g54 (n_120, B[8], n_117);
  nand g55 (n_122, n_118, n_119, n_120);
  xor g56 (n_121, A[8], B[8]);
  xor g57 (Z[8], n_117, n_121);
  nand g58 (n_123, A[9], B[9]);
  nand g59 (n_124, A[9], n_122);
  nand g60 (n_125, B[9], n_122);
  nand g61 (n_127, n_123, n_124, n_125);
  xor g62 (n_126, A[9], B[9]);
  xor g63 (Z[9], n_122, n_126);
  nand g64 (n_128, A[10], B[10]);
  nand g65 (n_129, A[10], n_127);
  nand g66 (n_130, B[10], n_127);
  nand g67 (n_132, n_128, n_129, n_130);
  xor g68 (n_131, A[10], B[10]);
  xor g69 (Z[10], n_127, n_131);
  nand g70 (n_133, A[11], B[11]);
  nand g71 (n_134, A[11], n_132);
  nand g72 (n_135, B[11], n_132);
  nand g73 (n_137, n_133, n_134, n_135);
  xor g74 (n_136, A[11], B[11]);
  xor g75 (Z[11], n_132, n_136);
  nand g76 (n_138, A[12], B[12]);
  nand g77 (n_139, A[12], n_137);
  nand g78 (n_140, B[12], n_137);
  nand g79 (n_142, n_138, n_139, n_140);
  xor g80 (n_141, A[12], B[12]);
  xor g81 (Z[12], n_137, n_141);
  nand g82 (n_143, A[13], B[13]);
  nand g83 (n_144, A[13], n_142);
  nand g84 (n_145, B[13], n_142);
  nand g85 (n_147, n_143, n_144, n_145);
  xor g86 (n_146, A[13], B[13]);
  xor g87 (Z[13], n_142, n_146);
  nand g88 (n_148, A[14], B[14]);
  nand g89 (n_149, A[14], n_147);
  nand g90 (n_150, B[14], n_147);
  nand g91 (n_152, n_148, n_149, n_150);
  xor g92 (n_151, A[14], B[14]);
  xor g93 (Z[14], n_147, n_151);
  nand g94 (n_153, A[15], B[15]);
  nand g95 (n_154, A[15], n_152);
  nand g96 (n_155, B[15], n_152);
  nand g97 (n_157, n_153, n_154, n_155);
  xor g98 (n_156, A[15], B[15]);
  xor g99 (Z[15], n_152, n_156);
  nand g100 (n_158, A[16], B[16]);
  nand g101 (n_159, A[16], n_157);
  nand g102 (n_160, B[16], n_157);
  nand g103 (n_162, n_158, n_159, n_160);
  xor g104 (n_161, A[16], B[16]);
  xor g105 (Z[16], n_157, n_161);
  nand g106 (n_163, A[17], B[17]);
  nand g107 (n_164, A[17], n_162);
  nand g108 (n_165, B[17], n_162);
  nand g109 (n_167, n_163, n_164, n_165);
  xor g110 (n_166, A[17], B[17]);
  xor g111 (Z[17], n_162, n_166);
  nand g112 (n_168, A[18], B[18]);
  nand g113 (n_169, A[18], n_167);
  nand g114 (n_170, B[18], n_167);
  nand g115 (n_172, n_168, n_169, n_170);
  xor g116 (n_171, A[18], B[18]);
  xor g117 (Z[18], n_167, n_171);
  nand g118 (n_173, A[19], B[19]);
  nand g119 (n_174, A[19], n_172);
  nand g120 (n_175, B[19], n_172);
  nand g121 (n_177, n_173, n_174, n_175);
  xor g122 (n_176, A[19], B[19]);
  xor g123 (Z[19], n_172, n_176);
  nand g124 (n_178, A[20], B[20]);
  nand g125 (n_179, A[20], n_177);
  nand g126 (n_180, B[20], n_177);
  nand g127 (n_182, n_178, n_179, n_180);
  xor g128 (n_181, A[20], B[20]);
  xor g129 (Z[20], n_177, n_181);
  nand g130 (n_183, A[21], B[21]);
  nand g131 (n_184, A[21], n_182);
  nand g132 (n_185, B[21], n_182);
  nand g133 (n_187, n_183, n_184, n_185);
  xor g134 (n_186, A[21], B[21]);
  xor g135 (Z[21], n_182, n_186);
  nand g136 (n_188, A[22], B[22]);
  nand g137 (n_189, A[22], n_187);
  nand g138 (n_190, B[22], n_187);
  nand g139 (n_192, n_188, n_189, n_190);
  xor g140 (n_191, A[22], B[22]);
  xor g141 (Z[22], n_187, n_191);
  xor g147 (Z[23], n_192, n_196);
  xor g149 (n_196, A[23], B[23]);
  or g150 (n_84, wc, n_79);
  not gc (wc, A[1]);
  or g151 (n_85, wc0, n_79);
  not gc0 (wc0, B[1]);
  xnor g152 (Z[1], n_79, n_86);
endmodule

module add_signed_3180_GENERIC(A, B, Z);
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  add_signed_3180_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3180_1_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  wire n_79, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_196;
  nand g4 (n_79, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_83, A[1], B[1]);
  nand g13 (n_87, n_83, n_84, n_85);
  xor g14 (n_86, A[1], B[1]);
  nand g16 (n_88, A[2], B[2]);
  nand g17 (n_89, A[2], n_87);
  nand g18 (n_90, B[2], n_87);
  nand g19 (n_92, n_88, n_89, n_90);
  xor g20 (n_91, A[2], B[2]);
  xor g21 (Z[2], n_87, n_91);
  nand g22 (n_93, A[3], B[3]);
  nand g23 (n_94, A[3], n_92);
  nand g24 (n_95, B[3], n_92);
  nand g25 (n_97, n_93, n_94, n_95);
  xor g26 (n_96, A[3], B[3]);
  xor g27 (Z[3], n_92, n_96);
  nand g28 (n_98, A[4], B[4]);
  nand g29 (n_99, A[4], n_97);
  nand g30 (n_100, B[4], n_97);
  nand g31 (n_102, n_98, n_99, n_100);
  xor g32 (n_101, A[4], B[4]);
  xor g33 (Z[4], n_97, n_101);
  nand g34 (n_103, A[5], B[5]);
  nand g35 (n_104, A[5], n_102);
  nand g36 (n_105, B[5], n_102);
  nand g37 (n_107, n_103, n_104, n_105);
  xor g38 (n_106, A[5], B[5]);
  xor g39 (Z[5], n_102, n_106);
  nand g40 (n_108, A[6], B[6]);
  nand g41 (n_109, A[6], n_107);
  nand g42 (n_110, B[6], n_107);
  nand g43 (n_112, n_108, n_109, n_110);
  xor g44 (n_111, A[6], B[6]);
  xor g45 (Z[6], n_107, n_111);
  nand g46 (n_113, A[7], B[7]);
  nand g47 (n_114, A[7], n_112);
  nand g48 (n_115, B[7], n_112);
  nand g49 (n_117, n_113, n_114, n_115);
  xor g50 (n_116, A[7], B[7]);
  xor g51 (Z[7], n_112, n_116);
  nand g52 (n_118, A[8], B[8]);
  nand g53 (n_119, A[8], n_117);
  nand g54 (n_120, B[8], n_117);
  nand g55 (n_122, n_118, n_119, n_120);
  xor g56 (n_121, A[8], B[8]);
  xor g57 (Z[8], n_117, n_121);
  nand g58 (n_123, A[9], B[9]);
  nand g59 (n_124, A[9], n_122);
  nand g60 (n_125, B[9], n_122);
  nand g61 (n_127, n_123, n_124, n_125);
  xor g62 (n_126, A[9], B[9]);
  xor g63 (Z[9], n_122, n_126);
  nand g64 (n_128, A[10], B[10]);
  nand g65 (n_129, A[10], n_127);
  nand g66 (n_130, B[10], n_127);
  nand g67 (n_132, n_128, n_129, n_130);
  xor g68 (n_131, A[10], B[10]);
  xor g69 (Z[10], n_127, n_131);
  nand g70 (n_133, A[11], B[11]);
  nand g71 (n_134, A[11], n_132);
  nand g72 (n_135, B[11], n_132);
  nand g73 (n_137, n_133, n_134, n_135);
  xor g74 (n_136, A[11], B[11]);
  xor g75 (Z[11], n_132, n_136);
  nand g76 (n_138, A[12], B[12]);
  nand g77 (n_139, A[12], n_137);
  nand g78 (n_140, B[12], n_137);
  nand g79 (n_142, n_138, n_139, n_140);
  xor g80 (n_141, A[12], B[12]);
  xor g81 (Z[12], n_137, n_141);
  nand g82 (n_143, A[13], B[13]);
  nand g83 (n_144, A[13], n_142);
  nand g84 (n_145, B[13], n_142);
  nand g85 (n_147, n_143, n_144, n_145);
  xor g86 (n_146, A[13], B[13]);
  xor g87 (Z[13], n_142, n_146);
  nand g88 (n_148, A[14], B[14]);
  nand g89 (n_149, A[14], n_147);
  nand g90 (n_150, B[14], n_147);
  nand g91 (n_152, n_148, n_149, n_150);
  xor g92 (n_151, A[14], B[14]);
  xor g93 (Z[14], n_147, n_151);
  nand g94 (n_153, A[15], B[15]);
  nand g95 (n_154, A[15], n_152);
  nand g96 (n_155, B[15], n_152);
  nand g97 (n_157, n_153, n_154, n_155);
  xor g98 (n_156, A[15], B[15]);
  xor g99 (Z[15], n_152, n_156);
  nand g100 (n_158, A[16], B[16]);
  nand g101 (n_159, A[16], n_157);
  nand g102 (n_160, B[16], n_157);
  nand g103 (n_162, n_158, n_159, n_160);
  xor g104 (n_161, A[16], B[16]);
  xor g105 (Z[16], n_157, n_161);
  nand g106 (n_163, A[17], B[17]);
  nand g107 (n_164, A[17], n_162);
  nand g108 (n_165, B[17], n_162);
  nand g109 (n_167, n_163, n_164, n_165);
  xor g110 (n_166, A[17], B[17]);
  xor g111 (Z[17], n_162, n_166);
  nand g112 (n_168, A[18], B[18]);
  nand g113 (n_169, A[18], n_167);
  nand g114 (n_170, B[18], n_167);
  nand g115 (n_172, n_168, n_169, n_170);
  xor g116 (n_171, A[18], B[18]);
  xor g117 (Z[18], n_167, n_171);
  nand g118 (n_173, A[19], B[19]);
  nand g119 (n_174, A[19], n_172);
  nand g120 (n_175, B[19], n_172);
  nand g121 (n_177, n_173, n_174, n_175);
  xor g122 (n_176, A[19], B[19]);
  xor g123 (Z[19], n_172, n_176);
  nand g124 (n_178, A[20], B[20]);
  nand g125 (n_179, A[20], n_177);
  nand g126 (n_180, B[20], n_177);
  nand g127 (n_182, n_178, n_179, n_180);
  xor g128 (n_181, A[20], B[20]);
  xor g129 (Z[20], n_177, n_181);
  nand g130 (n_183, A[21], B[21]);
  nand g131 (n_184, A[21], n_182);
  nand g132 (n_185, B[21], n_182);
  nand g133 (n_187, n_183, n_184, n_185);
  xor g134 (n_186, A[21], B[21]);
  xor g135 (Z[21], n_182, n_186);
  nand g136 (n_188, A[22], B[22]);
  nand g137 (n_189, A[22], n_187);
  nand g138 (n_190, B[22], n_187);
  nand g139 (n_192, n_188, n_189, n_190);
  xor g140 (n_191, A[22], B[22]);
  xor g141 (Z[22], n_187, n_191);
  xor g147 (Z[23], n_192, n_196);
  xor g149 (n_196, A[23], B[23]);
  or g150 (n_84, wc, n_79);
  not gc (wc, A[1]);
  or g151 (n_85, wc0, n_79);
  not gc0 (wc0, B[1]);
  xnor g152 (Z[1], n_79, n_86);
endmodule

module add_signed_3180_1_GENERIC(A, B, Z);
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  add_signed_3180_1_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3180_2_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  wire n_79, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_196;
  nand g4 (n_79, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_83, A[1], B[1]);
  nand g13 (n_87, n_83, n_84, n_85);
  xor g14 (n_86, A[1], B[1]);
  nand g16 (n_88, A[2], B[2]);
  nand g17 (n_89, A[2], n_87);
  nand g18 (n_90, B[2], n_87);
  nand g19 (n_92, n_88, n_89, n_90);
  xor g20 (n_91, A[2], B[2]);
  xor g21 (Z[2], n_87, n_91);
  nand g22 (n_93, A[3], B[3]);
  nand g23 (n_94, A[3], n_92);
  nand g24 (n_95, B[3], n_92);
  nand g25 (n_97, n_93, n_94, n_95);
  xor g26 (n_96, A[3], B[3]);
  xor g27 (Z[3], n_92, n_96);
  nand g28 (n_98, A[4], B[4]);
  nand g29 (n_99, A[4], n_97);
  nand g30 (n_100, B[4], n_97);
  nand g31 (n_102, n_98, n_99, n_100);
  xor g32 (n_101, A[4], B[4]);
  xor g33 (Z[4], n_97, n_101);
  nand g34 (n_103, A[5], B[5]);
  nand g35 (n_104, A[5], n_102);
  nand g36 (n_105, B[5], n_102);
  nand g37 (n_107, n_103, n_104, n_105);
  xor g38 (n_106, A[5], B[5]);
  xor g39 (Z[5], n_102, n_106);
  nand g40 (n_108, A[6], B[6]);
  nand g41 (n_109, A[6], n_107);
  nand g42 (n_110, B[6], n_107);
  nand g43 (n_112, n_108, n_109, n_110);
  xor g44 (n_111, A[6], B[6]);
  xor g45 (Z[6], n_107, n_111);
  nand g46 (n_113, A[7], B[7]);
  nand g47 (n_114, A[7], n_112);
  nand g48 (n_115, B[7], n_112);
  nand g49 (n_117, n_113, n_114, n_115);
  xor g50 (n_116, A[7], B[7]);
  xor g51 (Z[7], n_112, n_116);
  nand g52 (n_118, A[8], B[8]);
  nand g53 (n_119, A[8], n_117);
  nand g54 (n_120, B[8], n_117);
  nand g55 (n_122, n_118, n_119, n_120);
  xor g56 (n_121, A[8], B[8]);
  xor g57 (Z[8], n_117, n_121);
  nand g58 (n_123, A[9], B[9]);
  nand g59 (n_124, A[9], n_122);
  nand g60 (n_125, B[9], n_122);
  nand g61 (n_127, n_123, n_124, n_125);
  xor g62 (n_126, A[9], B[9]);
  xor g63 (Z[9], n_122, n_126);
  nand g64 (n_128, A[10], B[10]);
  nand g65 (n_129, A[10], n_127);
  nand g66 (n_130, B[10], n_127);
  nand g67 (n_132, n_128, n_129, n_130);
  xor g68 (n_131, A[10], B[10]);
  xor g69 (Z[10], n_127, n_131);
  nand g70 (n_133, A[11], B[11]);
  nand g71 (n_134, A[11], n_132);
  nand g72 (n_135, B[11], n_132);
  nand g73 (n_137, n_133, n_134, n_135);
  xor g74 (n_136, A[11], B[11]);
  xor g75 (Z[11], n_132, n_136);
  nand g76 (n_138, A[12], B[12]);
  nand g77 (n_139, A[12], n_137);
  nand g78 (n_140, B[12], n_137);
  nand g79 (n_142, n_138, n_139, n_140);
  xor g80 (n_141, A[12], B[12]);
  xor g81 (Z[12], n_137, n_141);
  nand g82 (n_143, A[13], B[13]);
  nand g83 (n_144, A[13], n_142);
  nand g84 (n_145, B[13], n_142);
  nand g85 (n_147, n_143, n_144, n_145);
  xor g86 (n_146, A[13], B[13]);
  xor g87 (Z[13], n_142, n_146);
  nand g88 (n_148, A[14], B[14]);
  nand g89 (n_149, A[14], n_147);
  nand g90 (n_150, B[14], n_147);
  nand g91 (n_152, n_148, n_149, n_150);
  xor g92 (n_151, A[14], B[14]);
  xor g93 (Z[14], n_147, n_151);
  nand g94 (n_153, A[15], B[15]);
  nand g95 (n_154, A[15], n_152);
  nand g96 (n_155, B[15], n_152);
  nand g97 (n_157, n_153, n_154, n_155);
  xor g98 (n_156, A[15], B[15]);
  xor g99 (Z[15], n_152, n_156);
  nand g100 (n_158, A[16], B[16]);
  nand g101 (n_159, A[16], n_157);
  nand g102 (n_160, B[16], n_157);
  nand g103 (n_162, n_158, n_159, n_160);
  xor g104 (n_161, A[16], B[16]);
  xor g105 (Z[16], n_157, n_161);
  nand g106 (n_163, A[17], B[17]);
  nand g107 (n_164, A[17], n_162);
  nand g108 (n_165, B[17], n_162);
  nand g109 (n_167, n_163, n_164, n_165);
  xor g110 (n_166, A[17], B[17]);
  xor g111 (Z[17], n_162, n_166);
  nand g112 (n_168, A[18], B[18]);
  nand g113 (n_169, A[18], n_167);
  nand g114 (n_170, B[18], n_167);
  nand g115 (n_172, n_168, n_169, n_170);
  xor g116 (n_171, A[18], B[18]);
  xor g117 (Z[18], n_167, n_171);
  nand g118 (n_173, A[19], B[19]);
  nand g119 (n_174, A[19], n_172);
  nand g120 (n_175, B[19], n_172);
  nand g121 (n_177, n_173, n_174, n_175);
  xor g122 (n_176, A[19], B[19]);
  xor g123 (Z[19], n_172, n_176);
  nand g124 (n_178, A[20], B[20]);
  nand g125 (n_179, A[20], n_177);
  nand g126 (n_180, B[20], n_177);
  nand g127 (n_182, n_178, n_179, n_180);
  xor g128 (n_181, A[20], B[20]);
  xor g129 (Z[20], n_177, n_181);
  nand g130 (n_183, A[21], B[21]);
  nand g131 (n_184, A[21], n_182);
  nand g132 (n_185, B[21], n_182);
  nand g133 (n_187, n_183, n_184, n_185);
  xor g134 (n_186, A[21], B[21]);
  xor g135 (Z[21], n_182, n_186);
  nand g136 (n_188, A[22], B[22]);
  nand g137 (n_189, A[22], n_187);
  nand g138 (n_190, B[22], n_187);
  nand g139 (n_192, n_188, n_189, n_190);
  xor g140 (n_191, A[22], B[22]);
  xor g141 (Z[22], n_187, n_191);
  xor g147 (Z[23], n_192, n_196);
  xor g149 (n_196, A[23], B[23]);
  or g150 (n_84, wc, n_79);
  not gc (wc, A[1]);
  or g151 (n_85, wc0, n_79);
  not gc0 (wc0, B[1]);
  xnor g152 (Z[1], n_79, n_86);
endmodule

module add_signed_3180_2_GENERIC(A, B, Z);
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  add_signed_3180_2_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_3180_3_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  wire n_79, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97;
  wire n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105;
  wire n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113;
  wire n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121;
  wire n_122, n_123, n_124, n_125, n_126, n_127, n_128, n_129;
  wire n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137;
  wire n_138, n_139, n_140, n_141, n_142, n_143, n_144, n_145;
  wire n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153;
  wire n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_196;
  nand g4 (n_79, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_83, A[1], B[1]);
  nand g13 (n_87, n_83, n_84, n_85);
  xor g14 (n_86, A[1], B[1]);
  nand g16 (n_88, A[2], B[2]);
  nand g17 (n_89, A[2], n_87);
  nand g18 (n_90, B[2], n_87);
  nand g19 (n_92, n_88, n_89, n_90);
  xor g20 (n_91, A[2], B[2]);
  xor g21 (Z[2], n_87, n_91);
  nand g22 (n_93, A[3], B[3]);
  nand g23 (n_94, A[3], n_92);
  nand g24 (n_95, B[3], n_92);
  nand g25 (n_97, n_93, n_94, n_95);
  xor g26 (n_96, A[3], B[3]);
  xor g27 (Z[3], n_92, n_96);
  nand g28 (n_98, A[4], B[4]);
  nand g29 (n_99, A[4], n_97);
  nand g30 (n_100, B[4], n_97);
  nand g31 (n_102, n_98, n_99, n_100);
  xor g32 (n_101, A[4], B[4]);
  xor g33 (Z[4], n_97, n_101);
  nand g34 (n_103, A[5], B[5]);
  nand g35 (n_104, A[5], n_102);
  nand g36 (n_105, B[5], n_102);
  nand g37 (n_107, n_103, n_104, n_105);
  xor g38 (n_106, A[5], B[5]);
  xor g39 (Z[5], n_102, n_106);
  nand g40 (n_108, A[6], B[6]);
  nand g41 (n_109, A[6], n_107);
  nand g42 (n_110, B[6], n_107);
  nand g43 (n_112, n_108, n_109, n_110);
  xor g44 (n_111, A[6], B[6]);
  xor g45 (Z[6], n_107, n_111);
  nand g46 (n_113, A[7], B[7]);
  nand g47 (n_114, A[7], n_112);
  nand g48 (n_115, B[7], n_112);
  nand g49 (n_117, n_113, n_114, n_115);
  xor g50 (n_116, A[7], B[7]);
  xor g51 (Z[7], n_112, n_116);
  nand g52 (n_118, A[8], B[8]);
  nand g53 (n_119, A[8], n_117);
  nand g54 (n_120, B[8], n_117);
  nand g55 (n_122, n_118, n_119, n_120);
  xor g56 (n_121, A[8], B[8]);
  xor g57 (Z[8], n_117, n_121);
  nand g58 (n_123, A[9], B[9]);
  nand g59 (n_124, A[9], n_122);
  nand g60 (n_125, B[9], n_122);
  nand g61 (n_127, n_123, n_124, n_125);
  xor g62 (n_126, A[9], B[9]);
  xor g63 (Z[9], n_122, n_126);
  nand g64 (n_128, A[10], B[10]);
  nand g65 (n_129, A[10], n_127);
  nand g66 (n_130, B[10], n_127);
  nand g67 (n_132, n_128, n_129, n_130);
  xor g68 (n_131, A[10], B[10]);
  xor g69 (Z[10], n_127, n_131);
  nand g70 (n_133, A[11], B[11]);
  nand g71 (n_134, A[11], n_132);
  nand g72 (n_135, B[11], n_132);
  nand g73 (n_137, n_133, n_134, n_135);
  xor g74 (n_136, A[11], B[11]);
  xor g75 (Z[11], n_132, n_136);
  nand g76 (n_138, A[12], B[12]);
  nand g77 (n_139, A[12], n_137);
  nand g78 (n_140, B[12], n_137);
  nand g79 (n_142, n_138, n_139, n_140);
  xor g80 (n_141, A[12], B[12]);
  xor g81 (Z[12], n_137, n_141);
  nand g82 (n_143, A[13], B[13]);
  nand g83 (n_144, A[13], n_142);
  nand g84 (n_145, B[13], n_142);
  nand g85 (n_147, n_143, n_144, n_145);
  xor g86 (n_146, A[13], B[13]);
  xor g87 (Z[13], n_142, n_146);
  nand g88 (n_148, A[14], B[14]);
  nand g89 (n_149, A[14], n_147);
  nand g90 (n_150, B[14], n_147);
  nand g91 (n_152, n_148, n_149, n_150);
  xor g92 (n_151, A[14], B[14]);
  xor g93 (Z[14], n_147, n_151);
  nand g94 (n_153, A[15], B[15]);
  nand g95 (n_154, A[15], n_152);
  nand g96 (n_155, B[15], n_152);
  nand g97 (n_157, n_153, n_154, n_155);
  xor g98 (n_156, A[15], B[15]);
  xor g99 (Z[15], n_152, n_156);
  nand g100 (n_158, A[16], B[16]);
  nand g101 (n_159, A[16], n_157);
  nand g102 (n_160, B[16], n_157);
  nand g103 (n_162, n_158, n_159, n_160);
  xor g104 (n_161, A[16], B[16]);
  xor g105 (Z[16], n_157, n_161);
  nand g106 (n_163, A[17], B[17]);
  nand g107 (n_164, A[17], n_162);
  nand g108 (n_165, B[17], n_162);
  nand g109 (n_167, n_163, n_164, n_165);
  xor g110 (n_166, A[17], B[17]);
  xor g111 (Z[17], n_162, n_166);
  nand g112 (n_168, A[18], B[18]);
  nand g113 (n_169, A[18], n_167);
  nand g114 (n_170, B[18], n_167);
  nand g115 (n_172, n_168, n_169, n_170);
  xor g116 (n_171, A[18], B[18]);
  xor g117 (Z[18], n_167, n_171);
  nand g118 (n_173, A[19], B[19]);
  nand g119 (n_174, A[19], n_172);
  nand g120 (n_175, B[19], n_172);
  nand g121 (n_177, n_173, n_174, n_175);
  xor g122 (n_176, A[19], B[19]);
  xor g123 (Z[19], n_172, n_176);
  nand g124 (n_178, A[20], B[20]);
  nand g125 (n_179, A[20], n_177);
  nand g126 (n_180, B[20], n_177);
  nand g127 (n_182, n_178, n_179, n_180);
  xor g128 (n_181, A[20], B[20]);
  xor g129 (Z[20], n_177, n_181);
  nand g130 (n_183, A[21], B[21]);
  nand g131 (n_184, A[21], n_182);
  nand g132 (n_185, B[21], n_182);
  nand g133 (n_187, n_183, n_184, n_185);
  xor g134 (n_186, A[21], B[21]);
  xor g135 (Z[21], n_182, n_186);
  nand g136 (n_188, A[22], B[22]);
  nand g137 (n_189, A[22], n_187);
  nand g138 (n_190, B[22], n_187);
  nand g139 (n_192, n_188, n_189, n_190);
  xor g140 (n_191, A[22], B[22]);
  xor g141 (Z[22], n_187, n_191);
  xor g147 (Z[23], n_192, n_196);
  xor g149 (n_196, A[23], B[23]);
  or g150 (n_84, wc, n_79);
  not gc (wc, A[1]);
  or g151 (n_85, wc0, n_79);
  not gc0 (wc0, B[1]);
  xnor g152 (Z[1], n_79, n_86);
endmodule

module add_signed_3180_3_GENERIC(A, B, Z);
  input [25:0] A, B;
  output [23:0] Z;
  wire [25:0] A, B;
  wire [23:0] Z;
  add_signed_3180_3_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_33_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [21:0] A, B;
  output [22:0] Z;
  wire [21:0] A, B;
  wire [22:0] Z;
  wire n_71, n_72, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180;
  not g3 (Z[22], n_71);
  nand g4 (n_72, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_77, A[1], B[1]);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_117, A[9], B[9]);
  nand g59 (n_118, A[9], n_116);
  nand g60 (n_119, B[9], n_116);
  nand g61 (n_121, n_117, n_118, n_119);
  xor g62 (n_120, A[9], B[9]);
  xor g63 (Z[9], n_116, n_120);
  nand g64 (n_122, A[10], B[10]);
  nand g65 (n_123, A[10], n_121);
  nand g66 (n_124, B[10], n_121);
  nand g67 (n_126, n_122, n_123, n_124);
  xor g68 (n_125, A[10], B[10]);
  xor g69 (Z[10], n_121, n_125);
  nand g70 (n_127, A[11], B[11]);
  nand g71 (n_128, A[11], n_126);
  nand g72 (n_129, B[11], n_126);
  nand g73 (n_131, n_127, n_128, n_129);
  xor g74 (n_130, A[11], B[11]);
  xor g75 (Z[11], n_126, n_130);
  nand g76 (n_132, A[12], B[12]);
  nand g77 (n_133, A[12], n_131);
  nand g78 (n_134, B[12], n_131);
  nand g79 (n_136, n_132, n_133, n_134);
  xor g80 (n_135, A[12], B[12]);
  xor g81 (Z[12], n_131, n_135);
  nand g82 (n_137, A[13], B[13]);
  nand g83 (n_138, A[13], n_136);
  nand g84 (n_139, B[13], n_136);
  nand g85 (n_141, n_137, n_138, n_139);
  xor g86 (n_140, A[13], B[13]);
  xor g87 (Z[13], n_136, n_140);
  nand g88 (n_142, A[14], B[14]);
  nand g89 (n_143, A[14], n_141);
  nand g90 (n_144, B[14], n_141);
  nand g91 (n_146, n_142, n_143, n_144);
  xor g92 (n_145, A[14], B[14]);
  xor g93 (Z[14], n_141, n_145);
  nand g94 (n_147, A[15], B[15]);
  nand g95 (n_148, A[15], n_146);
  nand g96 (n_149, B[15], n_146);
  nand g97 (n_151, n_147, n_148, n_149);
  xor g98 (n_150, A[15], B[15]);
  xor g99 (Z[15], n_146, n_150);
  nand g100 (n_152, A[16], B[16]);
  nand g101 (n_153, A[16], n_151);
  nand g102 (n_154, B[16], n_151);
  nand g103 (n_156, n_152, n_153, n_154);
  xor g104 (n_155, A[16], B[16]);
  xor g105 (Z[16], n_151, n_155);
  nand g106 (n_157, A[17], B[17]);
  nand g107 (n_158, A[17], n_156);
  nand g108 (n_159, B[17], n_156);
  nand g109 (n_161, n_157, n_158, n_159);
  xor g110 (n_160, A[17], B[17]);
  xor g111 (Z[17], n_156, n_160);
  nand g112 (n_162, A[18], B[18]);
  nand g113 (n_163, A[18], n_161);
  nand g114 (n_164, B[18], n_161);
  nand g115 (n_166, n_162, n_163, n_164);
  xor g116 (n_165, A[18], B[18]);
  xor g117 (Z[18], n_161, n_165);
  nand g118 (n_167, A[19], B[19]);
  nand g119 (n_168, A[19], n_166);
  nand g120 (n_169, B[19], n_166);
  nand g121 (n_171, n_167, n_168, n_169);
  xor g122 (n_170, A[19], B[19]);
  xor g123 (Z[19], n_166, n_170);
  nand g124 (n_172, A[20], B[20]);
  nand g125 (n_173, A[20], n_171);
  nand g126 (n_174, B[20], n_171);
  nand g127 (n_176, n_172, n_173, n_174);
  xor g128 (n_175, A[20], B[20]);
  xor g129 (Z[20], n_171, n_175);
  nand g133 (n_71, n_177, n_178, n_179);
  xor g135 (Z[21], n_176, n_180);
  or g137 (n_177, A[21], B[21]);
  xor g138 (n_180, A[21], B[21]);
  or g139 (n_78, wc, n_72);
  not gc (wc, A[1]);
  or g140 (n_79, wc0, n_72);
  not gc0 (wc0, B[1]);
  xnor g141 (Z[1], n_72, n_80);
  or g142 (n_178, A[21], wc1);
  not gc1 (wc1, n_176);
  or g143 (n_179, B[21], wc2);
  not gc2 (wc2, n_176);
endmodule

module add_signed_33_GENERIC(A, B, Z);
  input [21:0] A, B;
  output [22:0] Z;
  wire [21:0] A, B;
  wire [22:0] Z;
  add_signed_33_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_62_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [20:0] A, B;
  output [21:0] Z;
  wire [20:0] A, B;
  wire [21:0] Z;
  wire n_68, n_69, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172;
  not g3 (Z[21], n_68);
  nand g4 (n_69, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_74, A[1], B[1]);
  nand g13 (n_78, n_74, n_75, n_76);
  xor g14 (n_77, A[1], B[1]);
  nand g16 (n_79, A[2], B[2]);
  nand g17 (n_80, A[2], n_78);
  nand g18 (n_81, B[2], n_78);
  nand g19 (n_83, n_79, n_80, n_81);
  xor g20 (n_82, A[2], B[2]);
  xor g21 (Z[2], n_78, n_82);
  nand g22 (n_84, A[3], B[3]);
  nand g23 (n_85, A[3], n_83);
  nand g24 (n_86, B[3], n_83);
  nand g25 (n_88, n_84, n_85, n_86);
  xor g26 (n_87, A[3], B[3]);
  xor g27 (Z[3], n_83, n_87);
  nand g28 (n_89, A[4], B[4]);
  nand g29 (n_90, A[4], n_88);
  nand g30 (n_91, B[4], n_88);
  nand g31 (n_93, n_89, n_90, n_91);
  xor g32 (n_92, A[4], B[4]);
  xor g33 (Z[4], n_88, n_92);
  nand g34 (n_94, A[5], B[5]);
  nand g35 (n_95, A[5], n_93);
  nand g36 (n_96, B[5], n_93);
  nand g37 (n_98, n_94, n_95, n_96);
  xor g38 (n_97, A[5], B[5]);
  xor g39 (Z[5], n_93, n_97);
  nand g40 (n_99, A[6], B[6]);
  nand g41 (n_100, A[6], n_98);
  nand g42 (n_101, B[6], n_98);
  nand g43 (n_103, n_99, n_100, n_101);
  xor g44 (n_102, A[6], B[6]);
  xor g45 (Z[6], n_98, n_102);
  nand g46 (n_104, A[7], B[7]);
  nand g47 (n_105, A[7], n_103);
  nand g48 (n_106, B[7], n_103);
  nand g49 (n_108, n_104, n_105, n_106);
  xor g50 (n_107, A[7], B[7]);
  xor g51 (Z[7], n_103, n_107);
  nand g52 (n_109, A[8], B[8]);
  nand g53 (n_110, A[8], n_108);
  nand g54 (n_111, B[8], n_108);
  nand g55 (n_113, n_109, n_110, n_111);
  xor g56 (n_112, A[8], B[8]);
  xor g57 (Z[8], n_108, n_112);
  nand g58 (n_114, A[9], B[9]);
  nand g59 (n_115, A[9], n_113);
  nand g60 (n_116, B[9], n_113);
  nand g61 (n_118, n_114, n_115, n_116);
  xor g62 (n_117, A[9], B[9]);
  xor g63 (Z[9], n_113, n_117);
  nand g64 (n_119, A[10], B[10]);
  nand g65 (n_120, A[10], n_118);
  nand g66 (n_121, B[10], n_118);
  nand g67 (n_123, n_119, n_120, n_121);
  xor g68 (n_122, A[10], B[10]);
  xor g69 (Z[10], n_118, n_122);
  nand g70 (n_124, A[11], B[11]);
  nand g71 (n_125, A[11], n_123);
  nand g72 (n_126, B[11], n_123);
  nand g73 (n_128, n_124, n_125, n_126);
  xor g74 (n_127, A[11], B[11]);
  xor g75 (Z[11], n_123, n_127);
  nand g76 (n_129, A[12], B[12]);
  nand g77 (n_130, A[12], n_128);
  nand g78 (n_131, B[12], n_128);
  nand g79 (n_133, n_129, n_130, n_131);
  xor g80 (n_132, A[12], B[12]);
  xor g81 (Z[12], n_128, n_132);
  nand g82 (n_134, A[13], B[13]);
  nand g83 (n_135, A[13], n_133);
  nand g84 (n_136, B[13], n_133);
  nand g85 (n_138, n_134, n_135, n_136);
  xor g86 (n_137, A[13], B[13]);
  xor g87 (Z[13], n_133, n_137);
  nand g88 (n_139, A[14], B[14]);
  nand g89 (n_140, A[14], n_138);
  nand g90 (n_141, B[14], n_138);
  nand g91 (n_143, n_139, n_140, n_141);
  xor g92 (n_142, A[14], B[14]);
  xor g93 (Z[14], n_138, n_142);
  nand g94 (n_144, A[15], B[15]);
  nand g95 (n_145, A[15], n_143);
  nand g96 (n_146, B[15], n_143);
  nand g97 (n_148, n_144, n_145, n_146);
  xor g98 (n_147, A[15], B[15]);
  xor g99 (Z[15], n_143, n_147);
  nand g100 (n_149, A[16], B[16]);
  nand g101 (n_150, A[16], n_148);
  nand g102 (n_151, B[16], n_148);
  nand g103 (n_153, n_149, n_150, n_151);
  xor g104 (n_152, A[16], B[16]);
  xor g105 (Z[16], n_148, n_152);
  nand g106 (n_154, A[17], B[17]);
  nand g107 (n_155, A[17], n_153);
  nand g108 (n_156, B[17], n_153);
  nand g109 (n_158, n_154, n_155, n_156);
  xor g110 (n_157, A[17], B[17]);
  xor g111 (Z[17], n_153, n_157);
  nand g112 (n_159, A[18], B[18]);
  nand g113 (n_160, A[18], n_158);
  nand g114 (n_161, B[18], n_158);
  nand g115 (n_163, n_159, n_160, n_161);
  xor g116 (n_162, A[18], B[18]);
  xor g117 (Z[18], n_158, n_162);
  nand g118 (n_164, A[19], B[19]);
  nand g119 (n_165, A[19], n_163);
  nand g120 (n_166, B[19], n_163);
  nand g121 (n_168, n_164, n_165, n_166);
  xor g122 (n_167, A[19], B[19]);
  xor g123 (Z[19], n_163, n_167);
  nand g127 (n_68, n_169, n_170, n_171);
  xor g129 (Z[20], n_168, n_172);
  or g131 (n_169, A[20], B[20]);
  xor g132 (n_172, A[20], B[20]);
  or g133 (n_75, wc, n_69);
  not gc (wc, A[1]);
  or g134 (n_76, wc0, n_69);
  not gc0 (wc0, B[1]);
  xnor g135 (Z[1], n_69, n_77);
  or g136 (n_170, A[20], wc1);
  not gc1 (wc1, n_168);
  or g137 (n_171, B[20], wc2);
  not gc2 (wc2, n_168);
endmodule

module add_signed_62_GENERIC(A, B, Z);
  input [20:0] A, B;
  output [21:0] Z;
  wire [20:0] A, B;
  wire [21:0] Z;
  add_signed_62_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_65_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [21:0] A, B;
  output [22:0] Z;
  wire [21:0] A, B;
  wire [22:0] Z;
  wire n_71, n_72, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180;
  not g3 (Z[22], n_71);
  nand g4 (n_72, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_77, A[1], B[1]);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_117, A[9], B[9]);
  nand g59 (n_118, A[9], n_116);
  nand g60 (n_119, B[9], n_116);
  nand g61 (n_121, n_117, n_118, n_119);
  xor g62 (n_120, A[9], B[9]);
  xor g63 (Z[9], n_116, n_120);
  nand g64 (n_122, A[10], B[10]);
  nand g65 (n_123, A[10], n_121);
  nand g66 (n_124, B[10], n_121);
  nand g67 (n_126, n_122, n_123, n_124);
  xor g68 (n_125, A[10], B[10]);
  xor g69 (Z[10], n_121, n_125);
  nand g70 (n_127, A[11], B[11]);
  nand g71 (n_128, A[11], n_126);
  nand g72 (n_129, B[11], n_126);
  nand g73 (n_131, n_127, n_128, n_129);
  xor g74 (n_130, A[11], B[11]);
  xor g75 (Z[11], n_126, n_130);
  nand g76 (n_132, A[12], B[12]);
  nand g77 (n_133, A[12], n_131);
  nand g78 (n_134, B[12], n_131);
  nand g79 (n_136, n_132, n_133, n_134);
  xor g80 (n_135, A[12], B[12]);
  xor g81 (Z[12], n_131, n_135);
  nand g82 (n_137, A[13], B[13]);
  nand g83 (n_138, A[13], n_136);
  nand g84 (n_139, B[13], n_136);
  nand g85 (n_141, n_137, n_138, n_139);
  xor g86 (n_140, A[13], B[13]);
  xor g87 (Z[13], n_136, n_140);
  nand g88 (n_142, A[14], B[14]);
  nand g89 (n_143, A[14], n_141);
  nand g90 (n_144, B[14], n_141);
  nand g91 (n_146, n_142, n_143, n_144);
  xor g92 (n_145, A[14], B[14]);
  xor g93 (Z[14], n_141, n_145);
  nand g94 (n_147, A[15], B[15]);
  nand g95 (n_148, A[15], n_146);
  nand g96 (n_149, B[15], n_146);
  nand g97 (n_151, n_147, n_148, n_149);
  xor g98 (n_150, A[15], B[15]);
  xor g99 (Z[15], n_146, n_150);
  nand g100 (n_152, A[16], B[16]);
  nand g101 (n_153, A[16], n_151);
  nand g102 (n_154, B[16], n_151);
  nand g103 (n_156, n_152, n_153, n_154);
  xor g104 (n_155, A[16], B[16]);
  xor g105 (Z[16], n_151, n_155);
  nand g106 (n_157, A[17], B[17]);
  nand g107 (n_158, A[17], n_156);
  nand g108 (n_159, B[17], n_156);
  nand g109 (n_161, n_157, n_158, n_159);
  xor g110 (n_160, A[17], B[17]);
  xor g111 (Z[17], n_156, n_160);
  nand g112 (n_162, A[18], B[18]);
  nand g113 (n_163, A[18], n_161);
  nand g114 (n_164, B[18], n_161);
  nand g115 (n_166, n_162, n_163, n_164);
  xor g116 (n_165, A[18], B[18]);
  xor g117 (Z[18], n_161, n_165);
  nand g118 (n_167, A[19], B[19]);
  nand g119 (n_168, A[19], n_166);
  nand g120 (n_169, B[19], n_166);
  nand g121 (n_171, n_167, n_168, n_169);
  xor g122 (n_170, A[19], B[19]);
  xor g123 (Z[19], n_166, n_170);
  nand g124 (n_172, A[20], B[20]);
  nand g125 (n_173, A[20], n_171);
  nand g126 (n_174, B[20], n_171);
  nand g127 (n_176, n_172, n_173, n_174);
  xor g128 (n_175, A[20], B[20]);
  xor g129 (Z[20], n_171, n_175);
  nand g133 (n_71, n_177, n_178, n_179);
  xor g135 (Z[21], n_176, n_180);
  or g137 (n_177, A[21], B[21]);
  xor g138 (n_180, A[21], B[21]);
  or g139 (n_78, wc, n_72);
  not gc (wc, A[1]);
  or g140 (n_79, wc0, n_72);
  not gc0 (wc0, B[1]);
  xnor g141 (Z[1], n_72, n_80);
  or g142 (n_178, A[21], wc1);
  not gc1 (wc1, n_176);
  or g143 (n_179, B[21], wc2);
  not gc2 (wc2, n_176);
endmodule

module add_signed_65_GENERIC(A, B, Z);
  input [21:0] A, B;
  output [22:0] Z;
  wire [21:0] A, B;
  wire [22:0] Z;
  add_signed_65_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_6773_GENERIC_REAL(A, B, Z);
// synthesis_equation add_signed
  input [26:0] A, B;
  output [24:0] Z;
  wire [26:0] A, B;
  wire [24:0] Z;
  wire n_82, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_204;
  nand g4 (n_82, A[0], B[0]);
  xor g8 (Z[0], A[0], B[0]);
  nand g10 (n_86, A[1], B[1]);
  nand g13 (n_90, n_86, n_87, n_88);
  xor g14 (n_89, A[1], B[1]);
  nand g16 (n_91, A[2], B[2]);
  nand g17 (n_92, A[2], n_90);
  nand g18 (n_93, B[2], n_90);
  nand g19 (n_95, n_91, n_92, n_93);
  xor g20 (n_94, A[2], B[2]);
  xor g21 (Z[2], n_90, n_94);
  nand g22 (n_96, A[3], B[3]);
  nand g23 (n_97, A[3], n_95);
  nand g24 (n_98, B[3], n_95);
  nand g25 (n_100, n_96, n_97, n_98);
  xor g26 (n_99, A[3], B[3]);
  xor g27 (Z[3], n_95, n_99);
  nand g28 (n_101, A[4], B[4]);
  nand g29 (n_102, A[4], n_100);
  nand g30 (n_103, B[4], n_100);
  nand g31 (n_105, n_101, n_102, n_103);
  xor g32 (n_104, A[4], B[4]);
  xor g33 (Z[4], n_100, n_104);
  nand g34 (n_106, A[5], B[5]);
  nand g35 (n_107, A[5], n_105);
  nand g36 (n_108, B[5], n_105);
  nand g37 (n_110, n_106, n_107, n_108);
  xor g38 (n_109, A[5], B[5]);
  xor g39 (Z[5], n_105, n_109);
  nand g40 (n_111, A[6], B[6]);
  nand g41 (n_112, A[6], n_110);
  nand g42 (n_113, B[6], n_110);
  nand g43 (n_115, n_111, n_112, n_113);
  xor g44 (n_114, A[6], B[6]);
  xor g45 (Z[6], n_110, n_114);
  nand g46 (n_116, A[7], B[7]);
  nand g47 (n_117, A[7], n_115);
  nand g48 (n_118, B[7], n_115);
  nand g49 (n_120, n_116, n_117, n_118);
  xor g50 (n_119, A[7], B[7]);
  xor g51 (Z[7], n_115, n_119);
  nand g52 (n_121, A[8], B[8]);
  nand g53 (n_122, A[8], n_120);
  nand g54 (n_123, B[8], n_120);
  nand g55 (n_125, n_121, n_122, n_123);
  xor g56 (n_124, A[8], B[8]);
  xor g57 (Z[8], n_120, n_124);
  nand g58 (n_126, A[9], B[9]);
  nand g59 (n_127, A[9], n_125);
  nand g60 (n_128, B[9], n_125);
  nand g61 (n_130, n_126, n_127, n_128);
  xor g62 (n_129, A[9], B[9]);
  xor g63 (Z[9], n_125, n_129);
  nand g64 (n_131, A[10], B[10]);
  nand g65 (n_132, A[10], n_130);
  nand g66 (n_133, B[10], n_130);
  nand g67 (n_135, n_131, n_132, n_133);
  xor g68 (n_134, A[10], B[10]);
  xor g69 (Z[10], n_130, n_134);
  nand g70 (n_136, A[11], B[11]);
  nand g71 (n_137, A[11], n_135);
  nand g72 (n_138, B[11], n_135);
  nand g73 (n_140, n_136, n_137, n_138);
  xor g74 (n_139, A[11], B[11]);
  xor g75 (Z[11], n_135, n_139);
  nand g76 (n_141, A[12], B[12]);
  nand g77 (n_142, A[12], n_140);
  nand g78 (n_143, B[12], n_140);
  nand g79 (n_145, n_141, n_142, n_143);
  xor g80 (n_144, A[12], B[12]);
  xor g81 (Z[12], n_140, n_144);
  nand g82 (n_146, A[13], B[13]);
  nand g83 (n_147, A[13], n_145);
  nand g84 (n_148, B[13], n_145);
  nand g85 (n_150, n_146, n_147, n_148);
  xor g86 (n_149, A[13], B[13]);
  xor g87 (Z[13], n_145, n_149);
  nand g88 (n_151, A[14], B[14]);
  nand g89 (n_152, A[14], n_150);
  nand g90 (n_153, B[14], n_150);
  nand g91 (n_155, n_151, n_152, n_153);
  xor g92 (n_154, A[14], B[14]);
  xor g93 (Z[14], n_150, n_154);
  nand g94 (n_156, A[15], B[15]);
  nand g95 (n_157, A[15], n_155);
  nand g96 (n_158, B[15], n_155);
  nand g97 (n_160, n_156, n_157, n_158);
  xor g98 (n_159, A[15], B[15]);
  xor g99 (Z[15], n_155, n_159);
  nand g100 (n_161, A[16], B[16]);
  nand g101 (n_162, A[16], n_160);
  nand g102 (n_163, B[16], n_160);
  nand g103 (n_165, n_161, n_162, n_163);
  xor g104 (n_164, A[16], B[16]);
  xor g105 (Z[16], n_160, n_164);
  nand g106 (n_166, A[17], B[17]);
  nand g107 (n_167, A[17], n_165);
  nand g108 (n_168, B[17], n_165);
  nand g109 (n_170, n_166, n_167, n_168);
  xor g110 (n_169, A[17], B[17]);
  xor g111 (Z[17], n_165, n_169);
  nand g112 (n_171, A[18], B[18]);
  nand g113 (n_172, A[18], n_170);
  nand g114 (n_173, B[18], n_170);
  nand g115 (n_175, n_171, n_172, n_173);
  xor g116 (n_174, A[18], B[18]);
  xor g117 (Z[18], n_170, n_174);
  nand g118 (n_176, A[19], B[19]);
  nand g119 (n_177, A[19], n_175);
  nand g120 (n_178, B[19], n_175);
  nand g121 (n_180, n_176, n_177, n_178);
  xor g122 (n_179, A[19], B[19]);
  xor g123 (Z[19], n_175, n_179);
  nand g124 (n_181, A[20], B[20]);
  nand g125 (n_182, A[20], n_180);
  nand g126 (n_183, B[20], n_180);
  nand g127 (n_185, n_181, n_182, n_183);
  xor g128 (n_184, A[20], B[20]);
  xor g129 (Z[20], n_180, n_184);
  nand g130 (n_186, A[21], B[21]);
  nand g131 (n_187, A[21], n_185);
  nand g132 (n_188, B[21], n_185);
  nand g133 (n_190, n_186, n_187, n_188);
  xor g134 (n_189, A[21], B[21]);
  xor g135 (Z[21], n_185, n_189);
  nand g136 (n_191, A[22], B[22]);
  nand g137 (n_192, A[22], n_190);
  nand g138 (n_193, B[22], n_190);
  nand g139 (n_195, n_191, n_192, n_193);
  xor g140 (n_194, A[22], B[22]);
  xor g141 (Z[22], n_190, n_194);
  nand g142 (n_196, A[23], B[23]);
  nand g143 (n_197, A[23], n_195);
  nand g144 (n_198, B[23], n_195);
  nand g145 (n_200, n_196, n_197, n_198);
  xor g146 (n_199, A[23], B[23]);
  xor g147 (Z[23], n_195, n_199);
  xor g153 (Z[24], n_200, n_204);
  xor g155 (n_204, A[24], B[24]);
  or g156 (n_87, wc, n_82);
  not gc (wc, A[1]);
  or g157 (n_88, wc0, n_82);
  not gc0 (wc0, B[1]);
  xnor g158 (Z[1], n_82, n_89);
endmodule

module add_signed_6773_GENERIC(A, B, Z);
  input [26:0] A, B;
  output [24:0] Z;
  wire [26:0] A, B;
  wire [24:0] Z;
  add_signed_6773_GENERIC_REAL g1(.A (A), .B (B), .Z (Z));
endmodule

module add_signed_carry_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_signed_carry
  input [20:0] A, B;
  input CI;
  output [20:0] Z;
  wire [20:0] A, B;
  wire CI;
  wire [20:0] Z;
  wire n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_172;
  nand g4 (n_69, A[0], B[0]);
  nand g5 (n_70, A[0], CI);
  nand g6 (n_71, B[0], CI);
  nand g7 (n_73, n_69, n_70, n_71);
  xor g8 (n_72, A[0], B[0]);
  xor g9 (Z[0], CI, n_72);
  nand g10 (n_74, A[1], B[1]);
  nand g11 (n_75, A[1], n_73);
  nand g12 (n_76, B[1], n_73);
  nand g13 (n_78, n_74, n_75, n_76);
  xor g14 (n_77, A[1], B[1]);
  xor g15 (Z[1], n_73, n_77);
  nand g16 (n_79, A[2], B[2]);
  nand g17 (n_80, A[2], n_78);
  nand g18 (n_81, B[2], n_78);
  nand g19 (n_83, n_79, n_80, n_81);
  xor g20 (n_82, A[2], B[2]);
  xor g21 (Z[2], n_78, n_82);
  nand g22 (n_84, A[3], B[3]);
  nand g23 (n_85, A[3], n_83);
  nand g24 (n_86, B[3], n_83);
  nand g25 (n_88, n_84, n_85, n_86);
  xor g26 (n_87, A[3], B[3]);
  xor g27 (Z[3], n_83, n_87);
  nand g28 (n_89, A[4], B[4]);
  nand g29 (n_90, A[4], n_88);
  nand g30 (n_91, B[4], n_88);
  nand g31 (n_93, n_89, n_90, n_91);
  xor g32 (n_92, A[4], B[4]);
  xor g33 (Z[4], n_88, n_92);
  nand g34 (n_94, A[5], B[5]);
  nand g35 (n_95, A[5], n_93);
  nand g36 (n_96, B[5], n_93);
  nand g37 (n_98, n_94, n_95, n_96);
  xor g38 (n_97, A[5], B[5]);
  xor g39 (Z[5], n_93, n_97);
  nand g40 (n_99, A[6], B[6]);
  nand g41 (n_100, A[6], n_98);
  nand g42 (n_101, B[6], n_98);
  nand g43 (n_103, n_99, n_100, n_101);
  xor g44 (n_102, A[6], B[6]);
  xor g45 (Z[6], n_98, n_102);
  nand g46 (n_104, A[7], B[7]);
  nand g47 (n_105, A[7], n_103);
  nand g48 (n_106, B[7], n_103);
  nand g49 (n_108, n_104, n_105, n_106);
  xor g50 (n_107, A[7], B[7]);
  xor g51 (Z[7], n_103, n_107);
  nand g52 (n_109, A[8], B[8]);
  nand g53 (n_110, A[8], n_108);
  nand g54 (n_111, B[8], n_108);
  nand g55 (n_113, n_109, n_110, n_111);
  xor g56 (n_112, A[8], B[8]);
  xor g57 (Z[8], n_108, n_112);
  nand g58 (n_114, A[9], B[9]);
  nand g59 (n_115, A[9], n_113);
  nand g60 (n_116, B[9], n_113);
  nand g61 (n_118, n_114, n_115, n_116);
  xor g62 (n_117, A[9], B[9]);
  xor g63 (Z[9], n_113, n_117);
  nand g64 (n_119, A[10], B[10]);
  nand g65 (n_120, A[10], n_118);
  nand g66 (n_121, B[10], n_118);
  nand g67 (n_123, n_119, n_120, n_121);
  xor g68 (n_122, A[10], B[10]);
  xor g69 (Z[10], n_118, n_122);
  nand g70 (n_124, A[11], B[11]);
  nand g71 (n_125, A[11], n_123);
  nand g72 (n_126, B[11], n_123);
  nand g73 (n_128, n_124, n_125, n_126);
  xor g74 (n_127, A[11], B[11]);
  xor g75 (Z[11], n_123, n_127);
  nand g76 (n_129, A[12], B[12]);
  nand g77 (n_130, A[12], n_128);
  nand g78 (n_131, B[12], n_128);
  nand g79 (n_133, n_129, n_130, n_131);
  xor g80 (n_132, A[12], B[12]);
  xor g81 (Z[12], n_128, n_132);
  nand g82 (n_134, A[13], B[13]);
  nand g83 (n_135, A[13], n_133);
  nand g84 (n_136, B[13], n_133);
  nand g85 (n_138, n_134, n_135, n_136);
  xor g86 (n_137, A[13], B[13]);
  xor g87 (Z[13], n_133, n_137);
  nand g88 (n_139, A[14], B[14]);
  nand g89 (n_140, A[14], n_138);
  nand g90 (n_141, B[14], n_138);
  nand g91 (n_143, n_139, n_140, n_141);
  xor g92 (n_142, A[14], B[14]);
  xor g93 (Z[14], n_138, n_142);
  nand g94 (n_144, A[15], B[15]);
  nand g95 (n_145, A[15], n_143);
  nand g96 (n_146, B[15], n_143);
  nand g97 (n_148, n_144, n_145, n_146);
  xor g98 (n_147, A[15], B[15]);
  xor g99 (Z[15], n_143, n_147);
  nand g100 (n_149, A[16], B[16]);
  nand g101 (n_150, A[16], n_148);
  nand g102 (n_151, B[16], n_148);
  nand g103 (n_153, n_149, n_150, n_151);
  xor g104 (n_152, A[16], B[16]);
  xor g105 (Z[16], n_148, n_152);
  nand g106 (n_154, A[17], B[17]);
  nand g107 (n_155, A[17], n_153);
  nand g108 (n_156, B[17], n_153);
  nand g109 (n_158, n_154, n_155, n_156);
  xor g110 (n_157, A[17], B[17]);
  xor g111 (Z[17], n_153, n_157);
  nand g112 (n_159, A[18], B[18]);
  nand g113 (n_160, A[18], n_158);
  nand g114 (n_161, B[18], n_158);
  nand g115 (n_163, n_159, n_160, n_161);
  xor g116 (n_162, A[18], B[18]);
  xor g117 (Z[18], n_158, n_162);
  nand g118 (n_164, A[19], B[19]);
  nand g119 (n_165, A[19], n_163);
  nand g120 (n_166, B[19], n_163);
  nand g121 (n_168, n_164, n_165, n_166);
  xor g122 (n_167, A[19], B[19]);
  xor g123 (Z[19], n_163, n_167);
  xor g129 (Z[20], n_168, n_172);
  xor g130 (n_172, A[20], B[20]);
endmodule

module add_signed_carry_GENERIC(A, B, CI, Z);
  input [20:0] A, B;
  input CI;
  output [20:0] Z;
  wire [20:0] A, B;
  wire CI;
  wire [20:0] Z;
  add_signed_carry_GENERIC_REAL g1(.A ({A[19], A[19:0]}), .B ({B[19],
       B[19:0]}), .CI (CI), .Z (Z));
endmodule

module add_signed_carry_3209_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_signed_carry
  input [21:0] A, B;
  input CI;
  output [21:0] Z;
  wire [21:0] A, B;
  wire CI;
  wire [21:0] Z;
  wire n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_180;
  nand g4 (n_72, A[0], B[0]);
  nand g5 (n_73, A[0], CI);
  nand g6 (n_74, B[0], CI);
  nand g7 (n_76, n_72, n_73, n_74);
  xor g8 (n_75, A[0], B[0]);
  xor g9 (Z[0], CI, n_75);
  nand g10 (n_77, A[1], B[1]);
  nand g11 (n_78, A[1], n_76);
  nand g12 (n_79, B[1], n_76);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  xor g15 (Z[1], n_76, n_80);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_117, A[9], B[9]);
  nand g59 (n_118, A[9], n_116);
  nand g60 (n_119, B[9], n_116);
  nand g61 (n_121, n_117, n_118, n_119);
  xor g62 (n_120, A[9], B[9]);
  xor g63 (Z[9], n_116, n_120);
  nand g64 (n_122, A[10], B[10]);
  nand g65 (n_123, A[10], n_121);
  nand g66 (n_124, B[10], n_121);
  nand g67 (n_126, n_122, n_123, n_124);
  xor g68 (n_125, A[10], B[10]);
  xor g69 (Z[10], n_121, n_125);
  nand g70 (n_127, A[11], B[11]);
  nand g71 (n_128, A[11], n_126);
  nand g72 (n_129, B[11], n_126);
  nand g73 (n_131, n_127, n_128, n_129);
  xor g74 (n_130, A[11], B[11]);
  xor g75 (Z[11], n_126, n_130);
  nand g76 (n_132, A[12], B[12]);
  nand g77 (n_133, A[12], n_131);
  nand g78 (n_134, B[12], n_131);
  nand g79 (n_136, n_132, n_133, n_134);
  xor g80 (n_135, A[12], B[12]);
  xor g81 (Z[12], n_131, n_135);
  nand g82 (n_137, A[13], B[13]);
  nand g83 (n_138, A[13], n_136);
  nand g84 (n_139, B[13], n_136);
  nand g85 (n_141, n_137, n_138, n_139);
  xor g86 (n_140, A[13], B[13]);
  xor g87 (Z[13], n_136, n_140);
  nand g88 (n_142, A[14], B[14]);
  nand g89 (n_143, A[14], n_141);
  nand g90 (n_144, B[14], n_141);
  nand g91 (n_146, n_142, n_143, n_144);
  xor g92 (n_145, A[14], B[14]);
  xor g93 (Z[14], n_141, n_145);
  nand g94 (n_147, A[15], B[15]);
  nand g95 (n_148, A[15], n_146);
  nand g96 (n_149, B[15], n_146);
  nand g97 (n_151, n_147, n_148, n_149);
  xor g98 (n_150, A[15], B[15]);
  xor g99 (Z[15], n_146, n_150);
  nand g100 (n_152, A[16], B[16]);
  nand g101 (n_153, A[16], n_151);
  nand g102 (n_154, B[16], n_151);
  nand g103 (n_156, n_152, n_153, n_154);
  xor g104 (n_155, A[16], B[16]);
  xor g105 (Z[16], n_151, n_155);
  nand g106 (n_157, A[17], B[17]);
  nand g107 (n_158, A[17], n_156);
  nand g108 (n_159, B[17], n_156);
  nand g109 (n_161, n_157, n_158, n_159);
  xor g110 (n_160, A[17], B[17]);
  xor g111 (Z[17], n_156, n_160);
  nand g112 (n_162, A[18], B[18]);
  nand g113 (n_163, A[18], n_161);
  nand g114 (n_164, B[18], n_161);
  nand g115 (n_166, n_162, n_163, n_164);
  xor g116 (n_165, A[18], B[18]);
  xor g117 (Z[18], n_161, n_165);
  nand g118 (n_167, A[19], B[19]);
  nand g119 (n_168, A[19], n_166);
  nand g120 (n_169, B[19], n_166);
  nand g121 (n_171, n_167, n_168, n_169);
  xor g122 (n_170, A[19], B[19]);
  xor g123 (Z[19], n_166, n_170);
  nand g124 (n_172, A[20], B[20]);
  nand g125 (n_173, A[20], n_171);
  nand g126 (n_174, B[20], n_171);
  nand g127 (n_176, n_172, n_173, n_174);
  xor g128 (n_175, A[20], B[20]);
  xor g129 (Z[20], n_171, n_175);
  xor g135 (Z[21], n_176, n_180);
  xor g136 (n_180, A[21], B[21]);
endmodule

module add_signed_carry_3209_GENERIC(A, B, CI, Z);
  input [21:0] A, B;
  input CI;
  output [21:0] Z;
  wire [21:0] A, B;
  wire CI;
  wire [21:0] Z;
  add_signed_carry_3209_GENERIC_REAL g1(.A ({A[20], A[20:0]}), .B
       ({B[20], B[20:0]}), .CI (CI), .Z (Z));
endmodule

module add_signed_carry_3209_1_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_signed_carry
  input [21:0] A, B;
  input CI;
  output [21:0] Z;
  wire [21:0] A, B;
  wire CI;
  wire [21:0] Z;
  wire n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79;
  wire n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87;
  wire n_88, n_89, n_90, n_91, n_92, n_93, n_94, n_95;
  wire n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103;
  wire n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111;
  wire n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119;
  wire n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_180;
  nand g4 (n_72, A[0], B[0]);
  nand g5 (n_73, A[0], CI);
  nand g6 (n_74, B[0], CI);
  nand g7 (n_76, n_72, n_73, n_74);
  xor g8 (n_75, A[0], B[0]);
  xor g9 (Z[0], CI, n_75);
  nand g10 (n_77, A[1], B[1]);
  nand g11 (n_78, A[1], n_76);
  nand g12 (n_79, B[1], n_76);
  nand g13 (n_81, n_77, n_78, n_79);
  xor g14 (n_80, A[1], B[1]);
  xor g15 (Z[1], n_76, n_80);
  nand g16 (n_82, A[2], B[2]);
  nand g17 (n_83, A[2], n_81);
  nand g18 (n_84, B[2], n_81);
  nand g19 (n_86, n_82, n_83, n_84);
  xor g20 (n_85, A[2], B[2]);
  xor g21 (Z[2], n_81, n_85);
  nand g22 (n_87, A[3], B[3]);
  nand g23 (n_88, A[3], n_86);
  nand g24 (n_89, B[3], n_86);
  nand g25 (n_91, n_87, n_88, n_89);
  xor g26 (n_90, A[3], B[3]);
  xor g27 (Z[3], n_86, n_90);
  nand g28 (n_92, A[4], B[4]);
  nand g29 (n_93, A[4], n_91);
  nand g30 (n_94, B[4], n_91);
  nand g31 (n_96, n_92, n_93, n_94);
  xor g32 (n_95, A[4], B[4]);
  xor g33 (Z[4], n_91, n_95);
  nand g34 (n_97, A[5], B[5]);
  nand g35 (n_98, A[5], n_96);
  nand g36 (n_99, B[5], n_96);
  nand g37 (n_101, n_97, n_98, n_99);
  xor g38 (n_100, A[5], B[5]);
  xor g39 (Z[5], n_96, n_100);
  nand g40 (n_102, A[6], B[6]);
  nand g41 (n_103, A[6], n_101);
  nand g42 (n_104, B[6], n_101);
  nand g43 (n_106, n_102, n_103, n_104);
  xor g44 (n_105, A[6], B[6]);
  xor g45 (Z[6], n_101, n_105);
  nand g46 (n_107, A[7], B[7]);
  nand g47 (n_108, A[7], n_106);
  nand g48 (n_109, B[7], n_106);
  nand g49 (n_111, n_107, n_108, n_109);
  xor g50 (n_110, A[7], B[7]);
  xor g51 (Z[7], n_106, n_110);
  nand g52 (n_112, A[8], B[8]);
  nand g53 (n_113, A[8], n_111);
  nand g54 (n_114, B[8], n_111);
  nand g55 (n_116, n_112, n_113, n_114);
  xor g56 (n_115, A[8], B[8]);
  xor g57 (Z[8], n_111, n_115);
  nand g58 (n_117, A[9], B[9]);
  nand g59 (n_118, A[9], n_116);
  nand g60 (n_119, B[9], n_116);
  nand g61 (n_121, n_117, n_118, n_119);
  xor g62 (n_120, A[9], B[9]);
  xor g63 (Z[9], n_116, n_120);
  nand g64 (n_122, A[10], B[10]);
  nand g65 (n_123, A[10], n_121);
  nand g66 (n_124, B[10], n_121);
  nand g67 (n_126, n_122, n_123, n_124);
  xor g68 (n_125, A[10], B[10]);
  xor g69 (Z[10], n_121, n_125);
  nand g70 (n_127, A[11], B[11]);
  nand g71 (n_128, A[11], n_126);
  nand g72 (n_129, B[11], n_126);
  nand g73 (n_131, n_127, n_128, n_129);
  xor g74 (n_130, A[11], B[11]);
  xor g75 (Z[11], n_126, n_130);
  nand g76 (n_132, A[12], B[12]);
  nand g77 (n_133, A[12], n_131);
  nand g78 (n_134, B[12], n_131);
  nand g79 (n_136, n_132, n_133, n_134);
  xor g80 (n_135, A[12], B[12]);
  xor g81 (Z[12], n_131, n_135);
  nand g82 (n_137, A[13], B[13]);
  nand g83 (n_138, A[13], n_136);
  nand g84 (n_139, B[13], n_136);
  nand g85 (n_141, n_137, n_138, n_139);
  xor g86 (n_140, A[13], B[13]);
  xor g87 (Z[13], n_136, n_140);
  nand g88 (n_142, A[14], B[14]);
  nand g89 (n_143, A[14], n_141);
  nand g90 (n_144, B[14], n_141);
  nand g91 (n_146, n_142, n_143, n_144);
  xor g92 (n_145, A[14], B[14]);
  xor g93 (Z[14], n_141, n_145);
  nand g94 (n_147, A[15], B[15]);
  nand g95 (n_148, A[15], n_146);
  nand g96 (n_149, B[15], n_146);
  nand g97 (n_151, n_147, n_148, n_149);
  xor g98 (n_150, A[15], B[15]);
  xor g99 (Z[15], n_146, n_150);
  nand g100 (n_152, A[16], B[16]);
  nand g101 (n_153, A[16], n_151);
  nand g102 (n_154, B[16], n_151);
  nand g103 (n_156, n_152, n_153, n_154);
  xor g104 (n_155, A[16], B[16]);
  xor g105 (Z[16], n_151, n_155);
  nand g106 (n_157, A[17], B[17]);
  nand g107 (n_158, A[17], n_156);
  nand g108 (n_159, B[17], n_156);
  nand g109 (n_161, n_157, n_158, n_159);
  xor g110 (n_160, A[17], B[17]);
  xor g111 (Z[17], n_156, n_160);
  nand g112 (n_162, A[18], B[18]);
  nand g113 (n_163, A[18], n_161);
  nand g114 (n_164, B[18], n_161);
  nand g115 (n_166, n_162, n_163, n_164);
  xor g116 (n_165, A[18], B[18]);
  xor g117 (Z[18], n_161, n_165);
  nand g118 (n_167, A[19], B[19]);
  nand g119 (n_168, A[19], n_166);
  nand g120 (n_169, B[19], n_166);
  nand g121 (n_171, n_167, n_168, n_169);
  xor g122 (n_170, A[19], B[19]);
  xor g123 (Z[19], n_166, n_170);
  nand g124 (n_172, A[20], B[20]);
  nand g125 (n_173, A[20], n_171);
  nand g126 (n_174, B[20], n_171);
  nand g127 (n_176, n_172, n_173, n_174);
  xor g128 (n_175, A[20], B[20]);
  xor g129 (Z[20], n_171, n_175);
  xor g135 (Z[21], n_176, n_180);
  xor g136 (n_180, A[21], B[21]);
endmodule

module add_signed_carry_3209_1_GENERIC(A, B, CI, Z);
  input [21:0] A, B;
  input CI;
  output [21:0] Z;
  wire [21:0] A, B;
  wire CI;
  wire [21:0] Z;
  add_signed_carry_3209_1_GENERIC_REAL g1(.A ({A[20], A[20:0]}), .B
       ({B[20], B[20:0]}), .CI (CI), .Z (Z));
endmodule

module add_signed_carry_6718_GENERIC_REAL(A, B, CI, Z);
// synthesis_equation add_signed_carry
  input [22:0] A, B;
  input CI;
  output [22:0] Z;
  wire [22:0] A, B;
  wire CI;
  wire [22:0] Z;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_188;
  nand g4 (n_75, A[0], B[0]);
  nand g5 (n_76, A[0], CI);
  nand g6 (n_77, B[0], CI);
  nand g7 (n_79, n_75, n_76, n_77);
  xor g8 (n_78, A[0], B[0]);
  xor g9 (Z[0], CI, n_78);
  nand g10 (n_80, A[1], B[1]);
  nand g11 (n_81, A[1], n_79);
  nand g12 (n_82, B[1], n_79);
  nand g13 (n_84, n_80, n_81, n_82);
  xor g14 (n_83, A[1], B[1]);
  xor g15 (Z[1], n_79, n_83);
  nand g16 (n_85, A[2], B[2]);
  nand g17 (n_86, A[2], n_84);
  nand g18 (n_87, B[2], n_84);
  nand g19 (n_89, n_85, n_86, n_87);
  xor g20 (n_88, A[2], B[2]);
  xor g21 (Z[2], n_84, n_88);
  nand g22 (n_90, A[3], B[3]);
  nand g23 (n_91, A[3], n_89);
  nand g24 (n_92, B[3], n_89);
  nand g25 (n_94, n_90, n_91, n_92);
  xor g26 (n_93, A[3], B[3]);
  xor g27 (Z[3], n_89, n_93);
  nand g28 (n_95, A[4], B[4]);
  nand g29 (n_96, A[4], n_94);
  nand g30 (n_97, B[4], n_94);
  nand g31 (n_99, n_95, n_96, n_97);
  xor g32 (n_98, A[4], B[4]);
  xor g33 (Z[4], n_94, n_98);
  nand g34 (n_100, A[5], B[5]);
  nand g35 (n_101, A[5], n_99);
  nand g36 (n_102, B[5], n_99);
  nand g37 (n_104, n_100, n_101, n_102);
  xor g38 (n_103, A[5], B[5]);
  xor g39 (Z[5], n_99, n_103);
  nand g40 (n_105, A[6], B[6]);
  nand g41 (n_106, A[6], n_104);
  nand g42 (n_107, B[6], n_104);
  nand g43 (n_109, n_105, n_106, n_107);
  xor g44 (n_108, A[6], B[6]);
  xor g45 (Z[6], n_104, n_108);
  nand g46 (n_110, A[7], B[7]);
  nand g47 (n_111, A[7], n_109);
  nand g48 (n_112, B[7], n_109);
  nand g49 (n_114, n_110, n_111, n_112);
  xor g50 (n_113, A[7], B[7]);
  xor g51 (Z[7], n_109, n_113);
  nand g52 (n_115, A[8], B[8]);
  nand g53 (n_116, A[8], n_114);
  nand g54 (n_117, B[8], n_114);
  nand g55 (n_119, n_115, n_116, n_117);
  xor g56 (n_118, A[8], B[8]);
  xor g57 (Z[8], n_114, n_118);
  nand g58 (n_120, A[9], B[9]);
  nand g59 (n_121, A[9], n_119);
  nand g60 (n_122, B[9], n_119);
  nand g61 (n_124, n_120, n_121, n_122);
  xor g62 (n_123, A[9], B[9]);
  xor g63 (Z[9], n_119, n_123);
  nand g64 (n_125, A[10], B[10]);
  nand g65 (n_126, A[10], n_124);
  nand g66 (n_127, B[10], n_124);
  nand g67 (n_129, n_125, n_126, n_127);
  xor g68 (n_128, A[10], B[10]);
  xor g69 (Z[10], n_124, n_128);
  nand g70 (n_130, A[11], B[11]);
  nand g71 (n_131, A[11], n_129);
  nand g72 (n_132, B[11], n_129);
  nand g73 (n_134, n_130, n_131, n_132);
  xor g74 (n_133, A[11], B[11]);
  xor g75 (Z[11], n_129, n_133);
  nand g76 (n_135, A[12], B[12]);
  nand g77 (n_136, A[12], n_134);
  nand g78 (n_137, B[12], n_134);
  nand g79 (n_139, n_135, n_136, n_137);
  xor g80 (n_138, A[12], B[12]);
  xor g81 (Z[12], n_134, n_138);
  nand g82 (n_140, A[13], B[13]);
  nand g83 (n_141, A[13], n_139);
  nand g84 (n_142, B[13], n_139);
  nand g85 (n_144, n_140, n_141, n_142);
  xor g86 (n_143, A[13], B[13]);
  xor g87 (Z[13], n_139, n_143);
  nand g88 (n_145, A[14], B[14]);
  nand g89 (n_146, A[14], n_144);
  nand g90 (n_147, B[14], n_144);
  nand g91 (n_149, n_145, n_146, n_147);
  xor g92 (n_148, A[14], B[14]);
  xor g93 (Z[14], n_144, n_148);
  nand g94 (n_150, A[15], B[15]);
  nand g95 (n_151, A[15], n_149);
  nand g96 (n_152, B[15], n_149);
  nand g97 (n_154, n_150, n_151, n_152);
  xor g98 (n_153, A[15], B[15]);
  xor g99 (Z[15], n_149, n_153);
  nand g100 (n_155, A[16], B[16]);
  nand g101 (n_156, A[16], n_154);
  nand g102 (n_157, B[16], n_154);
  nand g103 (n_159, n_155, n_156, n_157);
  xor g104 (n_158, A[16], B[16]);
  xor g105 (Z[16], n_154, n_158);
  nand g106 (n_160, A[17], B[17]);
  nand g107 (n_161, A[17], n_159);
  nand g108 (n_162, B[17], n_159);
  nand g109 (n_164, n_160, n_161, n_162);
  xor g110 (n_163, A[17], B[17]);
  xor g111 (Z[17], n_159, n_163);
  nand g112 (n_165, A[18], B[18]);
  nand g113 (n_166, A[18], n_164);
  nand g114 (n_167, B[18], n_164);
  nand g115 (n_169, n_165, n_166, n_167);
  xor g116 (n_168, A[18], B[18]);
  xor g117 (Z[18], n_164, n_168);
  nand g118 (n_170, A[19], B[19]);
  nand g119 (n_171, A[19], n_169);
  nand g120 (n_172, B[19], n_169);
  nand g121 (n_174, n_170, n_171, n_172);
  xor g122 (n_173, A[19], B[19]);
  xor g123 (Z[19], n_169, n_173);
  nand g124 (n_175, A[20], B[20]);
  nand g125 (n_176, A[20], n_174);
  nand g126 (n_177, B[20], n_174);
  nand g127 (n_179, n_175, n_176, n_177);
  xor g128 (n_178, A[20], B[20]);
  xor g129 (Z[20], n_174, n_178);
  nand g130 (n_180, A[21], B[21]);
  nand g131 (n_181, A[21], n_179);
  nand g132 (n_182, B[21], n_179);
  nand g133 (n_184, n_180, n_181, n_182);
  xor g134 (n_183, A[21], B[21]);
  xor g135 (Z[21], n_179, n_183);
  xor g141 (Z[22], n_184, n_188);
  xor g142 (n_188, A[22], B[22]);
endmodule

module add_signed_carry_6718_GENERIC(A, B, CI, Z);
  input [22:0] A, B;
  input CI;
  output [22:0] Z;
  wire [22:0] A, B;
  wire CI;
  wire [22:0] Z;
  add_signed_carry_6718_GENERIC_REAL g1(.A ({A[21], A[21:0]}), .B
       ({B[21], B[21:0]}), .CI (CI), .Z (Z));
endmodule

module csa_tree_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 24'b0;"
  input [20:0] in_0, in_1, in_2;
  output [23:0] out_0, out_1;
  wire [20:0] in_0, in_1, in_2;
  wire [23:0] out_0, out_1;
  wire n_67, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_194;
  assign out_1[22] = 1'b0;
  assign out_1[23] = 1'b0;
  assign out_0[0] = in_1[0];
  assign out_0[22] = 1'b1;
  assign out_0[23] = 1'b1;
  xor g26 (out_1[0], in_0[0], in_2[0]);
  and g27 (out_0[1], in_0[0], in_2[0]);
  xor g28 (n_116, in_0[1], in_1[1]);
  xor g29 (out_1[1], n_116, in_2[1]);
  nand g30 (n_117, in_0[1], in_1[1]);
  nand g4 (n_118, in_2[1], in_1[1]);
  nand g5 (n_119, in_0[1], in_2[1]);
  nand g31 (out_0[2], n_117, n_118, n_119);
  xor g32 (n_120, in_0[2], in_1[2]);
  xor g33 (out_1[2], n_120, in_2[2]);
  nand g34 (n_121, in_0[2], in_1[2]);
  nand g35 (n_122, in_2[2], in_1[2]);
  nand g36 (n_123, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_121, n_122, n_123);
  xor g37 (n_124, in_0[3], in_1[3]);
  xor g38 (out_1[3], n_124, in_2[3]);
  nand g39 (n_125, in_0[3], in_1[3]);
  nand g40 (n_126, in_2[3], in_1[3]);
  nand g41 (n_127, in_0[3], in_2[3]);
  nand g42 (out_0[4], n_125, n_126, n_127);
  xor g43 (n_128, in_0[4], in_1[4]);
  xor g44 (out_1[4], n_128, in_2[4]);
  nand g45 (n_129, in_0[4], in_1[4]);
  nand g46 (n_130, in_2[4], in_1[4]);
  nand g47 (n_131, in_0[4], in_2[4]);
  nand g48 (out_0[5], n_129, n_130, n_131);
  xor g49 (n_132, in_0[5], in_1[5]);
  xor g50 (out_1[5], n_132, in_2[5]);
  nand g51 (n_133, in_0[5], in_1[5]);
  nand g52 (n_134, in_2[5], in_1[5]);
  nand g53 (n_135, in_0[5], in_2[5]);
  nand g54 (out_0[6], n_133, n_134, n_135);
  xor g55 (n_136, in_0[6], in_1[6]);
  xor g56 (out_1[6], n_136, in_2[6]);
  nand g57 (n_137, in_0[6], in_1[6]);
  nand g58 (n_138, in_2[6], in_1[6]);
  nand g59 (n_139, in_0[6], in_2[6]);
  nand g60 (out_0[7], n_137, n_138, n_139);
  xor g61 (n_140, in_0[7], in_1[7]);
  xor g62 (out_1[7], n_140, in_2[7]);
  nand g63 (n_141, in_0[7], in_1[7]);
  nand g64 (n_142, in_2[7], in_1[7]);
  nand g65 (n_143, in_0[7], in_2[7]);
  nand g66 (out_0[8], n_141, n_142, n_143);
  xor g67 (n_144, in_0[8], in_1[8]);
  xor g68 (out_1[8], n_144, in_2[8]);
  nand g69 (n_145, in_0[8], in_1[8]);
  nand g70 (n_146, in_2[8], in_1[8]);
  nand g71 (n_147, in_0[8], in_2[8]);
  nand g72 (out_0[9], n_145, n_146, n_147);
  xor g73 (n_148, in_0[9], in_1[9]);
  xor g74 (out_1[9], n_148, in_2[9]);
  nand g75 (n_149, in_0[9], in_1[9]);
  nand g76 (n_150, in_2[9], in_1[9]);
  nand g77 (n_151, in_0[9], in_2[9]);
  nand g78 (out_0[10], n_149, n_150, n_151);
  xor g79 (n_152, in_0[10], in_1[10]);
  xor g80 (out_1[10], n_152, in_2[10]);
  nand g81 (n_153, in_0[10], in_1[10]);
  nand g82 (n_154, in_2[10], in_1[10]);
  nand g83 (n_155, in_0[10], in_2[10]);
  nand g84 (out_0[11], n_153, n_154, n_155);
  xor g85 (n_156, in_0[11], in_1[11]);
  xor g86 (out_1[11], n_156, in_2[11]);
  nand g87 (n_157, in_0[11], in_1[11]);
  nand g88 (n_158, in_2[11], in_1[11]);
  nand g89 (n_159, in_0[11], in_2[11]);
  nand g90 (out_0[12], n_157, n_158, n_159);
  xor g91 (n_160, in_0[12], in_1[12]);
  xor g92 (out_1[12], n_160, in_2[12]);
  nand g93 (n_161, in_0[12], in_1[12]);
  nand g94 (n_162, in_2[12], in_1[12]);
  nand g95 (n_163, in_0[12], in_2[12]);
  nand g96 (out_0[13], n_161, n_162, n_163);
  xor g97 (n_164, in_0[13], in_1[13]);
  xor g98 (out_1[13], n_164, in_2[13]);
  nand g99 (n_165, in_0[13], in_1[13]);
  nand g100 (n_166, in_2[13], in_1[13]);
  nand g101 (n_167, in_0[13], in_2[13]);
  nand g102 (out_0[14], n_165, n_166, n_167);
  xor g103 (n_168, in_0[14], in_1[14]);
  xor g104 (out_1[14], n_168, in_2[14]);
  nand g105 (n_169, in_0[14], in_1[14]);
  nand g106 (n_170, in_2[14], in_1[14]);
  nand g107 (n_171, in_0[14], in_2[14]);
  nand g108 (out_0[15], n_169, n_170, n_171);
  xor g109 (n_172, in_0[15], in_1[15]);
  xor g110 (out_1[15], n_172, in_2[15]);
  nand g111 (n_173, in_0[15], in_1[15]);
  nand g112 (n_174, in_2[15], in_1[15]);
  nand g113 (n_175, in_0[15], in_2[15]);
  nand g114 (out_0[16], n_173, n_174, n_175);
  xor g115 (n_176, in_0[16], in_1[16]);
  xor g116 (out_1[16], n_176, in_2[16]);
  nand g117 (n_177, in_0[16], in_1[16]);
  nand g118 (n_178, in_2[16], in_1[16]);
  nand g119 (n_179, in_0[16], in_2[16]);
  nand g120 (out_0[17], n_177, n_178, n_179);
  xor g121 (n_180, in_0[17], in_1[17]);
  xor g122 (out_1[17], n_180, in_2[17]);
  nand g123 (n_181, in_0[17], in_1[17]);
  nand g124 (n_182, in_2[17], in_1[17]);
  nand g125 (n_183, in_0[17], in_2[17]);
  nand g126 (out_0[18], n_181, n_182, n_183);
  xor g127 (n_184, in_0[18], in_1[18]);
  xor g128 (out_1[18], n_184, in_2[18]);
  nand g129 (n_185, in_0[18], in_1[18]);
  nand g130 (n_186, in_2[18], in_1[18]);
  nand g131 (n_187, in_0[18], in_2[18]);
  nand g132 (out_0[19], n_185, n_186, n_187);
  xor g133 (n_188, in_0[19], in_1[19]);
  xor g134 (out_1[19], n_188, in_2[19]);
  nand g135 (n_189, in_0[19], in_1[19]);
  nand g136 (n_190, in_2[19], in_1[19]);
  nand g137 (n_191, in_0[19], in_2[19]);
  nand g138 (out_0[20], n_189, n_190, n_191);
  xor g142 (out_1[20], in_2[20], n_67);
  xor g147 (n_67, in_0[20], in_1[20]);
  nor g148 (out_0[21], in_0[20], in_1[20]);
  or g149 (n_194, in_2[20], wc);
  not gc (wc, n_67);
  or g151 (out_1[21], wc0, wc1, n_67);
  not gc1 (wc1, n_194);
  not gc0 (wc0, in_2[20]);
endmodule

module csa_tree_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [20:0] in_0, in_1, in_2;
  output [23:0] out_0, out_1;
  wire [20:0] in_0, in_1, in_2;
  wire [23:0] out_0, out_1;
  csa_tree_GENERIC_REAL g1(.in_0 ({in_0[19], in_0[19:0]}), .in_1
       ({in_1[19], in_1[19:0]}), .in_2 (in_2), .out_0 (out_0), .out_1
       (out_1));
endmodule

module csa_tree_3124_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 25'b0;"
  input [23:0] in_0, in_1;
  input [21:0] in_2;
  output [24:0] out_0, out_1;
  wire [23:0] in_0, in_1;
  wire [21:0] in_2;
  wire [24:0] out_0, out_1;
  wire n_70, n_74, n_75, n_79, n_80, n_131, n_132, n_133;
  wire n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141;
  wire n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149;
  wire n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157;
  wire n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_213, n_217, n_221;
  assign out_0[0] = in_1[0];
  xor g31 (out_1[0], in_0[0], in_2[0]);
  and g32 (out_0[1], in_0[0], in_2[0]);
  xor g33 (n_131, in_0[1], in_1[1]);
  xor g34 (out_1[1], n_131, in_2[1]);
  nand g35 (n_132, in_0[1], in_1[1]);
  nand g4 (n_133, in_2[1], in_1[1]);
  nand g5 (n_134, in_0[1], in_2[1]);
  nand g36 (out_0[2], n_132, n_133, n_134);
  xor g37 (n_135, in_0[2], in_1[2]);
  xor g38 (out_1[2], n_135, in_2[2]);
  nand g39 (n_136, in_0[2], in_1[2]);
  nand g40 (n_137, in_2[2], in_1[2]);
  nand g41 (n_138, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_136, n_137, n_138);
  xor g42 (n_139, in_0[3], in_1[3]);
  xor g43 (out_1[3], n_139, in_2[3]);
  nand g44 (n_140, in_0[3], in_1[3]);
  nand g45 (n_141, in_2[3], in_1[3]);
  nand g46 (n_142, in_0[3], in_2[3]);
  nand g47 (out_0[4], n_140, n_141, n_142);
  xor g48 (n_143, in_0[4], in_1[4]);
  xor g49 (out_1[4], n_143, in_2[4]);
  nand g50 (n_144, in_0[4], in_1[4]);
  nand g51 (n_145, in_2[4], in_1[4]);
  nand g52 (n_146, in_0[4], in_2[4]);
  nand g53 (out_0[5], n_144, n_145, n_146);
  xor g54 (n_147, in_0[5], in_1[5]);
  xor g55 (out_1[5], n_147, in_2[5]);
  nand g56 (n_148, in_0[5], in_1[5]);
  nand g57 (n_149, in_2[5], in_1[5]);
  nand g58 (n_150, in_0[5], in_2[5]);
  nand g59 (out_0[6], n_148, n_149, n_150);
  xor g60 (n_151, in_0[6], in_1[6]);
  xor g61 (out_1[6], n_151, in_2[6]);
  nand g62 (n_152, in_0[6], in_1[6]);
  nand g63 (n_153, in_2[6], in_1[6]);
  nand g64 (n_154, in_0[6], in_2[6]);
  nand g65 (out_0[7], n_152, n_153, n_154);
  xor g66 (n_155, in_0[7], in_1[7]);
  xor g67 (out_1[7], n_155, in_2[7]);
  nand g68 (n_156, in_0[7], in_1[7]);
  nand g69 (n_157, in_2[7], in_1[7]);
  nand g70 (n_158, in_0[7], in_2[7]);
  nand g71 (out_0[8], n_156, n_157, n_158);
  xor g72 (n_159, in_0[8], in_1[8]);
  xor g73 (out_1[8], n_159, in_2[8]);
  nand g74 (n_160, in_0[8], in_1[8]);
  nand g75 (n_161, in_2[8], in_1[8]);
  nand g76 (n_162, in_0[8], in_2[8]);
  nand g77 (out_0[9], n_160, n_161, n_162);
  xor g78 (n_163, in_0[9], in_1[9]);
  xor g79 (out_1[9], n_163, in_2[9]);
  nand g80 (n_164, in_0[9], in_1[9]);
  nand g81 (n_165, in_2[9], in_1[9]);
  nand g82 (n_166, in_0[9], in_2[9]);
  nand g83 (out_0[10], n_164, n_165, n_166);
  xor g84 (n_167, in_0[10], in_1[10]);
  xor g85 (out_1[10], n_167, in_2[10]);
  nand g86 (n_168, in_0[10], in_1[10]);
  nand g87 (n_169, in_2[10], in_1[10]);
  nand g88 (n_170, in_0[10], in_2[10]);
  nand g89 (out_0[11], n_168, n_169, n_170);
  xor g90 (n_171, in_0[11], in_1[11]);
  xor g91 (out_1[11], n_171, in_2[11]);
  nand g92 (n_172, in_0[11], in_1[11]);
  nand g93 (n_173, in_2[11], in_1[11]);
  nand g94 (n_174, in_0[11], in_2[11]);
  nand g95 (out_0[12], n_172, n_173, n_174);
  xor g96 (n_175, in_0[12], in_1[12]);
  xor g97 (out_1[12], n_175, in_2[12]);
  nand g98 (n_176, in_0[12], in_1[12]);
  nand g99 (n_177, in_2[12], in_1[12]);
  nand g100 (n_178, in_0[12], in_2[12]);
  nand g101 (out_0[13], n_176, n_177, n_178);
  xor g102 (n_179, in_0[13], in_1[13]);
  xor g103 (out_1[13], n_179, in_2[13]);
  nand g104 (n_180, in_0[13], in_1[13]);
  nand g105 (n_181, in_2[13], in_1[13]);
  nand g106 (n_182, in_0[13], in_2[13]);
  nand g107 (out_0[14], n_180, n_181, n_182);
  xor g108 (n_183, in_0[14], in_1[14]);
  xor g109 (out_1[14], n_183, in_2[14]);
  nand g110 (n_184, in_0[14], in_1[14]);
  nand g111 (n_185, in_2[14], in_1[14]);
  nand g112 (n_186, in_0[14], in_2[14]);
  nand g113 (out_0[15], n_184, n_185, n_186);
  xor g114 (n_187, in_0[15], in_1[15]);
  xor g115 (out_1[15], n_187, in_2[15]);
  nand g116 (n_188, in_0[15], in_1[15]);
  nand g117 (n_189, in_2[15], in_1[15]);
  nand g118 (n_190, in_0[15], in_2[15]);
  nand g119 (out_0[16], n_188, n_189, n_190);
  xor g120 (n_191, in_0[16], in_1[16]);
  xor g121 (out_1[16], n_191, in_2[16]);
  nand g122 (n_192, in_0[16], in_1[16]);
  nand g123 (n_193, in_2[16], in_1[16]);
  nand g124 (n_194, in_0[16], in_2[16]);
  nand g125 (out_0[17], n_192, n_193, n_194);
  xor g126 (n_195, in_0[17], in_1[17]);
  xor g127 (out_1[17], n_195, in_2[17]);
  nand g128 (n_196, in_0[17], in_1[17]);
  nand g129 (n_197, in_2[17], in_1[17]);
  nand g130 (n_198, in_0[17], in_2[17]);
  nand g131 (out_0[18], n_196, n_197, n_198);
  xor g132 (n_199, in_0[18], in_1[18]);
  xor g133 (out_1[18], n_199, in_2[18]);
  nand g134 (n_200, in_0[18], in_1[18]);
  nand g135 (n_201, in_2[18], in_1[18]);
  nand g136 (n_202, in_0[18], in_2[18]);
  nand g137 (out_0[19], n_200, n_201, n_202);
  xor g138 (n_203, in_0[19], in_1[19]);
  xor g139 (out_1[19], n_203, in_2[19]);
  nand g140 (n_204, in_0[19], in_1[19]);
  nand g141 (n_205, in_2[19], in_1[19]);
  nand g142 (n_206, in_0[19], in_2[19]);
  nand g143 (out_0[20], n_204, n_205, n_206);
  xor g144 (n_207, in_0[20], in_1[20]);
  xor g145 (out_1[20], n_207, in_2[20]);
  nand g146 (n_208, in_0[20], in_1[20]);
  nand g147 (n_209, in_2[20], in_1[20]);
  nand g148 (n_210, in_0[20], in_2[20]);
  nand g149 (out_0[21], n_208, n_209, n_210);
  xor g150 (n_70, in_0[21], in_1[21]);
  and g151 (n_75, in_0[21], in_1[21]);
  xor g153 (out_1[21], in_2[21], n_70);
  xor g158 (n_74, in_0[22], in_1[22]);
  and g159 (n_80, in_0[22], in_1[22]);
  nand g163 (n_217, n_75, n_74);
  nand g171 (n_221, n_80, n_79);
  or g174 (n_213, in_2[21], wc);
  not gc (wc, n_70);
  xor g178 (n_79, in_0[23], in_1[23]);
  nor g179 (out_0[24], in_0[23], in_1[23]);
  or g181 (out_0[22], wc0, wc1, n_70);
  not gc1 (wc1, n_213);
  not gc0 (wc0, in_2[21]);
  xnor g182 (out_1[22], n_75, n_74);
  or g183 (out_0[23], wc2, n_74, n_75);
  not gc2 (wc2, n_217);
  xnor g185 (out_1[23], n_80, n_79);
  or g186 (out_1[24], n_79, wc3, n_80);
  not gc3 (wc3, n_221);
endmodule

module csa_tree_3124_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [23:0] in_0, in_1;
  input [21:0] in_2;
  output [24:0] out_0, out_1;
  wire [23:0] in_0, in_1;
  wire [21:0] in_2;
  wire [24:0] out_0, out_1;
  csa_tree_3124_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_3152_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 26'b0;"
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  wire n_73, n_77, n_78, n_82, n_83, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_222, n_226, n_230;
  assign out_0[0] = in_1[0];
  xor g32 (out_1[0], in_0[0], in_2[0]);
  and g33 (out_0[1], in_0[0], in_2[0]);
  xor g34 (n_136, in_0[1], in_1[1]);
  xor g35 (out_1[1], n_136, in_2[1]);
  nand g36 (n_137, in_0[1], in_1[1]);
  nand g4 (n_138, in_2[1], in_1[1]);
  nand g5 (n_139, in_0[1], in_2[1]);
  nand g37 (out_0[2], n_137, n_138, n_139);
  xor g38 (n_140, in_0[2], in_1[2]);
  xor g39 (out_1[2], n_140, in_2[2]);
  nand g40 (n_141, in_0[2], in_1[2]);
  nand g41 (n_142, in_2[2], in_1[2]);
  nand g42 (n_143, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_141, n_142, n_143);
  xor g43 (n_144, in_0[3], in_1[3]);
  xor g44 (out_1[3], n_144, in_2[3]);
  nand g45 (n_145, in_0[3], in_1[3]);
  nand g46 (n_146, in_2[3], in_1[3]);
  nand g47 (n_147, in_0[3], in_2[3]);
  nand g48 (out_0[4], n_145, n_146, n_147);
  xor g49 (n_148, in_0[4], in_1[4]);
  xor g50 (out_1[4], n_148, in_2[4]);
  nand g51 (n_149, in_0[4], in_1[4]);
  nand g52 (n_150, in_2[4], in_1[4]);
  nand g53 (n_151, in_0[4], in_2[4]);
  nand g54 (out_0[5], n_149, n_150, n_151);
  xor g55 (n_152, in_0[5], in_1[5]);
  xor g56 (out_1[5], n_152, in_2[5]);
  nand g57 (n_153, in_0[5], in_1[5]);
  nand g58 (n_154, in_2[5], in_1[5]);
  nand g59 (n_155, in_0[5], in_2[5]);
  nand g60 (out_0[6], n_153, n_154, n_155);
  xor g61 (n_156, in_0[6], in_1[6]);
  xor g62 (out_1[6], n_156, in_2[6]);
  nand g63 (n_157, in_0[6], in_1[6]);
  nand g64 (n_158, in_2[6], in_1[6]);
  nand g65 (n_159, in_0[6], in_2[6]);
  nand g66 (out_0[7], n_157, n_158, n_159);
  xor g67 (n_160, in_0[7], in_1[7]);
  xor g68 (out_1[7], n_160, in_2[7]);
  nand g69 (n_161, in_0[7], in_1[7]);
  nand g70 (n_162, in_2[7], in_1[7]);
  nand g71 (n_163, in_0[7], in_2[7]);
  nand g72 (out_0[8], n_161, n_162, n_163);
  xor g73 (n_164, in_0[8], in_1[8]);
  xor g74 (out_1[8], n_164, in_2[8]);
  nand g75 (n_165, in_0[8], in_1[8]);
  nand g76 (n_166, in_2[8], in_1[8]);
  nand g77 (n_167, in_0[8], in_2[8]);
  nand g78 (out_0[9], n_165, n_166, n_167);
  xor g79 (n_168, in_0[9], in_1[9]);
  xor g80 (out_1[9], n_168, in_2[9]);
  nand g81 (n_169, in_0[9], in_1[9]);
  nand g82 (n_170, in_2[9], in_1[9]);
  nand g83 (n_171, in_0[9], in_2[9]);
  nand g84 (out_0[10], n_169, n_170, n_171);
  xor g85 (n_172, in_0[10], in_1[10]);
  xor g86 (out_1[10], n_172, in_2[10]);
  nand g87 (n_173, in_0[10], in_1[10]);
  nand g88 (n_174, in_2[10], in_1[10]);
  nand g89 (n_175, in_0[10], in_2[10]);
  nand g90 (out_0[11], n_173, n_174, n_175);
  xor g91 (n_176, in_0[11], in_1[11]);
  xor g92 (out_1[11], n_176, in_2[11]);
  nand g93 (n_177, in_0[11], in_1[11]);
  nand g94 (n_178, in_2[11], in_1[11]);
  nand g95 (n_179, in_0[11], in_2[11]);
  nand g96 (out_0[12], n_177, n_178, n_179);
  xor g97 (n_180, in_0[12], in_1[12]);
  xor g98 (out_1[12], n_180, in_2[12]);
  nand g99 (n_181, in_0[12], in_1[12]);
  nand g100 (n_182, in_2[12], in_1[12]);
  nand g101 (n_183, in_0[12], in_2[12]);
  nand g102 (out_0[13], n_181, n_182, n_183);
  xor g103 (n_184, in_0[13], in_1[13]);
  xor g104 (out_1[13], n_184, in_2[13]);
  nand g105 (n_185, in_0[13], in_1[13]);
  nand g106 (n_186, in_2[13], in_1[13]);
  nand g107 (n_187, in_0[13], in_2[13]);
  nand g108 (out_0[14], n_185, n_186, n_187);
  xor g109 (n_188, in_0[14], in_1[14]);
  xor g110 (out_1[14], n_188, in_2[14]);
  nand g111 (n_189, in_0[14], in_1[14]);
  nand g112 (n_190, in_2[14], in_1[14]);
  nand g113 (n_191, in_0[14], in_2[14]);
  nand g114 (out_0[15], n_189, n_190, n_191);
  xor g115 (n_192, in_0[15], in_1[15]);
  xor g116 (out_1[15], n_192, in_2[15]);
  nand g117 (n_193, in_0[15], in_1[15]);
  nand g118 (n_194, in_2[15], in_1[15]);
  nand g119 (n_195, in_0[15], in_2[15]);
  nand g120 (out_0[16], n_193, n_194, n_195);
  xor g121 (n_196, in_0[16], in_1[16]);
  xor g122 (out_1[16], n_196, in_2[16]);
  nand g123 (n_197, in_0[16], in_1[16]);
  nand g124 (n_198, in_2[16], in_1[16]);
  nand g125 (n_199, in_0[16], in_2[16]);
  nand g126 (out_0[17], n_197, n_198, n_199);
  xor g127 (n_200, in_0[17], in_1[17]);
  xor g128 (out_1[17], n_200, in_2[17]);
  nand g129 (n_201, in_0[17], in_1[17]);
  nand g130 (n_202, in_2[17], in_1[17]);
  nand g131 (n_203, in_0[17], in_2[17]);
  nand g132 (out_0[18], n_201, n_202, n_203);
  xor g133 (n_204, in_0[18], in_1[18]);
  xor g134 (out_1[18], n_204, in_2[18]);
  nand g135 (n_205, in_0[18], in_1[18]);
  nand g136 (n_206, in_2[18], in_1[18]);
  nand g137 (n_207, in_0[18], in_2[18]);
  nand g138 (out_0[19], n_205, n_206, n_207);
  xor g139 (n_208, in_0[19], in_1[19]);
  xor g140 (out_1[19], n_208, in_2[19]);
  nand g141 (n_209, in_0[19], in_1[19]);
  nand g142 (n_210, in_2[19], in_1[19]);
  nand g143 (n_211, in_0[19], in_2[19]);
  nand g144 (out_0[20], n_209, n_210, n_211);
  xor g145 (n_212, in_0[20], in_1[20]);
  xor g146 (out_1[20], n_212, in_2[20]);
  nand g147 (n_213, in_0[20], in_1[20]);
  nand g148 (n_214, in_2[20], in_1[20]);
  nand g149 (n_215, in_0[20], in_2[20]);
  nand g150 (out_0[21], n_213, n_214, n_215);
  xor g151 (n_216, in_0[21], in_1[21]);
  xor g152 (out_1[21], n_216, in_2[21]);
  nand g153 (n_217, in_0[21], in_1[21]);
  nand g154 (n_218, in_2[21], in_1[21]);
  nand g155 (n_219, in_0[21], in_2[21]);
  nand g156 (out_0[22], n_217, n_218, n_219);
  xor g157 (n_73, in_0[22], in_1[22]);
  and g158 (n_78, in_0[22], in_1[22]);
  xor g160 (out_1[22], in_2[22], n_73);
  xor g165 (n_77, in_0[23], in_1[23]);
  and g166 (n_83, in_0[23], in_1[23]);
  nand g170 (n_226, n_78, n_77);
  nand g178 (n_230, n_83, n_82);
  or g181 (n_222, in_2[22], wc);
  not gc (wc, n_73);
  xor g185 (n_82, in_0[24], in_1[24]);
  nor g186 (out_0[25], in_0[24], in_1[24]);
  or g188 (out_0[23], wc0, wc1, n_73);
  not gc1 (wc1, n_222);
  not gc0 (wc0, in_2[22]);
  xnor g189 (out_1[23], n_78, n_77);
  or g190 (out_0[24], wc2, n_77, n_78);
  not gc2 (wc2, n_226);
  xnor g192 (out_1[24], n_83, n_82);
  or g193 (out_1[25], n_82, wc3, n_83);
  not gc3 (wc3, n_230);
endmodule

module csa_tree_3152_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  csa_tree_3152_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_3152_1_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 26'b0;"
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  wire n_73, n_77, n_78, n_82, n_83, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_222, n_226, n_230;
  assign out_0[0] = in_1[0];
  xor g32 (out_1[0], in_0[0], in_2[0]);
  and g33 (out_0[1], in_0[0], in_2[0]);
  xor g34 (n_136, in_0[1], in_1[1]);
  xor g35 (out_1[1], n_136, in_2[1]);
  nand g36 (n_137, in_0[1], in_1[1]);
  nand g4 (n_138, in_2[1], in_1[1]);
  nand g5 (n_139, in_0[1], in_2[1]);
  nand g37 (out_0[2], n_137, n_138, n_139);
  xor g38 (n_140, in_0[2], in_1[2]);
  xor g39 (out_1[2], n_140, in_2[2]);
  nand g40 (n_141, in_0[2], in_1[2]);
  nand g41 (n_142, in_2[2], in_1[2]);
  nand g42 (n_143, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_141, n_142, n_143);
  xor g43 (n_144, in_0[3], in_1[3]);
  xor g44 (out_1[3], n_144, in_2[3]);
  nand g45 (n_145, in_0[3], in_1[3]);
  nand g46 (n_146, in_2[3], in_1[3]);
  nand g47 (n_147, in_0[3], in_2[3]);
  nand g48 (out_0[4], n_145, n_146, n_147);
  xor g49 (n_148, in_0[4], in_1[4]);
  xor g50 (out_1[4], n_148, in_2[4]);
  nand g51 (n_149, in_0[4], in_1[4]);
  nand g52 (n_150, in_2[4], in_1[4]);
  nand g53 (n_151, in_0[4], in_2[4]);
  nand g54 (out_0[5], n_149, n_150, n_151);
  xor g55 (n_152, in_0[5], in_1[5]);
  xor g56 (out_1[5], n_152, in_2[5]);
  nand g57 (n_153, in_0[5], in_1[5]);
  nand g58 (n_154, in_2[5], in_1[5]);
  nand g59 (n_155, in_0[5], in_2[5]);
  nand g60 (out_0[6], n_153, n_154, n_155);
  xor g61 (n_156, in_0[6], in_1[6]);
  xor g62 (out_1[6], n_156, in_2[6]);
  nand g63 (n_157, in_0[6], in_1[6]);
  nand g64 (n_158, in_2[6], in_1[6]);
  nand g65 (n_159, in_0[6], in_2[6]);
  nand g66 (out_0[7], n_157, n_158, n_159);
  xor g67 (n_160, in_0[7], in_1[7]);
  xor g68 (out_1[7], n_160, in_2[7]);
  nand g69 (n_161, in_0[7], in_1[7]);
  nand g70 (n_162, in_2[7], in_1[7]);
  nand g71 (n_163, in_0[7], in_2[7]);
  nand g72 (out_0[8], n_161, n_162, n_163);
  xor g73 (n_164, in_0[8], in_1[8]);
  xor g74 (out_1[8], n_164, in_2[8]);
  nand g75 (n_165, in_0[8], in_1[8]);
  nand g76 (n_166, in_2[8], in_1[8]);
  nand g77 (n_167, in_0[8], in_2[8]);
  nand g78 (out_0[9], n_165, n_166, n_167);
  xor g79 (n_168, in_0[9], in_1[9]);
  xor g80 (out_1[9], n_168, in_2[9]);
  nand g81 (n_169, in_0[9], in_1[9]);
  nand g82 (n_170, in_2[9], in_1[9]);
  nand g83 (n_171, in_0[9], in_2[9]);
  nand g84 (out_0[10], n_169, n_170, n_171);
  xor g85 (n_172, in_0[10], in_1[10]);
  xor g86 (out_1[10], n_172, in_2[10]);
  nand g87 (n_173, in_0[10], in_1[10]);
  nand g88 (n_174, in_2[10], in_1[10]);
  nand g89 (n_175, in_0[10], in_2[10]);
  nand g90 (out_0[11], n_173, n_174, n_175);
  xor g91 (n_176, in_0[11], in_1[11]);
  xor g92 (out_1[11], n_176, in_2[11]);
  nand g93 (n_177, in_0[11], in_1[11]);
  nand g94 (n_178, in_2[11], in_1[11]);
  nand g95 (n_179, in_0[11], in_2[11]);
  nand g96 (out_0[12], n_177, n_178, n_179);
  xor g97 (n_180, in_0[12], in_1[12]);
  xor g98 (out_1[12], n_180, in_2[12]);
  nand g99 (n_181, in_0[12], in_1[12]);
  nand g100 (n_182, in_2[12], in_1[12]);
  nand g101 (n_183, in_0[12], in_2[12]);
  nand g102 (out_0[13], n_181, n_182, n_183);
  xor g103 (n_184, in_0[13], in_1[13]);
  xor g104 (out_1[13], n_184, in_2[13]);
  nand g105 (n_185, in_0[13], in_1[13]);
  nand g106 (n_186, in_2[13], in_1[13]);
  nand g107 (n_187, in_0[13], in_2[13]);
  nand g108 (out_0[14], n_185, n_186, n_187);
  xor g109 (n_188, in_0[14], in_1[14]);
  xor g110 (out_1[14], n_188, in_2[14]);
  nand g111 (n_189, in_0[14], in_1[14]);
  nand g112 (n_190, in_2[14], in_1[14]);
  nand g113 (n_191, in_0[14], in_2[14]);
  nand g114 (out_0[15], n_189, n_190, n_191);
  xor g115 (n_192, in_0[15], in_1[15]);
  xor g116 (out_1[15], n_192, in_2[15]);
  nand g117 (n_193, in_0[15], in_1[15]);
  nand g118 (n_194, in_2[15], in_1[15]);
  nand g119 (n_195, in_0[15], in_2[15]);
  nand g120 (out_0[16], n_193, n_194, n_195);
  xor g121 (n_196, in_0[16], in_1[16]);
  xor g122 (out_1[16], n_196, in_2[16]);
  nand g123 (n_197, in_0[16], in_1[16]);
  nand g124 (n_198, in_2[16], in_1[16]);
  nand g125 (n_199, in_0[16], in_2[16]);
  nand g126 (out_0[17], n_197, n_198, n_199);
  xor g127 (n_200, in_0[17], in_1[17]);
  xor g128 (out_1[17], n_200, in_2[17]);
  nand g129 (n_201, in_0[17], in_1[17]);
  nand g130 (n_202, in_2[17], in_1[17]);
  nand g131 (n_203, in_0[17], in_2[17]);
  nand g132 (out_0[18], n_201, n_202, n_203);
  xor g133 (n_204, in_0[18], in_1[18]);
  xor g134 (out_1[18], n_204, in_2[18]);
  nand g135 (n_205, in_0[18], in_1[18]);
  nand g136 (n_206, in_2[18], in_1[18]);
  nand g137 (n_207, in_0[18], in_2[18]);
  nand g138 (out_0[19], n_205, n_206, n_207);
  xor g139 (n_208, in_0[19], in_1[19]);
  xor g140 (out_1[19], n_208, in_2[19]);
  nand g141 (n_209, in_0[19], in_1[19]);
  nand g142 (n_210, in_2[19], in_1[19]);
  nand g143 (n_211, in_0[19], in_2[19]);
  nand g144 (out_0[20], n_209, n_210, n_211);
  xor g145 (n_212, in_0[20], in_1[20]);
  xor g146 (out_1[20], n_212, in_2[20]);
  nand g147 (n_213, in_0[20], in_1[20]);
  nand g148 (n_214, in_2[20], in_1[20]);
  nand g149 (n_215, in_0[20], in_2[20]);
  nand g150 (out_0[21], n_213, n_214, n_215);
  xor g151 (n_216, in_0[21], in_1[21]);
  xor g152 (out_1[21], n_216, in_2[21]);
  nand g153 (n_217, in_0[21], in_1[21]);
  nand g154 (n_218, in_2[21], in_1[21]);
  nand g155 (n_219, in_0[21], in_2[21]);
  nand g156 (out_0[22], n_217, n_218, n_219);
  xor g157 (n_73, in_0[22], in_1[22]);
  and g158 (n_78, in_0[22], in_1[22]);
  xor g160 (out_1[22], in_2[22], n_73);
  xor g165 (n_77, in_0[23], in_1[23]);
  and g166 (n_83, in_0[23], in_1[23]);
  nand g170 (n_226, n_78, n_77);
  nand g178 (n_230, n_83, n_82);
  or g181 (n_222, in_2[22], wc);
  not gc (wc, n_73);
  xor g185 (n_82, in_0[24], in_1[24]);
  nor g186 (out_0[25], in_0[24], in_1[24]);
  or g188 (out_0[23], wc0, wc1, n_73);
  not gc1 (wc1, n_222);
  not gc0 (wc0, in_2[22]);
  xnor g189 (out_1[23], n_78, n_77);
  or g190 (out_0[24], wc2, n_77, n_78);
  not gc2 (wc2, n_226);
  xnor g192 (out_1[24], n_83, n_82);
  or g193 (out_1[25], n_82, wc3, n_83);
  not gc3 (wc3, n_230);
endmodule

module csa_tree_3152_1_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  csa_tree_3152_1_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_3152_2_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 26'b0;"
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  wire n_73, n_77, n_78, n_82, n_83, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162;
  wire n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170;
  wire n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178;
  wire n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_222, n_226, n_230;
  assign out_0[0] = in_1[0];
  xor g32 (out_1[0], in_0[0], in_2[0]);
  and g33 (out_0[1], in_0[0], in_2[0]);
  xor g34 (n_136, in_0[1], in_1[1]);
  xor g35 (out_1[1], n_136, in_2[1]);
  nand g36 (n_137, in_0[1], in_1[1]);
  nand g4 (n_138, in_2[1], in_1[1]);
  nand g5 (n_139, in_0[1], in_2[1]);
  nand g37 (out_0[2], n_137, n_138, n_139);
  xor g38 (n_140, in_0[2], in_1[2]);
  xor g39 (out_1[2], n_140, in_2[2]);
  nand g40 (n_141, in_0[2], in_1[2]);
  nand g41 (n_142, in_2[2], in_1[2]);
  nand g42 (n_143, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_141, n_142, n_143);
  xor g43 (n_144, in_0[3], in_1[3]);
  xor g44 (out_1[3], n_144, in_2[3]);
  nand g45 (n_145, in_0[3], in_1[3]);
  nand g46 (n_146, in_2[3], in_1[3]);
  nand g47 (n_147, in_0[3], in_2[3]);
  nand g48 (out_0[4], n_145, n_146, n_147);
  xor g49 (n_148, in_0[4], in_1[4]);
  xor g50 (out_1[4], n_148, in_2[4]);
  nand g51 (n_149, in_0[4], in_1[4]);
  nand g52 (n_150, in_2[4], in_1[4]);
  nand g53 (n_151, in_0[4], in_2[4]);
  nand g54 (out_0[5], n_149, n_150, n_151);
  xor g55 (n_152, in_0[5], in_1[5]);
  xor g56 (out_1[5], n_152, in_2[5]);
  nand g57 (n_153, in_0[5], in_1[5]);
  nand g58 (n_154, in_2[5], in_1[5]);
  nand g59 (n_155, in_0[5], in_2[5]);
  nand g60 (out_0[6], n_153, n_154, n_155);
  xor g61 (n_156, in_0[6], in_1[6]);
  xor g62 (out_1[6], n_156, in_2[6]);
  nand g63 (n_157, in_0[6], in_1[6]);
  nand g64 (n_158, in_2[6], in_1[6]);
  nand g65 (n_159, in_0[6], in_2[6]);
  nand g66 (out_0[7], n_157, n_158, n_159);
  xor g67 (n_160, in_0[7], in_1[7]);
  xor g68 (out_1[7], n_160, in_2[7]);
  nand g69 (n_161, in_0[7], in_1[7]);
  nand g70 (n_162, in_2[7], in_1[7]);
  nand g71 (n_163, in_0[7], in_2[7]);
  nand g72 (out_0[8], n_161, n_162, n_163);
  xor g73 (n_164, in_0[8], in_1[8]);
  xor g74 (out_1[8], n_164, in_2[8]);
  nand g75 (n_165, in_0[8], in_1[8]);
  nand g76 (n_166, in_2[8], in_1[8]);
  nand g77 (n_167, in_0[8], in_2[8]);
  nand g78 (out_0[9], n_165, n_166, n_167);
  xor g79 (n_168, in_0[9], in_1[9]);
  xor g80 (out_1[9], n_168, in_2[9]);
  nand g81 (n_169, in_0[9], in_1[9]);
  nand g82 (n_170, in_2[9], in_1[9]);
  nand g83 (n_171, in_0[9], in_2[9]);
  nand g84 (out_0[10], n_169, n_170, n_171);
  xor g85 (n_172, in_0[10], in_1[10]);
  xor g86 (out_1[10], n_172, in_2[10]);
  nand g87 (n_173, in_0[10], in_1[10]);
  nand g88 (n_174, in_2[10], in_1[10]);
  nand g89 (n_175, in_0[10], in_2[10]);
  nand g90 (out_0[11], n_173, n_174, n_175);
  xor g91 (n_176, in_0[11], in_1[11]);
  xor g92 (out_1[11], n_176, in_2[11]);
  nand g93 (n_177, in_0[11], in_1[11]);
  nand g94 (n_178, in_2[11], in_1[11]);
  nand g95 (n_179, in_0[11], in_2[11]);
  nand g96 (out_0[12], n_177, n_178, n_179);
  xor g97 (n_180, in_0[12], in_1[12]);
  xor g98 (out_1[12], n_180, in_2[12]);
  nand g99 (n_181, in_0[12], in_1[12]);
  nand g100 (n_182, in_2[12], in_1[12]);
  nand g101 (n_183, in_0[12], in_2[12]);
  nand g102 (out_0[13], n_181, n_182, n_183);
  xor g103 (n_184, in_0[13], in_1[13]);
  xor g104 (out_1[13], n_184, in_2[13]);
  nand g105 (n_185, in_0[13], in_1[13]);
  nand g106 (n_186, in_2[13], in_1[13]);
  nand g107 (n_187, in_0[13], in_2[13]);
  nand g108 (out_0[14], n_185, n_186, n_187);
  xor g109 (n_188, in_0[14], in_1[14]);
  xor g110 (out_1[14], n_188, in_2[14]);
  nand g111 (n_189, in_0[14], in_1[14]);
  nand g112 (n_190, in_2[14], in_1[14]);
  nand g113 (n_191, in_0[14], in_2[14]);
  nand g114 (out_0[15], n_189, n_190, n_191);
  xor g115 (n_192, in_0[15], in_1[15]);
  xor g116 (out_1[15], n_192, in_2[15]);
  nand g117 (n_193, in_0[15], in_1[15]);
  nand g118 (n_194, in_2[15], in_1[15]);
  nand g119 (n_195, in_0[15], in_2[15]);
  nand g120 (out_0[16], n_193, n_194, n_195);
  xor g121 (n_196, in_0[16], in_1[16]);
  xor g122 (out_1[16], n_196, in_2[16]);
  nand g123 (n_197, in_0[16], in_1[16]);
  nand g124 (n_198, in_2[16], in_1[16]);
  nand g125 (n_199, in_0[16], in_2[16]);
  nand g126 (out_0[17], n_197, n_198, n_199);
  xor g127 (n_200, in_0[17], in_1[17]);
  xor g128 (out_1[17], n_200, in_2[17]);
  nand g129 (n_201, in_0[17], in_1[17]);
  nand g130 (n_202, in_2[17], in_1[17]);
  nand g131 (n_203, in_0[17], in_2[17]);
  nand g132 (out_0[18], n_201, n_202, n_203);
  xor g133 (n_204, in_0[18], in_1[18]);
  xor g134 (out_1[18], n_204, in_2[18]);
  nand g135 (n_205, in_0[18], in_1[18]);
  nand g136 (n_206, in_2[18], in_1[18]);
  nand g137 (n_207, in_0[18], in_2[18]);
  nand g138 (out_0[19], n_205, n_206, n_207);
  xor g139 (n_208, in_0[19], in_1[19]);
  xor g140 (out_1[19], n_208, in_2[19]);
  nand g141 (n_209, in_0[19], in_1[19]);
  nand g142 (n_210, in_2[19], in_1[19]);
  nand g143 (n_211, in_0[19], in_2[19]);
  nand g144 (out_0[20], n_209, n_210, n_211);
  xor g145 (n_212, in_0[20], in_1[20]);
  xor g146 (out_1[20], n_212, in_2[20]);
  nand g147 (n_213, in_0[20], in_1[20]);
  nand g148 (n_214, in_2[20], in_1[20]);
  nand g149 (n_215, in_0[20], in_2[20]);
  nand g150 (out_0[21], n_213, n_214, n_215);
  xor g151 (n_216, in_0[21], in_1[21]);
  xor g152 (out_1[21], n_216, in_2[21]);
  nand g153 (n_217, in_0[21], in_1[21]);
  nand g154 (n_218, in_2[21], in_1[21]);
  nand g155 (n_219, in_0[21], in_2[21]);
  nand g156 (out_0[22], n_217, n_218, n_219);
  xor g157 (n_73, in_0[22], in_1[22]);
  and g158 (n_78, in_0[22], in_1[22]);
  xor g160 (out_1[22], in_2[22], n_73);
  xor g165 (n_77, in_0[23], in_1[23]);
  and g166 (n_83, in_0[23], in_1[23]);
  nand g170 (n_226, n_78, n_77);
  nand g178 (n_230, n_83, n_82);
  or g181 (n_222, in_2[22], wc);
  not gc (wc, n_73);
  xor g185 (n_82, in_0[24], in_1[24]);
  nor g186 (out_0[25], in_0[24], in_1[24]);
  or g188 (out_0[23], wc0, wc1, n_73);
  not gc1 (wc1, n_222);
  not gc0 (wc0, in_2[22]);
  xnor g189 (out_1[23], n_78, n_77);
  or g190 (out_0[24], wc2, n_77, n_78);
  not gc2 (wc2, n_226);
  xnor g192 (out_1[24], n_83, n_82);
  or g193 (out_1[25], n_82, wc3, n_83);
  not gc3 (wc3, n_230);
endmodule

module csa_tree_3152_2_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [24:0] in_0, in_1;
  input [22:0] in_2;
  output [25:0] out_0, out_1;
  wire [24:0] in_0, in_1;
  wire [22:0] in_2;
  wire [25:0] out_0, out_1;
  csa_tree_3152_2_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_3210_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 25'b0;"
  input [21:0] in_0, in_1, in_2;
  output [24:0] out_0, out_1;
  wire [21:0] in_0, in_1, in_2;
  wire [24:0] out_0, out_1;
  wire n_70, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_203;
  assign out_1[23] = 1'b0;
  assign out_1[24] = 1'b0;
  assign out_0[0] = in_1[0];
  assign out_0[23] = 1'b1;
  assign out_0[24] = 1'b1;
  xor g27 (out_1[0], in_0[0], in_2[0]);
  and g28 (out_0[1], in_0[0], in_2[0]);
  xor g29 (n_121, in_0[1], in_1[1]);
  xor g30 (out_1[1], n_121, in_2[1]);
  nand g31 (n_122, in_0[1], in_1[1]);
  nand g4 (n_123, in_2[1], in_1[1]);
  nand g5 (n_124, in_0[1], in_2[1]);
  nand g32 (out_0[2], n_122, n_123, n_124);
  xor g33 (n_125, in_0[2], in_1[2]);
  xor g34 (out_1[2], n_125, in_2[2]);
  nand g35 (n_126, in_0[2], in_1[2]);
  nand g36 (n_127, in_2[2], in_1[2]);
  nand g37 (n_128, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_126, n_127, n_128);
  xor g38 (n_129, in_0[3], in_1[3]);
  xor g39 (out_1[3], n_129, in_2[3]);
  nand g40 (n_130, in_0[3], in_1[3]);
  nand g41 (n_131, in_2[3], in_1[3]);
  nand g42 (n_132, in_0[3], in_2[3]);
  nand g43 (out_0[4], n_130, n_131, n_132);
  xor g44 (n_133, in_0[4], in_1[4]);
  xor g45 (out_1[4], n_133, in_2[4]);
  nand g46 (n_134, in_0[4], in_1[4]);
  nand g47 (n_135, in_2[4], in_1[4]);
  nand g48 (n_136, in_0[4], in_2[4]);
  nand g49 (out_0[5], n_134, n_135, n_136);
  xor g50 (n_137, in_0[5], in_1[5]);
  xor g51 (out_1[5], n_137, in_2[5]);
  nand g52 (n_138, in_0[5], in_1[5]);
  nand g53 (n_139, in_2[5], in_1[5]);
  nand g54 (n_140, in_0[5], in_2[5]);
  nand g55 (out_0[6], n_138, n_139, n_140);
  xor g56 (n_141, in_0[6], in_1[6]);
  xor g57 (out_1[6], n_141, in_2[6]);
  nand g58 (n_142, in_0[6], in_1[6]);
  nand g59 (n_143, in_2[6], in_1[6]);
  nand g60 (n_144, in_0[6], in_2[6]);
  nand g61 (out_0[7], n_142, n_143, n_144);
  xor g62 (n_145, in_0[7], in_1[7]);
  xor g63 (out_1[7], n_145, in_2[7]);
  nand g64 (n_146, in_0[7], in_1[7]);
  nand g65 (n_147, in_2[7], in_1[7]);
  nand g66 (n_148, in_0[7], in_2[7]);
  nand g67 (out_0[8], n_146, n_147, n_148);
  xor g68 (n_149, in_0[8], in_1[8]);
  xor g69 (out_1[8], n_149, in_2[8]);
  nand g70 (n_150, in_0[8], in_1[8]);
  nand g71 (n_151, in_2[8], in_1[8]);
  nand g72 (n_152, in_0[8], in_2[8]);
  nand g73 (out_0[9], n_150, n_151, n_152);
  xor g74 (n_153, in_0[9], in_1[9]);
  xor g75 (out_1[9], n_153, in_2[9]);
  nand g76 (n_154, in_0[9], in_1[9]);
  nand g77 (n_155, in_2[9], in_1[9]);
  nand g78 (n_156, in_0[9], in_2[9]);
  nand g79 (out_0[10], n_154, n_155, n_156);
  xor g80 (n_157, in_0[10], in_1[10]);
  xor g81 (out_1[10], n_157, in_2[10]);
  nand g82 (n_158, in_0[10], in_1[10]);
  nand g83 (n_159, in_2[10], in_1[10]);
  nand g84 (n_160, in_0[10], in_2[10]);
  nand g85 (out_0[11], n_158, n_159, n_160);
  xor g86 (n_161, in_0[11], in_1[11]);
  xor g87 (out_1[11], n_161, in_2[11]);
  nand g88 (n_162, in_0[11], in_1[11]);
  nand g89 (n_163, in_2[11], in_1[11]);
  nand g90 (n_164, in_0[11], in_2[11]);
  nand g91 (out_0[12], n_162, n_163, n_164);
  xor g92 (n_165, in_0[12], in_1[12]);
  xor g93 (out_1[12], n_165, in_2[12]);
  nand g94 (n_166, in_0[12], in_1[12]);
  nand g95 (n_167, in_2[12], in_1[12]);
  nand g96 (n_168, in_0[12], in_2[12]);
  nand g97 (out_0[13], n_166, n_167, n_168);
  xor g98 (n_169, in_0[13], in_1[13]);
  xor g99 (out_1[13], n_169, in_2[13]);
  nand g100 (n_170, in_0[13], in_1[13]);
  nand g101 (n_171, in_2[13], in_1[13]);
  nand g102 (n_172, in_0[13], in_2[13]);
  nand g103 (out_0[14], n_170, n_171, n_172);
  xor g104 (n_173, in_0[14], in_1[14]);
  xor g105 (out_1[14], n_173, in_2[14]);
  nand g106 (n_174, in_0[14], in_1[14]);
  nand g107 (n_175, in_2[14], in_1[14]);
  nand g108 (n_176, in_0[14], in_2[14]);
  nand g109 (out_0[15], n_174, n_175, n_176);
  xor g110 (n_177, in_0[15], in_1[15]);
  xor g111 (out_1[15], n_177, in_2[15]);
  nand g112 (n_178, in_0[15], in_1[15]);
  nand g113 (n_179, in_2[15], in_1[15]);
  nand g114 (n_180, in_0[15], in_2[15]);
  nand g115 (out_0[16], n_178, n_179, n_180);
  xor g116 (n_181, in_0[16], in_1[16]);
  xor g117 (out_1[16], n_181, in_2[16]);
  nand g118 (n_182, in_0[16], in_1[16]);
  nand g119 (n_183, in_2[16], in_1[16]);
  nand g120 (n_184, in_0[16], in_2[16]);
  nand g121 (out_0[17], n_182, n_183, n_184);
  xor g122 (n_185, in_0[17], in_1[17]);
  xor g123 (out_1[17], n_185, in_2[17]);
  nand g124 (n_186, in_0[17], in_1[17]);
  nand g125 (n_187, in_2[17], in_1[17]);
  nand g126 (n_188, in_0[17], in_2[17]);
  nand g127 (out_0[18], n_186, n_187, n_188);
  xor g128 (n_189, in_0[18], in_1[18]);
  xor g129 (out_1[18], n_189, in_2[18]);
  nand g130 (n_190, in_0[18], in_1[18]);
  nand g131 (n_191, in_2[18], in_1[18]);
  nand g132 (n_192, in_0[18], in_2[18]);
  nand g133 (out_0[19], n_190, n_191, n_192);
  xor g134 (n_193, in_0[19], in_1[19]);
  xor g135 (out_1[19], n_193, in_2[19]);
  nand g136 (n_194, in_0[19], in_1[19]);
  nand g137 (n_195, in_2[19], in_1[19]);
  nand g138 (n_196, in_0[19], in_2[19]);
  nand g139 (out_0[20], n_194, n_195, n_196);
  xor g140 (n_197, in_0[20], in_1[20]);
  xor g141 (out_1[20], n_197, in_2[20]);
  nand g142 (n_198, in_0[20], in_1[20]);
  nand g143 (n_199, in_2[20], in_1[20]);
  nand g144 (n_200, in_0[20], in_2[20]);
  nand g145 (out_0[21], n_198, n_199, n_200);
  xor g149 (out_1[21], in_2[21], n_70);
  xor g154 (n_70, in_0[21], in_1[21]);
  nor g155 (out_0[22], in_0[21], in_1[21]);
  or g156 (n_203, in_2[21], wc);
  not gc (wc, n_70);
  or g158 (out_1[22], wc0, wc1, n_70);
  not gc1 (wc1, n_203);
  not gc0 (wc0, in_2[21]);
endmodule

module csa_tree_3210_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [21:0] in_0, in_1, in_2;
  output [24:0] out_0, out_1;
  wire [21:0] in_0, in_1, in_2;
  wire [24:0] out_0, out_1;
  csa_tree_3210_GENERIC_REAL g1(.in_0 ({in_0[20], in_0[20:0]}), .in_1
       ({in_1[20], in_1[20:0]}), .in_2 (in_2), .out_0 (out_0), .out_1
       (out_1));
endmodule

module csa_tree_3210_1_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 25'b0;"
  input [21:0] in_0, in_1, in_2;
  output [24:0] out_0, out_1;
  wire [21:0] in_0, in_1, in_2;
  wire [24:0] out_0, out_1;
  wire n_70, n_121, n_122, n_123, n_124, n_125, n_126, n_127;
  wire n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135;
  wire n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_203;
  assign out_1[23] = 1'b0;
  assign out_1[24] = 1'b0;
  assign out_0[0] = in_1[0];
  assign out_0[23] = 1'b1;
  assign out_0[24] = 1'b1;
  xor g27 (out_1[0], in_0[0], in_2[0]);
  and g28 (out_0[1], in_0[0], in_2[0]);
  xor g29 (n_121, in_0[1], in_1[1]);
  xor g30 (out_1[1], n_121, in_2[1]);
  nand g31 (n_122, in_0[1], in_1[1]);
  nand g4 (n_123, in_2[1], in_1[1]);
  nand g5 (n_124, in_0[1], in_2[1]);
  nand g32 (out_0[2], n_122, n_123, n_124);
  xor g33 (n_125, in_0[2], in_1[2]);
  xor g34 (out_1[2], n_125, in_2[2]);
  nand g35 (n_126, in_0[2], in_1[2]);
  nand g36 (n_127, in_2[2], in_1[2]);
  nand g37 (n_128, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_126, n_127, n_128);
  xor g38 (n_129, in_0[3], in_1[3]);
  xor g39 (out_1[3], n_129, in_2[3]);
  nand g40 (n_130, in_0[3], in_1[3]);
  nand g41 (n_131, in_2[3], in_1[3]);
  nand g42 (n_132, in_0[3], in_2[3]);
  nand g43 (out_0[4], n_130, n_131, n_132);
  xor g44 (n_133, in_0[4], in_1[4]);
  xor g45 (out_1[4], n_133, in_2[4]);
  nand g46 (n_134, in_0[4], in_1[4]);
  nand g47 (n_135, in_2[4], in_1[4]);
  nand g48 (n_136, in_0[4], in_2[4]);
  nand g49 (out_0[5], n_134, n_135, n_136);
  xor g50 (n_137, in_0[5], in_1[5]);
  xor g51 (out_1[5], n_137, in_2[5]);
  nand g52 (n_138, in_0[5], in_1[5]);
  nand g53 (n_139, in_2[5], in_1[5]);
  nand g54 (n_140, in_0[5], in_2[5]);
  nand g55 (out_0[6], n_138, n_139, n_140);
  xor g56 (n_141, in_0[6], in_1[6]);
  xor g57 (out_1[6], n_141, in_2[6]);
  nand g58 (n_142, in_0[6], in_1[6]);
  nand g59 (n_143, in_2[6], in_1[6]);
  nand g60 (n_144, in_0[6], in_2[6]);
  nand g61 (out_0[7], n_142, n_143, n_144);
  xor g62 (n_145, in_0[7], in_1[7]);
  xor g63 (out_1[7], n_145, in_2[7]);
  nand g64 (n_146, in_0[7], in_1[7]);
  nand g65 (n_147, in_2[7], in_1[7]);
  nand g66 (n_148, in_0[7], in_2[7]);
  nand g67 (out_0[8], n_146, n_147, n_148);
  xor g68 (n_149, in_0[8], in_1[8]);
  xor g69 (out_1[8], n_149, in_2[8]);
  nand g70 (n_150, in_0[8], in_1[8]);
  nand g71 (n_151, in_2[8], in_1[8]);
  nand g72 (n_152, in_0[8], in_2[8]);
  nand g73 (out_0[9], n_150, n_151, n_152);
  xor g74 (n_153, in_0[9], in_1[9]);
  xor g75 (out_1[9], n_153, in_2[9]);
  nand g76 (n_154, in_0[9], in_1[9]);
  nand g77 (n_155, in_2[9], in_1[9]);
  nand g78 (n_156, in_0[9], in_2[9]);
  nand g79 (out_0[10], n_154, n_155, n_156);
  xor g80 (n_157, in_0[10], in_1[10]);
  xor g81 (out_1[10], n_157, in_2[10]);
  nand g82 (n_158, in_0[10], in_1[10]);
  nand g83 (n_159, in_2[10], in_1[10]);
  nand g84 (n_160, in_0[10], in_2[10]);
  nand g85 (out_0[11], n_158, n_159, n_160);
  xor g86 (n_161, in_0[11], in_1[11]);
  xor g87 (out_1[11], n_161, in_2[11]);
  nand g88 (n_162, in_0[11], in_1[11]);
  nand g89 (n_163, in_2[11], in_1[11]);
  nand g90 (n_164, in_0[11], in_2[11]);
  nand g91 (out_0[12], n_162, n_163, n_164);
  xor g92 (n_165, in_0[12], in_1[12]);
  xor g93 (out_1[12], n_165, in_2[12]);
  nand g94 (n_166, in_0[12], in_1[12]);
  nand g95 (n_167, in_2[12], in_1[12]);
  nand g96 (n_168, in_0[12], in_2[12]);
  nand g97 (out_0[13], n_166, n_167, n_168);
  xor g98 (n_169, in_0[13], in_1[13]);
  xor g99 (out_1[13], n_169, in_2[13]);
  nand g100 (n_170, in_0[13], in_1[13]);
  nand g101 (n_171, in_2[13], in_1[13]);
  nand g102 (n_172, in_0[13], in_2[13]);
  nand g103 (out_0[14], n_170, n_171, n_172);
  xor g104 (n_173, in_0[14], in_1[14]);
  xor g105 (out_1[14], n_173, in_2[14]);
  nand g106 (n_174, in_0[14], in_1[14]);
  nand g107 (n_175, in_2[14], in_1[14]);
  nand g108 (n_176, in_0[14], in_2[14]);
  nand g109 (out_0[15], n_174, n_175, n_176);
  xor g110 (n_177, in_0[15], in_1[15]);
  xor g111 (out_1[15], n_177, in_2[15]);
  nand g112 (n_178, in_0[15], in_1[15]);
  nand g113 (n_179, in_2[15], in_1[15]);
  nand g114 (n_180, in_0[15], in_2[15]);
  nand g115 (out_0[16], n_178, n_179, n_180);
  xor g116 (n_181, in_0[16], in_1[16]);
  xor g117 (out_1[16], n_181, in_2[16]);
  nand g118 (n_182, in_0[16], in_1[16]);
  nand g119 (n_183, in_2[16], in_1[16]);
  nand g120 (n_184, in_0[16], in_2[16]);
  nand g121 (out_0[17], n_182, n_183, n_184);
  xor g122 (n_185, in_0[17], in_1[17]);
  xor g123 (out_1[17], n_185, in_2[17]);
  nand g124 (n_186, in_0[17], in_1[17]);
  nand g125 (n_187, in_2[17], in_1[17]);
  nand g126 (n_188, in_0[17], in_2[17]);
  nand g127 (out_0[18], n_186, n_187, n_188);
  xor g128 (n_189, in_0[18], in_1[18]);
  xor g129 (out_1[18], n_189, in_2[18]);
  nand g130 (n_190, in_0[18], in_1[18]);
  nand g131 (n_191, in_2[18], in_1[18]);
  nand g132 (n_192, in_0[18], in_2[18]);
  nand g133 (out_0[19], n_190, n_191, n_192);
  xor g134 (n_193, in_0[19], in_1[19]);
  xor g135 (out_1[19], n_193, in_2[19]);
  nand g136 (n_194, in_0[19], in_1[19]);
  nand g137 (n_195, in_2[19], in_1[19]);
  nand g138 (n_196, in_0[19], in_2[19]);
  nand g139 (out_0[20], n_194, n_195, n_196);
  xor g140 (n_197, in_0[20], in_1[20]);
  xor g141 (out_1[20], n_197, in_2[20]);
  nand g142 (n_198, in_0[20], in_1[20]);
  nand g143 (n_199, in_2[20], in_1[20]);
  nand g144 (n_200, in_0[20], in_2[20]);
  nand g145 (out_0[21], n_198, n_199, n_200);
  xor g149 (out_1[21], in_2[21], n_70);
  xor g154 (n_70, in_0[21], in_1[21]);
  nor g155 (out_0[22], in_0[21], in_1[21]);
  or g156 (n_203, in_2[21], wc);
  not gc (wc, n_70);
  or g158 (out_1[22], wc0, wc1, n_70);
  not gc1 (wc1, n_203);
  not gc0 (wc0, in_2[21]);
endmodule

module csa_tree_3210_1_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [21:0] in_0, in_1, in_2;
  output [24:0] out_0, out_1;
  wire [21:0] in_0, in_1, in_2;
  wire [24:0] out_0, out_1;
  csa_tree_3210_1_GENERIC_REAL g1(.in_0 ({in_0[20], in_0[20:0]}), .in_1
       ({in_1[20], in_1[20:0]}), .in_2 (in_2), .out_0 (out_0), .out_1
       (out_1));
endmodule

module csa_tree_6719_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 26'b0;"
  input [22:0] in_0, in_1, in_2;
  output [25:0] out_0, out_1;
  wire [22:0] in_0, in_1, in_2;
  wire [25:0] out_0, out_1;
  wire n_73, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196;
  wire n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204;
  wire n_205, n_206, n_207, n_208, n_209, n_212;
  assign out_1[24] = 1'b0;
  assign out_1[25] = 1'b0;
  assign out_0[0] = in_1[0];
  assign out_0[24] = 1'b1;
  assign out_0[25] = 1'b1;
  xor g28 (out_1[0], in_0[0], in_2[0]);
  and g29 (out_0[1], in_0[0], in_2[0]);
  xor g30 (n_126, in_0[1], in_1[1]);
  xor g31 (out_1[1], n_126, in_2[1]);
  nand g32 (n_127, in_0[1], in_1[1]);
  nand g4 (n_128, in_2[1], in_1[1]);
  nand g5 (n_129, in_0[1], in_2[1]);
  nand g33 (out_0[2], n_127, n_128, n_129);
  xor g34 (n_130, in_0[2], in_1[2]);
  xor g35 (out_1[2], n_130, in_2[2]);
  nand g36 (n_131, in_0[2], in_1[2]);
  nand g37 (n_132, in_2[2], in_1[2]);
  nand g38 (n_133, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_131, n_132, n_133);
  xor g39 (n_134, in_0[3], in_1[3]);
  xor g40 (out_1[3], n_134, in_2[3]);
  nand g41 (n_135, in_0[3], in_1[3]);
  nand g42 (n_136, in_2[3], in_1[3]);
  nand g43 (n_137, in_0[3], in_2[3]);
  nand g44 (out_0[4], n_135, n_136, n_137);
  xor g45 (n_138, in_0[4], in_1[4]);
  xor g46 (out_1[4], n_138, in_2[4]);
  nand g47 (n_139, in_0[4], in_1[4]);
  nand g48 (n_140, in_2[4], in_1[4]);
  nand g49 (n_141, in_0[4], in_2[4]);
  nand g50 (out_0[5], n_139, n_140, n_141);
  xor g51 (n_142, in_0[5], in_1[5]);
  xor g52 (out_1[5], n_142, in_2[5]);
  nand g53 (n_143, in_0[5], in_1[5]);
  nand g54 (n_144, in_2[5], in_1[5]);
  nand g55 (n_145, in_0[5], in_2[5]);
  nand g56 (out_0[6], n_143, n_144, n_145);
  xor g57 (n_146, in_0[6], in_1[6]);
  xor g58 (out_1[6], n_146, in_2[6]);
  nand g59 (n_147, in_0[6], in_1[6]);
  nand g60 (n_148, in_2[6], in_1[6]);
  nand g61 (n_149, in_0[6], in_2[6]);
  nand g62 (out_0[7], n_147, n_148, n_149);
  xor g63 (n_150, in_0[7], in_1[7]);
  xor g64 (out_1[7], n_150, in_2[7]);
  nand g65 (n_151, in_0[7], in_1[7]);
  nand g66 (n_152, in_2[7], in_1[7]);
  nand g67 (n_153, in_0[7], in_2[7]);
  nand g68 (out_0[8], n_151, n_152, n_153);
  xor g69 (n_154, in_0[8], in_1[8]);
  xor g70 (out_1[8], n_154, in_2[8]);
  nand g71 (n_155, in_0[8], in_1[8]);
  nand g72 (n_156, in_2[8], in_1[8]);
  nand g73 (n_157, in_0[8], in_2[8]);
  nand g74 (out_0[9], n_155, n_156, n_157);
  xor g75 (n_158, in_0[9], in_1[9]);
  xor g76 (out_1[9], n_158, in_2[9]);
  nand g77 (n_159, in_0[9], in_1[9]);
  nand g78 (n_160, in_2[9], in_1[9]);
  nand g79 (n_161, in_0[9], in_2[9]);
  nand g80 (out_0[10], n_159, n_160, n_161);
  xor g81 (n_162, in_0[10], in_1[10]);
  xor g82 (out_1[10], n_162, in_2[10]);
  nand g83 (n_163, in_0[10], in_1[10]);
  nand g84 (n_164, in_2[10], in_1[10]);
  nand g85 (n_165, in_0[10], in_2[10]);
  nand g86 (out_0[11], n_163, n_164, n_165);
  xor g87 (n_166, in_0[11], in_1[11]);
  xor g88 (out_1[11], n_166, in_2[11]);
  nand g89 (n_167, in_0[11], in_1[11]);
  nand g90 (n_168, in_2[11], in_1[11]);
  nand g91 (n_169, in_0[11], in_2[11]);
  nand g92 (out_0[12], n_167, n_168, n_169);
  xor g93 (n_170, in_0[12], in_1[12]);
  xor g94 (out_1[12], n_170, in_2[12]);
  nand g95 (n_171, in_0[12], in_1[12]);
  nand g96 (n_172, in_2[12], in_1[12]);
  nand g97 (n_173, in_0[12], in_2[12]);
  nand g98 (out_0[13], n_171, n_172, n_173);
  xor g99 (n_174, in_0[13], in_1[13]);
  xor g100 (out_1[13], n_174, in_2[13]);
  nand g101 (n_175, in_0[13], in_1[13]);
  nand g102 (n_176, in_2[13], in_1[13]);
  nand g103 (n_177, in_0[13], in_2[13]);
  nand g104 (out_0[14], n_175, n_176, n_177);
  xor g105 (n_178, in_0[14], in_1[14]);
  xor g106 (out_1[14], n_178, in_2[14]);
  nand g107 (n_179, in_0[14], in_1[14]);
  nand g108 (n_180, in_2[14], in_1[14]);
  nand g109 (n_181, in_0[14], in_2[14]);
  nand g110 (out_0[15], n_179, n_180, n_181);
  xor g111 (n_182, in_0[15], in_1[15]);
  xor g112 (out_1[15], n_182, in_2[15]);
  nand g113 (n_183, in_0[15], in_1[15]);
  nand g114 (n_184, in_2[15], in_1[15]);
  nand g115 (n_185, in_0[15], in_2[15]);
  nand g116 (out_0[16], n_183, n_184, n_185);
  xor g117 (n_186, in_0[16], in_1[16]);
  xor g118 (out_1[16], n_186, in_2[16]);
  nand g119 (n_187, in_0[16], in_1[16]);
  nand g120 (n_188, in_2[16], in_1[16]);
  nand g121 (n_189, in_0[16], in_2[16]);
  nand g122 (out_0[17], n_187, n_188, n_189);
  xor g123 (n_190, in_0[17], in_1[17]);
  xor g124 (out_1[17], n_190, in_2[17]);
  nand g125 (n_191, in_0[17], in_1[17]);
  nand g126 (n_192, in_2[17], in_1[17]);
  nand g127 (n_193, in_0[17], in_2[17]);
  nand g128 (out_0[18], n_191, n_192, n_193);
  xor g129 (n_194, in_0[18], in_1[18]);
  xor g130 (out_1[18], n_194, in_2[18]);
  nand g131 (n_195, in_0[18], in_1[18]);
  nand g132 (n_196, in_2[18], in_1[18]);
  nand g133 (n_197, in_0[18], in_2[18]);
  nand g134 (out_0[19], n_195, n_196, n_197);
  xor g135 (n_198, in_0[19], in_1[19]);
  xor g136 (out_1[19], n_198, in_2[19]);
  nand g137 (n_199, in_0[19], in_1[19]);
  nand g138 (n_200, in_2[19], in_1[19]);
  nand g139 (n_201, in_0[19], in_2[19]);
  nand g140 (out_0[20], n_199, n_200, n_201);
  xor g141 (n_202, in_0[20], in_1[20]);
  xor g142 (out_1[20], n_202, in_2[20]);
  nand g143 (n_203, in_0[20], in_1[20]);
  nand g144 (n_204, in_2[20], in_1[20]);
  nand g145 (n_205, in_0[20], in_2[20]);
  nand g146 (out_0[21], n_203, n_204, n_205);
  xor g147 (n_206, in_0[21], in_1[21]);
  xor g148 (out_1[21], n_206, in_2[21]);
  nand g149 (n_207, in_0[21], in_1[21]);
  nand g150 (n_208, in_2[21], in_1[21]);
  nand g151 (n_209, in_0[21], in_2[21]);
  nand g152 (out_0[22], n_207, n_208, n_209);
  xor g156 (out_1[22], in_2[22], n_73);
  xor g161 (n_73, in_0[22], in_1[22]);
  nor g162 (out_0[23], in_0[22], in_1[22]);
  or g163 (n_212, in_2[22], wc);
  not gc (wc, n_73);
  or g165 (out_1[23], wc0, wc1, n_73);
  not gc1 (wc1, n_212);
  not gc0 (wc0, in_2[22]);
endmodule

module csa_tree_6719_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [22:0] in_0, in_1, in_2;
  output [25:0] out_0, out_1;
  wire [22:0] in_0, in_1, in_2;
  wire [25:0] out_0, out_1;
  csa_tree_6719_GENERIC_REAL g1(.in_0 ({in_0[21], in_0[21:0]}), .in_1
       ({in_1[21], in_1[21:0]}), .in_2 (in_2), .out_0 (out_0), .out_1
       (out_1));
endmodule

module csa_tree_6744_GENERIC_REAL(in_0, in_1, in_2, out_0, out_1);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ; assign out_1 = 27'b0;"
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [26:0] out_0, out_1;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [26:0] out_0, out_1;
  wire n_76, n_80, n_81, n_85, n_86, n_141, n_142, n_143;
  wire n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151;
  wire n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159;
  wire n_160, n_161, n_162, n_163, n_164, n_165, n_166, n_167;
  wire n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199;
  wire n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207;
  wire n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215;
  wire n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223;
  wire n_224, n_225, n_226, n_227, n_228, n_231, n_235, n_239;
  assign out_0[0] = in_1[0];
  xor g33 (out_1[0], in_0[0], in_2[0]);
  and g34 (out_0[1], in_0[0], in_2[0]);
  xor g35 (n_141, in_0[1], in_1[1]);
  xor g36 (out_1[1], n_141, in_2[1]);
  nand g37 (n_142, in_0[1], in_1[1]);
  nand g4 (n_143, in_2[1], in_1[1]);
  nand g5 (n_144, in_0[1], in_2[1]);
  nand g38 (out_0[2], n_142, n_143, n_144);
  xor g39 (n_145, in_0[2], in_1[2]);
  xor g40 (out_1[2], n_145, in_2[2]);
  nand g41 (n_146, in_0[2], in_1[2]);
  nand g42 (n_147, in_2[2], in_1[2]);
  nand g43 (n_148, in_0[2], in_2[2]);
  nand g6 (out_0[3], n_146, n_147, n_148);
  xor g44 (n_149, in_0[3], in_1[3]);
  xor g45 (out_1[3], n_149, in_2[3]);
  nand g46 (n_150, in_0[3], in_1[3]);
  nand g47 (n_151, in_2[3], in_1[3]);
  nand g48 (n_152, in_0[3], in_2[3]);
  nand g49 (out_0[4], n_150, n_151, n_152);
  xor g50 (n_153, in_0[4], in_1[4]);
  xor g51 (out_1[4], n_153, in_2[4]);
  nand g52 (n_154, in_0[4], in_1[4]);
  nand g53 (n_155, in_2[4], in_1[4]);
  nand g54 (n_156, in_0[4], in_2[4]);
  nand g55 (out_0[5], n_154, n_155, n_156);
  xor g56 (n_157, in_0[5], in_1[5]);
  xor g57 (out_1[5], n_157, in_2[5]);
  nand g58 (n_158, in_0[5], in_1[5]);
  nand g59 (n_159, in_2[5], in_1[5]);
  nand g60 (n_160, in_0[5], in_2[5]);
  nand g61 (out_0[6], n_158, n_159, n_160);
  xor g62 (n_161, in_0[6], in_1[6]);
  xor g63 (out_1[6], n_161, in_2[6]);
  nand g64 (n_162, in_0[6], in_1[6]);
  nand g65 (n_163, in_2[6], in_1[6]);
  nand g66 (n_164, in_0[6], in_2[6]);
  nand g67 (out_0[7], n_162, n_163, n_164);
  xor g68 (n_165, in_0[7], in_1[7]);
  xor g69 (out_1[7], n_165, in_2[7]);
  nand g70 (n_166, in_0[7], in_1[7]);
  nand g71 (n_167, in_2[7], in_1[7]);
  nand g72 (n_168, in_0[7], in_2[7]);
  nand g73 (out_0[8], n_166, n_167, n_168);
  xor g74 (n_169, in_0[8], in_1[8]);
  xor g75 (out_1[8], n_169, in_2[8]);
  nand g76 (n_170, in_0[8], in_1[8]);
  nand g77 (n_171, in_2[8], in_1[8]);
  nand g78 (n_172, in_0[8], in_2[8]);
  nand g79 (out_0[9], n_170, n_171, n_172);
  xor g80 (n_173, in_0[9], in_1[9]);
  xor g81 (out_1[9], n_173, in_2[9]);
  nand g82 (n_174, in_0[9], in_1[9]);
  nand g83 (n_175, in_2[9], in_1[9]);
  nand g84 (n_176, in_0[9], in_2[9]);
  nand g85 (out_0[10], n_174, n_175, n_176);
  xor g86 (n_177, in_0[10], in_1[10]);
  xor g87 (out_1[10], n_177, in_2[10]);
  nand g88 (n_178, in_0[10], in_1[10]);
  nand g89 (n_179, in_2[10], in_1[10]);
  nand g90 (n_180, in_0[10], in_2[10]);
  nand g91 (out_0[11], n_178, n_179, n_180);
  xor g92 (n_181, in_0[11], in_1[11]);
  xor g93 (out_1[11], n_181, in_2[11]);
  nand g94 (n_182, in_0[11], in_1[11]);
  nand g95 (n_183, in_2[11], in_1[11]);
  nand g96 (n_184, in_0[11], in_2[11]);
  nand g97 (out_0[12], n_182, n_183, n_184);
  xor g98 (n_185, in_0[12], in_1[12]);
  xor g99 (out_1[12], n_185, in_2[12]);
  nand g100 (n_186, in_0[12], in_1[12]);
  nand g101 (n_187, in_2[12], in_1[12]);
  nand g102 (n_188, in_0[12], in_2[12]);
  nand g103 (out_0[13], n_186, n_187, n_188);
  xor g104 (n_189, in_0[13], in_1[13]);
  xor g105 (out_1[13], n_189, in_2[13]);
  nand g106 (n_190, in_0[13], in_1[13]);
  nand g107 (n_191, in_2[13], in_1[13]);
  nand g108 (n_192, in_0[13], in_2[13]);
  nand g109 (out_0[14], n_190, n_191, n_192);
  xor g110 (n_193, in_0[14], in_1[14]);
  xor g111 (out_1[14], n_193, in_2[14]);
  nand g112 (n_194, in_0[14], in_1[14]);
  nand g113 (n_195, in_2[14], in_1[14]);
  nand g114 (n_196, in_0[14], in_2[14]);
  nand g115 (out_0[15], n_194, n_195, n_196);
  xor g116 (n_197, in_0[15], in_1[15]);
  xor g117 (out_1[15], n_197, in_2[15]);
  nand g118 (n_198, in_0[15], in_1[15]);
  nand g119 (n_199, in_2[15], in_1[15]);
  nand g120 (n_200, in_0[15], in_2[15]);
  nand g121 (out_0[16], n_198, n_199, n_200);
  xor g122 (n_201, in_0[16], in_1[16]);
  xor g123 (out_1[16], n_201, in_2[16]);
  nand g124 (n_202, in_0[16], in_1[16]);
  nand g125 (n_203, in_2[16], in_1[16]);
  nand g126 (n_204, in_0[16], in_2[16]);
  nand g127 (out_0[17], n_202, n_203, n_204);
  xor g128 (n_205, in_0[17], in_1[17]);
  xor g129 (out_1[17], n_205, in_2[17]);
  nand g130 (n_206, in_0[17], in_1[17]);
  nand g131 (n_207, in_2[17], in_1[17]);
  nand g132 (n_208, in_0[17], in_2[17]);
  nand g133 (out_0[18], n_206, n_207, n_208);
  xor g134 (n_209, in_0[18], in_1[18]);
  xor g135 (out_1[18], n_209, in_2[18]);
  nand g136 (n_210, in_0[18], in_1[18]);
  nand g137 (n_211, in_2[18], in_1[18]);
  nand g138 (n_212, in_0[18], in_2[18]);
  nand g139 (out_0[19], n_210, n_211, n_212);
  xor g140 (n_213, in_0[19], in_1[19]);
  xor g141 (out_1[19], n_213, in_2[19]);
  nand g142 (n_214, in_0[19], in_1[19]);
  nand g143 (n_215, in_2[19], in_1[19]);
  nand g144 (n_216, in_0[19], in_2[19]);
  nand g145 (out_0[20], n_214, n_215, n_216);
  xor g146 (n_217, in_0[20], in_1[20]);
  xor g147 (out_1[20], n_217, in_2[20]);
  nand g148 (n_218, in_0[20], in_1[20]);
  nand g149 (n_219, in_2[20], in_1[20]);
  nand g150 (n_220, in_0[20], in_2[20]);
  nand g151 (out_0[21], n_218, n_219, n_220);
  xor g152 (n_221, in_0[21], in_1[21]);
  xor g153 (out_1[21], n_221, in_2[21]);
  nand g154 (n_222, in_0[21], in_1[21]);
  nand g155 (n_223, in_2[21], in_1[21]);
  nand g156 (n_224, in_0[21], in_2[21]);
  nand g157 (out_0[22], n_222, n_223, n_224);
  xor g158 (n_225, in_0[22], in_1[22]);
  xor g159 (out_1[22], n_225, in_2[22]);
  nand g160 (n_226, in_0[22], in_1[22]);
  nand g161 (n_227, in_2[22], in_1[22]);
  nand g162 (n_228, in_0[22], in_2[22]);
  nand g163 (out_0[23], n_226, n_227, n_228);
  xor g164 (n_76, in_0[23], in_1[23]);
  and g165 (n_81, in_0[23], in_1[23]);
  xor g167 (out_1[23], in_2[23], n_76);
  xor g172 (n_80, in_0[24], in_1[24]);
  and g173 (n_86, in_0[24], in_1[24]);
  nand g177 (n_235, n_81, n_80);
  nand g185 (n_239, n_86, n_85);
  or g188 (n_231, in_2[23], wc);
  not gc (wc, n_76);
  xor g192 (n_85, in_0[25], in_1[25]);
  nor g193 (out_0[26], in_0[25], in_1[25]);
  or g195 (out_0[24], wc0, wc1, n_76);
  not gc1 (wc1, n_231);
  not gc0 (wc0, in_2[23]);
  xnor g196 (out_1[24], n_81, n_80);
  or g197 (out_0[25], wc2, n_80, n_81);
  not gc2 (wc2, n_235);
  xnor g199 (out_1[25], n_86, n_85);
  or g200 (out_1[26], n_85, wc3, n_86);
  not gc3 (wc3, n_239);
endmodule

module csa_tree_6744_GENERIC(in_0, in_1, in_2, out_0, out_1);
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [26:0] out_0, out_1;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [26:0] out_0, out_1;
  csa_tree_6744_GENERIC_REAL g1(.in_0 (in_0), .in_1 (in_1), .in_2
       (in_2), .out_0 (out_0), .out_1 (out_1));
endmodule

module csa_tree_add_178_36_group_6829_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_157, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_242, n_243;
  wire n_244, n_245, n_246, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_255, n_256, n_257, n_258, n_259, n_261, n_262;
  wire n_263, n_264, n_265, n_267, n_268, n_269, n_270, n_271;
  wire n_273, n_274, n_275, n_276, n_277, n_279, n_280, n_281;
  wire n_282, n_283, n_285, n_286, n_287, n_288, n_289, n_291;
  wire n_292, n_293, n_294, n_295, n_297, n_298, n_299, n_300;
  wire n_301, n_303, n_304, n_305, n_306, n_307, n_309, n_310;
  wire n_311, n_312, n_313, n_315, n_316, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_325, n_327, n_329, n_330, n_332;
  wire n_333, n_335, n_337, n_339, n_340, n_342, n_343, n_345;
  wire n_347, n_349, n_350, n_352, n_353, n_355, n_357, n_359;
  wire n_360, n_362, n_363, n_365, n_367, n_369, n_370, n_372;
  wire n_374, n_375, n_376, n_378, n_379, n_380, n_382, n_383;
  wire n_384, n_385, n_387, n_389, n_391, n_392, n_393, n_395;
  wire n_396, n_397, n_399, n_400, n_402, n_404, n_406, n_407;
  wire n_408, n_410, n_411, n_412, n_414, n_416, n_417, n_418;
  wire n_420, n_421, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_441, n_443, n_444, n_445, n_447;
  wire n_448, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_464, n_465;
  wire n_466, n_468, n_469, n_470, n_471, n_473, n_474, n_475;
  wire n_477, n_478, n_479, n_480, n_482, n_483, n_485, n_486;
  wire n_488, n_489, n_490, n_491, n_493, n_494, n_495, n_497;
  wire n_498, n_499, n_500, n_502, n_503, n_505, n_506, n_508;
  wire n_509, n_510, n_511, n_513, n_514, n_515, n_516, n_517;
  xor g26 (n_125, in_2[1], in_0[1]);
  and g2 (n_153, in_2[1], in_0[1]);
  xor g27 (n_157, in_2[2], n_153);
  xor g28 (n_149, n_157, in_0[2]);
  nand g3 (n_124, in_2[2], n_153);
  nand g29 (n_158, in_0[2], n_153);
  nand g30 (n_126, in_2[2], in_0[2]);
  nand g31 (n_123, n_124, n_158, n_126);
  xor g32 (n_159, in_2[3], in_0[3]);
  xor g33 (n_148, n_159, in_1[3]);
  nand g34 (n_160, in_2[3], in_0[3]);
  nand g4 (n_161, in_1[3], in_0[3]);
  nand g35 (n_162, in_2[3], in_1[3]);
  nand g36 (n_122, n_160, n_161, n_162);
  xor g37 (n_163, in_2[4], in_0[4]);
  xor g38 (n_147, n_163, in_1[4]);
  nand g39 (n_164, in_2[4], in_0[4]);
  nand g40 (n_165, in_1[4], in_0[4]);
  nand g5 (n_166, in_2[4], in_1[4]);
  nand g41 (n_121, n_164, n_165, n_166);
  xor g42 (n_167, in_2[5], in_0[5]);
  xor g43 (n_146, n_167, in_1[5]);
  nand g44 (n_168, in_2[5], in_0[5]);
  nand g45 (n_169, in_1[5], in_0[5]);
  nand g46 (n_170, in_2[5], in_1[5]);
  nand g6 (n_120, n_168, n_169, n_170);
  xor g47 (n_171, in_2[6], in_0[6]);
  xor g48 (n_145, n_171, in_1[6]);
  nand g49 (n_172, in_2[6], in_0[6]);
  nand g50 (n_173, in_1[6], in_0[6]);
  nand g51 (n_174, in_2[6], in_1[6]);
  nand g52 (n_119, n_172, n_173, n_174);
  xor g53 (n_175, in_2[7], in_0[7]);
  xor g54 (n_144, n_175, in_1[7]);
  nand g55 (n_176, in_2[7], in_0[7]);
  nand g56 (n_177, in_1[7], in_0[7]);
  nand g57 (n_178, in_2[7], in_1[7]);
  nand g58 (n_118, n_176, n_177, n_178);
  xor g59 (n_179, in_2[8], in_0[8]);
  xor g60 (n_143, n_179, in_1[8]);
  nand g61 (n_180, in_2[8], in_0[8]);
  nand g62 (n_181, in_1[8], in_0[8]);
  nand g63 (n_150, in_2[8], in_1[8]);
  nand g64 (n_117, n_180, n_181, n_150);
  xor g65 (n_151, in_2[9], in_0[9]);
  xor g66 (n_142, n_151, in_1[9]);
  nand g67 (n_152, in_2[9], in_0[9]);
  nand g68 (n_182, in_1[9], in_0[9]);
  nand g69 (n_183, in_2[9], in_1[9]);
  nand g70 (n_116, n_152, n_182, n_183);
  xor g71 (n_184, in_2[10], in_0[10]);
  xor g72 (n_141, n_184, in_1[10]);
  nand g73 (n_185, in_2[10], in_0[10]);
  nand g74 (n_186, in_1[10], in_0[10]);
  nand g75 (n_187, in_2[10], in_1[10]);
  nand g76 (n_115, n_185, n_186, n_187);
  xor g77 (n_188, in_2[11], in_0[11]);
  xor g78 (n_140, n_188, in_1[11]);
  nand g79 (n_189, in_2[11], in_0[11]);
  nand g80 (n_190, in_1[11], in_0[11]);
  nand g81 (n_191, in_2[11], in_1[11]);
  nand g82 (n_114, n_189, n_190, n_191);
  xor g83 (n_192, in_2[12], in_0[12]);
  xor g84 (n_139, n_192, in_1[12]);
  nand g85 (n_193, in_2[12], in_0[12]);
  nand g86 (n_194, in_1[12], in_0[12]);
  nand g87 (n_195, in_2[12], in_1[12]);
  nand g88 (n_113, n_193, n_194, n_195);
  xor g89 (n_196, in_2[13], in_0[13]);
  xor g90 (n_138, n_196, in_1[13]);
  nand g91 (n_197, in_2[13], in_0[13]);
  nand g92 (n_198, in_1[13], in_0[13]);
  nand g93 (n_199, in_2[13], in_1[13]);
  nand g94 (n_112, n_197, n_198, n_199);
  xor g95 (n_200, in_2[14], in_0[14]);
  xor g96 (n_137, n_200, in_1[14]);
  nand g97 (n_201, in_2[14], in_0[14]);
  nand g98 (n_202, in_1[14], in_0[14]);
  nand g99 (n_203, in_2[14], in_1[14]);
  nand g100 (n_111, n_201, n_202, n_203);
  xor g101 (n_204, in_2[15], in_0[15]);
  xor g102 (n_136, n_204, in_1[15]);
  nand g103 (n_205, in_2[15], in_0[15]);
  nand g104 (n_206, in_1[15], in_0[15]);
  nand g105 (n_207, in_2[15], in_1[15]);
  nand g106 (n_110, n_205, n_206, n_207);
  xor g107 (n_208, in_2[16], in_0[16]);
  xor g108 (n_135, n_208, in_1[16]);
  nand g109 (n_209, in_2[16], in_0[16]);
  nand g110 (n_210, in_1[16], in_0[16]);
  nand g111 (n_211, in_2[16], in_1[16]);
  nand g112 (n_109, n_209, n_210, n_211);
  xor g113 (n_212, in_2[17], in_0[17]);
  xor g114 (n_134, n_212, in_1[17]);
  nand g115 (n_213, in_2[17], in_0[17]);
  nand g116 (n_214, in_1[17], in_0[17]);
  nand g117 (n_215, in_2[17], in_1[17]);
  nand g118 (n_108, n_213, n_214, n_215);
  xor g119 (n_216, in_2[18], in_0[18]);
  xor g120 (n_133, n_216, in_1[18]);
  nand g121 (n_217, in_2[18], in_0[18]);
  nand g122 (n_218, in_1[18], in_0[18]);
  nand g123 (n_219, in_2[18], in_1[18]);
  nand g124 (n_107, n_217, n_218, n_219);
  xor g125 (n_220, in_2[19], in_0[19]);
  xor g126 (n_132, n_220, in_1[19]);
  nand g127 (n_221, in_2[19], in_0[19]);
  nand g128 (n_222, in_1[19], in_0[19]);
  nand g129 (n_223, in_2[19], in_1[19]);
  nand g130 (n_106, n_221, n_222, n_223);
  xor g131 (n_224, in_2[20], in_0[20]);
  xor g132 (n_131, n_224, in_1[20]);
  nand g133 (n_225, in_2[20], in_0[20]);
  nand g134 (n_226, in_1[20], in_0[20]);
  nand g135 (n_227, in_2[20], in_1[20]);
  nand g136 (n_105, n_225, n_226, n_227);
  xor g137 (n_228, in_2[21], in_0[21]);
  xor g138 (n_130, n_228, in_1[21]);
  nand g139 (n_229, in_2[21], in_0[21]);
  nand g140 (n_230, in_1[21], in_0[21]);
  nand g141 (n_231, in_2[21], in_1[21]);
  nand g142 (n_104, n_229, n_230, n_231);
  xor g143 (n_232, in_2[22], in_0[22]);
  xor g144 (n_129, n_232, in_1[22]);
  nand g145 (n_233, in_2[22], in_0[22]);
  nand g146 (n_234, in_1[22], in_0[22]);
  nand g147 (n_235, in_2[22], in_1[22]);
  nand g148 (n_128, n_233, n_234, n_235);
  xor g151 (n_236, in_2[23], in_1[23]);
  xor g152 (n_103, n_236, in_0[23]);
  nand g153 (n_237, in_2[23], in_1[23]);
  nand g154 (n_238, in_0[23], in_1[23]);
  nand g155 (n_239, in_2[23], in_0[23]);
  nand g156 (n_127, n_237, n_238, n_239);
  xor g159 (n_517, in_0[0], in_1[0]);
  nand g160 (n_242, in_0[0], in_1[0]);
  nand g161 (n_243, in_0[0], in_2[0]);
  nand g7 (n_244, in_1[0], in_2[0]);
  nand g8 (n_246, n_242, n_243, n_244);
  nor g9 (n_245, n_125, in_1[1]);
  nand g10 (n_248, n_125, in_1[1]);
  nor g11 (n_255, in_1[2], n_149);
  nand g12 (n_250, in_1[2], n_149);
  nor g13 (n_251, n_123, n_148);
  nand g14 (n_252, n_123, n_148);
  nor g15 (n_261, n_122, n_147);
  nand g16 (n_256, n_122, n_147);
  nor g17 (n_257, n_121, n_146);
  nand g18 (n_258, n_121, n_146);
  nor g19 (n_267, n_120, n_145);
  nand g20 (n_262, n_120, n_145);
  nor g21 (n_263, n_119, n_144);
  nand g22 (n_264, n_119, n_144);
  nor g23 (n_273, n_118, n_143);
  nand g24 (n_268, n_118, n_143);
  nor g25 (n_269, n_117, n_142);
  nand g162 (n_270, n_117, n_142);
  nor g163 (n_279, n_116, n_141);
  nand g164 (n_274, n_116, n_141);
  nor g165 (n_275, n_115, n_140);
  nand g166 (n_276, n_115, n_140);
  nor g167 (n_285, n_114, n_139);
  nand g168 (n_280, n_114, n_139);
  nor g169 (n_281, n_113, n_138);
  nand g170 (n_282, n_113, n_138);
  nor g171 (n_291, n_112, n_137);
  nand g172 (n_286, n_112, n_137);
  nor g173 (n_287, n_111, n_136);
  nand g174 (n_288, n_111, n_136);
  nor g175 (n_297, n_110, n_135);
  nand g176 (n_292, n_110, n_135);
  nor g177 (n_293, n_109, n_134);
  nand g178 (n_294, n_109, n_134);
  nor g179 (n_303, n_108, n_133);
  nand g180 (n_298, n_108, n_133);
  nor g181 (n_299, n_107, n_132);
  nand g182 (n_300, n_107, n_132);
  nor g183 (n_309, n_106, n_131);
  nand g184 (n_304, n_106, n_131);
  nor g185 (n_305, n_105, n_130);
  nand g186 (n_306, n_105, n_130);
  nor g187 (n_315, n_104, n_129);
  nand g188 (n_310, n_104, n_129);
  nor g189 (n_311, n_103, n_128);
  nand g190 (n_312, n_103, n_128);
  nand g195 (n_316, n_248, n_249);
  nor g196 (n_253, n_250, n_251);
  nor g199 (n_319, n_255, n_251);
  nor g200 (n_259, n_256, n_257);
  nor g203 (n_325, n_261, n_257);
  nor g204 (n_265, n_262, n_263);
  nor g207 (n_327, n_267, n_263);
  nor g208 (n_271, n_268, n_269);
  nor g211 (n_335, n_273, n_269);
  nor g212 (n_277, n_274, n_275);
  nor g215 (n_337, n_279, n_275);
  nor g216 (n_283, n_280, n_281);
  nor g219 (n_345, n_285, n_281);
  nor g220 (n_289, n_286, n_287);
  nor g223 (n_347, n_291, n_287);
  nor g224 (n_295, n_292, n_293);
  nor g227 (n_355, n_297, n_293);
  nor g228 (n_301, n_298, n_299);
  nor g231 (n_357, n_303, n_299);
  nor g232 (n_307, n_304, n_305);
  nor g235 (n_365, n_309, n_305);
  nor g236 (n_313, n_310, n_311);
  nor g239 (n_367, n_315, n_311);
  nand g242 (n_464, n_250, n_318);
  nand g243 (n_321, n_319, n_316);
  nand g244 (n_372, n_320, n_321);
  nor g245 (n_323, n_267, n_322);
  nand g254 (n_380, n_325, n_327);
  nor g255 (n_333, n_279, n_332);
  nand g264 (n_387, n_335, n_337);
  nor g265 (n_343, n_291, n_342);
  nand g274 (n_395, n_345, n_347);
  nor g275 (n_353, n_303, n_352);
  nand g284 (n_402, n_355, n_357);
  nor g285 (n_363, n_315, n_362);
  nand g294 (n_410, n_365, n_367);
  nand g297 (n_468, n_256, n_374);
  nand g298 (n_375, n_325, n_372);
  nand g299 (n_470, n_322, n_375);
  nand g302 (n_473, n_378, n_379);
  nand g305 (n_414, n_382, n_383);
  nor g306 (n_385, n_285, n_384);
  nor g309 (n_424, n_285, n_387);
  nor g315 (n_393, n_391, n_384);
  nor g318 (n_430, n_387, n_391);
  nor g319 (n_397, n_395, n_384);
  nor g322 (n_433, n_387, n_395);
  nor g323 (n_400, n_309, n_399);
  nor g326 (n_451, n_309, n_402);
  nor g332 (n_408, n_406, n_399);
  nor g335 (n_457, n_402, n_406);
  nor g336 (n_412, n_410, n_399);
  nor g339 (n_439, n_402, n_410);
  nand g342 (n_477, n_268, n_416);
  nand g343 (n_417, n_335, n_414);
  nand g344 (n_479, n_332, n_417);
  nand g347 (n_482, n_420, n_421);
  nand g350 (n_485, n_384, n_423);
  nand g351 (n_426, n_424, n_414);
  nand g352 (n_488, n_425, n_426);
  nand g353 (n_429, n_427, n_414);
  nand g354 (n_490, n_428, n_429);
  nand g355 (n_432, n_430, n_414);
  nand g356 (n_493, n_431, n_432);
  nand g357 (n_435, n_433, n_414);
  nand g358 (n_441, n_434, n_435);
  nand g362 (n_497, n_292, n_443);
  nand g363 (n_444, n_355, n_441);
  nand g364 (n_499, n_352, n_444);
  nand g367 (n_502, n_447, n_448);
  nand g370 (n_505, n_399, n_450);
  nand g371 (n_453, n_451, n_441);
  nand g372 (n_508, n_452, n_453);
  nand g373 (n_456, n_454, n_441);
  nand g374 (n_510, n_455, n_456);
  nand g375 (n_459, n_457, n_441);
  nand g376 (n_513, n_458, n_459);
  nand g377 (n_460, n_439, n_441);
  nand g378 (n_515, n_437, n_460);
  xnor g380 (out_0[1], n_246, n_461);
  xnor g382 (out_0[2], n_316, n_462);
  xnor g385 (out_0[3], n_464, n_465);
  xnor g387 (out_0[4], n_372, n_466);
  xnor g390 (out_0[5], n_468, n_469);
  xnor g392 (out_0[6], n_470, n_471);
  xnor g395 (out_0[7], n_473, n_474);
  xnor g397 (out_0[8], n_414, n_475);
  xnor g400 (out_0[9], n_477, n_478);
  xnor g402 (out_0[10], n_479, n_480);
  xnor g405 (out_0[11], n_482, n_483);
  xnor g408 (out_0[12], n_485, n_486);
  xnor g411 (out_0[13], n_488, n_489);
  xnor g413 (out_0[14], n_490, n_491);
  xnor g416 (out_0[15], n_493, n_494);
  xnor g418 (out_0[16], n_441, n_495);
  xnor g421 (out_0[17], n_497, n_498);
  xnor g423 (out_0[18], n_499, n_500);
  xnor g426 (out_0[19], n_502, n_503);
  xnor g429 (out_0[20], n_505, n_506);
  xnor g432 (out_0[21], n_508, n_509);
  xnor g434 (out_0[22], n_510, n_511);
  xnor g437 (out_0[23], n_513, n_514);
  xnor g439 (out_0[24], n_515, n_516);
  xor g440 (out_0[0], in_2[0], n_517);
  or g441 (n_249, n_245, wc);
  not gc (wc, n_246);
  or g442 (n_461, wc0, n_245);
  not gc0 (wc0, n_248);
  and g443 (n_322, wc1, n_258);
  not gc1 (wc1, n_259);
  and g444 (n_329, wc2, n_264);
  not gc2 (wc2, n_265);
  and g445 (n_332, wc3, n_270);
  not gc3 (wc3, n_271);
  and g446 (n_339, wc4, n_276);
  not gc4 (wc4, n_277);
  and g447 (n_342, wc5, n_282);
  not gc5 (wc5, n_283);
  and g448 (n_349, wc6, n_288);
  not gc6 (wc6, n_289);
  and g449 (n_352, wc7, n_294);
  not gc7 (wc7, n_295);
  and g450 (n_359, wc8, n_300);
  not gc8 (wc8, n_301);
  and g451 (n_362, wc9, n_306);
  not gc9 (wc9, n_307);
  or g452 (n_376, wc10, n_267);
  not gc10 (wc10, n_325);
  or g453 (n_418, wc11, n_279);
  not gc11 (wc11, n_335);
  or g454 (n_391, wc12, n_291);
  not gc12 (wc12, n_345);
  or g455 (n_445, wc13, n_303);
  not gc13 (wc13, n_355);
  or g456 (n_406, wc14, n_315);
  not gc14 (wc14, n_365);
  or g457 (n_466, wc15, n_261);
  not gc15 (wc15, n_256);
  or g458 (n_469, wc16, n_257);
  not gc16 (wc16, n_258);
  or g459 (n_471, wc17, n_267);
  not gc17 (wc17, n_262);
  or g460 (n_474, wc18, n_263);
  not gc18 (wc18, n_264);
  or g461 (n_475, wc19, n_273);
  not gc19 (wc19, n_268);
  or g462 (n_478, wc20, n_269);
  not gc20 (wc20, n_270);
  or g463 (n_480, wc21, n_279);
  not gc21 (wc21, n_274);
  or g464 (n_483, wc22, n_275);
  not gc22 (wc22, n_276);
  or g465 (n_486, wc23, n_285);
  not gc23 (wc23, n_280);
  or g466 (n_489, wc24, n_281);
  not gc24 (wc24, n_282);
  or g467 (n_491, wc25, n_291);
  not gc25 (wc25, n_286);
  or g468 (n_494, wc26, n_287);
  not gc26 (wc26, n_288);
  or g469 (n_495, wc27, n_297);
  not gc27 (wc27, n_292);
  or g470 (n_498, wc28, n_293);
  not gc28 (wc28, n_294);
  or g471 (n_500, wc29, n_303);
  not gc29 (wc29, n_298);
  or g472 (n_503, wc30, n_299);
  not gc30 (wc30, n_300);
  or g473 (n_506, wc31, n_309);
  not gc31 (wc31, n_304);
  or g474 (n_509, wc32, n_305);
  not gc32 (wc32, n_306);
  or g475 (n_511, wc33, n_315);
  not gc33 (wc33, n_310);
  and g476 (n_436, wc34, n_127);
  not gc34 (wc34, in_2[23]);
  or g477 (n_438, wc35, n_127);
  not gc35 (wc35, in_2[23]);
  and g478 (n_320, wc36, n_252);
  not gc36 (wc36, n_253);
  or g479 (n_318, wc37, n_255);
  not gc37 (wc37, n_316);
  and g480 (n_330, wc38, n_327);
  not gc38 (wc38, n_322);
  and g481 (n_340, wc39, n_337);
  not gc39 (wc39, n_332);
  and g482 (n_350, wc40, n_347);
  not gc40 (wc40, n_342);
  and g483 (n_360, wc41, n_357);
  not gc41 (wc41, n_352);
  and g484 (n_427, wc42, n_345);
  not gc42 (wc42, n_387);
  and g485 (n_454, wc43, n_365);
  not gc43 (wc43, n_402);
  or g486 (n_462, wc44, n_255);
  not gc44 (wc44, n_250);
  or g487 (n_465, wc45, n_251);
  not gc45 (wc45, n_252);
  and g488 (n_369, wc46, n_312);
  not gc46 (wc46, n_313);
  and g489 (n_378, wc47, n_262);
  not gc47 (wc47, n_323);
  and g490 (n_382, wc48, n_329);
  not gc48 (wc48, n_330);
  and g491 (n_420, wc49, n_274);
  not gc49 (wc49, n_333);
  and g492 (n_384, wc50, n_339);
  not gc50 (wc50, n_340);
  and g493 (n_392, wc51, n_286);
  not gc51 (wc51, n_343);
  and g494 (n_396, wc52, n_349);
  not gc52 (wc52, n_350);
  and g495 (n_447, wc53, n_298);
  not gc53 (wc53, n_353);
  and g496 (n_399, wc54, n_359);
  not gc54 (wc54, n_360);
  and g497 (n_407, wc55, n_310);
  not gc55 (wc55, n_363);
  or g498 (n_514, wc56, n_311);
  not gc56 (wc56, n_312);
  and g499 (n_370, wc57, n_367);
  not gc57 (wc57, n_362);
  or g500 (n_374, wc58, n_261);
  not gc58 (wc58, n_372);
  or g501 (n_379, n_376, wc59);
  not gc59 (wc59, n_372);
  or g502 (n_383, n_380, wc60);
  not gc60 (wc60, n_372);
  and g503 (n_389, wc61, n_345);
  not gc61 (wc61, n_384);
  and g504 (n_404, wc62, n_365);
  not gc62 (wc62, n_399);
  or g505 (n_516, wc63, n_436);
  not gc63 (wc63, n_438);
  and g506 (n_411, wc64, n_369);
  not gc64 (wc64, n_370);
  and g507 (n_425, wc65, n_280);
  not gc65 (wc65, n_385);
  and g508 (n_428, wc66, n_342);
  not gc66 (wc66, n_389);
  and g509 (n_431, n_392, wc67);
  not gc67 (wc67, n_393);
  and g510 (n_434, n_396, wc68);
  not gc68 (wc68, n_397);
  and g511 (n_452, wc69, n_304);
  not gc69 (wc69, n_400);
  and g512 (n_455, wc70, n_362);
  not gc70 (wc70, n_404);
  and g513 (n_458, n_407, wc71);
  not gc71 (wc71, n_408);
  or g514 (n_416, wc72, n_273);
  not gc72 (wc72, n_414);
  or g515 (n_421, n_418, wc73);
  not gc73 (wc73, n_414);
  or g516 (n_423, wc74, n_387);
  not gc74 (wc74, n_414);
  and g517 (n_437, n_411, wc75);
  not gc75 (wc75, n_412);
  or g518 (n_443, wc76, n_297);
  not gc76 (wc76, n_441);
  or g519 (n_448, n_445, wc77);
  not gc77 (wc77, n_441);
  or g520 (n_450, wc78, n_402);
  not gc78 (wc78, n_441);
endmodule

module csa_tree_add_178_36_group_6829_GENERIC(in_0, in_1, in_2, out_0);
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  csa_tree_add_178_36_group_6829_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_181_36_group_6825_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_242, n_243;
  wire n_244, n_245, n_246, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_255, n_256, n_257, n_258, n_259, n_261, n_262;
  wire n_263, n_264, n_265, n_267, n_268, n_269, n_270, n_271;
  wire n_273, n_274, n_275, n_276, n_277, n_279, n_280, n_281;
  wire n_282, n_283, n_285, n_286, n_287, n_288, n_289, n_291;
  wire n_292, n_293, n_294, n_295, n_297, n_298, n_299, n_300;
  wire n_301, n_303, n_304, n_305, n_306, n_307, n_309, n_310;
  wire n_311, n_312, n_313, n_315, n_316, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_325, n_327, n_329, n_330, n_332;
  wire n_333, n_335, n_337, n_339, n_340, n_342, n_343, n_345;
  wire n_347, n_349, n_350, n_352, n_353, n_355, n_357, n_359;
  wire n_360, n_362, n_363, n_365, n_367, n_369, n_370, n_372;
  wire n_374, n_375, n_376, n_378, n_379, n_380, n_382, n_383;
  wire n_384, n_385, n_387, n_389, n_391, n_392, n_393, n_395;
  wire n_396, n_397, n_399, n_400, n_402, n_404, n_406, n_407;
  wire n_408, n_410, n_411, n_412, n_414, n_416, n_417, n_418;
  wire n_420, n_421, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_441, n_443, n_444, n_445, n_447;
  wire n_448, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_464, n_465;
  wire n_466, n_468, n_469, n_470, n_471, n_473, n_474, n_475;
  wire n_477, n_478, n_479, n_480, n_482, n_483, n_485, n_486;
  wire n_488, n_489, n_490, n_491, n_493, n_494, n_495, n_497;
  wire n_498, n_499, n_500, n_502, n_503, n_505, n_506, n_508;
  wire n_509, n_510, n_511, n_513, n_514, n_515, n_516, n_517;
  xor g26 (n_125, in_2[1], in_0[1]);
  and g2 (n_153, in_2[1], in_0[1]);
  xor g27 (n_123, in_2[2], n_153);
  xor g28 (n_149, n_123, in_0[2]);
  nand g3 (n_124, in_2[2], n_153);
  nand g29 (n_158, in_0[2], n_153);
  nand g30 (n_126, in_2[2], in_0[2]);
  nand g31 (n_154, n_124, n_158, n_126);
  xor g32 (n_159, in_2[3], in_0[3]);
  xor g33 (n_148, n_159, n_154);
  nand g34 (n_160, in_2[3], in_0[3]);
  nand g4 (n_161, n_154, in_0[3]);
  nand g35 (n_162, in_2[3], n_154);
  nand g36 (n_122, n_160, n_161, n_162);
  xor g37 (n_163, in_2[4], in_0[4]);
  xor g38 (n_147, n_163, in_1[4]);
  nand g39 (n_164, in_2[4], in_0[4]);
  nand g40 (n_165, in_1[4], in_0[4]);
  nand g5 (n_166, in_2[4], in_1[4]);
  nand g41 (n_121, n_164, n_165, n_166);
  xor g42 (n_167, in_2[5], in_0[5]);
  xor g43 (n_146, n_167, in_1[5]);
  nand g44 (n_168, in_2[5], in_0[5]);
  nand g45 (n_169, in_1[5], in_0[5]);
  nand g46 (n_170, in_2[5], in_1[5]);
  nand g6 (n_120, n_168, n_169, n_170);
  xor g47 (n_171, in_2[6], in_0[6]);
  xor g48 (n_145, n_171, in_1[6]);
  nand g49 (n_172, in_2[6], in_0[6]);
  nand g50 (n_173, in_1[6], in_0[6]);
  nand g51 (n_174, in_2[6], in_1[6]);
  nand g52 (n_119, n_172, n_173, n_174);
  xor g53 (n_175, in_2[7], in_0[7]);
  xor g54 (n_144, n_175, in_1[7]);
  nand g55 (n_176, in_2[7], in_0[7]);
  nand g56 (n_177, in_1[7], in_0[7]);
  nand g57 (n_178, in_2[7], in_1[7]);
  nand g58 (n_118, n_176, n_177, n_178);
  xor g59 (n_179, in_2[8], in_0[8]);
  xor g60 (n_143, n_179, in_1[8]);
  nand g61 (n_180, in_2[8], in_0[8]);
  nand g62 (n_181, in_1[8], in_0[8]);
  nand g63 (n_150, in_2[8], in_1[8]);
  nand g64 (n_117, n_180, n_181, n_150);
  xor g65 (n_151, in_2[9], in_0[9]);
  xor g66 (n_142, n_151, in_1[9]);
  nand g67 (n_152, in_2[9], in_0[9]);
  nand g68 (n_182, in_1[9], in_0[9]);
  nand g69 (n_183, in_2[9], in_1[9]);
  nand g70 (n_116, n_152, n_182, n_183);
  xor g71 (n_184, in_2[10], in_0[10]);
  xor g72 (n_141, n_184, in_1[10]);
  nand g73 (n_185, in_2[10], in_0[10]);
  nand g74 (n_186, in_1[10], in_0[10]);
  nand g75 (n_187, in_2[10], in_1[10]);
  nand g76 (n_115, n_185, n_186, n_187);
  xor g77 (n_188, in_2[11], in_0[11]);
  xor g78 (n_140, n_188, in_1[11]);
  nand g79 (n_189, in_2[11], in_0[11]);
  nand g80 (n_190, in_1[11], in_0[11]);
  nand g81 (n_191, in_2[11], in_1[11]);
  nand g82 (n_114, n_189, n_190, n_191);
  xor g83 (n_192, in_2[12], in_0[12]);
  xor g84 (n_139, n_192, in_1[12]);
  nand g85 (n_193, in_2[12], in_0[12]);
  nand g86 (n_194, in_1[12], in_0[12]);
  nand g87 (n_195, in_2[12], in_1[12]);
  nand g88 (n_113, n_193, n_194, n_195);
  xor g89 (n_196, in_2[13], in_0[13]);
  xor g90 (n_138, n_196, in_1[13]);
  nand g91 (n_197, in_2[13], in_0[13]);
  nand g92 (n_198, in_1[13], in_0[13]);
  nand g93 (n_199, in_2[13], in_1[13]);
  nand g94 (n_112, n_197, n_198, n_199);
  xor g95 (n_200, in_2[14], in_0[14]);
  xor g96 (n_137, n_200, in_1[14]);
  nand g97 (n_201, in_2[14], in_0[14]);
  nand g98 (n_202, in_1[14], in_0[14]);
  nand g99 (n_203, in_2[14], in_1[14]);
  nand g100 (n_111, n_201, n_202, n_203);
  xor g101 (n_204, in_2[15], in_0[15]);
  xor g102 (n_136, n_204, in_1[15]);
  nand g103 (n_205, in_2[15], in_0[15]);
  nand g104 (n_206, in_1[15], in_0[15]);
  nand g105 (n_207, in_2[15], in_1[15]);
  nand g106 (n_110, n_205, n_206, n_207);
  xor g107 (n_208, in_2[16], in_0[16]);
  xor g108 (n_135, n_208, in_1[16]);
  nand g109 (n_209, in_2[16], in_0[16]);
  nand g110 (n_210, in_1[16], in_0[16]);
  nand g111 (n_211, in_2[16], in_1[16]);
  nand g112 (n_109, n_209, n_210, n_211);
  xor g113 (n_212, in_2[17], in_0[17]);
  xor g114 (n_134, n_212, in_1[17]);
  nand g115 (n_213, in_2[17], in_0[17]);
  nand g116 (n_214, in_1[17], in_0[17]);
  nand g117 (n_215, in_2[17], in_1[17]);
  nand g118 (n_108, n_213, n_214, n_215);
  xor g119 (n_216, in_2[18], in_0[18]);
  xor g120 (n_133, n_216, in_1[18]);
  nand g121 (n_217, in_2[18], in_0[18]);
  nand g122 (n_218, in_1[18], in_0[18]);
  nand g123 (n_219, in_2[18], in_1[18]);
  nand g124 (n_107, n_217, n_218, n_219);
  xor g125 (n_220, in_2[19], in_0[19]);
  xor g126 (n_132, n_220, in_1[19]);
  nand g127 (n_221, in_2[19], in_0[19]);
  nand g128 (n_222, in_1[19], in_0[19]);
  nand g129 (n_223, in_2[19], in_1[19]);
  nand g130 (n_106, n_221, n_222, n_223);
  xor g131 (n_224, in_2[20], in_0[20]);
  xor g132 (n_131, n_224, in_1[20]);
  nand g133 (n_225, in_2[20], in_0[20]);
  nand g134 (n_226, in_1[20], in_0[20]);
  nand g135 (n_227, in_2[20], in_1[20]);
  nand g136 (n_105, n_225, n_226, n_227);
  xor g137 (n_228, in_2[21], in_0[21]);
  xor g138 (n_130, n_228, in_1[21]);
  nand g139 (n_229, in_2[21], in_0[21]);
  nand g140 (n_230, in_1[21], in_0[21]);
  nand g141 (n_231, in_2[21], in_1[21]);
  nand g142 (n_104, n_229, n_230, n_231);
  xor g143 (n_232, in_2[22], in_0[22]);
  xor g144 (n_129, n_232, in_1[22]);
  nand g145 (n_233, in_2[22], in_0[22]);
  nand g146 (n_234, in_1[22], in_0[22]);
  nand g147 (n_235, in_2[22], in_1[22]);
  nand g148 (n_103, n_233, n_234, n_235);
  xor g151 (n_236, in_2[23], in_1[23]);
  xor g152 (n_128, n_236, in_0[23]);
  nand g153 (n_237, in_2[23], in_1[23]);
  nand g154 (n_238, in_0[23], in_1[23]);
  nand g155 (n_239, in_2[23], in_0[23]);
  nand g156 (n_127, n_237, n_238, n_239);
  xor g159 (n_517, in_1[0], in_0[0]);
  nand g160 (n_242, in_1[0], in_0[0]);
  nand g161 (n_243, in_1[0], in_2[0]);
  nand g7 (n_244, in_0[0], in_2[0]);
  nand g8 (n_246, n_242, n_243, n_244);
  nor g9 (n_245, n_125, in_1[1]);
  nand g10 (n_248, n_125, in_1[1]);
  nor g11 (n_255, in_1[2], n_149);
  nand g12 (n_250, in_1[2], n_149);
  nor g13 (n_251, in_1[3], n_148);
  nand g14 (n_252, in_1[3], n_148);
  nor g15 (n_261, n_122, n_147);
  nand g16 (n_256, n_122, n_147);
  nor g17 (n_257, n_121, n_146);
  nand g18 (n_258, n_121, n_146);
  nor g19 (n_267, n_120, n_145);
  nand g20 (n_262, n_120, n_145);
  nor g21 (n_263, n_119, n_144);
  nand g22 (n_264, n_119, n_144);
  nor g23 (n_273, n_118, n_143);
  nand g24 (n_268, n_118, n_143);
  nor g25 (n_269, n_117, n_142);
  nand g162 (n_270, n_117, n_142);
  nor g163 (n_279, n_116, n_141);
  nand g164 (n_274, n_116, n_141);
  nor g165 (n_275, n_115, n_140);
  nand g166 (n_276, n_115, n_140);
  nor g167 (n_285, n_114, n_139);
  nand g168 (n_280, n_114, n_139);
  nor g169 (n_281, n_113, n_138);
  nand g170 (n_282, n_113, n_138);
  nor g171 (n_291, n_112, n_137);
  nand g172 (n_286, n_112, n_137);
  nor g173 (n_287, n_111, n_136);
  nand g174 (n_288, n_111, n_136);
  nor g175 (n_297, n_110, n_135);
  nand g176 (n_292, n_110, n_135);
  nor g177 (n_293, n_109, n_134);
  nand g178 (n_294, n_109, n_134);
  nor g179 (n_303, n_108, n_133);
  nand g180 (n_298, n_108, n_133);
  nor g181 (n_299, n_107, n_132);
  nand g182 (n_300, n_107, n_132);
  nor g183 (n_309, n_106, n_131);
  nand g184 (n_304, n_106, n_131);
  nor g185 (n_305, n_105, n_130);
  nand g186 (n_306, n_105, n_130);
  nor g187 (n_315, n_104, n_129);
  nand g188 (n_310, n_104, n_129);
  nor g189 (n_311, n_103, n_128);
  nand g190 (n_312, n_103, n_128);
  nand g195 (n_316, n_248, n_249);
  nor g196 (n_253, n_250, n_251);
  nor g199 (n_319, n_255, n_251);
  nor g200 (n_259, n_256, n_257);
  nor g203 (n_325, n_261, n_257);
  nor g204 (n_265, n_262, n_263);
  nor g207 (n_327, n_267, n_263);
  nor g208 (n_271, n_268, n_269);
  nor g211 (n_335, n_273, n_269);
  nor g212 (n_277, n_274, n_275);
  nor g215 (n_337, n_279, n_275);
  nor g216 (n_283, n_280, n_281);
  nor g219 (n_345, n_285, n_281);
  nor g220 (n_289, n_286, n_287);
  nor g223 (n_347, n_291, n_287);
  nor g224 (n_295, n_292, n_293);
  nor g227 (n_355, n_297, n_293);
  nor g228 (n_301, n_298, n_299);
  nor g231 (n_357, n_303, n_299);
  nor g232 (n_307, n_304, n_305);
  nor g235 (n_365, n_309, n_305);
  nor g236 (n_313, n_310, n_311);
  nor g239 (n_367, n_315, n_311);
  nand g242 (n_464, n_250, n_318);
  nand g243 (n_321, n_319, n_316);
  nand g244 (n_372, n_320, n_321);
  nor g245 (n_323, n_267, n_322);
  nand g254 (n_380, n_325, n_327);
  nor g255 (n_333, n_279, n_332);
  nand g264 (n_387, n_335, n_337);
  nor g265 (n_343, n_291, n_342);
  nand g274 (n_395, n_345, n_347);
  nor g275 (n_353, n_303, n_352);
  nand g284 (n_402, n_355, n_357);
  nor g285 (n_363, n_315, n_362);
  nand g294 (n_410, n_365, n_367);
  nand g297 (n_468, n_256, n_374);
  nand g298 (n_375, n_325, n_372);
  nand g299 (n_470, n_322, n_375);
  nand g302 (n_473, n_378, n_379);
  nand g305 (n_414, n_382, n_383);
  nor g306 (n_385, n_285, n_384);
  nor g309 (n_424, n_285, n_387);
  nor g315 (n_393, n_391, n_384);
  nor g318 (n_430, n_387, n_391);
  nor g319 (n_397, n_395, n_384);
  nor g322 (n_433, n_387, n_395);
  nor g323 (n_400, n_309, n_399);
  nor g326 (n_451, n_309, n_402);
  nor g332 (n_408, n_406, n_399);
  nor g335 (n_457, n_402, n_406);
  nor g336 (n_412, n_410, n_399);
  nor g339 (n_439, n_402, n_410);
  nand g342 (n_477, n_268, n_416);
  nand g343 (n_417, n_335, n_414);
  nand g344 (n_479, n_332, n_417);
  nand g347 (n_482, n_420, n_421);
  nand g350 (n_485, n_384, n_423);
  nand g351 (n_426, n_424, n_414);
  nand g352 (n_488, n_425, n_426);
  nand g353 (n_429, n_427, n_414);
  nand g354 (n_490, n_428, n_429);
  nand g355 (n_432, n_430, n_414);
  nand g356 (n_493, n_431, n_432);
  nand g357 (n_435, n_433, n_414);
  nand g358 (n_441, n_434, n_435);
  nand g362 (n_497, n_292, n_443);
  nand g363 (n_444, n_355, n_441);
  nand g364 (n_499, n_352, n_444);
  nand g367 (n_502, n_447, n_448);
  nand g370 (n_505, n_399, n_450);
  nand g371 (n_453, n_451, n_441);
  nand g372 (n_508, n_452, n_453);
  nand g373 (n_456, n_454, n_441);
  nand g374 (n_510, n_455, n_456);
  nand g375 (n_459, n_457, n_441);
  nand g376 (n_513, n_458, n_459);
  nand g377 (n_460, n_439, n_441);
  nand g378 (n_515, n_437, n_460);
  xnor g380 (out_0[1], n_246, n_461);
  xnor g382 (out_0[2], n_316, n_462);
  xnor g385 (out_0[3], n_464, n_465);
  xnor g387 (out_0[4], n_372, n_466);
  xnor g390 (out_0[5], n_468, n_469);
  xnor g392 (out_0[6], n_470, n_471);
  xnor g395 (out_0[7], n_473, n_474);
  xnor g397 (out_0[8], n_414, n_475);
  xnor g400 (out_0[9], n_477, n_478);
  xnor g402 (out_0[10], n_479, n_480);
  xnor g405 (out_0[11], n_482, n_483);
  xnor g408 (out_0[12], n_485, n_486);
  xnor g411 (out_0[13], n_488, n_489);
  xnor g413 (out_0[14], n_490, n_491);
  xnor g416 (out_0[15], n_493, n_494);
  xnor g418 (out_0[16], n_441, n_495);
  xnor g421 (out_0[17], n_497, n_498);
  xnor g423 (out_0[18], n_499, n_500);
  xnor g426 (out_0[19], n_502, n_503);
  xnor g429 (out_0[20], n_505, n_506);
  xnor g432 (out_0[21], n_508, n_509);
  xnor g434 (out_0[22], n_510, n_511);
  xnor g437 (out_0[23], n_513, n_514);
  xnor g439 (out_0[24], n_515, n_516);
  xor g440 (out_0[0], in_2[0], n_517);
  or g441 (n_249, n_245, wc);
  not gc (wc, n_246);
  or g442 (n_461, wc0, n_245);
  not gc0 (wc0, n_248);
  and g443 (n_329, wc1, n_264);
  not gc1 (wc1, n_265);
  and g444 (n_332, wc2, n_270);
  not gc2 (wc2, n_271);
  and g445 (n_339, wc3, n_276);
  not gc3 (wc3, n_277);
  and g446 (n_342, wc4, n_282);
  not gc4 (wc4, n_283);
  and g447 (n_349, wc5, n_288);
  not gc5 (wc5, n_289);
  and g448 (n_352, wc6, n_294);
  not gc6 (wc6, n_295);
  and g449 (n_359, wc7, n_300);
  not gc7 (wc7, n_301);
  and g450 (n_362, wc8, n_306);
  not gc8 (wc8, n_307);
  or g451 (n_418, wc9, n_279);
  not gc9 (wc9, n_335);
  or g452 (n_391, wc10, n_291);
  not gc10 (wc10, n_345);
  or g453 (n_445, wc11, n_303);
  not gc11 (wc11, n_355);
  or g454 (n_406, wc12, n_315);
  not gc12 (wc12, n_365);
  or g455 (n_469, wc13, n_257);
  not gc13 (wc13, n_258);
  or g456 (n_471, wc14, n_267);
  not gc14 (wc14, n_262);
  or g457 (n_474, wc15, n_263);
  not gc15 (wc15, n_264);
  or g458 (n_475, wc16, n_273);
  not gc16 (wc16, n_268);
  or g459 (n_478, wc17, n_269);
  not gc17 (wc17, n_270);
  or g460 (n_480, wc18, n_279);
  not gc18 (wc18, n_274);
  or g461 (n_483, wc19, n_275);
  not gc19 (wc19, n_276);
  or g462 (n_486, wc20, n_285);
  not gc20 (wc20, n_280);
  or g463 (n_489, wc21, n_281);
  not gc21 (wc21, n_282);
  or g464 (n_491, wc22, n_291);
  not gc22 (wc22, n_286);
  or g465 (n_494, wc23, n_287);
  not gc23 (wc23, n_288);
  or g466 (n_495, wc24, n_297);
  not gc24 (wc24, n_292);
  or g467 (n_498, wc25, n_293);
  not gc25 (wc25, n_294);
  or g468 (n_500, wc26, n_303);
  not gc26 (wc26, n_298);
  or g469 (n_503, wc27, n_299);
  not gc27 (wc27, n_300);
  or g470 (n_506, wc28, n_309);
  not gc28 (wc28, n_304);
  or g471 (n_509, wc29, n_305);
  not gc29 (wc29, n_306);
  or g472 (n_511, wc30, n_315);
  not gc30 (wc30, n_310);
  and g473 (n_436, wc31, n_127);
  not gc31 (wc31, in_2[23]);
  or g474 (n_438, wc32, n_127);
  not gc32 (wc32, in_2[23]);
  or g475 (n_318, wc33, n_255);
  not gc33 (wc33, n_316);
  and g476 (n_340, wc34, n_337);
  not gc34 (wc34, n_332);
  and g477 (n_350, wc35, n_347);
  not gc35 (wc35, n_342);
  and g478 (n_360, wc36, n_357);
  not gc36 (wc36, n_352);
  and g479 (n_427, wc37, n_345);
  not gc37 (wc37, n_387);
  and g480 (n_454, wc38, n_365);
  not gc38 (wc38, n_402);
  or g481 (n_462, wc39, n_255);
  not gc39 (wc39, n_250);
  and g482 (n_320, wc40, n_252);
  not gc40 (wc40, n_253);
  and g483 (n_369, wc41, n_312);
  not gc41 (wc41, n_313);
  and g484 (n_420, wc42, n_274);
  not gc42 (wc42, n_333);
  and g485 (n_384, wc43, n_339);
  not gc43 (wc43, n_340);
  and g486 (n_392, wc44, n_286);
  not gc44 (wc44, n_343);
  and g487 (n_396, wc45, n_349);
  not gc45 (wc45, n_350);
  and g488 (n_447, wc46, n_298);
  not gc46 (wc46, n_353);
  and g489 (n_399, wc47, n_359);
  not gc47 (wc47, n_360);
  and g490 (n_407, wc48, n_310);
  not gc48 (wc48, n_363);
  or g491 (n_465, wc49, n_251);
  not gc49 (wc49, n_252);
  or g492 (n_514, wc50, n_311);
  not gc50 (wc50, n_312);
  and g493 (n_322, wc51, n_258);
  not gc51 (wc51, n_259);
  or g494 (n_376, wc52, n_267);
  not gc52 (wc52, n_325);
  and g495 (n_370, wc53, n_367);
  not gc53 (wc53, n_362);
  and g496 (n_389, wc54, n_345);
  not gc54 (wc54, n_384);
  and g497 (n_404, wc55, n_365);
  not gc55 (wc55, n_399);
  or g498 (n_466, wc56, n_261);
  not gc56 (wc56, n_256);
  or g499 (n_516, wc57, n_436);
  not gc57 (wc57, n_438);
  and g500 (n_330, wc58, n_327);
  not gc58 (wc58, n_322);
  and g501 (n_411, wc59, n_369);
  not gc59 (wc59, n_370);
  or g502 (n_374, wc60, n_261);
  not gc60 (wc60, n_372);
  and g503 (n_425, wc61, n_280);
  not gc61 (wc61, n_385);
  and g504 (n_428, wc62, n_342);
  not gc62 (wc62, n_389);
  and g505 (n_431, n_392, wc63);
  not gc63 (wc63, n_393);
  and g506 (n_434, n_396, wc64);
  not gc64 (wc64, n_397);
  and g507 (n_452, wc65, n_304);
  not gc65 (wc65, n_400);
  and g508 (n_455, wc66, n_362);
  not gc66 (wc66, n_404);
  and g509 (n_458, n_407, wc67);
  not gc67 (wc67, n_408);
  and g510 (n_378, wc68, n_262);
  not gc68 (wc68, n_323);
  and g511 (n_382, wc69, n_329);
  not gc69 (wc69, n_330);
  or g512 (n_379, n_376, wc70);
  not gc70 (wc70, n_372);
  or g513 (n_383, n_380, wc71);
  not gc71 (wc71, n_372);
  and g514 (n_437, n_411, wc72);
  not gc72 (wc72, n_412);
  or g515 (n_416, wc73, n_273);
  not gc73 (wc73, n_414);
  or g516 (n_421, n_418, wc74);
  not gc74 (wc74, n_414);
  or g517 (n_423, wc75, n_387);
  not gc75 (wc75, n_414);
  or g518 (n_443, wc76, n_297);
  not gc76 (wc76, n_441);
  or g519 (n_448, n_445, wc77);
  not gc77 (wc77, n_441);
  or g520 (n_450, wc78, n_402);
  not gc78 (wc78, n_441);
endmodule

module csa_tree_add_181_36_group_6825_GENERIC(in_0, in_1, in_2, out_0);
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  csa_tree_add_181_36_group_6825_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_255_42_group_6823_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [20:0] in_0, in_1, in_2, in_3, in_4;
  output [23:0] out_0;
  wire [20:0] in_0, in_1, in_2, in_3, in_4;
  wire [23:0] out_0;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213;
  wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_250, n_256, n_257, n_258;
  wire n_259, n_260, n_263, n_265, n_266, n_267, n_268, n_269;
  wire n_270, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_285;
  wire n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_294, n_295, n_296, n_297, n_298, n_299, n_300, n_301;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317;
  wire n_318, n_319, n_320, n_321, n_322, n_323, n_324, n_325;
  wire n_326, n_327, n_328, n_329, n_330, n_331, n_332, n_333;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349;
  wire n_350, n_351, n_352, n_353, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373;
  wire n_374, n_375, n_376, n_377, n_378, n_379, n_380, n_381;
  wire n_382, n_383, n_384, n_385, n_386, n_387, n_388, n_389;
  wire n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397;
  wire n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405;
  wire n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413;
  wire n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421;
  wire n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429;
  wire n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437;
  wire n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445;
  wire n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453;
  wire n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461;
  wire n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477;
  wire n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485;
  wire n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_496, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_508, n_509, n_510, n_511, n_512, n_514, n_515;
  wire n_516, n_517, n_518, n_519, n_521, n_522, n_523, n_524;
  wire n_525, n_527, n_528, n_529, n_530, n_531, n_533, n_534;
  wire n_535, n_536, n_537, n_539, n_540, n_541, n_542, n_543;
  wire n_545, n_546, n_547, n_548, n_549, n_551, n_552, n_553;
  wire n_554, n_555, n_557, n_558, n_559, n_560, n_561, n_563;
  wire n_564, n_565, n_566, n_567, n_569, n_570, n_571, n_572;
  wire n_573, n_575, n_576, n_579, n_580, n_581, n_582, n_583;
  wire n_584, n_585, n_586, n_588, n_590, n_592, n_593, n_595;
  wire n_596, n_598, n_600, n_602, n_603, n_605, n_606, n_608;
  wire n_610, n_612, n_613, n_615, n_616, n_618, n_620, n_622;
  wire n_623, n_625, n_626, n_628, n_630, n_632, n_633, n_634;
  wire n_636, n_637, n_638, n_640, n_641, n_642, n_643, n_645;
  wire n_647, n_649, n_650, n_651, n_653, n_654, n_655, n_657;
  wire n_658, n_660, n_662, n_664, n_665, n_666, n_668, n_670;
  wire n_671, n_672, n_674, n_675, n_677, n_678, n_679, n_680;
  wire n_681, n_682, n_683, n_684, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_692, n_693, n_694, n_696, n_697, n_699;
  wire n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_712, n_713, n_714, n_716, n_717;
  wire n_718, n_719, n_721, n_722, n_723, n_725, n_726, n_727;
  wire n_728, n_730, n_731, n_733, n_734, n_736, n_737, n_738;
  wire n_739, n_741, n_742, n_743, n_745, n_746, n_747, n_748;
  wire n_750, n_751, n_753, n_754, n_756, n_757, n_758, n_759;
  wire n_761, n_763;
  xor g69 (n_266, in_0[0], in_4[0]);
  xor g70 (n_177, n_266, in_3[0]);
  nand g71 (n_267, in_0[0], in_4[0]);
  nand g72 (n_268, in_3[0], in_4[0]);
  nand g73 (n_269, in_0[0], in_3[0]);
  nand g6 (n_179, n_267, n_268, n_269);
  xor g74 (n_270, in_0[1], in_1[1]);
  xor g75 (n_152, n_270, in_4[1]);
  nand g76 (n_271, in_0[1], in_1[1]);
  nand g77 (n_272, in_4[1], in_1[1]);
  nand g78 (n_273, in_0[1], in_4[1]);
  nand g79 (n_181, n_271, n_272, n_273);
  xor g80 (n_274, in_3[1], in_2[1]);
  xor g81 (n_176, n_274, n_179);
  nand g82 (n_275, in_3[1], in_2[1]);
  nand g83 (n_276, n_179, in_2[1]);
  nand g84 (n_277, in_3[1], n_179);
  nand g85 (n_151, n_275, n_276, n_277);
  xor g86 (n_180, in_0[2], in_1[2]);
  and g87 (n_183, in_0[2], in_1[2]);
  xor g88 (n_278, in_3[2], in_4[2]);
  xor g89 (n_182, n_278, in_2[2]);
  nand g90 (n_279, in_3[2], in_4[2]);
  nand g91 (n_280, in_2[2], in_4[2]);
  nand g92 (n_281, in_3[2], in_2[2]);
  nand g93 (n_184, n_279, n_280, n_281);
  xor g94 (n_282, n_180, n_181);
  xor g95 (n_175, n_282, n_182);
  nand g96 (n_283, n_180, n_181);
  nand g97 (n_284, n_182, n_181);
  nand g98 (n_285, n_180, n_182);
  nand g99 (n_150, n_283, n_284, n_285);
  xor g100 (n_286, in_0[3], in_1[3]);
  xor g101 (n_185, n_286, in_3[3]);
  nand g102 (n_287, in_0[3], in_1[3]);
  nand g103 (n_288, in_3[3], in_1[3]);
  nand g104 (n_289, in_0[3], in_3[3]);
  nand g105 (n_187, n_287, n_288, n_289);
  xor g106 (n_290, in_4[3], in_2[3]);
  xor g107 (n_186, n_290, n_183);
  nand g108 (n_291, in_4[3], in_2[3]);
  nand g109 (n_292, n_183, in_2[3]);
  nand g110 (n_293, in_4[3], n_183);
  nand g111 (n_189, n_291, n_292, n_293);
  xor g112 (n_294, n_184, n_185);
  xor g113 (n_174, n_294, n_186);
  nand g114 (n_295, n_184, n_185);
  nand g115 (n_296, n_186, n_185);
  nand g116 (n_297, n_184, n_186);
  nand g117 (n_149, n_295, n_296, n_297);
  xor g118 (n_298, in_0[4], in_1[4]);
  xor g119 (n_188, n_298, in_3[4]);
  nand g120 (n_299, in_0[4], in_1[4]);
  nand g121 (n_300, in_3[4], in_1[4]);
  nand g122 (n_301, in_0[4], in_3[4]);
  nand g123 (n_191, n_299, n_300, n_301);
  xor g124 (n_302, in_4[4], in_2[4]);
  xor g125 (n_190, n_302, n_187);
  nand g126 (n_303, in_4[4], in_2[4]);
  nand g127 (n_304, n_187, in_2[4]);
  nand g128 (n_305, in_4[4], n_187);
  nand g129 (n_194, n_303, n_304, n_305);
  xor g130 (n_306, n_188, n_189);
  xor g131 (n_173, n_306, n_190);
  nand g132 (n_307, n_188, n_189);
  nand g133 (n_308, n_190, n_189);
  nand g134 (n_309, n_188, n_190);
  nand g135 (n_148, n_307, n_308, n_309);
  xor g136 (n_310, in_0[5], in_1[5]);
  xor g137 (n_192, n_310, in_3[5]);
  nand g138 (n_311, in_0[5], in_1[5]);
  nand g139 (n_312, in_3[5], in_1[5]);
  nand g140 (n_313, in_0[5], in_3[5]);
  nand g141 (n_195, n_311, n_312, n_313);
  xor g142 (n_314, in_4[5], in_2[5]);
  xor g143 (n_193, n_314, n_191);
  nand g144 (n_315, in_4[5], in_2[5]);
  nand g145 (n_316, n_191, in_2[5]);
  nand g146 (n_317, in_4[5], n_191);
  nand g147 (n_198, n_315, n_316, n_317);
  xor g148 (n_318, n_192, n_193);
  xor g149 (n_172, n_318, n_194);
  nand g150 (n_319, n_192, n_193);
  nand g151 (n_320, n_194, n_193);
  nand g152 (n_321, n_192, n_194);
  nand g153 (n_147, n_319, n_320, n_321);
  xor g154 (n_322, in_0[6], in_1[6]);
  xor g155 (n_196, n_322, in_3[6]);
  nand g156 (n_323, in_0[6], in_1[6]);
  nand g157 (n_324, in_3[6], in_1[6]);
  nand g158 (n_325, in_0[6], in_3[6]);
  nand g159 (n_199, n_323, n_324, n_325);
  xor g160 (n_326, in_4[6], in_2[6]);
  xor g161 (n_197, n_326, n_195);
  nand g162 (n_327, in_4[6], in_2[6]);
  nand g163 (n_328, n_195, in_2[6]);
  nand g164 (n_329, in_4[6], n_195);
  nand g165 (n_202, n_327, n_328, n_329);
  xor g166 (n_330, n_196, n_197);
  xor g167 (n_171, n_330, n_198);
  nand g168 (n_331, n_196, n_197);
  nand g169 (n_332, n_198, n_197);
  nand g170 (n_333, n_196, n_198);
  nand g171 (n_146, n_331, n_332, n_333);
  xor g172 (n_334, in_0[7], in_1[7]);
  xor g173 (n_200, n_334, in_3[7]);
  nand g174 (n_335, in_0[7], in_1[7]);
  nand g175 (n_336, in_3[7], in_1[7]);
  nand g176 (n_337, in_0[7], in_3[7]);
  nand g177 (n_203, n_335, n_336, n_337);
  xor g178 (n_338, in_4[7], in_2[7]);
  xor g179 (n_201, n_338, n_199);
  nand g180 (n_339, in_4[7], in_2[7]);
  nand g181 (n_340, n_199, in_2[7]);
  nand g182 (n_341, in_4[7], n_199);
  nand g183 (n_206, n_339, n_340, n_341);
  xor g184 (n_342, n_200, n_201);
  xor g185 (n_170, n_342, n_202);
  nand g186 (n_343, n_200, n_201);
  nand g187 (n_344, n_202, n_201);
  nand g188 (n_345, n_200, n_202);
  nand g189 (n_145, n_343, n_344, n_345);
  xor g190 (n_346, in_0[8], in_1[8]);
  xor g191 (n_204, n_346, in_3[8]);
  nand g192 (n_347, in_0[8], in_1[8]);
  nand g193 (n_348, in_3[8], in_1[8]);
  nand g194 (n_349, in_0[8], in_3[8]);
  nand g195 (n_207, n_347, n_348, n_349);
  xor g196 (n_350, in_4[8], in_2[8]);
  xor g197 (n_205, n_350, n_203);
  nand g198 (n_351, in_4[8], in_2[8]);
  nand g199 (n_352, n_203, in_2[8]);
  nand g200 (n_353, in_4[8], n_203);
  nand g201 (n_210, n_351, n_352, n_353);
  xor g202 (n_354, n_204, n_205);
  xor g203 (n_169, n_354, n_206);
  nand g204 (n_355, n_204, n_205);
  nand g205 (n_356, n_206, n_205);
  nand g206 (n_357, n_204, n_206);
  nand g207 (n_144, n_355, n_356, n_357);
  xor g208 (n_358, in_0[9], in_1[9]);
  xor g209 (n_208, n_358, in_3[9]);
  nand g210 (n_359, in_0[9], in_1[9]);
  nand g211 (n_360, in_3[9], in_1[9]);
  nand g212 (n_361, in_0[9], in_3[9]);
  nand g213 (n_211, n_359, n_360, n_361);
  xor g214 (n_362, in_4[9], in_2[9]);
  xor g215 (n_209, n_362, n_207);
  nand g216 (n_363, in_4[9], in_2[9]);
  nand g217 (n_364, n_207, in_2[9]);
  nand g218 (n_365, in_4[9], n_207);
  nand g219 (n_214, n_363, n_364, n_365);
  xor g220 (n_366, n_208, n_209);
  xor g221 (n_168, n_366, n_210);
  nand g222 (n_367, n_208, n_209);
  nand g223 (n_368, n_210, n_209);
  nand g224 (n_369, n_208, n_210);
  nand g225 (n_143, n_367, n_368, n_369);
  xor g226 (n_370, in_0[10], in_1[10]);
  xor g227 (n_212, n_370, in_3[10]);
  nand g228 (n_371, in_0[10], in_1[10]);
  nand g229 (n_372, in_3[10], in_1[10]);
  nand g230 (n_373, in_0[10], in_3[10]);
  nand g231 (n_215, n_371, n_372, n_373);
  xor g232 (n_374, in_4[10], in_2[10]);
  xor g233 (n_213, n_374, n_211);
  nand g234 (n_375, in_4[10], in_2[10]);
  nand g235 (n_376, n_211, in_2[10]);
  nand g236 (n_377, in_4[10], n_211);
  nand g237 (n_218, n_375, n_376, n_377);
  xor g238 (n_378, n_212, n_213);
  xor g239 (n_167, n_378, n_214);
  nand g240 (n_379, n_212, n_213);
  nand g241 (n_380, n_214, n_213);
  nand g242 (n_381, n_212, n_214);
  nand g243 (n_142, n_379, n_380, n_381);
  xor g244 (n_382, in_0[11], in_1[11]);
  xor g245 (n_216, n_382, in_3[11]);
  nand g246 (n_383, in_0[11], in_1[11]);
  nand g247 (n_384, in_3[11], in_1[11]);
  nand g248 (n_385, in_0[11], in_3[11]);
  nand g249 (n_219, n_383, n_384, n_385);
  xor g250 (n_386, in_4[11], in_2[11]);
  xor g251 (n_217, n_386, n_215);
  nand g252 (n_387, in_4[11], in_2[11]);
  nand g253 (n_388, n_215, in_2[11]);
  nand g254 (n_389, in_4[11], n_215);
  nand g255 (n_222, n_387, n_388, n_389);
  xor g256 (n_390, n_216, n_217);
  xor g257 (n_166, n_390, n_218);
  nand g258 (n_391, n_216, n_217);
  nand g259 (n_392, n_218, n_217);
  nand g260 (n_393, n_216, n_218);
  nand g261 (n_141, n_391, n_392, n_393);
  xor g262 (n_394, in_0[12], in_1[12]);
  xor g263 (n_220, n_394, in_3[12]);
  nand g264 (n_395, in_0[12], in_1[12]);
  nand g265 (n_396, in_3[12], in_1[12]);
  nand g266 (n_397, in_0[12], in_3[12]);
  nand g267 (n_223, n_395, n_396, n_397);
  xor g268 (n_398, in_4[12], in_2[12]);
  xor g269 (n_221, n_398, n_219);
  nand g270 (n_399, in_4[12], in_2[12]);
  nand g271 (n_400, n_219, in_2[12]);
  nand g272 (n_401, in_4[12], n_219);
  nand g273 (n_226, n_399, n_400, n_401);
  xor g274 (n_402, n_220, n_221);
  xor g275 (n_165, n_402, n_222);
  nand g276 (n_403, n_220, n_221);
  nand g277 (n_404, n_222, n_221);
  nand g278 (n_405, n_220, n_222);
  nand g279 (n_140, n_403, n_404, n_405);
  xor g280 (n_406, in_0[13], in_1[13]);
  xor g281 (n_224, n_406, in_3[13]);
  nand g282 (n_407, in_0[13], in_1[13]);
  nand g283 (n_408, in_3[13], in_1[13]);
  nand g284 (n_409, in_0[13], in_3[13]);
  nand g285 (n_227, n_407, n_408, n_409);
  xor g286 (n_410, in_4[13], in_2[13]);
  xor g287 (n_225, n_410, n_223);
  nand g288 (n_411, in_4[13], in_2[13]);
  nand g289 (n_412, n_223, in_2[13]);
  nand g290 (n_413, in_4[13], n_223);
  nand g291 (n_230, n_411, n_412, n_413);
  xor g292 (n_414, n_224, n_225);
  xor g293 (n_164, n_414, n_226);
  nand g294 (n_415, n_224, n_225);
  nand g295 (n_416, n_226, n_225);
  nand g296 (n_417, n_224, n_226);
  nand g297 (n_139, n_415, n_416, n_417);
  xor g298 (n_418, in_0[14], in_1[14]);
  xor g299 (n_228, n_418, in_3[14]);
  nand g300 (n_419, in_0[14], in_1[14]);
  nand g301 (n_420, in_3[14], in_1[14]);
  nand g302 (n_421, in_0[14], in_3[14]);
  nand g303 (n_231, n_419, n_420, n_421);
  xor g304 (n_422, in_4[14], in_2[14]);
  xor g305 (n_229, n_422, n_227);
  nand g306 (n_423, in_4[14], in_2[14]);
  nand g307 (n_424, n_227, in_2[14]);
  nand g308 (n_425, in_4[14], n_227);
  nand g309 (n_234, n_423, n_424, n_425);
  xor g310 (n_426, n_228, n_229);
  xor g311 (n_163, n_426, n_230);
  nand g312 (n_427, n_228, n_229);
  nand g313 (n_428, n_230, n_229);
  nand g314 (n_429, n_228, n_230);
  nand g315 (n_138, n_427, n_428, n_429);
  xor g316 (n_430, in_0[15], in_1[15]);
  xor g317 (n_232, n_430, in_3[15]);
  nand g318 (n_431, in_0[15], in_1[15]);
  nand g319 (n_432, in_3[15], in_1[15]);
  nand g320 (n_433, in_0[15], in_3[15]);
  nand g321 (n_235, n_431, n_432, n_433);
  xor g322 (n_434, in_4[15], in_2[15]);
  xor g323 (n_233, n_434, n_231);
  nand g324 (n_435, in_4[15], in_2[15]);
  nand g325 (n_436, n_231, in_2[15]);
  nand g326 (n_437, in_4[15], n_231);
  nand g327 (n_238, n_435, n_436, n_437);
  xor g328 (n_438, n_232, n_233);
  xor g329 (n_162, n_438, n_234);
  nand g330 (n_439, n_232, n_233);
  nand g331 (n_440, n_234, n_233);
  nand g332 (n_441, n_232, n_234);
  nand g333 (n_137, n_439, n_440, n_441);
  xor g334 (n_442, in_0[16], in_1[16]);
  xor g335 (n_236, n_442, in_3[16]);
  nand g336 (n_443, in_0[16], in_1[16]);
  nand g337 (n_444, in_3[16], in_1[16]);
  nand g338 (n_445, in_0[16], in_3[16]);
  nand g339 (n_239, n_443, n_444, n_445);
  xor g340 (n_446, in_4[16], in_2[16]);
  xor g341 (n_237, n_446, n_235);
  nand g342 (n_447, in_4[16], in_2[16]);
  nand g343 (n_448, n_235, in_2[16]);
  nand g344 (n_449, in_4[16], n_235);
  nand g345 (n_242, n_447, n_448, n_449);
  xor g346 (n_450, n_236, n_237);
  xor g347 (n_161, n_450, n_238);
  nand g348 (n_451, n_236, n_237);
  nand g349 (n_452, n_238, n_237);
  nand g350 (n_453, n_236, n_238);
  nand g351 (n_136, n_451, n_452, n_453);
  xor g352 (n_454, in_0[17], in_1[17]);
  xor g353 (n_240, n_454, in_3[17]);
  nand g354 (n_455, in_0[17], in_1[17]);
  nand g355 (n_456, in_3[17], in_1[17]);
  nand g356 (n_457, in_0[17], in_3[17]);
  nand g357 (n_243, n_455, n_456, n_457);
  xor g358 (n_458, in_4[17], in_2[17]);
  xor g359 (n_241, n_458, n_239);
  nand g360 (n_459, in_4[17], in_2[17]);
  nand g361 (n_460, n_239, in_2[17]);
  nand g362 (n_461, in_4[17], n_239);
  nand g363 (n_246, n_459, n_460, n_461);
  xor g364 (n_462, n_240, n_241);
  xor g365 (n_160, n_462, n_242);
  nand g366 (n_463, n_240, n_241);
  nand g367 (n_464, n_242, n_241);
  nand g368 (n_465, n_240, n_242);
  nand g369 (n_135, n_463, n_464, n_465);
  xor g370 (n_466, in_0[18], in_1[18]);
  xor g371 (n_244, n_466, in_3[18]);
  nand g372 (n_467, in_0[18], in_1[18]);
  nand g373 (n_468, in_3[18], in_1[18]);
  nand g374 (n_469, in_0[18], in_3[18]);
  nand g375 (n_247, n_467, n_468, n_469);
  xor g376 (n_470, in_4[18], in_2[18]);
  xor g377 (n_245, n_470, n_243);
  nand g378 (n_471, in_4[18], in_2[18]);
  nand g379 (n_472, n_243, in_2[18]);
  nand g380 (n_473, in_4[18], n_243);
  nand g381 (n_250, n_471, n_472, n_473);
  xor g382 (n_474, n_244, n_245);
  xor g383 (n_159, n_474, n_246);
  nand g384 (n_475, n_244, n_245);
  nand g385 (n_476, n_246, n_245);
  nand g386 (n_477, n_244, n_246);
  nand g387 (n_134, n_475, n_476, n_477);
  xor g388 (n_478, in_0[19], in_1[19]);
  xor g389 (n_248, n_478, in_3[19]);
  nand g390 (n_479, in_0[19], in_1[19]);
  nand g391 (n_480, in_3[19], in_1[19]);
  nand g392 (n_481, in_0[19], in_3[19]);
  nand g393 (n_257, n_479, n_480, n_481);
  xor g394 (n_482, in_4[19], in_2[19]);
  xor g395 (n_249, n_482, n_247);
  nand g396 (n_483, in_4[19], in_2[19]);
  nand g397 (n_484, n_247, in_2[19]);
  nand g398 (n_485, in_4[19], n_247);
  nand g399 (n_260, n_483, n_484, n_485);
  xor g400 (n_486, n_248, n_249);
  xor g401 (n_158, n_486, n_250);
  nand g402 (n_487, n_248, n_249);
  nand g403 (n_488, n_250, n_249);
  nand g404 (n_489, n_248, n_250);
  nand g405 (n_133, n_487, n_488, n_489);
  nand g413 (n_263, n_491, n_492, n_493);
  nand g417 (n_496, n_257, n_256);
  xor g420 (n_498, n_258, n_259);
  xor g421 (n_157, n_498, n_260);
  nand g422 (n_499, n_258, n_259);
  nand g423 (n_500, n_260, n_259);
  nand g424 (n_501, n_258, n_260);
  nand g425 (n_132, n_499, n_500, n_501);
  xor g429 (n_156, n_502, n_265);
  nand g432 (n_505, n_263, n_265);
  nand g433 (n_155, n_503, n_504, n_505);
  xor g436 (n_763, in_1[0], n_177);
  nand g437 (n_508, in_1[0], n_177);
  nand g438 (n_509, in_1[0], in_2[0]);
  nand g7 (n_510, n_177, in_2[0]);
  nand g8 (n_512, n_508, n_509, n_510);
  nor g9 (n_511, n_152, n_176);
  nand g10 (n_514, n_152, n_176);
  nor g11 (n_521, n_151, n_175);
  nand g12 (n_516, n_151, n_175);
  nor g13 (n_517, n_150, n_174);
  nand g14 (n_518, n_150, n_174);
  nor g15 (n_527, n_149, n_173);
  nand g16 (n_522, n_149, n_173);
  nor g17 (n_523, n_148, n_172);
  nand g18 (n_524, n_148, n_172);
  nor g19 (n_533, n_147, n_171);
  nand g20 (n_528, n_147, n_171);
  nor g21 (n_529, n_146, n_170);
  nand g22 (n_530, n_146, n_170);
  nor g23 (n_539, n_145, n_169);
  nand g24 (n_534, n_145, n_169);
  nor g25 (n_535, n_144, n_168);
  nand g26 (n_536, n_144, n_168);
  nor g27 (n_545, n_143, n_167);
  nand g28 (n_540, n_143, n_167);
  nor g29 (n_541, n_142, n_166);
  nand g30 (n_542, n_142, n_166);
  nor g31 (n_551, n_141, n_165);
  nand g32 (n_546, n_141, n_165);
  nor g33 (n_547, n_140, n_164);
  nand g34 (n_548, n_140, n_164);
  nor g35 (n_557, n_139, n_163);
  nand g36 (n_552, n_139, n_163);
  nor g37 (n_553, n_138, n_162);
  nand g38 (n_554, n_138, n_162);
  nor g39 (n_563, n_137, n_161);
  nand g40 (n_558, n_137, n_161);
  nor g41 (n_559, n_136, n_160);
  nand g42 (n_560, n_136, n_160);
  nor g43 (n_569, n_135, n_159);
  nand g44 (n_564, n_135, n_159);
  nor g45 (n_565, n_134, n_158);
  nand g46 (n_566, n_134, n_158);
  nor g47 (n_575, n_133, n_157);
  nand g48 (n_570, n_133, n_157);
  nor g49 (n_571, n_132, n_156);
  nand g50 (n_572, n_132, n_156);
  nor g51 (n_579, n_131, n_155);
  nand g52 (n_576, n_131, n_155);
  nand g57 (n_580, n_514, n_515);
  nor g58 (n_519, n_516, n_517);
  nor g61 (n_582, n_521, n_517);
  nor g62 (n_525, n_522, n_523);
  nor g65 (n_588, n_527, n_523);
  nor g66 (n_531, n_528, n_529);
  nor g439 (n_590, n_533, n_529);
  nor g440 (n_537, n_534, n_535);
  nor g443 (n_598, n_539, n_535);
  nor g444 (n_543, n_540, n_541);
  nor g447 (n_600, n_545, n_541);
  nor g448 (n_549, n_546, n_547);
  nor g451 (n_608, n_551, n_547);
  nor g452 (n_555, n_552, n_553);
  nor g455 (n_610, n_557, n_553);
  nor g456 (n_561, n_558, n_559);
  nor g459 (n_618, n_563, n_559);
  nor g460 (n_567, n_564, n_565);
  nor g463 (n_620, n_569, n_565);
  nor g464 (n_573, n_570, n_571);
  nor g467 (n_628, n_575, n_571);
  nand g470 (n_712, n_516, n_581);
  nand g471 (n_584, n_582, n_580);
  nand g472 (n_630, n_583, n_584);
  nor g473 (n_586, n_533, n_585);
  nand g482 (n_638, n_588, n_590);
  nor g483 (n_596, n_545, n_595);
  nand g492 (n_645, n_598, n_600);
  nor g493 (n_606, n_557, n_605);
  nand g502 (n_653, n_608, n_610);
  nor g503 (n_616, n_569, n_615);
  nand g512 (n_660, n_618, n_620);
  nor g513 (n_626, n_579, n_625);
  nand g520 (n_716, n_522, n_632);
  nand g521 (n_633, n_588, n_630);
  nand g522 (n_718, n_585, n_633);
  nand g525 (n_721, n_636, n_637);
  nand g528 (n_668, n_640, n_641);
  nor g529 (n_643, n_551, n_642);
  nor g532 (n_678, n_551, n_645);
  nor g538 (n_651, n_649, n_642);
  nor g541 (n_684, n_645, n_649);
  nor g542 (n_655, n_653, n_642);
  nor g545 (n_687, n_645, n_653);
  nor g546 (n_658, n_575, n_657);
  nor g549 (n_700, n_575, n_660);
  nor g555 (n_666, n_664, n_657);
  nor g558 (n_706, n_660, n_664);
  nand g561 (n_725, n_534, n_670);
  nand g562 (n_671, n_598, n_668);
  nand g563 (n_727, n_595, n_671);
  nand g566 (n_730, n_674, n_675);
  nand g569 (n_733, n_642, n_677);
  nand g570 (n_680, n_678, n_668);
  nand g571 (n_736, n_679, n_680);
  nand g572 (n_683, n_681, n_668);
  nand g573 (n_738, n_682, n_683);
  nand g574 (n_686, n_684, n_668);
  nand g575 (n_741, n_685, n_686);
  nand g576 (n_689, n_687, n_668);
  nand g577 (n_690, n_688, n_689);
  nand g580 (n_745, n_558, n_692);
  nand g581 (n_693, n_618, n_690);
  nand g582 (n_747, n_615, n_693);
  nand g585 (n_750, n_696, n_697);
  nand g588 (n_753, n_657, n_699);
  nand g589 (n_702, n_700, n_690);
  nand g590 (n_756, n_701, n_702);
  nand g591 (n_705, n_703, n_690);
  nand g592 (n_758, n_704, n_705);
  nand g593 (n_708, n_706, n_690);
  nand g594 (n_761, n_707, n_708);
  xnor g596 (out_0[1], n_512, n_709);
  xnor g598 (out_0[2], n_580, n_710);
  xnor g601 (out_0[3], n_712, n_713);
  xnor g603 (out_0[4], n_630, n_714);
  xnor g606 (out_0[5], n_716, n_717);
  xnor g608 (out_0[6], n_718, n_719);
  xnor g611 (out_0[7], n_721, n_722);
  xnor g613 (out_0[8], n_668, n_723);
  xnor g616 (out_0[9], n_725, n_726);
  xnor g618 (out_0[10], n_727, n_728);
  xnor g621 (out_0[11], n_730, n_731);
  xnor g624 (out_0[12], n_733, n_734);
  xnor g627 (out_0[13], n_736, n_737);
  xnor g629 (out_0[14], n_738, n_739);
  xnor g632 (out_0[15], n_741, n_742);
  xnor g634 (out_0[16], n_690, n_743);
  xnor g637 (out_0[17], n_745, n_746);
  xnor g639 (out_0[18], n_747, n_748);
  xnor g642 (out_0[19], n_750, n_751);
  xnor g645 (out_0[20], n_753, n_754);
  xnor g648 (out_0[21], n_756, n_757);
  xnor g650 (out_0[22], n_758, n_759);
  xor g654 (out_0[0], in_2[0], n_763);
  xor g655 (n_256, in_0[20], in_1[20]);
  nor g656 (n_131, in_0[20], in_1[20]);
  xor g657 (n_490, in_3[20], in_4[20]);
  or g658 (n_491, in_3[20], in_4[20]);
  or g659 (n_492, in_2[20], in_4[20]);
  or g660 (n_493, in_2[20], in_3[20]);
  xnor g661 (n_258, n_490, in_2[20]);
  xnor g665 (n_259, n_257, n_256);
  or g666 (n_265, n_256, wc, n_257);
  not gc (wc, n_496);
  xnor g667 (n_502, n_263, n_131);
  or g668 (n_503, n_131, wc0);
  not gc0 (wc0, n_263);
  or g669 (n_504, wc1, n_131);
  not gc1 (wc1, n_265);
  or g670 (n_515, n_511, wc2);
  not gc2 (wc2, n_512);
  or g671 (n_709, wc3, n_511);
  not gc3 (wc3, n_514);
  and g672 (n_583, wc4, n_518);
  not gc4 (wc4, n_519);
  or g673 (n_710, wc5, n_521);
  not gc5 (wc5, n_516);
  or g674 (n_713, wc6, n_517);
  not gc6 (wc6, n_518);
  and g675 (n_585, wc7, n_524);
  not gc7 (wc7, n_525);
  or g676 (n_581, wc8, n_521);
  not gc8 (wc8, n_580);
  or g677 (n_714, wc9, n_527);
  not gc9 (wc9, n_522);
  or g678 (n_717, wc10, n_523);
  not gc10 (wc10, n_524);
  and g679 (n_592, wc11, n_530);
  not gc11 (wc11, n_531);
  and g680 (n_595, wc12, n_536);
  not gc12 (wc12, n_537);
  and g681 (n_602, wc13, n_542);
  not gc13 (wc13, n_543);
  and g682 (n_605, wc14, n_548);
  not gc14 (wc14, n_549);
  and g683 (n_612, wc15, n_554);
  not gc15 (wc15, n_555);
  and g684 (n_615, wc16, n_560);
  not gc16 (wc16, n_561);
  and g685 (n_622, wc17, n_566);
  not gc17 (wc17, n_567);
  and g686 (n_625, wc18, n_572);
  not gc18 (wc18, n_573);
  or g687 (n_634, wc19, n_533);
  not gc19 (wc19, n_588);
  or g688 (n_672, wc20, n_545);
  not gc20 (wc20, n_598);
  or g689 (n_649, wc21, n_557);
  not gc21 (wc21, n_608);
  or g690 (n_694, wc22, n_569);
  not gc22 (wc22, n_618);
  or g691 (n_664, wc23, n_579);
  not gc23 (wc23, n_628);
  or g692 (n_719, wc24, n_533);
  not gc24 (wc24, n_528);
  or g693 (n_722, wc25, n_529);
  not gc25 (wc25, n_530);
  or g694 (n_723, wc26, n_539);
  not gc26 (wc26, n_534);
  or g695 (n_726, wc27, n_535);
  not gc27 (wc27, n_536);
  or g696 (n_728, wc28, n_545);
  not gc28 (wc28, n_540);
  or g697 (n_731, wc29, n_541);
  not gc29 (wc29, n_542);
  or g698 (n_734, wc30, n_551);
  not gc30 (wc30, n_546);
  or g699 (n_737, wc31, n_547);
  not gc31 (wc31, n_548);
  or g700 (n_739, wc32, n_557);
  not gc32 (wc32, n_552);
  or g701 (n_742, wc33, n_553);
  not gc33 (wc33, n_554);
  or g702 (n_743, wc34, n_563);
  not gc34 (wc34, n_558);
  or g703 (n_746, wc35, n_559);
  not gc35 (wc35, n_560);
  or g704 (n_748, wc36, n_569);
  not gc36 (wc36, n_564);
  or g705 (n_751, wc37, n_565);
  not gc37 (wc37, n_566);
  or g706 (n_754, wc38, n_575);
  not gc38 (wc38, n_570);
  or g707 (n_757, wc39, n_571);
  not gc39 (wc39, n_572);
  or g708 (n_759, wc40, n_579);
  not gc40 (wc40, n_576);
  and g709 (n_636, wc41, n_528);
  not gc41 (wc41, n_586);
  and g710 (n_593, wc42, n_590);
  not gc42 (wc42, n_585);
  and g711 (n_603, wc43, n_600);
  not gc43 (wc43, n_595);
  and g712 (n_613, wc44, n_610);
  not gc44 (wc44, n_605);
  and g713 (n_623, wc45, n_620);
  not gc45 (wc45, n_615);
  or g714 (n_632, wc46, n_527);
  not gc46 (wc46, n_630);
  and g715 (n_681, wc47, n_608);
  not gc47 (wc47, n_645);
  and g716 (n_703, wc48, n_628);
  not gc48 (wc48, n_660);
  and g717 (n_640, wc49, n_592);
  not gc49 (wc49, n_593);
  and g718 (n_674, wc50, n_540);
  not gc50 (wc50, n_596);
  and g719 (n_642, wc51, n_602);
  not gc51 (wc51, n_603);
  and g720 (n_650, wc52, n_552);
  not gc52 (wc52, n_606);
  and g721 (n_654, wc53, n_612);
  not gc53 (wc53, n_613);
  and g722 (n_696, wc54, n_564);
  not gc54 (wc54, n_616);
  and g723 (n_657, wc55, n_622);
  not gc55 (wc55, n_623);
  and g724 (n_665, wc56, n_576);
  not gc56 (wc56, n_626);
  or g725 (n_637, n_634, wc57);
  not gc57 (wc57, n_630);
  or g726 (n_641, n_638, wc58);
  not gc58 (wc58, n_630);
  and g727 (n_647, wc59, n_608);
  not gc59 (wc59, n_642);
  and g728 (n_662, wc60, n_628);
  not gc60 (wc60, n_657);
  and g729 (n_679, wc61, n_546);
  not gc61 (wc61, n_643);
  and g730 (n_682, wc62, n_605);
  not gc62 (wc62, n_647);
  and g731 (n_685, n_650, wc63);
  not gc63 (wc63, n_651);
  and g732 (n_688, n_654, wc64);
  not gc64 (wc64, n_655);
  and g733 (n_701, wc65, n_570);
  not gc65 (wc65, n_658);
  and g734 (n_704, wc66, n_625);
  not gc66 (wc66, n_662);
  and g735 (n_707, n_665, wc67);
  not gc67 (wc67, n_666);
  or g736 (n_670, wc68, n_539);
  not gc68 (wc68, n_668);
  or g737 (n_675, n_672, wc69);
  not gc69 (wc69, n_668);
  or g738 (n_677, wc70, n_645);
  not gc70 (wc70, n_668);
  or g739 (n_692, wc71, n_563);
  not gc71 (wc71, n_690);
  or g740 (n_697, n_694, wc72);
  not gc72 (wc72, n_690);
  or g741 (n_699, wc73, n_660);
  not gc73 (wc73, n_690);
  not g742 (out_0[23], n_761);
endmodule

module csa_tree_add_255_42_group_6823_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [20:0] in_0, in_1, in_2, in_3, in_4;
  output [23:0] out_0;
  wire [20:0] in_0, in_1, in_2, in_3, in_4;
  wire [23:0] out_0;
  csa_tree_add_255_42_group_6823_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_284_36_group_6827_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  wire n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110;
  wire n_111, n_112, n_113, n_114, n_115, n_116, n_117, n_118;
  wire n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_158, n_159, n_160, n_161;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201;
  wire n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209;
  wire n_210, n_211, n_212, n_213, n_214, n_215, n_216, n_217;
  wire n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225;
  wire n_226, n_227, n_228, n_229, n_230, n_231, n_232, n_233;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_242, n_243;
  wire n_244, n_245, n_246, n_248, n_249, n_250, n_251, n_252;
  wire n_253, n_255, n_256, n_257, n_258, n_259, n_261, n_262;
  wire n_263, n_264, n_265, n_267, n_268, n_269, n_270, n_271;
  wire n_273, n_274, n_275, n_276, n_277, n_279, n_280, n_281;
  wire n_282, n_283, n_285, n_286, n_287, n_288, n_289, n_291;
  wire n_292, n_293, n_294, n_295, n_297, n_298, n_299, n_300;
  wire n_301, n_303, n_304, n_305, n_306, n_307, n_309, n_310;
  wire n_311, n_312, n_313, n_315, n_316, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_325, n_327, n_329, n_330, n_332;
  wire n_333, n_335, n_337, n_339, n_340, n_342, n_343, n_345;
  wire n_347, n_349, n_350, n_352, n_353, n_355, n_357, n_359;
  wire n_360, n_362, n_363, n_365, n_367, n_369, n_370, n_372;
  wire n_374, n_375, n_376, n_378, n_379, n_380, n_382, n_383;
  wire n_384, n_385, n_387, n_389, n_391, n_392, n_393, n_395;
  wire n_396, n_397, n_399, n_400, n_402, n_404, n_406, n_407;
  wire n_408, n_410, n_411, n_412, n_414, n_416, n_417, n_418;
  wire n_420, n_421, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_441, n_443, n_444, n_445, n_447;
  wire n_448, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_464, n_465;
  wire n_466, n_468, n_469, n_470, n_471, n_473, n_474, n_475;
  wire n_477, n_478, n_479, n_480, n_482, n_483, n_485, n_486;
  wire n_488, n_489, n_490, n_491, n_493, n_494, n_495, n_497;
  wire n_498, n_499, n_500, n_502, n_503, n_505, n_506, n_508;
  wire n_509, n_510, n_511, n_513, n_514, n_515, n_516, n_517;
  xor g26 (n_125, in_2[1], in_0[1]);
  and g2 (n_153, in_2[1], in_0[1]);
  xor g27 (n_123, in_2[2], n_153);
  xor g28 (n_149, n_123, in_0[2]);
  nand g3 (n_124, in_2[2], n_153);
  nand g29 (n_158, in_0[2], n_153);
  nand g30 (n_126, in_2[2], in_0[2]);
  nand g31 (n_154, n_124, n_158, n_126);
  xor g32 (n_159, in_2[3], in_0[3]);
  xor g33 (n_148, n_159, n_154);
  nand g34 (n_160, in_2[3], in_0[3]);
  nand g4 (n_161, n_154, in_0[3]);
  nand g35 (n_162, in_2[3], n_154);
  nand g36 (n_122, n_160, n_161, n_162);
  xor g37 (n_163, in_2[4], in_0[4]);
  xor g38 (n_147, n_163, in_1[4]);
  nand g39 (n_164, in_2[4], in_0[4]);
  nand g40 (n_165, in_1[4], in_0[4]);
  nand g5 (n_166, in_2[4], in_1[4]);
  nand g41 (n_121, n_164, n_165, n_166);
  xor g42 (n_167, in_2[5], in_0[5]);
  xor g43 (n_146, n_167, in_1[5]);
  nand g44 (n_168, in_2[5], in_0[5]);
  nand g45 (n_169, in_1[5], in_0[5]);
  nand g46 (n_170, in_2[5], in_1[5]);
  nand g6 (n_120, n_168, n_169, n_170);
  xor g47 (n_171, in_2[6], in_0[6]);
  xor g48 (n_145, n_171, in_1[6]);
  nand g49 (n_172, in_2[6], in_0[6]);
  nand g50 (n_173, in_1[6], in_0[6]);
  nand g51 (n_174, in_2[6], in_1[6]);
  nand g52 (n_119, n_172, n_173, n_174);
  xor g53 (n_175, in_2[7], in_0[7]);
  xor g54 (n_144, n_175, in_1[7]);
  nand g55 (n_176, in_2[7], in_0[7]);
  nand g56 (n_177, in_1[7], in_0[7]);
  nand g57 (n_178, in_2[7], in_1[7]);
  nand g58 (n_118, n_176, n_177, n_178);
  xor g59 (n_179, in_2[8], in_0[8]);
  xor g60 (n_143, n_179, in_1[8]);
  nand g61 (n_180, in_2[8], in_0[8]);
  nand g62 (n_181, in_1[8], in_0[8]);
  nand g63 (n_150, in_2[8], in_1[8]);
  nand g64 (n_117, n_180, n_181, n_150);
  xor g65 (n_151, in_2[9], in_0[9]);
  xor g66 (n_142, n_151, in_1[9]);
  nand g67 (n_152, in_2[9], in_0[9]);
  nand g68 (n_182, in_1[9], in_0[9]);
  nand g69 (n_183, in_2[9], in_1[9]);
  nand g70 (n_116, n_152, n_182, n_183);
  xor g71 (n_184, in_2[10], in_0[10]);
  xor g72 (n_141, n_184, in_1[10]);
  nand g73 (n_185, in_2[10], in_0[10]);
  nand g74 (n_186, in_1[10], in_0[10]);
  nand g75 (n_187, in_2[10], in_1[10]);
  nand g76 (n_115, n_185, n_186, n_187);
  xor g77 (n_188, in_2[11], in_0[11]);
  xor g78 (n_140, n_188, in_1[11]);
  nand g79 (n_189, in_2[11], in_0[11]);
  nand g80 (n_190, in_1[11], in_0[11]);
  nand g81 (n_191, in_2[11], in_1[11]);
  nand g82 (n_114, n_189, n_190, n_191);
  xor g83 (n_192, in_2[12], in_0[12]);
  xor g84 (n_139, n_192, in_1[12]);
  nand g85 (n_193, in_2[12], in_0[12]);
  nand g86 (n_194, in_1[12], in_0[12]);
  nand g87 (n_195, in_2[12], in_1[12]);
  nand g88 (n_113, n_193, n_194, n_195);
  xor g89 (n_196, in_2[13], in_0[13]);
  xor g90 (n_138, n_196, in_1[13]);
  nand g91 (n_197, in_2[13], in_0[13]);
  nand g92 (n_198, in_1[13], in_0[13]);
  nand g93 (n_199, in_2[13], in_1[13]);
  nand g94 (n_112, n_197, n_198, n_199);
  xor g95 (n_200, in_2[14], in_0[14]);
  xor g96 (n_137, n_200, in_1[14]);
  nand g97 (n_201, in_2[14], in_0[14]);
  nand g98 (n_202, in_1[14], in_0[14]);
  nand g99 (n_203, in_2[14], in_1[14]);
  nand g100 (n_111, n_201, n_202, n_203);
  xor g101 (n_204, in_2[15], in_0[15]);
  xor g102 (n_136, n_204, in_1[15]);
  nand g103 (n_205, in_2[15], in_0[15]);
  nand g104 (n_206, in_1[15], in_0[15]);
  nand g105 (n_207, in_2[15], in_1[15]);
  nand g106 (n_110, n_205, n_206, n_207);
  xor g107 (n_208, in_2[16], in_0[16]);
  xor g108 (n_135, n_208, in_1[16]);
  nand g109 (n_209, in_2[16], in_0[16]);
  nand g110 (n_210, in_1[16], in_0[16]);
  nand g111 (n_211, in_2[16], in_1[16]);
  nand g112 (n_109, n_209, n_210, n_211);
  xor g113 (n_212, in_2[17], in_0[17]);
  xor g114 (n_134, n_212, in_1[17]);
  nand g115 (n_213, in_2[17], in_0[17]);
  nand g116 (n_214, in_1[17], in_0[17]);
  nand g117 (n_215, in_2[17], in_1[17]);
  nand g118 (n_108, n_213, n_214, n_215);
  xor g119 (n_216, in_2[18], in_0[18]);
  xor g120 (n_133, n_216, in_1[18]);
  nand g121 (n_217, in_2[18], in_0[18]);
  nand g122 (n_218, in_1[18], in_0[18]);
  nand g123 (n_219, in_2[18], in_1[18]);
  nand g124 (n_107, n_217, n_218, n_219);
  xor g125 (n_220, in_2[19], in_0[19]);
  xor g126 (n_132, n_220, in_1[19]);
  nand g127 (n_221, in_2[19], in_0[19]);
  nand g128 (n_222, in_1[19], in_0[19]);
  nand g129 (n_223, in_2[19], in_1[19]);
  nand g130 (n_106, n_221, n_222, n_223);
  xor g131 (n_224, in_2[20], in_0[20]);
  xor g132 (n_131, n_224, in_1[20]);
  nand g133 (n_225, in_2[20], in_0[20]);
  nand g134 (n_226, in_1[20], in_0[20]);
  nand g135 (n_227, in_2[20], in_1[20]);
  nand g136 (n_105, n_225, n_226, n_227);
  xor g137 (n_228, in_2[21], in_0[21]);
  xor g138 (n_130, n_228, in_1[21]);
  nand g139 (n_229, in_2[21], in_0[21]);
  nand g140 (n_230, in_1[21], in_0[21]);
  nand g141 (n_231, in_2[21], in_1[21]);
  nand g142 (n_104, n_229, n_230, n_231);
  xor g143 (n_232, in_2[22], in_0[22]);
  xor g144 (n_129, n_232, in_1[22]);
  nand g145 (n_233, in_2[22], in_0[22]);
  nand g146 (n_234, in_1[22], in_0[22]);
  nand g147 (n_235, in_2[22], in_1[22]);
  nand g148 (n_103, n_233, n_234, n_235);
  xor g151 (n_236, in_2[23], in_1[23]);
  xor g152 (n_128, n_236, in_0[23]);
  nand g153 (n_237, in_2[23], in_1[23]);
  nand g154 (n_238, in_0[23], in_1[23]);
  nand g155 (n_239, in_2[23], in_0[23]);
  nand g156 (n_127, n_237, n_238, n_239);
  xor g159 (n_517, in_1[0], in_0[0]);
  nand g160 (n_242, in_1[0], in_0[0]);
  nand g161 (n_243, in_1[0], in_2[0]);
  nand g7 (n_244, in_0[0], in_2[0]);
  nand g8 (n_246, n_242, n_243, n_244);
  nor g9 (n_245, n_125, in_1[1]);
  nand g10 (n_248, n_125, in_1[1]);
  nor g11 (n_255, in_1[2], n_149);
  nand g12 (n_250, in_1[2], n_149);
  nor g13 (n_251, in_1[3], n_148);
  nand g14 (n_252, in_1[3], n_148);
  nor g15 (n_261, n_122, n_147);
  nand g16 (n_256, n_122, n_147);
  nor g17 (n_257, n_121, n_146);
  nand g18 (n_258, n_121, n_146);
  nor g19 (n_267, n_120, n_145);
  nand g20 (n_262, n_120, n_145);
  nor g21 (n_263, n_119, n_144);
  nand g22 (n_264, n_119, n_144);
  nor g23 (n_273, n_118, n_143);
  nand g24 (n_268, n_118, n_143);
  nor g25 (n_269, n_117, n_142);
  nand g162 (n_270, n_117, n_142);
  nor g163 (n_279, n_116, n_141);
  nand g164 (n_274, n_116, n_141);
  nor g165 (n_275, n_115, n_140);
  nand g166 (n_276, n_115, n_140);
  nor g167 (n_285, n_114, n_139);
  nand g168 (n_280, n_114, n_139);
  nor g169 (n_281, n_113, n_138);
  nand g170 (n_282, n_113, n_138);
  nor g171 (n_291, n_112, n_137);
  nand g172 (n_286, n_112, n_137);
  nor g173 (n_287, n_111, n_136);
  nand g174 (n_288, n_111, n_136);
  nor g175 (n_297, n_110, n_135);
  nand g176 (n_292, n_110, n_135);
  nor g177 (n_293, n_109, n_134);
  nand g178 (n_294, n_109, n_134);
  nor g179 (n_303, n_108, n_133);
  nand g180 (n_298, n_108, n_133);
  nor g181 (n_299, n_107, n_132);
  nand g182 (n_300, n_107, n_132);
  nor g183 (n_309, n_106, n_131);
  nand g184 (n_304, n_106, n_131);
  nor g185 (n_305, n_105, n_130);
  nand g186 (n_306, n_105, n_130);
  nor g187 (n_315, n_104, n_129);
  nand g188 (n_310, n_104, n_129);
  nor g189 (n_311, n_103, n_128);
  nand g190 (n_312, n_103, n_128);
  nand g195 (n_316, n_248, n_249);
  nor g196 (n_253, n_250, n_251);
  nor g199 (n_319, n_255, n_251);
  nor g200 (n_259, n_256, n_257);
  nor g203 (n_325, n_261, n_257);
  nor g204 (n_265, n_262, n_263);
  nor g207 (n_327, n_267, n_263);
  nor g208 (n_271, n_268, n_269);
  nor g211 (n_335, n_273, n_269);
  nor g212 (n_277, n_274, n_275);
  nor g215 (n_337, n_279, n_275);
  nor g216 (n_283, n_280, n_281);
  nor g219 (n_345, n_285, n_281);
  nor g220 (n_289, n_286, n_287);
  nor g223 (n_347, n_291, n_287);
  nor g224 (n_295, n_292, n_293);
  nor g227 (n_355, n_297, n_293);
  nor g228 (n_301, n_298, n_299);
  nor g231 (n_357, n_303, n_299);
  nor g232 (n_307, n_304, n_305);
  nor g235 (n_365, n_309, n_305);
  nor g236 (n_313, n_310, n_311);
  nor g239 (n_367, n_315, n_311);
  nand g242 (n_464, n_250, n_318);
  nand g243 (n_321, n_319, n_316);
  nand g244 (n_372, n_320, n_321);
  nor g245 (n_323, n_267, n_322);
  nand g254 (n_380, n_325, n_327);
  nor g255 (n_333, n_279, n_332);
  nand g264 (n_387, n_335, n_337);
  nor g265 (n_343, n_291, n_342);
  nand g274 (n_395, n_345, n_347);
  nor g275 (n_353, n_303, n_352);
  nand g284 (n_402, n_355, n_357);
  nor g285 (n_363, n_315, n_362);
  nand g294 (n_410, n_365, n_367);
  nand g297 (n_468, n_256, n_374);
  nand g298 (n_375, n_325, n_372);
  nand g299 (n_470, n_322, n_375);
  nand g302 (n_473, n_378, n_379);
  nand g305 (n_414, n_382, n_383);
  nor g306 (n_385, n_285, n_384);
  nor g309 (n_424, n_285, n_387);
  nor g315 (n_393, n_391, n_384);
  nor g318 (n_430, n_387, n_391);
  nor g319 (n_397, n_395, n_384);
  nor g322 (n_433, n_387, n_395);
  nor g323 (n_400, n_309, n_399);
  nor g326 (n_451, n_309, n_402);
  nor g332 (n_408, n_406, n_399);
  nor g335 (n_457, n_402, n_406);
  nor g336 (n_412, n_410, n_399);
  nor g339 (n_439, n_402, n_410);
  nand g342 (n_477, n_268, n_416);
  nand g343 (n_417, n_335, n_414);
  nand g344 (n_479, n_332, n_417);
  nand g347 (n_482, n_420, n_421);
  nand g350 (n_485, n_384, n_423);
  nand g351 (n_426, n_424, n_414);
  nand g352 (n_488, n_425, n_426);
  nand g353 (n_429, n_427, n_414);
  nand g354 (n_490, n_428, n_429);
  nand g355 (n_432, n_430, n_414);
  nand g356 (n_493, n_431, n_432);
  nand g357 (n_435, n_433, n_414);
  nand g358 (n_441, n_434, n_435);
  nand g362 (n_497, n_292, n_443);
  nand g363 (n_444, n_355, n_441);
  nand g364 (n_499, n_352, n_444);
  nand g367 (n_502, n_447, n_448);
  nand g370 (n_505, n_399, n_450);
  nand g371 (n_453, n_451, n_441);
  nand g372 (n_508, n_452, n_453);
  nand g373 (n_456, n_454, n_441);
  nand g374 (n_510, n_455, n_456);
  nand g375 (n_459, n_457, n_441);
  nand g376 (n_513, n_458, n_459);
  nand g377 (n_460, n_439, n_441);
  nand g378 (n_515, n_437, n_460);
  xnor g380 (out_0[1], n_246, n_461);
  xnor g382 (out_0[2], n_316, n_462);
  xnor g385 (out_0[3], n_464, n_465);
  xnor g387 (out_0[4], n_372, n_466);
  xnor g390 (out_0[5], n_468, n_469);
  xnor g392 (out_0[6], n_470, n_471);
  xnor g395 (out_0[7], n_473, n_474);
  xnor g397 (out_0[8], n_414, n_475);
  xnor g400 (out_0[9], n_477, n_478);
  xnor g402 (out_0[10], n_479, n_480);
  xnor g405 (out_0[11], n_482, n_483);
  xnor g408 (out_0[12], n_485, n_486);
  xnor g411 (out_0[13], n_488, n_489);
  xnor g413 (out_0[14], n_490, n_491);
  xnor g416 (out_0[15], n_493, n_494);
  xnor g418 (out_0[16], n_441, n_495);
  xnor g421 (out_0[17], n_497, n_498);
  xnor g423 (out_0[18], n_499, n_500);
  xnor g426 (out_0[19], n_502, n_503);
  xnor g429 (out_0[20], n_505, n_506);
  xnor g432 (out_0[21], n_508, n_509);
  xnor g434 (out_0[22], n_510, n_511);
  xnor g437 (out_0[23], n_513, n_514);
  xnor g439 (out_0[24], n_515, n_516);
  xor g440 (out_0[0], in_2[0], n_517);
  or g441 (n_249, n_245, wc);
  not gc (wc, n_246);
  or g442 (n_461, wc0, n_245);
  not gc0 (wc0, n_248);
  and g443 (n_329, wc1, n_264);
  not gc1 (wc1, n_265);
  and g444 (n_332, wc2, n_270);
  not gc2 (wc2, n_271);
  and g445 (n_339, wc3, n_276);
  not gc3 (wc3, n_277);
  and g446 (n_342, wc4, n_282);
  not gc4 (wc4, n_283);
  and g447 (n_349, wc5, n_288);
  not gc5 (wc5, n_289);
  and g448 (n_352, wc6, n_294);
  not gc6 (wc6, n_295);
  and g449 (n_359, wc7, n_300);
  not gc7 (wc7, n_301);
  and g450 (n_362, wc8, n_306);
  not gc8 (wc8, n_307);
  or g451 (n_418, wc9, n_279);
  not gc9 (wc9, n_335);
  or g452 (n_391, wc10, n_291);
  not gc10 (wc10, n_345);
  or g453 (n_445, wc11, n_303);
  not gc11 (wc11, n_355);
  or g454 (n_406, wc12, n_315);
  not gc12 (wc12, n_365);
  or g455 (n_469, wc13, n_257);
  not gc13 (wc13, n_258);
  or g456 (n_471, wc14, n_267);
  not gc14 (wc14, n_262);
  or g457 (n_474, wc15, n_263);
  not gc15 (wc15, n_264);
  or g458 (n_475, wc16, n_273);
  not gc16 (wc16, n_268);
  or g459 (n_478, wc17, n_269);
  not gc17 (wc17, n_270);
  or g460 (n_480, wc18, n_279);
  not gc18 (wc18, n_274);
  or g461 (n_483, wc19, n_275);
  not gc19 (wc19, n_276);
  or g462 (n_486, wc20, n_285);
  not gc20 (wc20, n_280);
  or g463 (n_489, wc21, n_281);
  not gc21 (wc21, n_282);
  or g464 (n_491, wc22, n_291);
  not gc22 (wc22, n_286);
  or g465 (n_494, wc23, n_287);
  not gc23 (wc23, n_288);
  or g466 (n_495, wc24, n_297);
  not gc24 (wc24, n_292);
  or g467 (n_498, wc25, n_293);
  not gc25 (wc25, n_294);
  or g468 (n_500, wc26, n_303);
  not gc26 (wc26, n_298);
  or g469 (n_503, wc27, n_299);
  not gc27 (wc27, n_300);
  or g470 (n_506, wc28, n_309);
  not gc28 (wc28, n_304);
  or g471 (n_509, wc29, n_305);
  not gc29 (wc29, n_306);
  or g472 (n_511, wc30, n_315);
  not gc30 (wc30, n_310);
  and g473 (n_436, wc31, n_127);
  not gc31 (wc31, in_2[23]);
  or g474 (n_438, wc32, n_127);
  not gc32 (wc32, in_2[23]);
  or g475 (n_318, wc33, n_255);
  not gc33 (wc33, n_316);
  and g476 (n_340, wc34, n_337);
  not gc34 (wc34, n_332);
  and g477 (n_350, wc35, n_347);
  not gc35 (wc35, n_342);
  and g478 (n_360, wc36, n_357);
  not gc36 (wc36, n_352);
  and g479 (n_427, wc37, n_345);
  not gc37 (wc37, n_387);
  and g480 (n_454, wc38, n_365);
  not gc38 (wc38, n_402);
  or g481 (n_462, wc39, n_255);
  not gc39 (wc39, n_250);
  and g482 (n_320, wc40, n_252);
  not gc40 (wc40, n_253);
  and g483 (n_369, wc41, n_312);
  not gc41 (wc41, n_313);
  and g484 (n_420, wc42, n_274);
  not gc42 (wc42, n_333);
  and g485 (n_384, wc43, n_339);
  not gc43 (wc43, n_340);
  and g486 (n_392, wc44, n_286);
  not gc44 (wc44, n_343);
  and g487 (n_396, wc45, n_349);
  not gc45 (wc45, n_350);
  and g488 (n_447, wc46, n_298);
  not gc46 (wc46, n_353);
  and g489 (n_399, wc47, n_359);
  not gc47 (wc47, n_360);
  and g490 (n_407, wc48, n_310);
  not gc48 (wc48, n_363);
  or g491 (n_465, wc49, n_251);
  not gc49 (wc49, n_252);
  or g492 (n_514, wc50, n_311);
  not gc50 (wc50, n_312);
  and g493 (n_322, wc51, n_258);
  not gc51 (wc51, n_259);
  or g494 (n_376, wc52, n_267);
  not gc52 (wc52, n_325);
  and g495 (n_370, wc53, n_367);
  not gc53 (wc53, n_362);
  and g496 (n_389, wc54, n_345);
  not gc54 (wc54, n_384);
  and g497 (n_404, wc55, n_365);
  not gc55 (wc55, n_399);
  or g498 (n_466, wc56, n_261);
  not gc56 (wc56, n_256);
  or g499 (n_516, wc57, n_436);
  not gc57 (wc57, n_438);
  and g500 (n_330, wc58, n_327);
  not gc58 (wc58, n_322);
  and g501 (n_411, wc59, n_369);
  not gc59 (wc59, n_370);
  or g502 (n_374, wc60, n_261);
  not gc60 (wc60, n_372);
  and g503 (n_425, wc61, n_280);
  not gc61 (wc61, n_385);
  and g504 (n_428, wc62, n_342);
  not gc62 (wc62, n_389);
  and g505 (n_431, n_392, wc63);
  not gc63 (wc63, n_393);
  and g506 (n_434, n_396, wc64);
  not gc64 (wc64, n_397);
  and g507 (n_452, wc65, n_304);
  not gc65 (wc65, n_400);
  and g508 (n_455, wc66, n_362);
  not gc66 (wc66, n_404);
  and g509 (n_458, n_407, wc67);
  not gc67 (wc67, n_408);
  and g510 (n_378, wc68, n_262);
  not gc68 (wc68, n_323);
  and g511 (n_382, wc69, n_329);
  not gc69 (wc69, n_330);
  or g512 (n_379, n_376, wc70);
  not gc70 (wc70, n_372);
  or g513 (n_383, n_380, wc71);
  not gc71 (wc71, n_372);
  and g514 (n_437, n_411, wc72);
  not gc72 (wc72, n_412);
  or g515 (n_416, wc73, n_273);
  not gc73 (wc73, n_414);
  or g516 (n_421, n_418, wc74);
  not gc74 (wc74, n_414);
  or g517 (n_423, wc75, n_387);
  not gc75 (wc75, n_414);
  or g518 (n_443, wc76, n_297);
  not gc76 (wc76, n_441);
  or g519 (n_448, n_445, wc77);
  not gc77 (wc77, n_441);
  or g520 (n_450, wc78, n_402);
  not gc78 (wc78, n_441);
endmodule

module csa_tree_add_284_36_group_6827_GENERIC(in_0, in_1, in_2, out_0);
  input [25:0] in_0, in_1;
  input [23:0] in_2;
  output [24:0] out_0;
  wire [25:0] in_0, in_1;
  wire [23:0] in_2;
  wire [24:0] out_0;
  csa_tree_add_284_36_group_6827_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_287_40_group_6803_GENERIC_REAL(in_0, in_1, in_2,
     out_0);
// synthesis_equation "assign out_0 = ( ( $signed(in_0) + $signed(in_1) ) + $signed(in_2) )  ;"
  input [26:0] in_0, in_1;
  input [24:0] in_2;
  output [25:0] out_0;
  wire [26:0] in_0, in_1;
  wire [24:0] in_2;
  wire [25:0] out_0;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130;
  wire n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138;
  wire n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146;
  wire n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154;
  wire n_155, n_156, n_157, n_158, n_159, n_160, n_164, n_165;
  wire n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173;
  wire n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181;
  wire n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
  wire n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197;
  wire n_198, n_199, n_200, n_201, n_202, n_203, n_204, n_205;
  wire n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213;
  wire n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221;
  wire n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229;
  wire n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245;
  wire n_246, n_247, n_248, n_249, n_252, n_253, n_254, n_255;
  wire n_256, n_258, n_259, n_260, n_261, n_262, n_263, n_265;
  wire n_266, n_267, n_268, n_269, n_271, n_272, n_273, n_274;
  wire n_275, n_277, n_278, n_279, n_280, n_281, n_283, n_284;
  wire n_285, n_286, n_287, n_289, n_290, n_291, n_292, n_293;
  wire n_295, n_296, n_297, n_298, n_299, n_301, n_302, n_303;
  wire n_304, n_305, n_307, n_308, n_309, n_310, n_311, n_313;
  wire n_314, n_315, n_316, n_317, n_319, n_320, n_321, n_322;
  wire n_323, n_325, n_326, n_327, n_328, n_329, n_330, n_332;
  wire n_333, n_334, n_335, n_336, n_337, n_339, n_341, n_343;
  wire n_344, n_346, n_347, n_349, n_351, n_353, n_354, n_356;
  wire n_357, n_359, n_361, n_363, n_364, n_366, n_367, n_369;
  wire n_371, n_373, n_374, n_376, n_377, n_379, n_381, n_383;
  wire n_384, n_386, n_388, n_389, n_390, n_392, n_393, n_394;
  wire n_396, n_397, n_398, n_399, n_401, n_403, n_405, n_406;
  wire n_407, n_409, n_410, n_411, n_413, n_414, n_416, n_418;
  wire n_420, n_421, n_422, n_424, n_425, n_426, n_428, n_430;
  wire n_431, n_432, n_434, n_435, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_453, n_455, n_457, n_458, n_459;
  wire n_461, n_462, n_464, n_465, n_466, n_467, n_468, n_469;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_477, n_478;
  wire n_479, n_480, n_482, n_483, n_484, n_486, n_487, n_488;
  wire n_489, n_491, n_492, n_493, n_495, n_496, n_497, n_498;
  wire n_500, n_501, n_503, n_504, n_506, n_507, n_508, n_509;
  wire n_511, n_512, n_513, n_515, n_516, n_517, n_518, n_520;
  wire n_521, n_523, n_524, n_526, n_527, n_528, n_529, n_531;
  wire n_532, n_533, n_534, n_536, n_537, n_538;
  xor g27 (n_130, in_2[1], in_0[1]);
  and g2 (n_159, in_2[1], in_0[1]);
  xor g28 (n_128, in_2[2], n_159);
  xor g29 (n_155, n_128, in_0[2]);
  nand g3 (n_129, in_2[2], n_159);
  nand g30 (n_164, in_0[2], n_159);
  nand g31 (n_131, in_2[2], in_0[2]);
  nand g32 (n_160, n_129, n_164, n_131);
  xor g33 (n_165, in_2[3], in_0[3]);
  xor g34 (n_154, n_165, n_160);
  nand g35 (n_166, in_2[3], in_0[3]);
  nand g4 (n_167, n_160, in_0[3]);
  nand g36 (n_168, in_2[3], n_160);
  nand g37 (n_127, n_166, n_167, n_168);
  xor g38 (n_169, in_2[4], in_0[4]);
  xor g39 (n_153, n_169, in_1[4]);
  nand g40 (n_170, in_2[4], in_0[4]);
  nand g41 (n_171, in_1[4], in_0[4]);
  nand g5 (n_172, in_2[4], in_1[4]);
  nand g42 (n_126, n_170, n_171, n_172);
  xor g43 (n_173, in_2[5], in_0[5]);
  xor g44 (n_152, n_173, in_1[5]);
  nand g45 (n_174, in_2[5], in_0[5]);
  nand g46 (n_175, in_1[5], in_0[5]);
  nand g47 (n_176, in_2[5], in_1[5]);
  nand g6 (n_125, n_174, n_175, n_176);
  xor g48 (n_177, in_2[6], in_0[6]);
  xor g49 (n_151, n_177, in_1[6]);
  nand g50 (n_178, in_2[6], in_0[6]);
  nand g51 (n_179, in_1[6], in_0[6]);
  nand g52 (n_180, in_2[6], in_1[6]);
  nand g53 (n_124, n_178, n_179, n_180);
  xor g54 (n_181, in_2[7], in_0[7]);
  xor g55 (n_150, n_181, in_1[7]);
  nand g56 (n_182, in_2[7], in_0[7]);
  nand g57 (n_183, in_1[7], in_0[7]);
  nand g58 (n_184, in_2[7], in_1[7]);
  nand g59 (n_123, n_182, n_183, n_184);
  xor g60 (n_185, in_2[8], in_0[8]);
  xor g61 (n_149, n_185, in_1[8]);
  nand g62 (n_186, in_2[8], in_0[8]);
  nand g63 (n_187, in_1[8], in_0[8]);
  nand g64 (n_188, in_2[8], in_1[8]);
  nand g65 (n_122, n_186, n_187, n_188);
  xor g66 (n_156, in_2[9], in_0[9]);
  xor g67 (n_148, n_156, in_1[9]);
  nand g68 (n_157, in_2[9], in_0[9]);
  nand g69 (n_158, in_1[9], in_0[9]);
  nand g70 (n_189, in_2[9], in_1[9]);
  nand g71 (n_121, n_157, n_158, n_189);
  xor g72 (n_190, in_2[10], in_0[10]);
  xor g73 (n_147, n_190, in_1[10]);
  nand g74 (n_191, in_2[10], in_0[10]);
  nand g75 (n_192, in_1[10], in_0[10]);
  nand g76 (n_193, in_2[10], in_1[10]);
  nand g77 (n_120, n_191, n_192, n_193);
  xor g78 (n_194, in_2[11], in_0[11]);
  xor g79 (n_146, n_194, in_1[11]);
  nand g80 (n_195, in_2[11], in_0[11]);
  nand g81 (n_196, in_1[11], in_0[11]);
  nand g82 (n_197, in_2[11], in_1[11]);
  nand g83 (n_119, n_195, n_196, n_197);
  xor g84 (n_198, in_2[12], in_0[12]);
  xor g85 (n_145, n_198, in_1[12]);
  nand g86 (n_199, in_2[12], in_0[12]);
  nand g87 (n_200, in_1[12], in_0[12]);
  nand g88 (n_201, in_2[12], in_1[12]);
  nand g89 (n_118, n_199, n_200, n_201);
  xor g90 (n_202, in_2[13], in_0[13]);
  xor g91 (n_144, n_202, in_1[13]);
  nand g92 (n_203, in_2[13], in_0[13]);
  nand g93 (n_204, in_1[13], in_0[13]);
  nand g94 (n_205, in_2[13], in_1[13]);
  nand g95 (n_117, n_203, n_204, n_205);
  xor g96 (n_206, in_2[14], in_0[14]);
  xor g97 (n_143, n_206, in_1[14]);
  nand g98 (n_207, in_2[14], in_0[14]);
  nand g99 (n_208, in_1[14], in_0[14]);
  nand g100 (n_209, in_2[14], in_1[14]);
  nand g101 (n_116, n_207, n_208, n_209);
  xor g102 (n_210, in_2[15], in_0[15]);
  xor g103 (n_142, n_210, in_1[15]);
  nand g104 (n_211, in_2[15], in_0[15]);
  nand g105 (n_212, in_1[15], in_0[15]);
  nand g106 (n_213, in_2[15], in_1[15]);
  nand g107 (n_115, n_211, n_212, n_213);
  xor g108 (n_214, in_2[16], in_0[16]);
  xor g109 (n_141, n_214, in_1[16]);
  nand g110 (n_215, in_2[16], in_0[16]);
  nand g111 (n_216, in_1[16], in_0[16]);
  nand g112 (n_217, in_2[16], in_1[16]);
  nand g113 (n_114, n_215, n_216, n_217);
  xor g114 (n_218, in_2[17], in_0[17]);
  xor g115 (n_140, n_218, in_1[17]);
  nand g116 (n_219, in_2[17], in_0[17]);
  nand g117 (n_220, in_1[17], in_0[17]);
  nand g118 (n_221, in_2[17], in_1[17]);
  nand g119 (n_113, n_219, n_220, n_221);
  xor g120 (n_222, in_2[18], in_0[18]);
  xor g121 (n_139, n_222, in_1[18]);
  nand g122 (n_223, in_2[18], in_0[18]);
  nand g123 (n_224, in_1[18], in_0[18]);
  nand g124 (n_225, in_2[18], in_1[18]);
  nand g125 (n_112, n_223, n_224, n_225);
  xor g126 (n_226, in_2[19], in_0[19]);
  xor g127 (n_138, n_226, in_1[19]);
  nand g128 (n_227, in_2[19], in_0[19]);
  nand g129 (n_228, in_1[19], in_0[19]);
  nand g130 (n_229, in_2[19], in_1[19]);
  nand g131 (n_111, n_227, n_228, n_229);
  xor g132 (n_230, in_2[20], in_0[20]);
  xor g133 (n_137, n_230, in_1[20]);
  nand g134 (n_231, in_2[20], in_0[20]);
  nand g135 (n_232, in_1[20], in_0[20]);
  nand g136 (n_233, in_2[20], in_1[20]);
  nand g137 (n_110, n_231, n_232, n_233);
  xor g138 (n_234, in_2[21], in_0[21]);
  xor g139 (n_136, n_234, in_1[21]);
  nand g140 (n_235, in_2[21], in_0[21]);
  nand g141 (n_236, in_1[21], in_0[21]);
  nand g142 (n_237, in_2[21], in_1[21]);
  nand g143 (n_109, n_235, n_236, n_237);
  xor g144 (n_238, in_2[22], in_0[22]);
  xor g145 (n_135, n_238, in_1[22]);
  nand g146 (n_239, in_2[22], in_0[22]);
  nand g147 (n_240, in_1[22], in_0[22]);
  nand g148 (n_241, in_2[22], in_1[22]);
  nand g149 (n_108, n_239, n_240, n_241);
  xor g150 (n_242, in_2[23], in_0[23]);
  xor g151 (n_134, n_242, in_1[23]);
  nand g152 (n_243, in_2[23], in_0[23]);
  nand g153 (n_244, in_1[23], in_0[23]);
  nand g154 (n_245, in_2[23], in_1[23]);
  nand g155 (n_133, n_243, n_244, n_245);
  xor g158 (n_246, in_2[24], in_1[24]);
  xor g159 (n_107, n_246, in_0[24]);
  nand g160 (n_247, in_2[24], in_1[24]);
  nand g161 (n_248, in_0[24], in_1[24]);
  nand g162 (n_249, in_2[24], in_0[24]);
  nand g163 (n_132, n_247, n_248, n_249);
  xor g166 (n_538, in_1[0], in_0[0]);
  nand g167 (n_252, in_1[0], in_0[0]);
  nand g168 (n_253, in_1[0], in_2[0]);
  nand g7 (n_254, in_0[0], in_2[0]);
  nand g8 (n_256, n_252, n_253, n_254);
  nor g9 (n_255, n_130, in_1[1]);
  nand g10 (n_258, n_130, in_1[1]);
  nor g11 (n_265, in_1[2], n_155);
  nand g12 (n_260, in_1[2], n_155);
  nor g13 (n_261, in_1[3], n_154);
  nand g14 (n_262, in_1[3], n_154);
  nor g15 (n_271, n_127, n_153);
  nand g16 (n_266, n_127, n_153);
  nor g17 (n_267, n_126, n_152);
  nand g18 (n_268, n_126, n_152);
  nor g19 (n_277, n_125, n_151);
  nand g20 (n_272, n_125, n_151);
  nor g21 (n_273, n_124, n_150);
  nand g22 (n_274, n_124, n_150);
  nor g23 (n_283, n_123, n_149);
  nand g24 (n_278, n_123, n_149);
  nor g25 (n_279, n_122, n_148);
  nand g26 (n_280, n_122, n_148);
  nor g169 (n_289, n_121, n_147);
  nand g170 (n_284, n_121, n_147);
  nor g171 (n_285, n_120, n_146);
  nand g172 (n_286, n_120, n_146);
  nor g173 (n_295, n_119, n_145);
  nand g174 (n_290, n_119, n_145);
  nor g175 (n_291, n_118, n_144);
  nand g176 (n_292, n_118, n_144);
  nor g177 (n_301, n_117, n_143);
  nand g178 (n_296, n_117, n_143);
  nor g179 (n_297, n_116, n_142);
  nand g180 (n_298, n_116, n_142);
  nor g181 (n_307, n_115, n_141);
  nand g182 (n_302, n_115, n_141);
  nor g183 (n_303, n_114, n_140);
  nand g184 (n_304, n_114, n_140);
  nor g185 (n_313, n_113, n_139);
  nand g186 (n_308, n_113, n_139);
  nor g187 (n_309, n_112, n_138);
  nand g188 (n_310, n_112, n_138);
  nor g189 (n_319, n_111, n_137);
  nand g190 (n_314, n_111, n_137);
  nor g191 (n_315, n_110, n_136);
  nand g192 (n_316, n_110, n_136);
  nor g193 (n_325, n_109, n_135);
  nand g194 (n_320, n_109, n_135);
  nor g195 (n_321, n_108, n_134);
  nand g196 (n_322, n_108, n_134);
  nor g197 (n_329, n_107, n_133);
  nand g198 (n_326, n_107, n_133);
  nand g203 (n_330, n_258, n_259);
  nor g204 (n_263, n_260, n_261);
  nor g207 (n_333, n_265, n_261);
  nor g208 (n_269, n_266, n_267);
  nor g211 (n_339, n_271, n_267);
  nor g212 (n_275, n_272, n_273);
  nor g215 (n_341, n_277, n_273);
  nor g216 (n_281, n_278, n_279);
  nor g219 (n_349, n_283, n_279);
  nor g220 (n_287, n_284, n_285);
  nor g223 (n_351, n_289, n_285);
  nor g224 (n_293, n_290, n_291);
  nor g227 (n_359, n_295, n_291);
  nor g228 (n_299, n_296, n_297);
  nor g231 (n_361, n_301, n_297);
  nor g232 (n_305, n_302, n_303);
  nor g235 (n_369, n_307, n_303);
  nor g236 (n_311, n_308, n_309);
  nor g239 (n_371, n_313, n_309);
  nor g240 (n_317, n_314, n_315);
  nor g243 (n_379, n_319, n_315);
  nor g244 (n_323, n_320, n_321);
  nor g247 (n_381, n_325, n_321);
  nand g250 (n_482, n_260, n_332);
  nand g251 (n_335, n_333, n_330);
  nand g252 (n_386, n_334, n_335);
  nor g253 (n_337, n_277, n_336);
  nand g262 (n_394, n_339, n_341);
  nor g263 (n_347, n_289, n_346);
  nand g272 (n_401, n_349, n_351);
  nor g273 (n_357, n_301, n_356);
  nand g282 (n_409, n_359, n_361);
  nor g283 (n_367, n_313, n_366);
  nand g292 (n_416, n_369, n_371);
  nor g293 (n_377, n_325, n_376);
  nand g302 (n_424, n_379, n_381);
  nand g305 (n_486, n_266, n_388);
  nand g306 (n_389, n_339, n_386);
  nand g307 (n_488, n_336, n_389);
  nand g310 (n_491, n_392, n_393);
  nand g313 (n_428, n_396, n_397);
  nor g314 (n_399, n_295, n_398);
  nor g317 (n_438, n_295, n_401);
  nor g323 (n_407, n_405, n_398);
  nor g326 (n_444, n_401, n_405);
  nor g327 (n_411, n_409, n_398);
  nor g330 (n_447, n_401, n_409);
  nor g331 (n_414, n_319, n_413);
  nor g334 (n_465, n_319, n_416);
  nor g340 (n_422, n_420, n_413);
  nor g343 (n_471, n_416, n_420);
  nor g344 (n_426, n_424, n_413);
  nor g347 (n_453, n_416, n_424);
  nand g350 (n_495, n_278, n_430);
  nand g351 (n_431, n_349, n_428);
  nand g352 (n_497, n_346, n_431);
  nand g355 (n_500, n_434, n_435);
  nand g358 (n_503, n_398, n_437);
  nand g359 (n_440, n_438, n_428);
  nand g360 (n_506, n_439, n_440);
  nand g361 (n_443, n_441, n_428);
  nand g362 (n_508, n_442, n_443);
  nand g363 (n_446, n_444, n_428);
  nand g364 (n_511, n_445, n_446);
  nand g365 (n_449, n_447, n_428);
  nand g366 (n_455, n_448, n_449);
  nor g367 (n_451, n_329, n_450);
  nand g374 (n_515, n_302, n_457);
  nand g375 (n_458, n_369, n_455);
  nand g376 (n_517, n_366, n_458);
  nand g379 (n_520, n_461, n_462);
  nand g382 (n_523, n_413, n_464);
  nand g383 (n_467, n_465, n_455);
  nand g384 (n_526, n_466, n_467);
  nand g385 (n_470, n_468, n_455);
  nand g386 (n_528, n_469, n_470);
  nand g387 (n_473, n_471, n_455);
  nand g388 (n_531, n_472, n_473);
  nand g389 (n_474, n_453, n_455);
  nand g390 (n_533, n_450, n_474);
  nand g393 (n_536, n_477, n_478);
  xnor g395 (out_0[1], n_256, n_479);
  xnor g397 (out_0[2], n_330, n_480);
  xnor g400 (out_0[3], n_482, n_483);
  xnor g402 (out_0[4], n_386, n_484);
  xnor g405 (out_0[5], n_486, n_487);
  xnor g407 (out_0[6], n_488, n_489);
  xnor g410 (out_0[7], n_491, n_492);
  xnor g412 (out_0[8], n_428, n_493);
  xnor g415 (out_0[9], n_495, n_496);
  xnor g417 (out_0[10], n_497, n_498);
  xnor g420 (out_0[11], n_500, n_501);
  xnor g423 (out_0[12], n_503, n_504);
  xnor g426 (out_0[13], n_506, n_507);
  xnor g428 (out_0[14], n_508, n_509);
  xnor g431 (out_0[15], n_511, n_512);
  xnor g433 (out_0[16], n_455, n_513);
  xnor g436 (out_0[17], n_515, n_516);
  xnor g438 (out_0[18], n_517, n_518);
  xnor g441 (out_0[19], n_520, n_521);
  xnor g444 (out_0[20], n_523, n_524);
  xnor g447 (out_0[21], n_526, n_527);
  xnor g449 (out_0[22], n_528, n_529);
  xnor g452 (out_0[23], n_531, n_532);
  xnor g454 (out_0[24], n_533, n_534);
  xnor g457 (out_0[25], n_536, n_537);
  xor g458 (out_0[0], in_2[0], n_538);
  or g459 (n_259, n_255, wc);
  not gc (wc, n_256);
  or g460 (n_479, wc0, n_255);
  not gc0 (wc0, n_258);
  and g461 (n_343, wc1, n_274);
  not gc1 (wc1, n_275);
  and g462 (n_346, wc2, n_280);
  not gc2 (wc2, n_281);
  and g463 (n_353, wc3, n_286);
  not gc3 (wc3, n_287);
  and g464 (n_356, wc4, n_292);
  not gc4 (wc4, n_293);
  and g465 (n_363, wc5, n_298);
  not gc5 (wc5, n_299);
  and g466 (n_366, wc6, n_304);
  not gc6 (wc6, n_305);
  and g467 (n_373, wc7, n_310);
  not gc7 (wc7, n_311);
  and g468 (n_376, wc8, n_316);
  not gc8 (wc8, n_317);
  and g469 (n_383, wc9, n_322);
  not gc9 (wc9, n_323);
  or g470 (n_432, wc10, n_289);
  not gc10 (wc10, n_349);
  or g471 (n_405, wc11, n_301);
  not gc11 (wc11, n_359);
  or g472 (n_459, wc12, n_313);
  not gc12 (wc12, n_369);
  or g473 (n_420, wc13, n_325);
  not gc13 (wc13, n_379);
  or g474 (n_487, wc14, n_267);
  not gc14 (wc14, n_268);
  or g475 (n_489, wc15, n_277);
  not gc15 (wc15, n_272);
  or g476 (n_492, wc16, n_273);
  not gc16 (wc16, n_274);
  or g477 (n_493, wc17, n_283);
  not gc17 (wc17, n_278);
  or g478 (n_496, wc18, n_279);
  not gc18 (wc18, n_280);
  or g479 (n_498, wc19, n_289);
  not gc19 (wc19, n_284);
  or g480 (n_501, wc20, n_285);
  not gc20 (wc20, n_286);
  or g481 (n_504, wc21, n_295);
  not gc21 (wc21, n_290);
  or g482 (n_507, wc22, n_291);
  not gc22 (wc22, n_292);
  or g483 (n_509, wc23, n_301);
  not gc23 (wc23, n_296);
  or g484 (n_512, wc24, n_297);
  not gc24 (wc24, n_298);
  or g485 (n_513, wc25, n_307);
  not gc25 (wc25, n_302);
  or g486 (n_516, wc26, n_303);
  not gc26 (wc26, n_304);
  or g487 (n_518, wc27, n_313);
  not gc27 (wc27, n_308);
  or g488 (n_521, wc28, n_309);
  not gc28 (wc28, n_310);
  or g489 (n_524, wc29, n_319);
  not gc29 (wc29, n_314);
  or g490 (n_527, wc30, n_315);
  not gc30 (wc30, n_316);
  or g491 (n_529, wc31, n_325);
  not gc31 (wc31, n_320);
  or g492 (n_532, wc32, n_321);
  not gc32 (wc32, n_322);
  and g493 (n_327, wc33, n_132);
  not gc33 (wc33, in_2[24]);
  or g494 (n_328, wc34, n_132);
  not gc34 (wc34, in_2[24]);
  or g495 (n_332, wc35, n_265);
  not gc35 (wc35, n_330);
  and g496 (n_354, wc36, n_351);
  not gc36 (wc36, n_346);
  and g497 (n_364, wc37, n_361);
  not gc37 (wc37, n_356);
  and g498 (n_374, wc38, n_371);
  not gc38 (wc38, n_366);
  and g499 (n_384, wc39, n_381);
  not gc39 (wc39, n_376);
  and g500 (n_441, wc40, n_359);
  not gc40 (wc40, n_401);
  and g501 (n_468, wc41, n_379);
  not gc41 (wc41, n_416);
  or g502 (n_480, wc42, n_265);
  not gc42 (wc42, n_260);
  and g503 (n_334, wc43, n_262);
  not gc43 (wc43, n_263);
  and g504 (n_434, wc44, n_284);
  not gc44 (wc44, n_347);
  and g505 (n_398, wc45, n_353);
  not gc45 (wc45, n_354);
  and g506 (n_406, wc46, n_296);
  not gc46 (wc46, n_357);
  and g507 (n_410, wc47, n_363);
  not gc47 (wc47, n_364);
  and g508 (n_461, wc48, n_308);
  not gc48 (wc48, n_367);
  and g509 (n_413, wc49, n_373);
  not gc49 (wc49, n_374);
  and g510 (n_421, wc50, n_320);
  not gc50 (wc50, n_377);
  and g511 (n_425, wc51, n_383);
  not gc51 (wc51, n_384);
  or g512 (n_475, wc52, n_329);
  not gc52 (wc52, n_453);
  or g513 (n_483, wc53, n_261);
  not gc53 (wc53, n_262);
  or g514 (n_534, wc54, n_329);
  not gc54 (wc54, n_326);
  and g515 (n_336, wc55, n_268);
  not gc55 (wc55, n_269);
  or g516 (n_390, wc56, n_277);
  not gc56 (wc56, n_339);
  and g517 (n_403, wc57, n_359);
  not gc57 (wc57, n_398);
  and g518 (n_418, wc58, n_379);
  not gc58 (wc58, n_413);
  or g519 (n_484, wc59, n_271);
  not gc59 (wc59, n_266);
  or g520 (n_537, wc60, n_327);
  not gc60 (wc60, n_328);
  and g521 (n_344, wc61, n_341);
  not gc61 (wc61, n_336);
  or g522 (n_388, wc62, n_271);
  not gc62 (wc62, n_386);
  and g523 (n_439, wc63, n_290);
  not gc63 (wc63, n_399);
  and g524 (n_442, wc64, n_356);
  not gc64 (wc64, n_403);
  and g525 (n_445, n_406, wc65);
  not gc65 (wc65, n_407);
  and g526 (n_448, n_410, wc66);
  not gc66 (wc66, n_411);
  and g527 (n_466, wc67, n_314);
  not gc67 (wc67, n_414);
  and g528 (n_469, wc68, n_376);
  not gc68 (wc68, n_418);
  and g529 (n_472, n_421, wc69);
  not gc69 (wc69, n_422);
  and g530 (n_450, n_425, wc70);
  not gc70 (wc70, n_426);
  and g531 (n_392, wc71, n_272);
  not gc71 (wc71, n_337);
  and g532 (n_396, wc72, n_343);
  not gc72 (wc72, n_344);
  or g533 (n_393, n_390, wc73);
  not gc73 (wc73, n_386);
  or g534 (n_397, n_394, wc74);
  not gc74 (wc74, n_386);
  and g535 (n_477, wc75, n_326);
  not gc75 (wc75, n_451);
  or g536 (n_430, wc76, n_283);
  not gc76 (wc76, n_428);
  or g537 (n_435, n_432, wc77);
  not gc77 (wc77, n_428);
  or g538 (n_437, wc78, n_401);
  not gc78 (wc78, n_428);
  or g539 (n_457, wc79, n_307);
  not gc79 (wc79, n_455);
  or g540 (n_462, n_459, wc80);
  not gc80 (wc80, n_455);
  or g541 (n_464, wc81, n_416);
  not gc81 (wc81, n_455);
  or g542 (n_478, n_475, wc82);
  not gc82 (wc82, n_455);
endmodule

module csa_tree_add_287_40_group_6803_GENERIC(in_0, in_1, in_2, out_0);
  input [26:0] in_0, in_1;
  input [24:0] in_2;
  output [25:0] out_0;
  wire [26:0] in_0, in_1;
  wire [24:0] in_2;
  wire [25:0] out_0;
  csa_tree_add_287_40_group_6803_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .out_0 (out_0));
endmodule

module csa_tree_add_329_38_group_6821_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_329_38_group_6821_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_329_38_group_6821_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_402_38_group_6813_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_402_38_group_6813_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_402_38_group_6813_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_475_38_group_6815_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_475_38_group_6815_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_475_38_group_6815_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_548_38_group_6817_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_548_38_group_6817_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_548_38_group_6817_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_621_38_group_6819_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_621_38_group_6819_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_621_38_group_6819_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_694_38_group_6811_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  wire n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169;
  wire n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_194;
  wire n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234;
  wire n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242;
  wire n_243, n_244, n_245, n_246, n_247, n_248, n_249, n_250;
  wire n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258;
  wire n_259, n_260, n_261, n_262, n_268, n_269, n_270, n_271;
  wire n_272, n_275, n_277, n_278, n_279, n_280, n_281, n_282;
  wire n_283, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_294, n_295, n_296, n_297, n_298;
  wire n_299, n_300, n_301, n_302, n_303, n_304, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330;
  wire n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_346;
  wire n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362;
  wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434;
  wire n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442;
  wire n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450;
  wire n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_520, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_532, n_533, n_534, n_535;
  wire n_536, n_538, n_539, n_540, n_541, n_542, n_543, n_545;
  wire n_546, n_547, n_548, n_549, n_551, n_552, n_553, n_554;
  wire n_555, n_557, n_558, n_559, n_560, n_561, n_563, n_564;
  wire n_565, n_566, n_567, n_569, n_570, n_571, n_572, n_573;
  wire n_575, n_576, n_577, n_578, n_579, n_581, n_582, n_583;
  wire n_584, n_585, n_587, n_588, n_589, n_590, n_591, n_593;
  wire n_594, n_595, n_596, n_597, n_599, n_600, n_601, n_602;
  wire n_603, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_614, n_616, n_618, n_619, n_621, n_622, n_624, n_626;
  wire n_628, n_629, n_631, n_632, n_634, n_636, n_638, n_639;
  wire n_641, n_642, n_644, n_646, n_648, n_649, n_651, n_652;
  wire n_654, n_656, n_658, n_659, n_661, n_663, n_664, n_665;
  wire n_667, n_668, n_669, n_671, n_672, n_673, n_674, n_676;
  wire n_678, n_680, n_681, n_682, n_684, n_685, n_686, n_688;
  wire n_689, n_691, n_693, n_695, n_696, n_697, n_699, n_700;
  wire n_701, n_703, n_705, n_706, n_707, n_709, n_710, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_719, n_720;
  wire n_721, n_722, n_723, n_724, n_726, n_728, n_730, n_732;
  wire n_733, n_734, n_736, n_737, n_739, n_740, n_741, n_742;
  wire n_743, n_744, n_745, n_746, n_747, n_748, n_749, n_750;
  wire n_751, n_753, n_754, n_755, n_757, n_758, n_759, n_760;
  wire n_762, n_763, n_764, n_766, n_767, n_768, n_769, n_771;
  wire n_772, n_774, n_775, n_777, n_778, n_779, n_780, n_782;
  wire n_783, n_784, n_786, n_787, n_788, n_789, n_791, n_792;
  wire n_794, n_795, n_797, n_798, n_799, n_800, n_802, n_803;
  wire n_804, n_806;
  xor g72 (n_278, in_0[0], in_4[0]);
  xor g73 (n_185, n_278, in_3[0]);
  nand g74 (n_279, in_0[0], in_4[0]);
  nand g75 (n_280, in_3[0], in_4[0]);
  nand g76 (n_281, in_0[0], in_3[0]);
  nand g6 (n_187, n_279, n_280, n_281);
  xor g77 (n_282, in_0[1], in_1[1]);
  xor g78 (n_159, n_282, in_4[1]);
  nand g79 (n_283, in_0[1], in_1[1]);
  nand g80 (n_284, in_4[1], in_1[1]);
  nand g81 (n_285, in_0[1], in_4[1]);
  nand g82 (n_189, n_283, n_284, n_285);
  xor g83 (n_286, in_3[1], in_2[1]);
  xor g84 (n_184, n_286, n_187);
  nand g85 (n_287, in_3[1], in_2[1]);
  nand g86 (n_288, n_187, in_2[1]);
  nand g87 (n_289, in_3[1], n_187);
  nand g88 (n_158, n_287, n_288, n_289);
  xor g89 (n_188, in_0[2], in_1[2]);
  and g90 (n_191, in_0[2], in_1[2]);
  xor g91 (n_290, in_3[2], in_4[2]);
  xor g92 (n_190, n_290, in_2[2]);
  nand g93 (n_291, in_3[2], in_4[2]);
  nand g94 (n_292, in_2[2], in_4[2]);
  nand g95 (n_293, in_3[2], in_2[2]);
  nand g96 (n_192, n_291, n_292, n_293);
  xor g97 (n_294, n_188, n_189);
  xor g98 (n_183, n_294, n_190);
  nand g99 (n_295, n_188, n_189);
  nand g100 (n_296, n_190, n_189);
  nand g101 (n_297, n_188, n_190);
  nand g102 (n_157, n_295, n_296, n_297);
  xor g103 (n_298, in_0[3], in_1[3]);
  xor g104 (n_193, n_298, in_3[3]);
  nand g105 (n_299, in_0[3], in_1[3]);
  nand g106 (n_300, in_3[3], in_1[3]);
  nand g107 (n_301, in_0[3], in_3[3]);
  nand g108 (n_195, n_299, n_300, n_301);
  xor g109 (n_302, in_4[3], in_2[3]);
  xor g110 (n_194, n_302, n_191);
  nand g111 (n_303, in_4[3], in_2[3]);
  nand g112 (n_304, n_191, in_2[3]);
  nand g113 (n_305, in_4[3], n_191);
  nand g114 (n_197, n_303, n_304, n_305);
  xor g115 (n_306, n_192, n_193);
  xor g116 (n_182, n_306, n_194);
  nand g117 (n_307, n_192, n_193);
  nand g118 (n_308, n_194, n_193);
  nand g119 (n_309, n_192, n_194);
  nand g120 (n_156, n_307, n_308, n_309);
  xor g121 (n_310, in_0[4], in_1[4]);
  xor g122 (n_196, n_310, in_3[4]);
  nand g123 (n_311, in_0[4], in_1[4]);
  nand g124 (n_312, in_3[4], in_1[4]);
  nand g125 (n_313, in_0[4], in_3[4]);
  nand g126 (n_199, n_311, n_312, n_313);
  xor g127 (n_314, in_4[4], in_2[4]);
  xor g128 (n_198, n_314, n_195);
  nand g129 (n_315, in_4[4], in_2[4]);
  nand g130 (n_316, n_195, in_2[4]);
  nand g131 (n_317, in_4[4], n_195);
  nand g132 (n_202, n_315, n_316, n_317);
  xor g133 (n_318, n_196, n_197);
  xor g134 (n_181, n_318, n_198);
  nand g135 (n_319, n_196, n_197);
  nand g136 (n_320, n_198, n_197);
  nand g137 (n_321, n_196, n_198);
  nand g138 (n_155, n_319, n_320, n_321);
  xor g139 (n_322, in_0[5], in_1[5]);
  xor g140 (n_200, n_322, in_3[5]);
  nand g141 (n_323, in_0[5], in_1[5]);
  nand g142 (n_324, in_3[5], in_1[5]);
  nand g143 (n_325, in_0[5], in_3[5]);
  nand g144 (n_203, n_323, n_324, n_325);
  xor g145 (n_326, in_4[5], in_2[5]);
  xor g146 (n_201, n_326, n_199);
  nand g147 (n_327, in_4[5], in_2[5]);
  nand g148 (n_328, n_199, in_2[5]);
  nand g149 (n_329, in_4[5], n_199);
  nand g150 (n_206, n_327, n_328, n_329);
  xor g151 (n_330, n_200, n_201);
  xor g152 (n_180, n_330, n_202);
  nand g153 (n_331, n_200, n_201);
  nand g154 (n_332, n_202, n_201);
  nand g155 (n_333, n_200, n_202);
  nand g156 (n_154, n_331, n_332, n_333);
  xor g157 (n_334, in_0[6], in_1[6]);
  xor g158 (n_204, n_334, in_3[6]);
  nand g159 (n_335, in_0[6], in_1[6]);
  nand g160 (n_336, in_3[6], in_1[6]);
  nand g161 (n_337, in_0[6], in_3[6]);
  nand g162 (n_207, n_335, n_336, n_337);
  xor g163 (n_338, in_4[6], in_2[6]);
  xor g164 (n_205, n_338, n_203);
  nand g165 (n_339, in_4[6], in_2[6]);
  nand g166 (n_340, n_203, in_2[6]);
  nand g167 (n_341, in_4[6], n_203);
  nand g168 (n_210, n_339, n_340, n_341);
  xor g169 (n_342, n_204, n_205);
  xor g170 (n_179, n_342, n_206);
  nand g171 (n_343, n_204, n_205);
  nand g172 (n_344, n_206, n_205);
  nand g173 (n_345, n_204, n_206);
  nand g174 (n_153, n_343, n_344, n_345);
  xor g175 (n_346, in_0[7], in_1[7]);
  xor g176 (n_208, n_346, in_3[7]);
  nand g177 (n_347, in_0[7], in_1[7]);
  nand g178 (n_348, in_3[7], in_1[7]);
  nand g179 (n_349, in_0[7], in_3[7]);
  nand g180 (n_211, n_347, n_348, n_349);
  xor g181 (n_350, in_4[7], in_2[7]);
  xor g182 (n_209, n_350, n_207);
  nand g183 (n_351, in_4[7], in_2[7]);
  nand g184 (n_352, n_207, in_2[7]);
  nand g185 (n_353, in_4[7], n_207);
  nand g186 (n_214, n_351, n_352, n_353);
  xor g187 (n_354, n_208, n_209);
  xor g188 (n_178, n_354, n_210);
  nand g189 (n_355, n_208, n_209);
  nand g190 (n_356, n_210, n_209);
  nand g191 (n_357, n_208, n_210);
  nand g192 (n_152, n_355, n_356, n_357);
  xor g193 (n_358, in_0[8], in_1[8]);
  xor g194 (n_212, n_358, in_3[8]);
  nand g195 (n_359, in_0[8], in_1[8]);
  nand g196 (n_360, in_3[8], in_1[8]);
  nand g197 (n_361, in_0[8], in_3[8]);
  nand g198 (n_215, n_359, n_360, n_361);
  xor g199 (n_362, in_4[8], in_2[8]);
  xor g200 (n_213, n_362, n_211);
  nand g201 (n_363, in_4[8], in_2[8]);
  nand g202 (n_364, n_211, in_2[8]);
  nand g203 (n_365, in_4[8], n_211);
  nand g204 (n_218, n_363, n_364, n_365);
  xor g205 (n_366, n_212, n_213);
  xor g206 (n_177, n_366, n_214);
  nand g207 (n_367, n_212, n_213);
  nand g208 (n_368, n_214, n_213);
  nand g209 (n_369, n_212, n_214);
  nand g210 (n_151, n_367, n_368, n_369);
  xor g211 (n_370, in_0[9], in_1[9]);
  xor g212 (n_216, n_370, in_3[9]);
  nand g213 (n_371, in_0[9], in_1[9]);
  nand g214 (n_372, in_3[9], in_1[9]);
  nand g215 (n_373, in_0[9], in_3[9]);
  nand g216 (n_219, n_371, n_372, n_373);
  xor g217 (n_374, in_4[9], in_2[9]);
  xor g218 (n_217, n_374, n_215);
  nand g219 (n_375, in_4[9], in_2[9]);
  nand g220 (n_376, n_215, in_2[9]);
  nand g221 (n_377, in_4[9], n_215);
  nand g222 (n_222, n_375, n_376, n_377);
  xor g223 (n_378, n_216, n_217);
  xor g224 (n_176, n_378, n_218);
  nand g225 (n_379, n_216, n_217);
  nand g226 (n_380, n_218, n_217);
  nand g227 (n_381, n_216, n_218);
  nand g228 (n_150, n_379, n_380, n_381);
  xor g229 (n_382, in_0[10], in_1[10]);
  xor g230 (n_220, n_382, in_3[10]);
  nand g231 (n_383, in_0[10], in_1[10]);
  nand g232 (n_384, in_3[10], in_1[10]);
  nand g233 (n_385, in_0[10], in_3[10]);
  nand g234 (n_223, n_383, n_384, n_385);
  xor g235 (n_386, in_4[10], in_2[10]);
  xor g236 (n_221, n_386, n_219);
  nand g237 (n_387, in_4[10], in_2[10]);
  nand g238 (n_388, n_219, in_2[10]);
  nand g239 (n_389, in_4[10], n_219);
  nand g240 (n_226, n_387, n_388, n_389);
  xor g241 (n_390, n_220, n_221);
  xor g242 (n_175, n_390, n_222);
  nand g243 (n_391, n_220, n_221);
  nand g244 (n_392, n_222, n_221);
  nand g245 (n_393, n_220, n_222);
  nand g246 (n_149, n_391, n_392, n_393);
  xor g247 (n_394, in_0[11], in_1[11]);
  xor g248 (n_224, n_394, in_3[11]);
  nand g249 (n_395, in_0[11], in_1[11]);
  nand g250 (n_396, in_3[11], in_1[11]);
  nand g251 (n_397, in_0[11], in_3[11]);
  nand g252 (n_227, n_395, n_396, n_397);
  xor g253 (n_398, in_4[11], in_2[11]);
  xor g254 (n_225, n_398, n_223);
  nand g255 (n_399, in_4[11], in_2[11]);
  nand g256 (n_400, n_223, in_2[11]);
  nand g257 (n_401, in_4[11], n_223);
  nand g258 (n_230, n_399, n_400, n_401);
  xor g259 (n_402, n_224, n_225);
  xor g260 (n_174, n_402, n_226);
  nand g261 (n_403, n_224, n_225);
  nand g262 (n_404, n_226, n_225);
  nand g263 (n_405, n_224, n_226);
  nand g264 (n_148, n_403, n_404, n_405);
  xor g265 (n_406, in_0[12], in_1[12]);
  xor g266 (n_228, n_406, in_3[12]);
  nand g267 (n_407, in_0[12], in_1[12]);
  nand g268 (n_408, in_3[12], in_1[12]);
  nand g269 (n_409, in_0[12], in_3[12]);
  nand g270 (n_231, n_407, n_408, n_409);
  xor g271 (n_410, in_4[12], in_2[12]);
  xor g272 (n_229, n_410, n_227);
  nand g273 (n_411, in_4[12], in_2[12]);
  nand g274 (n_412, n_227, in_2[12]);
  nand g275 (n_413, in_4[12], n_227);
  nand g276 (n_234, n_411, n_412, n_413);
  xor g277 (n_414, n_228, n_229);
  xor g278 (n_173, n_414, n_230);
  nand g279 (n_415, n_228, n_229);
  nand g280 (n_416, n_230, n_229);
  nand g281 (n_417, n_228, n_230);
  nand g282 (n_147, n_415, n_416, n_417);
  xor g283 (n_418, in_0[13], in_1[13]);
  xor g284 (n_232, n_418, in_3[13]);
  nand g285 (n_419, in_0[13], in_1[13]);
  nand g286 (n_420, in_3[13], in_1[13]);
  nand g287 (n_421, in_0[13], in_3[13]);
  nand g288 (n_235, n_419, n_420, n_421);
  xor g289 (n_422, in_4[13], in_2[13]);
  xor g290 (n_233, n_422, n_231);
  nand g291 (n_423, in_4[13], in_2[13]);
  nand g292 (n_424, n_231, in_2[13]);
  nand g293 (n_425, in_4[13], n_231);
  nand g294 (n_238, n_423, n_424, n_425);
  xor g295 (n_426, n_232, n_233);
  xor g296 (n_172, n_426, n_234);
  nand g297 (n_427, n_232, n_233);
  nand g298 (n_428, n_234, n_233);
  nand g299 (n_429, n_232, n_234);
  nand g300 (n_146, n_427, n_428, n_429);
  xor g301 (n_430, in_0[14], in_1[14]);
  xor g302 (n_236, n_430, in_3[14]);
  nand g303 (n_431, in_0[14], in_1[14]);
  nand g304 (n_432, in_3[14], in_1[14]);
  nand g305 (n_433, in_0[14], in_3[14]);
  nand g306 (n_239, n_431, n_432, n_433);
  xor g307 (n_434, in_4[14], in_2[14]);
  xor g308 (n_237, n_434, n_235);
  nand g309 (n_435, in_4[14], in_2[14]);
  nand g310 (n_436, n_235, in_2[14]);
  nand g311 (n_437, in_4[14], n_235);
  nand g312 (n_242, n_435, n_436, n_437);
  xor g313 (n_438, n_236, n_237);
  xor g314 (n_171, n_438, n_238);
  nand g315 (n_439, n_236, n_237);
  nand g316 (n_440, n_238, n_237);
  nand g317 (n_441, n_236, n_238);
  nand g318 (n_145, n_439, n_440, n_441);
  xor g319 (n_442, in_0[15], in_1[15]);
  xor g320 (n_240, n_442, in_3[15]);
  nand g321 (n_443, in_0[15], in_1[15]);
  nand g322 (n_444, in_3[15], in_1[15]);
  nand g323 (n_445, in_0[15], in_3[15]);
  nand g324 (n_243, n_443, n_444, n_445);
  xor g325 (n_446, in_4[15], in_2[15]);
  xor g326 (n_241, n_446, n_239);
  nand g327 (n_447, in_4[15], in_2[15]);
  nand g328 (n_448, n_239, in_2[15]);
  nand g329 (n_449, in_4[15], n_239);
  nand g330 (n_246, n_447, n_448, n_449);
  xor g331 (n_450, n_240, n_241);
  xor g332 (n_170, n_450, n_242);
  nand g333 (n_451, n_240, n_241);
  nand g334 (n_452, n_242, n_241);
  nand g335 (n_453, n_240, n_242);
  nand g336 (n_144, n_451, n_452, n_453);
  xor g337 (n_454, in_0[16], in_1[16]);
  xor g338 (n_244, n_454, in_3[16]);
  nand g339 (n_455, in_0[16], in_1[16]);
  nand g340 (n_456, in_3[16], in_1[16]);
  nand g341 (n_457, in_0[16], in_3[16]);
  nand g342 (n_247, n_455, n_456, n_457);
  xor g343 (n_458, in_4[16], in_2[16]);
  xor g344 (n_245, n_458, n_243);
  nand g345 (n_459, in_4[16], in_2[16]);
  nand g346 (n_460, n_243, in_2[16]);
  nand g347 (n_461, in_4[16], n_243);
  nand g348 (n_250, n_459, n_460, n_461);
  xor g349 (n_462, n_244, n_245);
  xor g350 (n_169, n_462, n_246);
  nand g351 (n_463, n_244, n_245);
  nand g352 (n_464, n_246, n_245);
  nand g353 (n_465, n_244, n_246);
  nand g354 (n_143, n_463, n_464, n_465);
  xor g355 (n_466, in_0[17], in_1[17]);
  xor g356 (n_248, n_466, in_3[17]);
  nand g357 (n_467, in_0[17], in_1[17]);
  nand g358 (n_468, in_3[17], in_1[17]);
  nand g359 (n_469, in_0[17], in_3[17]);
  nand g360 (n_251, n_467, n_468, n_469);
  xor g361 (n_470, in_4[17], in_2[17]);
  xor g362 (n_249, n_470, n_247);
  nand g363 (n_471, in_4[17], in_2[17]);
  nand g364 (n_472, n_247, in_2[17]);
  nand g365 (n_473, in_4[17], n_247);
  nand g366 (n_254, n_471, n_472, n_473);
  xor g367 (n_474, n_248, n_249);
  xor g368 (n_168, n_474, n_250);
  nand g369 (n_475, n_248, n_249);
  nand g370 (n_476, n_250, n_249);
  nand g371 (n_477, n_248, n_250);
  nand g372 (n_142, n_475, n_476, n_477);
  xor g373 (n_478, in_0[18], in_1[18]);
  xor g374 (n_252, n_478, in_3[18]);
  nand g375 (n_479, in_0[18], in_1[18]);
  nand g376 (n_480, in_3[18], in_1[18]);
  nand g377 (n_481, in_0[18], in_3[18]);
  nand g378 (n_255, n_479, n_480, n_481);
  xor g379 (n_482, in_4[18], in_2[18]);
  xor g380 (n_253, n_482, n_251);
  nand g381 (n_483, in_4[18], in_2[18]);
  nand g382 (n_484, n_251, in_2[18]);
  nand g383 (n_485, in_4[18], n_251);
  nand g384 (n_258, n_483, n_484, n_485);
  xor g385 (n_486, n_252, n_253);
  xor g386 (n_167, n_486, n_254);
  nand g387 (n_487, n_252, n_253);
  nand g388 (n_488, n_254, n_253);
  nand g389 (n_489, n_252, n_254);
  nand g390 (n_141, n_487, n_488, n_489);
  xor g391 (n_490, in_0[19], in_1[19]);
  xor g392 (n_256, n_490, in_3[19]);
  nand g393 (n_491, in_0[19], in_1[19]);
  nand g394 (n_492, in_3[19], in_1[19]);
  nand g395 (n_493, in_0[19], in_3[19]);
  nand g396 (n_259, n_491, n_492, n_493);
  xor g397 (n_494, in_4[19], in_2[19]);
  xor g398 (n_257, n_494, n_255);
  nand g399 (n_495, in_4[19], in_2[19]);
  nand g400 (n_496, n_255, in_2[19]);
  nand g401 (n_497, in_4[19], n_255);
  nand g402 (n_262, n_495, n_496, n_497);
  xor g403 (n_498, n_256, n_257);
  xor g404 (n_166, n_498, n_258);
  nand g405 (n_499, n_256, n_257);
  nand g406 (n_500, n_258, n_257);
  nand g407 (n_501, n_256, n_258);
  nand g408 (n_140, n_499, n_500, n_501);
  xor g409 (n_502, in_0[20], in_1[20]);
  xor g410 (n_260, n_502, in_3[20]);
  nand g411 (n_503, in_0[20], in_1[20]);
  nand g412 (n_504, in_3[20], in_1[20]);
  nand g413 (n_505, in_0[20], in_3[20]);
  nand g414 (n_269, n_503, n_504, n_505);
  xor g415 (n_506, in_4[20], in_2[20]);
  xor g416 (n_261, n_506, n_259);
  nand g417 (n_507, in_4[20], in_2[20]);
  nand g418 (n_508, n_259, in_2[20]);
  nand g419 (n_509, in_4[20], n_259);
  nand g420 (n_272, n_507, n_508, n_509);
  xor g421 (n_510, n_260, n_261);
  xor g422 (n_165, n_510, n_262);
  nand g423 (n_511, n_260, n_261);
  nand g424 (n_512, n_262, n_261);
  nand g425 (n_513, n_260, n_262);
  nand g426 (n_139, n_511, n_512, n_513);
  nand g434 (n_275, n_515, n_516, n_517);
  nand g438 (n_520, n_269, n_268);
  xor g441 (n_522, n_270, n_271);
  xor g442 (n_164, n_522, n_272);
  nand g443 (n_523, n_270, n_271);
  nand g444 (n_524, n_272, n_271);
  nand g445 (n_525, n_270, n_272);
  nand g446 (n_138, n_523, n_524, n_525);
  xor g450 (n_163, n_526, n_277);
  nand g453 (n_529, n_275, n_277);
  nand g454 (n_162, n_527, n_528, n_529);
  xor g457 (n_806, in_1[0], n_185);
  nand g458 (n_532, in_1[0], n_185);
  nand g459 (n_533, in_1[0], in_2[0]);
  nand g7 (n_534, n_185, in_2[0]);
  nand g8 (n_536, n_532, n_533, n_534);
  nor g9 (n_535, n_159, n_184);
  nand g10 (n_538, n_159, n_184);
  nor g11 (n_545, n_158, n_183);
  nand g12 (n_540, n_158, n_183);
  nor g13 (n_541, n_157, n_182);
  nand g14 (n_542, n_157, n_182);
  nor g15 (n_551, n_156, n_181);
  nand g16 (n_546, n_156, n_181);
  nor g17 (n_547, n_155, n_180);
  nand g18 (n_548, n_155, n_180);
  nor g19 (n_557, n_154, n_179);
  nand g20 (n_552, n_154, n_179);
  nor g21 (n_553, n_153, n_178);
  nand g22 (n_554, n_153, n_178);
  nor g23 (n_563, n_152, n_177);
  nand g24 (n_558, n_152, n_177);
  nor g25 (n_559, n_151, n_176);
  nand g26 (n_560, n_151, n_176);
  nor g27 (n_569, n_150, n_175);
  nand g28 (n_564, n_150, n_175);
  nor g29 (n_565, n_149, n_174);
  nand g30 (n_566, n_149, n_174);
  nor g31 (n_575, n_148, n_173);
  nand g32 (n_570, n_148, n_173);
  nor g33 (n_571, n_147, n_172);
  nand g34 (n_572, n_147, n_172);
  nor g35 (n_581, n_146, n_171);
  nand g36 (n_576, n_146, n_171);
  nor g37 (n_577, n_145, n_170);
  nand g38 (n_578, n_145, n_170);
  nor g39 (n_587, n_144, n_169);
  nand g40 (n_582, n_144, n_169);
  nor g41 (n_583, n_143, n_168);
  nand g42 (n_584, n_143, n_168);
  nor g43 (n_593, n_142, n_167);
  nand g44 (n_588, n_142, n_167);
  nor g45 (n_589, n_141, n_166);
  nand g46 (n_590, n_141, n_166);
  nor g47 (n_599, n_140, n_165);
  nand g48 (n_594, n_140, n_165);
  nor g49 (n_595, n_139, n_164);
  nand g50 (n_596, n_139, n_164);
  nor g51 (n_605, n_138, n_163);
  nand g52 (n_600, n_138, n_163);
  nor g53 (n_601, n_137, n_162);
  nand g54 (n_602, n_137, n_162);
  nand g59 (n_606, n_538, n_539);
  nor g60 (n_543, n_540, n_541);
  nor g63 (n_609, n_545, n_541);
  nor g64 (n_549, n_546, n_547);
  nor g67 (n_614, n_551, n_547);
  nor g68 (n_555, n_552, n_553);
  nor g71 (n_616, n_557, n_553);
  nor g460 (n_561, n_558, n_559);
  nor g463 (n_624, n_563, n_559);
  nor g464 (n_567, n_564, n_565);
  nor g467 (n_626, n_569, n_565);
  nor g468 (n_573, n_570, n_571);
  nor g471 (n_634, n_575, n_571);
  nor g472 (n_579, n_576, n_577);
  nor g475 (n_636, n_581, n_577);
  nor g476 (n_585, n_582, n_583);
  nor g479 (n_644, n_587, n_583);
  nor g480 (n_591, n_588, n_589);
  nor g483 (n_646, n_593, n_589);
  nor g484 (n_597, n_594, n_595);
  nor g487 (n_654, n_599, n_595);
  nor g488 (n_603, n_600, n_601);
  nor g491 (n_656, n_605, n_601);
  nand g494 (n_753, n_540, n_608);
  nand g495 (n_160, n_609, n_606);
  nand g496 (n_661, n_610, n_160);
  nor g497 (n_612, n_557, n_611);
  nand g506 (n_669, n_614, n_616);
  nor g507 (n_622, n_569, n_621);
  nand g516 (n_676, n_624, n_626);
  nor g517 (n_632, n_581, n_631);
  nand g526 (n_684, n_634, n_636);
  nor g527 (n_642, n_593, n_641);
  nand g536 (n_691, n_644, n_646);
  nor g537 (n_652, n_605, n_651);
  nand g546 (n_699, n_654, n_656);
  nand g549 (n_757, n_546, n_663);
  nand g550 (n_664, n_614, n_661);
  nand g551 (n_759, n_611, n_664);
  nand g554 (n_762, n_667, n_668);
  nand g557 (n_703, n_671, n_672);
  nor g558 (n_674, n_575, n_673);
  nor g561 (n_713, n_575, n_676);
  nor g567 (n_682, n_680, n_673);
  nor g570 (n_719, n_676, n_680);
  nor g571 (n_686, n_684, n_673);
  nor g574 (n_722, n_676, n_684);
  nor g575 (n_689, n_599, n_688);
  nor g578 (n_740, n_599, n_691);
  nor g584 (n_697, n_695, n_688);
  nor g587 (n_746, n_691, n_695);
  nor g588 (n_701, n_699, n_688);
  nor g591 (n_728, n_691, n_699);
  nand g594 (n_766, n_558, n_705);
  nand g595 (n_706, n_624, n_703);
  nand g596 (n_768, n_621, n_706);
  nand g599 (n_771, n_709, n_710);
  nand g602 (n_774, n_673, n_712);
  nand g603 (n_715, n_713, n_703);
  nand g604 (n_777, n_714, n_715);
  nand g605 (n_718, n_716, n_703);
  nand g606 (n_779, n_717, n_718);
  nand g607 (n_721, n_719, n_703);
  nand g608 (n_782, n_720, n_721);
  nand g609 (n_724, n_722, n_703);
  nand g610 (n_730, n_723, n_724);
  nand g614 (n_786, n_582, n_732);
  nand g615 (n_733, n_644, n_730);
  nand g616 (n_788, n_641, n_733);
  nand g619 (n_791, n_736, n_737);
  nand g622 (n_794, n_688, n_739);
  nand g623 (n_742, n_740, n_730);
  nand g624 (n_797, n_741, n_742);
  nand g625 (n_745, n_743, n_730);
  nand g626 (n_799, n_744, n_745);
  nand g627 (n_748, n_746, n_730);
  nand g628 (n_802, n_747, n_748);
  nand g629 (n_749, n_728, n_730);
  nand g630 (n_804, n_726, n_749);
  xnor g632 (out_0[1], n_536, n_750);
  xnor g634 (out_0[2], n_606, n_751);
  xnor g637 (out_0[3], n_753, n_754);
  xnor g639 (out_0[4], n_661, n_755);
  xnor g642 (out_0[5], n_757, n_758);
  xnor g644 (out_0[6], n_759, n_760);
  xnor g647 (out_0[7], n_762, n_763);
  xnor g649 (out_0[8], n_703, n_764);
  xnor g652 (out_0[9], n_766, n_767);
  xnor g654 (out_0[10], n_768, n_769);
  xnor g657 (out_0[11], n_771, n_772);
  xnor g660 (out_0[12], n_774, n_775);
  xnor g663 (out_0[13], n_777, n_778);
  xnor g665 (out_0[14], n_779, n_780);
  xnor g668 (out_0[15], n_782, n_783);
  xnor g670 (out_0[16], n_730, n_784);
  xnor g673 (out_0[17], n_786, n_787);
  xnor g675 (out_0[18], n_788, n_789);
  xnor g678 (out_0[19], n_791, n_792);
  xnor g681 (out_0[20], n_794, n_795);
  xnor g684 (out_0[21], n_797, n_798);
  xnor g686 (out_0[22], n_799, n_800);
  xnor g689 (out_0[23], n_802, n_803);
  xor g692 (out_0[0], in_2[0], n_806);
  xor g693 (n_268, in_0[21], in_1[21]);
  nor g694 (n_137, in_0[21], in_1[21]);
  xor g695 (n_514, in_3[21], in_4[21]);
  or g696 (n_515, in_3[21], in_4[21]);
  or g697 (n_516, in_2[21], in_4[21]);
  or g698 (n_517, in_2[21], in_3[21]);
  xnor g699 (n_270, n_514, in_2[21]);
  xnor g703 (n_271, n_269, n_268);
  or g704 (n_277, n_268, wc, n_269);
  not gc (wc, n_520);
  xnor g705 (n_526, n_275, n_137);
  or g706 (n_527, n_137, wc0);
  not gc0 (wc0, n_275);
  or g707 (n_528, wc1, n_137);
  not gc1 (wc1, n_277);
  or g708 (n_539, n_535, wc2);
  not gc2 (wc2, n_536);
  or g709 (n_750, wc3, n_535);
  not gc3 (wc3, n_538);
  and g710 (n_610, wc4, n_542);
  not gc4 (wc4, n_543);
  or g711 (n_751, wc5, n_545);
  not gc5 (wc5, n_540);
  or g712 (n_754, wc6, n_541);
  not gc6 (wc6, n_542);
  and g713 (n_611, wc7, n_548);
  not gc7 (wc7, n_549);
  or g714 (n_608, wc8, n_545);
  not gc8 (wc8, n_606);
  or g715 (n_755, wc9, n_551);
  not gc9 (wc9, n_546);
  or g716 (n_758, wc10, n_547);
  not gc10 (wc10, n_548);
  and g717 (n_618, wc11, n_554);
  not gc11 (wc11, n_555);
  and g718 (n_621, wc12, n_560);
  not gc12 (wc12, n_561);
  and g719 (n_628, wc13, n_566);
  not gc13 (wc13, n_567);
  and g720 (n_631, wc14, n_572);
  not gc14 (wc14, n_573);
  and g721 (n_638, wc15, n_578);
  not gc15 (wc15, n_579);
  and g722 (n_641, wc16, n_584);
  not gc16 (wc16, n_585);
  and g723 (n_648, wc17, n_590);
  not gc17 (wc17, n_591);
  and g724 (n_651, wc18, n_596);
  not gc18 (wc18, n_597);
  and g725 (n_658, wc19, n_602);
  not gc19 (wc19, n_603);
  or g726 (n_665, wc20, n_557);
  not gc20 (wc20, n_614);
  or g727 (n_707, wc21, n_569);
  not gc21 (wc21, n_624);
  or g728 (n_680, wc22, n_581);
  not gc22 (wc22, n_634);
  or g729 (n_734, wc23, n_593);
  not gc23 (wc23, n_644);
  or g730 (n_695, wc24, n_605);
  not gc24 (wc24, n_654);
  or g731 (n_760, wc25, n_557);
  not gc25 (wc25, n_552);
  or g732 (n_763, wc26, n_553);
  not gc26 (wc26, n_554);
  or g733 (n_764, wc27, n_563);
  not gc27 (wc27, n_558);
  or g734 (n_767, wc28, n_559);
  not gc28 (wc28, n_560);
  or g735 (n_769, wc29, n_569);
  not gc29 (wc29, n_564);
  or g736 (n_772, wc30, n_565);
  not gc30 (wc30, n_566);
  or g737 (n_775, wc31, n_575);
  not gc31 (wc31, n_570);
  or g738 (n_778, wc32, n_571);
  not gc32 (wc32, n_572);
  or g739 (n_780, wc33, n_581);
  not gc33 (wc33, n_576);
  or g740 (n_783, wc34, n_577);
  not gc34 (wc34, n_578);
  or g741 (n_784, wc35, n_587);
  not gc35 (wc35, n_582);
  or g742 (n_787, wc36, n_583);
  not gc36 (wc36, n_584);
  or g743 (n_789, wc37, n_593);
  not gc37 (wc37, n_588);
  or g744 (n_792, wc38, n_589);
  not gc38 (wc38, n_590);
  or g745 (n_795, wc39, n_599);
  not gc39 (wc39, n_594);
  or g746 (n_798, wc40, n_595);
  not gc40 (wc40, n_596);
  or g747 (n_800, wc41, n_605);
  not gc41 (wc41, n_600);
  or g748 (n_803, wc42, n_601);
  not gc42 (wc42, n_602);
  and g749 (n_667, wc43, n_552);
  not gc43 (wc43, n_612);
  and g750 (n_619, wc44, n_616);
  not gc44 (wc44, n_611);
  and g751 (n_629, wc45, n_626);
  not gc45 (wc45, n_621);
  and g752 (n_639, wc46, n_636);
  not gc46 (wc46, n_631);
  and g753 (n_649, wc47, n_646);
  not gc47 (wc47, n_641);
  and g754 (n_659, wc48, n_656);
  not gc48 (wc48, n_651);
  or g755 (n_663, wc49, n_551);
  not gc49 (wc49, n_661);
  and g756 (n_716, wc50, n_634);
  not gc50 (wc50, n_676);
  and g757 (n_743, wc51, n_654);
  not gc51 (wc51, n_691);
  and g758 (n_671, wc52, n_618);
  not gc52 (wc52, n_619);
  and g759 (n_709, wc53, n_564);
  not gc53 (wc53, n_622);
  and g760 (n_673, wc54, n_628);
  not gc54 (wc54, n_629);
  and g761 (n_681, wc55, n_576);
  not gc55 (wc55, n_632);
  and g762 (n_685, wc56, n_638);
  not gc56 (wc56, n_639);
  and g763 (n_736, wc57, n_588);
  not gc57 (wc57, n_642);
  and g764 (n_688, wc58, n_648);
  not gc58 (wc58, n_649);
  and g765 (n_696, wc59, n_600);
  not gc59 (wc59, n_652);
  and g766 (n_700, wc60, n_658);
  not gc60 (wc60, n_659);
  or g767 (n_668, n_665, wc61);
  not gc61 (wc61, n_661);
  or g768 (n_672, n_669, wc62);
  not gc62 (wc62, n_661);
  and g769 (n_678, wc63, n_634);
  not gc63 (wc63, n_673);
  and g770 (n_693, wc64, n_654);
  not gc64 (wc64, n_688);
  and g771 (n_714, wc65, n_570);
  not gc65 (wc65, n_674);
  and g772 (n_717, wc66, n_631);
  not gc66 (wc66, n_678);
  and g773 (n_720, n_681, wc67);
  not gc67 (wc67, n_682);
  and g774 (n_723, n_685, wc68);
  not gc68 (wc68, n_686);
  and g775 (n_741, wc69, n_594);
  not gc69 (wc69, n_689);
  and g776 (n_744, wc70, n_651);
  not gc70 (wc70, n_693);
  and g777 (n_747, n_696, wc71);
  not gc71 (wc71, n_697);
  and g778 (n_726, n_700, wc72);
  not gc72 (wc72, n_701);
  or g779 (n_705, wc73, n_563);
  not gc73 (wc73, n_703);
  or g780 (n_710, n_707, wc74);
  not gc74 (wc74, n_703);
  or g781 (n_712, wc75, n_676);
  not gc75 (wc75, n_703);
  or g782 (n_732, wc76, n_587);
  not gc76 (wc76, n_730);
  or g783 (n_737, n_734, wc77);
  not gc77 (wc77, n_730);
  or g784 (n_739, wc78, n_691);
  not gc78 (wc78, n_730);
  not g785 (out_0[24], n_804);
endmodule

module csa_tree_add_694_38_group_6811_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [21:0] in_0, in_1, in_2, in_3, in_4;
  output [24:0] out_0;
  wire [21:0] in_0, in_1, in_2, in_3, in_4;
  wire [24:0] out_0;
  csa_tree_add_694_38_group_6811_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_767_44_group_6809_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_280, n_281, n_282, n_283, n_284, n_287;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_544, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_556, n_557;
  wire n_558, n_559, n_560, n_562, n_563, n_564, n_565, n_566;
  wire n_567, n_569, n_570, n_571, n_572, n_573, n_575, n_576;
  wire n_577, n_578, n_579, n_581, n_582, n_583, n_584, n_585;
  wire n_587, n_588, n_589, n_590, n_591, n_593, n_594, n_595;
  wire n_596, n_597, n_599, n_600, n_601, n_602, n_603, n_605;
  wire n_606, n_607, n_608, n_609, n_611, n_612, n_613, n_614;
  wire n_615, n_617, n_618, n_619, n_620, n_621, n_623, n_624;
  wire n_625, n_626, n_627, n_629, n_630, n_633, n_634, n_636;
  wire n_637, n_638, n_639, n_640, n_642, n_644, n_646, n_647;
  wire n_649, n_650, n_652, n_654, n_656, n_657, n_659, n_660;
  wire n_662, n_664, n_666, n_667, n_669, n_670, n_672, n_674;
  wire n_676, n_677, n_679, n_680, n_682, n_684, n_686, n_687;
  wire n_689, n_691, n_692, n_693, n_695, n_696, n_697, n_699;
  wire n_700, n_701, n_702, n_704, n_706, n_708, n_709, n_710;
  wire n_712, n_713, n_714, n_716, n_717, n_719, n_721, n_723;
  wire n_724, n_725, n_727, n_728, n_729, n_731, n_733, n_734;
  wire n_735, n_737, n_738, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_756, n_758, n_760, n_761, n_762, n_764;
  wire n_765, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_780, n_781, n_782;
  wire n_783, n_785, n_786, n_787, n_789, n_790, n_791, n_792;
  wire n_794, n_795, n_796, n_798, n_799, n_800, n_801, n_803;
  wire n_804, n_806, n_807, n_809, n_810, n_811, n_812, n_814;
  wire n_815, n_816, n_818, n_819, n_820, n_821, n_823, n_824;
  wire n_826, n_827, n_829, n_830, n_831, n_832, n_834, n_835;
  wire n_836, n_837, n_839, n_841;
  xor g75 (n_290, in_0[0], in_4[0]);
  xor g76 (n_193, n_290, in_3[0]);
  nand g77 (n_291, in_0[0], in_4[0]);
  nand g78 (n_292, in_3[0], in_4[0]);
  nand g79 (n_293, in_0[0], in_3[0]);
  nand g6 (n_195, n_291, n_292, n_293);
  xor g80 (n_294, in_0[1], in_1[1]);
  xor g81 (n_166, n_294, in_4[1]);
  nand g82 (n_295, in_0[1], in_1[1]);
  nand g83 (n_296, in_4[1], in_1[1]);
  nand g84 (n_297, in_0[1], in_4[1]);
  nand g85 (n_197, n_295, n_296, n_297);
  xor g86 (n_298, in_3[1], in_2[1]);
  xor g87 (n_192, n_298, n_195);
  nand g88 (n_299, in_3[1], in_2[1]);
  nand g89 (n_300, n_195, in_2[1]);
  nand g90 (n_301, in_3[1], n_195);
  nand g91 (n_165, n_299, n_300, n_301);
  xor g92 (n_196, in_0[2], in_1[2]);
  and g93 (n_199, in_0[2], in_1[2]);
  xor g94 (n_302, in_3[2], in_4[2]);
  xor g95 (n_198, n_302, in_2[2]);
  nand g96 (n_303, in_3[2], in_4[2]);
  nand g97 (n_304, in_2[2], in_4[2]);
  nand g98 (n_305, in_3[2], in_2[2]);
  nand g99 (n_200, n_303, n_304, n_305);
  xor g100 (n_306, n_196, n_197);
  xor g101 (n_191, n_306, n_198);
  nand g102 (n_307, n_196, n_197);
  nand g103 (n_308, n_198, n_197);
  nand g104 (n_309, n_196, n_198);
  nand g105 (n_164, n_307, n_308, n_309);
  xor g106 (n_310, in_0[3], in_1[3]);
  xor g107 (n_201, n_310, in_3[3]);
  nand g108 (n_311, in_0[3], in_1[3]);
  nand g109 (n_312, in_3[3], in_1[3]);
  nand g110 (n_313, in_0[3], in_3[3]);
  nand g111 (n_203, n_311, n_312, n_313);
  xor g112 (n_314, in_4[3], in_2[3]);
  xor g113 (n_202, n_314, n_199);
  nand g114 (n_315, in_4[3], in_2[3]);
  nand g115 (n_316, n_199, in_2[3]);
  nand g116 (n_317, in_4[3], n_199);
  nand g117 (n_205, n_315, n_316, n_317);
  xor g118 (n_318, n_200, n_201);
  xor g119 (n_190, n_318, n_202);
  nand g120 (n_319, n_200, n_201);
  nand g121 (n_320, n_202, n_201);
  nand g122 (n_321, n_200, n_202);
  nand g123 (n_163, n_319, n_320, n_321);
  xor g124 (n_322, in_0[4], in_1[4]);
  xor g125 (n_204, n_322, in_3[4]);
  nand g126 (n_323, in_0[4], in_1[4]);
  nand g127 (n_324, in_3[4], in_1[4]);
  nand g128 (n_325, in_0[4], in_3[4]);
  nand g129 (n_207, n_323, n_324, n_325);
  xor g130 (n_326, in_4[4], in_2[4]);
  xor g131 (n_206, n_326, n_203);
  nand g132 (n_327, in_4[4], in_2[4]);
  nand g133 (n_328, n_203, in_2[4]);
  nand g134 (n_329, in_4[4], n_203);
  nand g135 (n_210, n_327, n_328, n_329);
  xor g136 (n_330, n_204, n_205);
  xor g137 (n_189, n_330, n_206);
  nand g138 (n_331, n_204, n_205);
  nand g139 (n_332, n_206, n_205);
  nand g140 (n_333, n_204, n_206);
  nand g141 (n_162, n_331, n_332, n_333);
  xor g142 (n_334, in_0[5], in_1[5]);
  xor g143 (n_208, n_334, in_3[5]);
  nand g144 (n_335, in_0[5], in_1[5]);
  nand g145 (n_336, in_3[5], in_1[5]);
  nand g146 (n_337, in_0[5], in_3[5]);
  nand g147 (n_211, n_335, n_336, n_337);
  xor g148 (n_338, in_4[5], in_2[5]);
  xor g149 (n_209, n_338, n_207);
  nand g150 (n_339, in_4[5], in_2[5]);
  nand g151 (n_340, n_207, in_2[5]);
  nand g152 (n_341, in_4[5], n_207);
  nand g153 (n_214, n_339, n_340, n_341);
  xor g154 (n_342, n_208, n_209);
  xor g155 (n_188, n_342, n_210);
  nand g156 (n_343, n_208, n_209);
  nand g157 (n_344, n_210, n_209);
  nand g158 (n_345, n_208, n_210);
  nand g159 (n_161, n_343, n_344, n_345);
  xor g160 (n_346, in_0[6], in_1[6]);
  xor g161 (n_212, n_346, in_3[6]);
  nand g162 (n_347, in_0[6], in_1[6]);
  nand g163 (n_348, in_3[6], in_1[6]);
  nand g164 (n_349, in_0[6], in_3[6]);
  nand g165 (n_215, n_347, n_348, n_349);
  xor g166 (n_350, in_4[6], in_2[6]);
  xor g167 (n_213, n_350, n_211);
  nand g168 (n_351, in_4[6], in_2[6]);
  nand g169 (n_352, n_211, in_2[6]);
  nand g170 (n_353, in_4[6], n_211);
  nand g171 (n_218, n_351, n_352, n_353);
  xor g172 (n_354, n_212, n_213);
  xor g173 (n_187, n_354, n_214);
  nand g174 (n_355, n_212, n_213);
  nand g175 (n_356, n_214, n_213);
  nand g176 (n_357, n_212, n_214);
  nand g177 (n_160, n_355, n_356, n_357);
  xor g178 (n_358, in_0[7], in_1[7]);
  xor g179 (n_216, n_358, in_3[7]);
  nand g180 (n_359, in_0[7], in_1[7]);
  nand g181 (n_360, in_3[7], in_1[7]);
  nand g182 (n_361, in_0[7], in_3[7]);
  nand g183 (n_219, n_359, n_360, n_361);
  xor g184 (n_362, in_4[7], in_2[7]);
  xor g185 (n_217, n_362, n_215);
  nand g186 (n_363, in_4[7], in_2[7]);
  nand g187 (n_364, n_215, in_2[7]);
  nand g188 (n_365, in_4[7], n_215);
  nand g189 (n_222, n_363, n_364, n_365);
  xor g190 (n_366, n_216, n_217);
  xor g191 (n_186, n_366, n_218);
  nand g192 (n_367, n_216, n_217);
  nand g193 (n_368, n_218, n_217);
  nand g194 (n_369, n_216, n_218);
  nand g195 (n_159, n_367, n_368, n_369);
  xor g196 (n_370, in_0[8], in_1[8]);
  xor g197 (n_220, n_370, in_3[8]);
  nand g198 (n_371, in_0[8], in_1[8]);
  nand g199 (n_372, in_3[8], in_1[8]);
  nand g200 (n_373, in_0[8], in_3[8]);
  nand g201 (n_223, n_371, n_372, n_373);
  xor g202 (n_374, in_4[8], in_2[8]);
  xor g203 (n_221, n_374, n_219);
  nand g204 (n_375, in_4[8], in_2[8]);
  nand g205 (n_376, n_219, in_2[8]);
  nand g206 (n_377, in_4[8], n_219);
  nand g207 (n_226, n_375, n_376, n_377);
  xor g208 (n_378, n_220, n_221);
  xor g209 (n_185, n_378, n_222);
  nand g210 (n_379, n_220, n_221);
  nand g211 (n_380, n_222, n_221);
  nand g212 (n_381, n_220, n_222);
  nand g213 (n_158, n_379, n_380, n_381);
  xor g214 (n_382, in_0[9], in_1[9]);
  xor g215 (n_224, n_382, in_3[9]);
  nand g216 (n_383, in_0[9], in_1[9]);
  nand g217 (n_384, in_3[9], in_1[9]);
  nand g218 (n_385, in_0[9], in_3[9]);
  nand g219 (n_227, n_383, n_384, n_385);
  xor g220 (n_386, in_4[9], in_2[9]);
  xor g221 (n_225, n_386, n_223);
  nand g222 (n_387, in_4[9], in_2[9]);
  nand g223 (n_388, n_223, in_2[9]);
  nand g224 (n_389, in_4[9], n_223);
  nand g225 (n_230, n_387, n_388, n_389);
  xor g226 (n_390, n_224, n_225);
  xor g227 (n_184, n_390, n_226);
  nand g228 (n_391, n_224, n_225);
  nand g229 (n_392, n_226, n_225);
  nand g230 (n_393, n_224, n_226);
  nand g231 (n_157, n_391, n_392, n_393);
  xor g232 (n_394, in_0[10], in_1[10]);
  xor g233 (n_228, n_394, in_3[10]);
  nand g234 (n_395, in_0[10], in_1[10]);
  nand g235 (n_396, in_3[10], in_1[10]);
  nand g236 (n_397, in_0[10], in_3[10]);
  nand g237 (n_231, n_395, n_396, n_397);
  xor g238 (n_398, in_4[10], in_2[10]);
  xor g239 (n_229, n_398, n_227);
  nand g240 (n_399, in_4[10], in_2[10]);
  nand g241 (n_400, n_227, in_2[10]);
  nand g242 (n_401, in_4[10], n_227);
  nand g243 (n_234, n_399, n_400, n_401);
  xor g244 (n_402, n_228, n_229);
  xor g245 (n_183, n_402, n_230);
  nand g246 (n_403, n_228, n_229);
  nand g247 (n_404, n_230, n_229);
  nand g248 (n_405, n_228, n_230);
  nand g249 (n_156, n_403, n_404, n_405);
  xor g250 (n_406, in_0[11], in_1[11]);
  xor g251 (n_232, n_406, in_3[11]);
  nand g252 (n_407, in_0[11], in_1[11]);
  nand g253 (n_408, in_3[11], in_1[11]);
  nand g254 (n_409, in_0[11], in_3[11]);
  nand g255 (n_235, n_407, n_408, n_409);
  xor g256 (n_410, in_4[11], in_2[11]);
  xor g257 (n_233, n_410, n_231);
  nand g258 (n_411, in_4[11], in_2[11]);
  nand g259 (n_412, n_231, in_2[11]);
  nand g260 (n_413, in_4[11], n_231);
  nand g261 (n_238, n_411, n_412, n_413);
  xor g262 (n_414, n_232, n_233);
  xor g263 (n_182, n_414, n_234);
  nand g264 (n_415, n_232, n_233);
  nand g265 (n_416, n_234, n_233);
  nand g266 (n_417, n_232, n_234);
  nand g267 (n_155, n_415, n_416, n_417);
  xor g268 (n_418, in_0[12], in_1[12]);
  xor g269 (n_236, n_418, in_3[12]);
  nand g270 (n_419, in_0[12], in_1[12]);
  nand g271 (n_420, in_3[12], in_1[12]);
  nand g272 (n_421, in_0[12], in_3[12]);
  nand g273 (n_239, n_419, n_420, n_421);
  xor g274 (n_422, in_4[12], in_2[12]);
  xor g275 (n_237, n_422, n_235);
  nand g276 (n_423, in_4[12], in_2[12]);
  nand g277 (n_424, n_235, in_2[12]);
  nand g278 (n_425, in_4[12], n_235);
  nand g279 (n_242, n_423, n_424, n_425);
  xor g280 (n_426, n_236, n_237);
  xor g281 (n_181, n_426, n_238);
  nand g282 (n_427, n_236, n_237);
  nand g283 (n_428, n_238, n_237);
  nand g284 (n_429, n_236, n_238);
  nand g285 (n_154, n_427, n_428, n_429);
  xor g286 (n_430, in_0[13], in_1[13]);
  xor g287 (n_240, n_430, in_3[13]);
  nand g288 (n_431, in_0[13], in_1[13]);
  nand g289 (n_432, in_3[13], in_1[13]);
  nand g290 (n_433, in_0[13], in_3[13]);
  nand g291 (n_243, n_431, n_432, n_433);
  xor g292 (n_434, in_4[13], in_2[13]);
  xor g293 (n_241, n_434, n_239);
  nand g294 (n_435, in_4[13], in_2[13]);
  nand g295 (n_436, n_239, in_2[13]);
  nand g296 (n_437, in_4[13], n_239);
  nand g297 (n_246, n_435, n_436, n_437);
  xor g298 (n_438, n_240, n_241);
  xor g299 (n_180, n_438, n_242);
  nand g300 (n_439, n_240, n_241);
  nand g301 (n_440, n_242, n_241);
  nand g302 (n_441, n_240, n_242);
  nand g303 (n_153, n_439, n_440, n_441);
  xor g304 (n_442, in_0[14], in_1[14]);
  xor g305 (n_244, n_442, in_3[14]);
  nand g306 (n_443, in_0[14], in_1[14]);
  nand g307 (n_444, in_3[14], in_1[14]);
  nand g308 (n_445, in_0[14], in_3[14]);
  nand g309 (n_247, n_443, n_444, n_445);
  xor g310 (n_446, in_4[14], in_2[14]);
  xor g311 (n_245, n_446, n_243);
  nand g312 (n_447, in_4[14], in_2[14]);
  nand g313 (n_448, n_243, in_2[14]);
  nand g314 (n_449, in_4[14], n_243);
  nand g315 (n_250, n_447, n_448, n_449);
  xor g316 (n_450, n_244, n_245);
  xor g317 (n_179, n_450, n_246);
  nand g318 (n_451, n_244, n_245);
  nand g319 (n_452, n_246, n_245);
  nand g320 (n_453, n_244, n_246);
  nand g321 (n_152, n_451, n_452, n_453);
  xor g322 (n_454, in_0[15], in_1[15]);
  xor g323 (n_248, n_454, in_3[15]);
  nand g324 (n_455, in_0[15], in_1[15]);
  nand g325 (n_456, in_3[15], in_1[15]);
  nand g326 (n_457, in_0[15], in_3[15]);
  nand g327 (n_251, n_455, n_456, n_457);
  xor g328 (n_458, in_4[15], in_2[15]);
  xor g329 (n_249, n_458, n_247);
  nand g330 (n_459, in_4[15], in_2[15]);
  nand g331 (n_460, n_247, in_2[15]);
  nand g332 (n_461, in_4[15], n_247);
  nand g333 (n_254, n_459, n_460, n_461);
  xor g334 (n_462, n_248, n_249);
  xor g335 (n_178, n_462, n_250);
  nand g336 (n_463, n_248, n_249);
  nand g337 (n_464, n_250, n_249);
  nand g338 (n_465, n_248, n_250);
  nand g339 (n_151, n_463, n_464, n_465);
  xor g340 (n_466, in_0[16], in_1[16]);
  xor g341 (n_252, n_466, in_3[16]);
  nand g342 (n_467, in_0[16], in_1[16]);
  nand g343 (n_468, in_3[16], in_1[16]);
  nand g344 (n_469, in_0[16], in_3[16]);
  nand g345 (n_255, n_467, n_468, n_469);
  xor g346 (n_470, in_4[16], in_2[16]);
  xor g347 (n_253, n_470, n_251);
  nand g348 (n_471, in_4[16], in_2[16]);
  nand g349 (n_472, n_251, in_2[16]);
  nand g350 (n_473, in_4[16], n_251);
  nand g351 (n_258, n_471, n_472, n_473);
  xor g352 (n_474, n_252, n_253);
  xor g353 (n_177, n_474, n_254);
  nand g354 (n_475, n_252, n_253);
  nand g355 (n_476, n_254, n_253);
  nand g356 (n_477, n_252, n_254);
  nand g357 (n_150, n_475, n_476, n_477);
  xor g358 (n_478, in_0[17], in_1[17]);
  xor g359 (n_256, n_478, in_3[17]);
  nand g360 (n_479, in_0[17], in_1[17]);
  nand g361 (n_480, in_3[17], in_1[17]);
  nand g362 (n_481, in_0[17], in_3[17]);
  nand g363 (n_259, n_479, n_480, n_481);
  xor g364 (n_482, in_4[17], in_2[17]);
  xor g365 (n_257, n_482, n_255);
  nand g366 (n_483, in_4[17], in_2[17]);
  nand g367 (n_484, n_255, in_2[17]);
  nand g368 (n_485, in_4[17], n_255);
  nand g369 (n_262, n_483, n_484, n_485);
  xor g370 (n_486, n_256, n_257);
  xor g371 (n_176, n_486, n_258);
  nand g372 (n_487, n_256, n_257);
  nand g373 (n_488, n_258, n_257);
  nand g374 (n_489, n_256, n_258);
  nand g375 (n_149, n_487, n_488, n_489);
  xor g376 (n_490, in_0[18], in_1[18]);
  xor g377 (n_260, n_490, in_3[18]);
  nand g378 (n_491, in_0[18], in_1[18]);
  nand g379 (n_492, in_3[18], in_1[18]);
  nand g380 (n_493, in_0[18], in_3[18]);
  nand g381 (n_263, n_491, n_492, n_493);
  xor g382 (n_494, in_4[18], in_2[18]);
  xor g383 (n_261, n_494, n_259);
  nand g384 (n_495, in_4[18], in_2[18]);
  nand g385 (n_496, n_259, in_2[18]);
  nand g386 (n_497, in_4[18], n_259);
  nand g387 (n_266, n_495, n_496, n_497);
  xor g388 (n_498, n_260, n_261);
  xor g389 (n_175, n_498, n_262);
  nand g390 (n_499, n_260, n_261);
  nand g391 (n_500, n_262, n_261);
  nand g392 (n_501, n_260, n_262);
  nand g393 (n_148, n_499, n_500, n_501);
  xor g394 (n_502, in_0[19], in_1[19]);
  xor g395 (n_264, n_502, in_3[19]);
  nand g396 (n_503, in_0[19], in_1[19]);
  nand g397 (n_504, in_3[19], in_1[19]);
  nand g398 (n_505, in_0[19], in_3[19]);
  nand g399 (n_267, n_503, n_504, n_505);
  xor g400 (n_506, in_4[19], in_2[19]);
  xor g401 (n_265, n_506, n_263);
  nand g402 (n_507, in_4[19], in_2[19]);
  nand g403 (n_508, n_263, in_2[19]);
  nand g404 (n_509, in_4[19], n_263);
  nand g405 (n_270, n_507, n_508, n_509);
  xor g406 (n_510, n_264, n_265);
  xor g407 (n_174, n_510, n_266);
  nand g408 (n_511, n_264, n_265);
  nand g409 (n_512, n_266, n_265);
  nand g410 (n_513, n_264, n_266);
  nand g411 (n_147, n_511, n_512, n_513);
  xor g412 (n_514, in_0[20], in_1[20]);
  xor g413 (n_268, n_514, in_3[20]);
  nand g414 (n_515, in_0[20], in_1[20]);
  nand g415 (n_516, in_3[20], in_1[20]);
  nand g416 (n_517, in_0[20], in_3[20]);
  nand g417 (n_271, n_515, n_516, n_517);
  xor g418 (n_518, in_4[20], in_2[20]);
  xor g419 (n_269, n_518, n_267);
  nand g420 (n_519, in_4[20], in_2[20]);
  nand g421 (n_520, n_267, in_2[20]);
  nand g422 (n_521, in_4[20], n_267);
  nand g423 (n_274, n_519, n_520, n_521);
  xor g424 (n_522, n_268, n_269);
  xor g425 (n_173, n_522, n_270);
  nand g426 (n_523, n_268, n_269);
  nand g427 (n_524, n_270, n_269);
  nand g428 (n_525, n_268, n_270);
  nand g429 (n_146, n_523, n_524, n_525);
  xor g430 (n_526, in_0[21], in_1[21]);
  xor g431 (n_272, n_526, in_3[21]);
  nand g432 (n_527, in_0[21], in_1[21]);
  nand g433 (n_528, in_3[21], in_1[21]);
  nand g434 (n_529, in_0[21], in_3[21]);
  nand g435 (n_281, n_527, n_528, n_529);
  xor g436 (n_530, in_4[21], in_2[21]);
  xor g437 (n_273, n_530, n_271);
  nand g438 (n_531, in_4[21], in_2[21]);
  nand g439 (n_532, n_271, in_2[21]);
  nand g440 (n_533, in_4[21], n_271);
  nand g441 (n_284, n_531, n_532, n_533);
  xor g442 (n_534, n_272, n_273);
  xor g443 (n_172, n_534, n_274);
  nand g444 (n_535, n_272, n_273);
  nand g445 (n_536, n_274, n_273);
  nand g446 (n_537, n_272, n_274);
  nand g447 (n_145, n_535, n_536, n_537);
  nand g455 (n_287, n_539, n_540, n_541);
  nand g459 (n_544, n_281, n_280);
  xor g462 (n_546, n_282, n_283);
  xor g463 (n_171, n_546, n_284);
  nand g464 (n_547, n_282, n_283);
  nand g465 (n_548, n_284, n_283);
  nand g466 (n_549, n_282, n_284);
  nand g467 (n_144, n_547, n_548, n_549);
  xor g471 (n_170, n_550, n_289);
  nand g474 (n_553, n_287, n_289);
  nand g475 (n_169, n_551, n_552, n_553);
  xor g478 (n_841, in_1[0], n_193);
  nand g479 (n_556, in_1[0], n_193);
  nand g480 (n_557, in_1[0], in_2[0]);
  nand g7 (n_558, n_193, in_2[0]);
  nand g8 (n_560, n_556, n_557, n_558);
  nor g9 (n_559, n_166, n_192);
  nand g10 (n_562, n_166, n_192);
  nor g11 (n_569, n_165, n_191);
  nand g12 (n_564, n_165, n_191);
  nor g13 (n_565, n_164, n_190);
  nand g14 (n_566, n_164, n_190);
  nor g15 (n_575, n_163, n_189);
  nand g16 (n_570, n_163, n_189);
  nor g17 (n_571, n_162, n_188);
  nand g18 (n_572, n_162, n_188);
  nor g19 (n_581, n_161, n_187);
  nand g20 (n_576, n_161, n_187);
  nor g21 (n_577, n_160, n_186);
  nand g22 (n_578, n_160, n_186);
  nor g23 (n_587, n_159, n_185);
  nand g24 (n_582, n_159, n_185);
  nor g25 (n_583, n_158, n_184);
  nand g26 (n_584, n_158, n_184);
  nor g27 (n_593, n_157, n_183);
  nand g28 (n_588, n_157, n_183);
  nor g29 (n_589, n_156, n_182);
  nand g30 (n_590, n_156, n_182);
  nor g31 (n_599, n_155, n_181);
  nand g32 (n_594, n_155, n_181);
  nor g33 (n_595, n_154, n_180);
  nand g34 (n_596, n_154, n_180);
  nor g35 (n_605, n_153, n_179);
  nand g36 (n_600, n_153, n_179);
  nor g37 (n_601, n_152, n_178);
  nand g38 (n_602, n_152, n_178);
  nor g39 (n_611, n_151, n_177);
  nand g40 (n_606, n_151, n_177);
  nor g41 (n_607, n_150, n_176);
  nand g42 (n_608, n_150, n_176);
  nor g43 (n_617, n_149, n_175);
  nand g44 (n_612, n_149, n_175);
  nor g45 (n_613, n_148, n_174);
  nand g46 (n_614, n_148, n_174);
  nor g47 (n_623, n_147, n_173);
  nand g48 (n_618, n_147, n_173);
  nor g49 (n_619, n_146, n_172);
  nand g50 (n_620, n_146, n_172);
  nor g51 (n_629, n_145, n_171);
  nand g52 (n_624, n_145, n_171);
  nor g53 (n_625, n_144, n_170);
  nand g54 (n_626, n_144, n_170);
  nor g55 (n_633, n_143, n_169);
  nand g56 (n_630, n_143, n_169);
  nand g61 (n_634, n_562, n_563);
  nor g62 (n_567, n_564, n_565);
  nor g65 (n_167, n_569, n_565);
  nor g66 (n_573, n_570, n_571);
  nor g69 (n_642, n_575, n_571);
  nor g70 (n_579, n_576, n_577);
  nor g73 (n_644, n_581, n_577);
  nor g74 (n_585, n_582, n_583);
  nor g483 (n_652, n_587, n_583);
  nor g484 (n_591, n_588, n_589);
  nor g487 (n_654, n_593, n_589);
  nor g488 (n_597, n_594, n_595);
  nor g491 (n_662, n_599, n_595);
  nor g492 (n_603, n_600, n_601);
  nor g495 (n_664, n_605, n_601);
  nor g496 (n_609, n_606, n_607);
  nor g499 (n_672, n_611, n_607);
  nor g500 (n_615, n_612, n_613);
  nor g503 (n_674, n_617, n_613);
  nor g504 (n_621, n_618, n_619);
  nor g507 (n_682, n_623, n_619);
  nor g508 (n_627, n_624, n_625);
  nor g511 (n_684, n_629, n_625);
  nand g514 (n_785, n_564, n_636);
  nand g515 (n_638, n_167, n_634);
  nand g516 (n_689, n_637, n_638);
  nor g517 (n_640, n_581, n_639);
  nand g526 (n_697, n_642, n_644);
  nor g527 (n_650, n_593, n_649);
  nand g536 (n_704, n_652, n_654);
  nor g537 (n_660, n_605, n_659);
  nand g546 (n_712, n_662, n_664);
  nor g547 (n_670, n_617, n_669);
  nand g556 (n_719, n_672, n_674);
  nor g557 (n_680, n_629, n_679);
  nand g566 (n_727, n_682, n_684);
  nand g569 (n_789, n_570, n_691);
  nand g570 (n_692, n_642, n_689);
  nand g571 (n_791, n_639, n_692);
  nand g574 (n_794, n_695, n_696);
  nand g577 (n_731, n_699, n_700);
  nor g578 (n_702, n_599, n_701);
  nor g581 (n_741, n_599, n_704);
  nor g587 (n_710, n_708, n_701);
  nor g590 (n_747, n_704, n_708);
  nor g591 (n_714, n_712, n_701);
  nor g594 (n_750, n_704, n_712);
  nor g595 (n_717, n_623, n_716);
  nor g598 (n_768, n_623, n_719);
  nor g604 (n_725, n_723, n_716);
  nor g607 (n_774, n_719, n_723);
  nor g608 (n_729, n_727, n_716);
  nor g611 (n_756, n_719, n_727);
  nand g614 (n_798, n_582, n_733);
  nand g615 (n_734, n_652, n_731);
  nand g616 (n_800, n_649, n_734);
  nand g619 (n_803, n_737, n_738);
  nand g622 (n_806, n_701, n_740);
  nand g623 (n_743, n_741, n_731);
  nand g624 (n_809, n_742, n_743);
  nand g625 (n_746, n_744, n_731);
  nand g626 (n_811, n_745, n_746);
  nand g627 (n_749, n_747, n_731);
  nand g628 (n_814, n_748, n_749);
  nand g629 (n_752, n_750, n_731);
  nand g630 (n_758, n_751, n_752);
  nor g631 (n_754, n_633, n_753);
  nand g638 (n_818, n_606, n_760);
  nand g639 (n_761, n_672, n_758);
  nand g640 (n_820, n_669, n_761);
  nand g643 (n_823, n_764, n_765);
  nand g646 (n_826, n_716, n_767);
  nand g647 (n_770, n_768, n_758);
  nand g648 (n_829, n_769, n_770);
  nand g649 (n_773, n_771, n_758);
  nand g650 (n_831, n_772, n_773);
  nand g651 (n_776, n_774, n_758);
  nand g652 (n_834, n_775, n_776);
  nand g653 (n_777, n_756, n_758);
  nand g654 (n_836, n_753, n_777);
  nand g657 (n_839, n_780, n_781);
  xnor g659 (out_0[1], n_560, n_782);
  xnor g661 (out_0[2], n_634, n_783);
  xnor g664 (out_0[3], n_785, n_786);
  xnor g666 (out_0[4], n_689, n_787);
  xnor g669 (out_0[5], n_789, n_790);
  xnor g671 (out_0[6], n_791, n_792);
  xnor g674 (out_0[7], n_794, n_795);
  xnor g676 (out_0[8], n_731, n_796);
  xnor g679 (out_0[9], n_798, n_799);
  xnor g681 (out_0[10], n_800, n_801);
  xnor g684 (out_0[11], n_803, n_804);
  xnor g687 (out_0[12], n_806, n_807);
  xnor g690 (out_0[13], n_809, n_810);
  xnor g692 (out_0[14], n_811, n_812);
  xnor g695 (out_0[15], n_814, n_815);
  xnor g697 (out_0[16], n_758, n_816);
  xnor g700 (out_0[17], n_818, n_819);
  xnor g702 (out_0[18], n_820, n_821);
  xnor g705 (out_0[19], n_823, n_824);
  xnor g708 (out_0[20], n_826, n_827);
  xnor g711 (out_0[21], n_829, n_830);
  xnor g713 (out_0[22], n_831, n_832);
  xnor g716 (out_0[23], n_834, n_835);
  xnor g718 (out_0[24], n_836, n_837);
  xor g722 (out_0[0], in_2[0], n_841);
  xor g723 (n_280, in_0[22], in_1[22]);
  nor g724 (n_143, in_0[22], in_1[22]);
  xor g725 (n_538, in_3[22], in_4[22]);
  or g726 (n_539, in_3[22], in_4[22]);
  or g727 (n_540, in_2[22], in_4[22]);
  or g728 (n_541, in_2[22], in_3[22]);
  xnor g729 (n_282, n_538, in_2[22]);
  xnor g733 (n_283, n_281, n_280);
  or g734 (n_289, n_280, wc, n_281);
  not gc (wc, n_544);
  xnor g735 (n_550, n_287, n_143);
  or g736 (n_551, n_143, wc0);
  not gc0 (wc0, n_287);
  or g737 (n_552, wc1, n_143);
  not gc1 (wc1, n_289);
  or g738 (n_563, n_559, wc2);
  not gc2 (wc2, n_560);
  or g739 (n_782, wc3, n_559);
  not gc3 (wc3, n_562);
  and g740 (n_637, wc4, n_566);
  not gc4 (wc4, n_567);
  or g741 (n_783, wc5, n_569);
  not gc5 (wc5, n_564);
  or g742 (n_786, wc6, n_565);
  not gc6 (wc6, n_566);
  and g743 (n_639, wc7, n_572);
  not gc7 (wc7, n_573);
  or g744 (n_636, wc8, n_569);
  not gc8 (wc8, n_634);
  or g745 (n_787, wc9, n_575);
  not gc9 (wc9, n_570);
  or g746 (n_790, wc10, n_571);
  not gc10 (wc10, n_572);
  and g747 (n_646, wc11, n_578);
  not gc11 (wc11, n_579);
  and g748 (n_649, wc12, n_584);
  not gc12 (wc12, n_585);
  and g749 (n_656, wc13, n_590);
  not gc13 (wc13, n_591);
  and g750 (n_659, wc14, n_596);
  not gc14 (wc14, n_597);
  and g751 (n_666, wc15, n_602);
  not gc15 (wc15, n_603);
  and g752 (n_669, wc16, n_608);
  not gc16 (wc16, n_609);
  and g753 (n_676, wc17, n_614);
  not gc17 (wc17, n_615);
  and g754 (n_679, wc18, n_620);
  not gc18 (wc18, n_621);
  and g755 (n_686, wc19, n_626);
  not gc19 (wc19, n_627);
  or g756 (n_693, wc20, n_581);
  not gc20 (wc20, n_642);
  or g757 (n_735, wc21, n_593);
  not gc21 (wc21, n_652);
  or g758 (n_708, wc22, n_605);
  not gc22 (wc22, n_662);
  or g759 (n_762, wc23, n_617);
  not gc23 (wc23, n_672);
  or g760 (n_723, wc24, n_629);
  not gc24 (wc24, n_682);
  or g761 (n_792, wc25, n_581);
  not gc25 (wc25, n_576);
  or g762 (n_795, wc26, n_577);
  not gc26 (wc26, n_578);
  or g763 (n_796, wc27, n_587);
  not gc27 (wc27, n_582);
  or g764 (n_799, wc28, n_583);
  not gc28 (wc28, n_584);
  or g765 (n_801, wc29, n_593);
  not gc29 (wc29, n_588);
  or g766 (n_804, wc30, n_589);
  not gc30 (wc30, n_590);
  or g767 (n_807, wc31, n_599);
  not gc31 (wc31, n_594);
  or g768 (n_810, wc32, n_595);
  not gc32 (wc32, n_596);
  or g769 (n_812, wc33, n_605);
  not gc33 (wc33, n_600);
  or g770 (n_815, wc34, n_601);
  not gc34 (wc34, n_602);
  or g771 (n_816, wc35, n_611);
  not gc35 (wc35, n_606);
  or g772 (n_819, wc36, n_607);
  not gc36 (wc36, n_608);
  or g773 (n_821, wc37, n_617);
  not gc37 (wc37, n_612);
  or g774 (n_824, wc38, n_613);
  not gc38 (wc38, n_614);
  or g775 (n_827, wc39, n_623);
  not gc39 (wc39, n_618);
  or g776 (n_830, wc40, n_619);
  not gc40 (wc40, n_620);
  or g777 (n_832, wc41, n_629);
  not gc41 (wc41, n_624);
  or g778 (n_835, wc42, n_625);
  not gc42 (wc42, n_626);
  or g779 (n_837, wc43, n_633);
  not gc43 (wc43, n_630);
  and g780 (n_695, wc44, n_576);
  not gc44 (wc44, n_640);
  and g781 (n_647, wc45, n_644);
  not gc45 (wc45, n_639);
  and g782 (n_657, wc46, n_654);
  not gc46 (wc46, n_649);
  and g783 (n_667, wc47, n_664);
  not gc47 (wc47, n_659);
  and g784 (n_677, wc48, n_674);
  not gc48 (wc48, n_669);
  and g785 (n_687, wc49, n_684);
  not gc49 (wc49, n_679);
  or g786 (n_691, wc50, n_575);
  not gc50 (wc50, n_689);
  and g787 (n_744, wc51, n_662);
  not gc51 (wc51, n_704);
  and g788 (n_771, wc52, n_682);
  not gc52 (wc52, n_719);
  and g789 (n_699, wc53, n_646);
  not gc53 (wc53, n_647);
  and g790 (n_737, wc54, n_588);
  not gc54 (wc54, n_650);
  and g791 (n_701, wc55, n_656);
  not gc55 (wc55, n_657);
  and g792 (n_709, wc56, n_600);
  not gc56 (wc56, n_660);
  and g793 (n_713, wc57, n_666);
  not gc57 (wc57, n_667);
  and g794 (n_764, wc58, n_612);
  not gc58 (wc58, n_670);
  and g795 (n_716, wc59, n_676);
  not gc59 (wc59, n_677);
  and g796 (n_724, wc60, n_624);
  not gc60 (wc60, n_680);
  and g797 (n_728, wc61, n_686);
  not gc61 (wc61, n_687);
  or g798 (n_696, n_693, wc62);
  not gc62 (wc62, n_689);
  or g799 (n_700, n_697, wc63);
  not gc63 (wc63, n_689);
  or g800 (n_778, wc64, n_633);
  not gc64 (wc64, n_756);
  and g801 (n_706, wc65, n_662);
  not gc65 (wc65, n_701);
  and g802 (n_721, wc66, n_682);
  not gc66 (wc66, n_716);
  and g803 (n_742, wc67, n_594);
  not gc67 (wc67, n_702);
  and g804 (n_745, wc68, n_659);
  not gc68 (wc68, n_706);
  and g805 (n_748, n_709, wc69);
  not gc69 (wc69, n_710);
  and g806 (n_751, n_713, wc70);
  not gc70 (wc70, n_714);
  and g807 (n_769, wc71, n_618);
  not gc71 (wc71, n_717);
  and g808 (n_772, wc72, n_679);
  not gc72 (wc72, n_721);
  and g809 (n_775, n_724, wc73);
  not gc73 (wc73, n_725);
  and g810 (n_753, n_728, wc74);
  not gc74 (wc74, n_729);
  or g811 (n_733, wc75, n_587);
  not gc75 (wc75, n_731);
  or g812 (n_738, n_735, wc76);
  not gc76 (wc76, n_731);
  or g813 (n_740, wc77, n_704);
  not gc77 (wc77, n_731);
  and g814 (n_780, wc78, n_630);
  not gc78 (wc78, n_754);
  or g815 (n_760, wc79, n_611);
  not gc79 (wc79, n_758);
  or g816 (n_765, n_762, wc80);
  not gc80 (wc80, n_758);
  or g817 (n_767, wc81, n_719);
  not gc81 (wc81, n_758);
  or g818 (n_781, n_778, wc82);
  not gc82 (wc82, n_758);
  not g819 (out_0[25], n_839);
endmodule

module csa_tree_add_767_44_group_6809_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  csa_tree_add_767_44_group_6809_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_841_44_group_6807_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_280, n_281, n_282, n_283, n_284, n_287;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_544, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_556, n_557;
  wire n_558, n_559, n_560, n_562, n_563, n_564, n_565, n_566;
  wire n_567, n_569, n_570, n_571, n_572, n_573, n_575, n_576;
  wire n_577, n_578, n_579, n_581, n_582, n_583, n_584, n_585;
  wire n_587, n_588, n_589, n_590, n_591, n_593, n_594, n_595;
  wire n_596, n_597, n_599, n_600, n_601, n_602, n_603, n_605;
  wire n_606, n_607, n_608, n_609, n_611, n_612, n_613, n_614;
  wire n_615, n_617, n_618, n_619, n_620, n_621, n_623, n_624;
  wire n_625, n_626, n_627, n_629, n_630, n_633, n_634, n_636;
  wire n_637, n_638, n_639, n_640, n_642, n_644, n_646, n_647;
  wire n_649, n_650, n_652, n_654, n_656, n_657, n_659, n_660;
  wire n_662, n_664, n_666, n_667, n_669, n_670, n_672, n_674;
  wire n_676, n_677, n_679, n_680, n_682, n_684, n_686, n_687;
  wire n_689, n_691, n_692, n_693, n_695, n_696, n_697, n_699;
  wire n_700, n_701, n_702, n_704, n_706, n_708, n_709, n_710;
  wire n_712, n_713, n_714, n_716, n_717, n_719, n_721, n_723;
  wire n_724, n_725, n_727, n_728, n_729, n_731, n_733, n_734;
  wire n_735, n_737, n_738, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_756, n_758, n_760, n_761, n_762, n_764;
  wire n_765, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_780, n_781, n_782;
  wire n_783, n_785, n_786, n_787, n_789, n_790, n_791, n_792;
  wire n_794, n_795, n_796, n_798, n_799, n_800, n_801, n_803;
  wire n_804, n_806, n_807, n_809, n_810, n_811, n_812, n_814;
  wire n_815, n_816, n_818, n_819, n_820, n_821, n_823, n_824;
  wire n_826, n_827, n_829, n_830, n_831, n_832, n_834, n_835;
  wire n_836, n_837, n_839, n_841;
  xor g75 (n_290, in_0[0], in_4[0]);
  xor g76 (n_193, n_290, in_3[0]);
  nand g77 (n_291, in_0[0], in_4[0]);
  nand g78 (n_292, in_3[0], in_4[0]);
  nand g79 (n_293, in_0[0], in_3[0]);
  nand g6 (n_195, n_291, n_292, n_293);
  xor g80 (n_294, in_0[1], in_1[1]);
  xor g81 (n_166, n_294, in_4[1]);
  nand g82 (n_295, in_0[1], in_1[1]);
  nand g83 (n_296, in_4[1], in_1[1]);
  nand g84 (n_297, in_0[1], in_4[1]);
  nand g85 (n_197, n_295, n_296, n_297);
  xor g86 (n_298, in_3[1], in_2[1]);
  xor g87 (n_192, n_298, n_195);
  nand g88 (n_299, in_3[1], in_2[1]);
  nand g89 (n_300, n_195, in_2[1]);
  nand g90 (n_301, in_3[1], n_195);
  nand g91 (n_165, n_299, n_300, n_301);
  xor g92 (n_196, in_0[2], in_1[2]);
  and g93 (n_199, in_0[2], in_1[2]);
  xor g94 (n_302, in_3[2], in_4[2]);
  xor g95 (n_198, n_302, in_2[2]);
  nand g96 (n_303, in_3[2], in_4[2]);
  nand g97 (n_304, in_2[2], in_4[2]);
  nand g98 (n_305, in_3[2], in_2[2]);
  nand g99 (n_200, n_303, n_304, n_305);
  xor g100 (n_306, n_196, n_197);
  xor g101 (n_191, n_306, n_198);
  nand g102 (n_307, n_196, n_197);
  nand g103 (n_308, n_198, n_197);
  nand g104 (n_309, n_196, n_198);
  nand g105 (n_164, n_307, n_308, n_309);
  xor g106 (n_310, in_0[3], in_1[3]);
  xor g107 (n_201, n_310, in_3[3]);
  nand g108 (n_311, in_0[3], in_1[3]);
  nand g109 (n_312, in_3[3], in_1[3]);
  nand g110 (n_313, in_0[3], in_3[3]);
  nand g111 (n_203, n_311, n_312, n_313);
  xor g112 (n_314, in_4[3], in_2[3]);
  xor g113 (n_202, n_314, n_199);
  nand g114 (n_315, in_4[3], in_2[3]);
  nand g115 (n_316, n_199, in_2[3]);
  nand g116 (n_317, in_4[3], n_199);
  nand g117 (n_205, n_315, n_316, n_317);
  xor g118 (n_318, n_200, n_201);
  xor g119 (n_190, n_318, n_202);
  nand g120 (n_319, n_200, n_201);
  nand g121 (n_320, n_202, n_201);
  nand g122 (n_321, n_200, n_202);
  nand g123 (n_163, n_319, n_320, n_321);
  xor g124 (n_322, in_0[4], in_1[4]);
  xor g125 (n_204, n_322, in_3[4]);
  nand g126 (n_323, in_0[4], in_1[4]);
  nand g127 (n_324, in_3[4], in_1[4]);
  nand g128 (n_325, in_0[4], in_3[4]);
  nand g129 (n_207, n_323, n_324, n_325);
  xor g130 (n_326, in_4[4], in_2[4]);
  xor g131 (n_206, n_326, n_203);
  nand g132 (n_327, in_4[4], in_2[4]);
  nand g133 (n_328, n_203, in_2[4]);
  nand g134 (n_329, in_4[4], n_203);
  nand g135 (n_210, n_327, n_328, n_329);
  xor g136 (n_330, n_204, n_205);
  xor g137 (n_189, n_330, n_206);
  nand g138 (n_331, n_204, n_205);
  nand g139 (n_332, n_206, n_205);
  nand g140 (n_333, n_204, n_206);
  nand g141 (n_162, n_331, n_332, n_333);
  xor g142 (n_334, in_0[5], in_1[5]);
  xor g143 (n_208, n_334, in_3[5]);
  nand g144 (n_335, in_0[5], in_1[5]);
  nand g145 (n_336, in_3[5], in_1[5]);
  nand g146 (n_337, in_0[5], in_3[5]);
  nand g147 (n_211, n_335, n_336, n_337);
  xor g148 (n_338, in_4[5], in_2[5]);
  xor g149 (n_209, n_338, n_207);
  nand g150 (n_339, in_4[5], in_2[5]);
  nand g151 (n_340, n_207, in_2[5]);
  nand g152 (n_341, in_4[5], n_207);
  nand g153 (n_214, n_339, n_340, n_341);
  xor g154 (n_342, n_208, n_209);
  xor g155 (n_188, n_342, n_210);
  nand g156 (n_343, n_208, n_209);
  nand g157 (n_344, n_210, n_209);
  nand g158 (n_345, n_208, n_210);
  nand g159 (n_161, n_343, n_344, n_345);
  xor g160 (n_346, in_0[6], in_1[6]);
  xor g161 (n_212, n_346, in_3[6]);
  nand g162 (n_347, in_0[6], in_1[6]);
  nand g163 (n_348, in_3[6], in_1[6]);
  nand g164 (n_349, in_0[6], in_3[6]);
  nand g165 (n_215, n_347, n_348, n_349);
  xor g166 (n_350, in_4[6], in_2[6]);
  xor g167 (n_213, n_350, n_211);
  nand g168 (n_351, in_4[6], in_2[6]);
  nand g169 (n_352, n_211, in_2[6]);
  nand g170 (n_353, in_4[6], n_211);
  nand g171 (n_218, n_351, n_352, n_353);
  xor g172 (n_354, n_212, n_213);
  xor g173 (n_187, n_354, n_214);
  nand g174 (n_355, n_212, n_213);
  nand g175 (n_356, n_214, n_213);
  nand g176 (n_357, n_212, n_214);
  nand g177 (n_160, n_355, n_356, n_357);
  xor g178 (n_358, in_0[7], in_1[7]);
  xor g179 (n_216, n_358, in_3[7]);
  nand g180 (n_359, in_0[7], in_1[7]);
  nand g181 (n_360, in_3[7], in_1[7]);
  nand g182 (n_361, in_0[7], in_3[7]);
  nand g183 (n_219, n_359, n_360, n_361);
  xor g184 (n_362, in_4[7], in_2[7]);
  xor g185 (n_217, n_362, n_215);
  nand g186 (n_363, in_4[7], in_2[7]);
  nand g187 (n_364, n_215, in_2[7]);
  nand g188 (n_365, in_4[7], n_215);
  nand g189 (n_222, n_363, n_364, n_365);
  xor g190 (n_366, n_216, n_217);
  xor g191 (n_186, n_366, n_218);
  nand g192 (n_367, n_216, n_217);
  nand g193 (n_368, n_218, n_217);
  nand g194 (n_369, n_216, n_218);
  nand g195 (n_159, n_367, n_368, n_369);
  xor g196 (n_370, in_0[8], in_1[8]);
  xor g197 (n_220, n_370, in_3[8]);
  nand g198 (n_371, in_0[8], in_1[8]);
  nand g199 (n_372, in_3[8], in_1[8]);
  nand g200 (n_373, in_0[8], in_3[8]);
  nand g201 (n_223, n_371, n_372, n_373);
  xor g202 (n_374, in_4[8], in_2[8]);
  xor g203 (n_221, n_374, n_219);
  nand g204 (n_375, in_4[8], in_2[8]);
  nand g205 (n_376, n_219, in_2[8]);
  nand g206 (n_377, in_4[8], n_219);
  nand g207 (n_226, n_375, n_376, n_377);
  xor g208 (n_378, n_220, n_221);
  xor g209 (n_185, n_378, n_222);
  nand g210 (n_379, n_220, n_221);
  nand g211 (n_380, n_222, n_221);
  nand g212 (n_381, n_220, n_222);
  nand g213 (n_158, n_379, n_380, n_381);
  xor g214 (n_382, in_0[9], in_1[9]);
  xor g215 (n_224, n_382, in_3[9]);
  nand g216 (n_383, in_0[9], in_1[9]);
  nand g217 (n_384, in_3[9], in_1[9]);
  nand g218 (n_385, in_0[9], in_3[9]);
  nand g219 (n_227, n_383, n_384, n_385);
  xor g220 (n_386, in_4[9], in_2[9]);
  xor g221 (n_225, n_386, n_223);
  nand g222 (n_387, in_4[9], in_2[9]);
  nand g223 (n_388, n_223, in_2[9]);
  nand g224 (n_389, in_4[9], n_223);
  nand g225 (n_230, n_387, n_388, n_389);
  xor g226 (n_390, n_224, n_225);
  xor g227 (n_184, n_390, n_226);
  nand g228 (n_391, n_224, n_225);
  nand g229 (n_392, n_226, n_225);
  nand g230 (n_393, n_224, n_226);
  nand g231 (n_157, n_391, n_392, n_393);
  xor g232 (n_394, in_0[10], in_1[10]);
  xor g233 (n_228, n_394, in_3[10]);
  nand g234 (n_395, in_0[10], in_1[10]);
  nand g235 (n_396, in_3[10], in_1[10]);
  nand g236 (n_397, in_0[10], in_3[10]);
  nand g237 (n_231, n_395, n_396, n_397);
  xor g238 (n_398, in_4[10], in_2[10]);
  xor g239 (n_229, n_398, n_227);
  nand g240 (n_399, in_4[10], in_2[10]);
  nand g241 (n_400, n_227, in_2[10]);
  nand g242 (n_401, in_4[10], n_227);
  nand g243 (n_234, n_399, n_400, n_401);
  xor g244 (n_402, n_228, n_229);
  xor g245 (n_183, n_402, n_230);
  nand g246 (n_403, n_228, n_229);
  nand g247 (n_404, n_230, n_229);
  nand g248 (n_405, n_228, n_230);
  nand g249 (n_156, n_403, n_404, n_405);
  xor g250 (n_406, in_0[11], in_1[11]);
  xor g251 (n_232, n_406, in_3[11]);
  nand g252 (n_407, in_0[11], in_1[11]);
  nand g253 (n_408, in_3[11], in_1[11]);
  nand g254 (n_409, in_0[11], in_3[11]);
  nand g255 (n_235, n_407, n_408, n_409);
  xor g256 (n_410, in_4[11], in_2[11]);
  xor g257 (n_233, n_410, n_231);
  nand g258 (n_411, in_4[11], in_2[11]);
  nand g259 (n_412, n_231, in_2[11]);
  nand g260 (n_413, in_4[11], n_231);
  nand g261 (n_238, n_411, n_412, n_413);
  xor g262 (n_414, n_232, n_233);
  xor g263 (n_182, n_414, n_234);
  nand g264 (n_415, n_232, n_233);
  nand g265 (n_416, n_234, n_233);
  nand g266 (n_417, n_232, n_234);
  nand g267 (n_155, n_415, n_416, n_417);
  xor g268 (n_418, in_0[12], in_1[12]);
  xor g269 (n_236, n_418, in_3[12]);
  nand g270 (n_419, in_0[12], in_1[12]);
  nand g271 (n_420, in_3[12], in_1[12]);
  nand g272 (n_421, in_0[12], in_3[12]);
  nand g273 (n_239, n_419, n_420, n_421);
  xor g274 (n_422, in_4[12], in_2[12]);
  xor g275 (n_237, n_422, n_235);
  nand g276 (n_423, in_4[12], in_2[12]);
  nand g277 (n_424, n_235, in_2[12]);
  nand g278 (n_425, in_4[12], n_235);
  nand g279 (n_242, n_423, n_424, n_425);
  xor g280 (n_426, n_236, n_237);
  xor g281 (n_181, n_426, n_238);
  nand g282 (n_427, n_236, n_237);
  nand g283 (n_428, n_238, n_237);
  nand g284 (n_429, n_236, n_238);
  nand g285 (n_154, n_427, n_428, n_429);
  xor g286 (n_430, in_0[13], in_1[13]);
  xor g287 (n_240, n_430, in_3[13]);
  nand g288 (n_431, in_0[13], in_1[13]);
  nand g289 (n_432, in_3[13], in_1[13]);
  nand g290 (n_433, in_0[13], in_3[13]);
  nand g291 (n_243, n_431, n_432, n_433);
  xor g292 (n_434, in_4[13], in_2[13]);
  xor g293 (n_241, n_434, n_239);
  nand g294 (n_435, in_4[13], in_2[13]);
  nand g295 (n_436, n_239, in_2[13]);
  nand g296 (n_437, in_4[13], n_239);
  nand g297 (n_246, n_435, n_436, n_437);
  xor g298 (n_438, n_240, n_241);
  xor g299 (n_180, n_438, n_242);
  nand g300 (n_439, n_240, n_241);
  nand g301 (n_440, n_242, n_241);
  nand g302 (n_441, n_240, n_242);
  nand g303 (n_153, n_439, n_440, n_441);
  xor g304 (n_442, in_0[14], in_1[14]);
  xor g305 (n_244, n_442, in_3[14]);
  nand g306 (n_443, in_0[14], in_1[14]);
  nand g307 (n_444, in_3[14], in_1[14]);
  nand g308 (n_445, in_0[14], in_3[14]);
  nand g309 (n_247, n_443, n_444, n_445);
  xor g310 (n_446, in_4[14], in_2[14]);
  xor g311 (n_245, n_446, n_243);
  nand g312 (n_447, in_4[14], in_2[14]);
  nand g313 (n_448, n_243, in_2[14]);
  nand g314 (n_449, in_4[14], n_243);
  nand g315 (n_250, n_447, n_448, n_449);
  xor g316 (n_450, n_244, n_245);
  xor g317 (n_179, n_450, n_246);
  nand g318 (n_451, n_244, n_245);
  nand g319 (n_452, n_246, n_245);
  nand g320 (n_453, n_244, n_246);
  nand g321 (n_152, n_451, n_452, n_453);
  xor g322 (n_454, in_0[15], in_1[15]);
  xor g323 (n_248, n_454, in_3[15]);
  nand g324 (n_455, in_0[15], in_1[15]);
  nand g325 (n_456, in_3[15], in_1[15]);
  nand g326 (n_457, in_0[15], in_3[15]);
  nand g327 (n_251, n_455, n_456, n_457);
  xor g328 (n_458, in_4[15], in_2[15]);
  xor g329 (n_249, n_458, n_247);
  nand g330 (n_459, in_4[15], in_2[15]);
  nand g331 (n_460, n_247, in_2[15]);
  nand g332 (n_461, in_4[15], n_247);
  nand g333 (n_254, n_459, n_460, n_461);
  xor g334 (n_462, n_248, n_249);
  xor g335 (n_178, n_462, n_250);
  nand g336 (n_463, n_248, n_249);
  nand g337 (n_464, n_250, n_249);
  nand g338 (n_465, n_248, n_250);
  nand g339 (n_151, n_463, n_464, n_465);
  xor g340 (n_466, in_0[16], in_1[16]);
  xor g341 (n_252, n_466, in_3[16]);
  nand g342 (n_467, in_0[16], in_1[16]);
  nand g343 (n_468, in_3[16], in_1[16]);
  nand g344 (n_469, in_0[16], in_3[16]);
  nand g345 (n_255, n_467, n_468, n_469);
  xor g346 (n_470, in_4[16], in_2[16]);
  xor g347 (n_253, n_470, n_251);
  nand g348 (n_471, in_4[16], in_2[16]);
  nand g349 (n_472, n_251, in_2[16]);
  nand g350 (n_473, in_4[16], n_251);
  nand g351 (n_258, n_471, n_472, n_473);
  xor g352 (n_474, n_252, n_253);
  xor g353 (n_177, n_474, n_254);
  nand g354 (n_475, n_252, n_253);
  nand g355 (n_476, n_254, n_253);
  nand g356 (n_477, n_252, n_254);
  nand g357 (n_150, n_475, n_476, n_477);
  xor g358 (n_478, in_0[17], in_1[17]);
  xor g359 (n_256, n_478, in_3[17]);
  nand g360 (n_479, in_0[17], in_1[17]);
  nand g361 (n_480, in_3[17], in_1[17]);
  nand g362 (n_481, in_0[17], in_3[17]);
  nand g363 (n_259, n_479, n_480, n_481);
  xor g364 (n_482, in_4[17], in_2[17]);
  xor g365 (n_257, n_482, n_255);
  nand g366 (n_483, in_4[17], in_2[17]);
  nand g367 (n_484, n_255, in_2[17]);
  nand g368 (n_485, in_4[17], n_255);
  nand g369 (n_262, n_483, n_484, n_485);
  xor g370 (n_486, n_256, n_257);
  xor g371 (n_176, n_486, n_258);
  nand g372 (n_487, n_256, n_257);
  nand g373 (n_488, n_258, n_257);
  nand g374 (n_489, n_256, n_258);
  nand g375 (n_149, n_487, n_488, n_489);
  xor g376 (n_490, in_0[18], in_1[18]);
  xor g377 (n_260, n_490, in_3[18]);
  nand g378 (n_491, in_0[18], in_1[18]);
  nand g379 (n_492, in_3[18], in_1[18]);
  nand g380 (n_493, in_0[18], in_3[18]);
  nand g381 (n_263, n_491, n_492, n_493);
  xor g382 (n_494, in_4[18], in_2[18]);
  xor g383 (n_261, n_494, n_259);
  nand g384 (n_495, in_4[18], in_2[18]);
  nand g385 (n_496, n_259, in_2[18]);
  nand g386 (n_497, in_4[18], n_259);
  nand g387 (n_266, n_495, n_496, n_497);
  xor g388 (n_498, n_260, n_261);
  xor g389 (n_175, n_498, n_262);
  nand g390 (n_499, n_260, n_261);
  nand g391 (n_500, n_262, n_261);
  nand g392 (n_501, n_260, n_262);
  nand g393 (n_148, n_499, n_500, n_501);
  xor g394 (n_502, in_0[19], in_1[19]);
  xor g395 (n_264, n_502, in_3[19]);
  nand g396 (n_503, in_0[19], in_1[19]);
  nand g397 (n_504, in_3[19], in_1[19]);
  nand g398 (n_505, in_0[19], in_3[19]);
  nand g399 (n_267, n_503, n_504, n_505);
  xor g400 (n_506, in_4[19], in_2[19]);
  xor g401 (n_265, n_506, n_263);
  nand g402 (n_507, in_4[19], in_2[19]);
  nand g403 (n_508, n_263, in_2[19]);
  nand g404 (n_509, in_4[19], n_263);
  nand g405 (n_270, n_507, n_508, n_509);
  xor g406 (n_510, n_264, n_265);
  xor g407 (n_174, n_510, n_266);
  nand g408 (n_511, n_264, n_265);
  nand g409 (n_512, n_266, n_265);
  nand g410 (n_513, n_264, n_266);
  nand g411 (n_147, n_511, n_512, n_513);
  xor g412 (n_514, in_0[20], in_1[20]);
  xor g413 (n_268, n_514, in_3[20]);
  nand g414 (n_515, in_0[20], in_1[20]);
  nand g415 (n_516, in_3[20], in_1[20]);
  nand g416 (n_517, in_0[20], in_3[20]);
  nand g417 (n_271, n_515, n_516, n_517);
  xor g418 (n_518, in_4[20], in_2[20]);
  xor g419 (n_269, n_518, n_267);
  nand g420 (n_519, in_4[20], in_2[20]);
  nand g421 (n_520, n_267, in_2[20]);
  nand g422 (n_521, in_4[20], n_267);
  nand g423 (n_274, n_519, n_520, n_521);
  xor g424 (n_522, n_268, n_269);
  xor g425 (n_173, n_522, n_270);
  nand g426 (n_523, n_268, n_269);
  nand g427 (n_524, n_270, n_269);
  nand g428 (n_525, n_268, n_270);
  nand g429 (n_146, n_523, n_524, n_525);
  xor g430 (n_526, in_0[21], in_1[21]);
  xor g431 (n_272, n_526, in_3[21]);
  nand g432 (n_527, in_0[21], in_1[21]);
  nand g433 (n_528, in_3[21], in_1[21]);
  nand g434 (n_529, in_0[21], in_3[21]);
  nand g435 (n_281, n_527, n_528, n_529);
  xor g436 (n_530, in_4[21], in_2[21]);
  xor g437 (n_273, n_530, n_271);
  nand g438 (n_531, in_4[21], in_2[21]);
  nand g439 (n_532, n_271, in_2[21]);
  nand g440 (n_533, in_4[21], n_271);
  nand g441 (n_284, n_531, n_532, n_533);
  xor g442 (n_534, n_272, n_273);
  xor g443 (n_172, n_534, n_274);
  nand g444 (n_535, n_272, n_273);
  nand g445 (n_536, n_274, n_273);
  nand g446 (n_537, n_272, n_274);
  nand g447 (n_145, n_535, n_536, n_537);
  nand g455 (n_287, n_539, n_540, n_541);
  nand g459 (n_544, n_281, n_280);
  xor g462 (n_546, n_282, n_283);
  xor g463 (n_171, n_546, n_284);
  nand g464 (n_547, n_282, n_283);
  nand g465 (n_548, n_284, n_283);
  nand g466 (n_549, n_282, n_284);
  nand g467 (n_144, n_547, n_548, n_549);
  xor g471 (n_170, n_550, n_289);
  nand g474 (n_553, n_287, n_289);
  nand g475 (n_169, n_551, n_552, n_553);
  xor g478 (n_841, in_1[0], n_193);
  nand g479 (n_556, in_1[0], n_193);
  nand g480 (n_557, in_1[0], in_2[0]);
  nand g7 (n_558, n_193, in_2[0]);
  nand g8 (n_560, n_556, n_557, n_558);
  nor g9 (n_559, n_166, n_192);
  nand g10 (n_562, n_166, n_192);
  nor g11 (n_569, n_165, n_191);
  nand g12 (n_564, n_165, n_191);
  nor g13 (n_565, n_164, n_190);
  nand g14 (n_566, n_164, n_190);
  nor g15 (n_575, n_163, n_189);
  nand g16 (n_570, n_163, n_189);
  nor g17 (n_571, n_162, n_188);
  nand g18 (n_572, n_162, n_188);
  nor g19 (n_581, n_161, n_187);
  nand g20 (n_576, n_161, n_187);
  nor g21 (n_577, n_160, n_186);
  nand g22 (n_578, n_160, n_186);
  nor g23 (n_587, n_159, n_185);
  nand g24 (n_582, n_159, n_185);
  nor g25 (n_583, n_158, n_184);
  nand g26 (n_584, n_158, n_184);
  nor g27 (n_593, n_157, n_183);
  nand g28 (n_588, n_157, n_183);
  nor g29 (n_589, n_156, n_182);
  nand g30 (n_590, n_156, n_182);
  nor g31 (n_599, n_155, n_181);
  nand g32 (n_594, n_155, n_181);
  nor g33 (n_595, n_154, n_180);
  nand g34 (n_596, n_154, n_180);
  nor g35 (n_605, n_153, n_179);
  nand g36 (n_600, n_153, n_179);
  nor g37 (n_601, n_152, n_178);
  nand g38 (n_602, n_152, n_178);
  nor g39 (n_611, n_151, n_177);
  nand g40 (n_606, n_151, n_177);
  nor g41 (n_607, n_150, n_176);
  nand g42 (n_608, n_150, n_176);
  nor g43 (n_617, n_149, n_175);
  nand g44 (n_612, n_149, n_175);
  nor g45 (n_613, n_148, n_174);
  nand g46 (n_614, n_148, n_174);
  nor g47 (n_623, n_147, n_173);
  nand g48 (n_618, n_147, n_173);
  nor g49 (n_619, n_146, n_172);
  nand g50 (n_620, n_146, n_172);
  nor g51 (n_629, n_145, n_171);
  nand g52 (n_624, n_145, n_171);
  nor g53 (n_625, n_144, n_170);
  nand g54 (n_626, n_144, n_170);
  nor g55 (n_633, n_143, n_169);
  nand g56 (n_630, n_143, n_169);
  nand g61 (n_634, n_562, n_563);
  nor g62 (n_567, n_564, n_565);
  nor g65 (n_167, n_569, n_565);
  nor g66 (n_573, n_570, n_571);
  nor g69 (n_642, n_575, n_571);
  nor g70 (n_579, n_576, n_577);
  nor g73 (n_644, n_581, n_577);
  nor g74 (n_585, n_582, n_583);
  nor g483 (n_652, n_587, n_583);
  nor g484 (n_591, n_588, n_589);
  nor g487 (n_654, n_593, n_589);
  nor g488 (n_597, n_594, n_595);
  nor g491 (n_662, n_599, n_595);
  nor g492 (n_603, n_600, n_601);
  nor g495 (n_664, n_605, n_601);
  nor g496 (n_609, n_606, n_607);
  nor g499 (n_672, n_611, n_607);
  nor g500 (n_615, n_612, n_613);
  nor g503 (n_674, n_617, n_613);
  nor g504 (n_621, n_618, n_619);
  nor g507 (n_682, n_623, n_619);
  nor g508 (n_627, n_624, n_625);
  nor g511 (n_684, n_629, n_625);
  nand g514 (n_785, n_564, n_636);
  nand g515 (n_638, n_167, n_634);
  nand g516 (n_689, n_637, n_638);
  nor g517 (n_640, n_581, n_639);
  nand g526 (n_697, n_642, n_644);
  nor g527 (n_650, n_593, n_649);
  nand g536 (n_704, n_652, n_654);
  nor g537 (n_660, n_605, n_659);
  nand g546 (n_712, n_662, n_664);
  nor g547 (n_670, n_617, n_669);
  nand g556 (n_719, n_672, n_674);
  nor g557 (n_680, n_629, n_679);
  nand g566 (n_727, n_682, n_684);
  nand g569 (n_789, n_570, n_691);
  nand g570 (n_692, n_642, n_689);
  nand g571 (n_791, n_639, n_692);
  nand g574 (n_794, n_695, n_696);
  nand g577 (n_731, n_699, n_700);
  nor g578 (n_702, n_599, n_701);
  nor g581 (n_741, n_599, n_704);
  nor g587 (n_710, n_708, n_701);
  nor g590 (n_747, n_704, n_708);
  nor g591 (n_714, n_712, n_701);
  nor g594 (n_750, n_704, n_712);
  nor g595 (n_717, n_623, n_716);
  nor g598 (n_768, n_623, n_719);
  nor g604 (n_725, n_723, n_716);
  nor g607 (n_774, n_719, n_723);
  nor g608 (n_729, n_727, n_716);
  nor g611 (n_756, n_719, n_727);
  nand g614 (n_798, n_582, n_733);
  nand g615 (n_734, n_652, n_731);
  nand g616 (n_800, n_649, n_734);
  nand g619 (n_803, n_737, n_738);
  nand g622 (n_806, n_701, n_740);
  nand g623 (n_743, n_741, n_731);
  nand g624 (n_809, n_742, n_743);
  nand g625 (n_746, n_744, n_731);
  nand g626 (n_811, n_745, n_746);
  nand g627 (n_749, n_747, n_731);
  nand g628 (n_814, n_748, n_749);
  nand g629 (n_752, n_750, n_731);
  nand g630 (n_758, n_751, n_752);
  nor g631 (n_754, n_633, n_753);
  nand g638 (n_818, n_606, n_760);
  nand g639 (n_761, n_672, n_758);
  nand g640 (n_820, n_669, n_761);
  nand g643 (n_823, n_764, n_765);
  nand g646 (n_826, n_716, n_767);
  nand g647 (n_770, n_768, n_758);
  nand g648 (n_829, n_769, n_770);
  nand g649 (n_773, n_771, n_758);
  nand g650 (n_831, n_772, n_773);
  nand g651 (n_776, n_774, n_758);
  nand g652 (n_834, n_775, n_776);
  nand g653 (n_777, n_756, n_758);
  nand g654 (n_836, n_753, n_777);
  nand g657 (n_839, n_780, n_781);
  xnor g659 (out_0[1], n_560, n_782);
  xnor g661 (out_0[2], n_634, n_783);
  xnor g664 (out_0[3], n_785, n_786);
  xnor g666 (out_0[4], n_689, n_787);
  xnor g669 (out_0[5], n_789, n_790);
  xnor g671 (out_0[6], n_791, n_792);
  xnor g674 (out_0[7], n_794, n_795);
  xnor g676 (out_0[8], n_731, n_796);
  xnor g679 (out_0[9], n_798, n_799);
  xnor g681 (out_0[10], n_800, n_801);
  xnor g684 (out_0[11], n_803, n_804);
  xnor g687 (out_0[12], n_806, n_807);
  xnor g690 (out_0[13], n_809, n_810);
  xnor g692 (out_0[14], n_811, n_812);
  xnor g695 (out_0[15], n_814, n_815);
  xnor g697 (out_0[16], n_758, n_816);
  xnor g700 (out_0[17], n_818, n_819);
  xnor g702 (out_0[18], n_820, n_821);
  xnor g705 (out_0[19], n_823, n_824);
  xnor g708 (out_0[20], n_826, n_827);
  xnor g711 (out_0[21], n_829, n_830);
  xnor g713 (out_0[22], n_831, n_832);
  xnor g716 (out_0[23], n_834, n_835);
  xnor g718 (out_0[24], n_836, n_837);
  xor g722 (out_0[0], in_2[0], n_841);
  xor g723 (n_280, in_0[22], in_1[22]);
  nor g724 (n_143, in_0[22], in_1[22]);
  xor g725 (n_538, in_3[22], in_4[22]);
  or g726 (n_539, in_3[22], in_4[22]);
  or g727 (n_540, in_2[22], in_4[22]);
  or g728 (n_541, in_2[22], in_3[22]);
  xnor g729 (n_282, n_538, in_2[22]);
  xnor g733 (n_283, n_281, n_280);
  or g734 (n_289, n_280, wc, n_281);
  not gc (wc, n_544);
  xnor g735 (n_550, n_287, n_143);
  or g736 (n_551, n_143, wc0);
  not gc0 (wc0, n_287);
  or g737 (n_552, wc1, n_143);
  not gc1 (wc1, n_289);
  or g738 (n_563, n_559, wc2);
  not gc2 (wc2, n_560);
  or g739 (n_782, wc3, n_559);
  not gc3 (wc3, n_562);
  and g740 (n_637, wc4, n_566);
  not gc4 (wc4, n_567);
  or g741 (n_783, wc5, n_569);
  not gc5 (wc5, n_564);
  or g742 (n_786, wc6, n_565);
  not gc6 (wc6, n_566);
  and g743 (n_639, wc7, n_572);
  not gc7 (wc7, n_573);
  or g744 (n_636, wc8, n_569);
  not gc8 (wc8, n_634);
  or g745 (n_787, wc9, n_575);
  not gc9 (wc9, n_570);
  or g746 (n_790, wc10, n_571);
  not gc10 (wc10, n_572);
  and g747 (n_646, wc11, n_578);
  not gc11 (wc11, n_579);
  and g748 (n_649, wc12, n_584);
  not gc12 (wc12, n_585);
  and g749 (n_656, wc13, n_590);
  not gc13 (wc13, n_591);
  and g750 (n_659, wc14, n_596);
  not gc14 (wc14, n_597);
  and g751 (n_666, wc15, n_602);
  not gc15 (wc15, n_603);
  and g752 (n_669, wc16, n_608);
  not gc16 (wc16, n_609);
  and g753 (n_676, wc17, n_614);
  not gc17 (wc17, n_615);
  and g754 (n_679, wc18, n_620);
  not gc18 (wc18, n_621);
  and g755 (n_686, wc19, n_626);
  not gc19 (wc19, n_627);
  or g756 (n_693, wc20, n_581);
  not gc20 (wc20, n_642);
  or g757 (n_735, wc21, n_593);
  not gc21 (wc21, n_652);
  or g758 (n_708, wc22, n_605);
  not gc22 (wc22, n_662);
  or g759 (n_762, wc23, n_617);
  not gc23 (wc23, n_672);
  or g760 (n_723, wc24, n_629);
  not gc24 (wc24, n_682);
  or g761 (n_792, wc25, n_581);
  not gc25 (wc25, n_576);
  or g762 (n_795, wc26, n_577);
  not gc26 (wc26, n_578);
  or g763 (n_796, wc27, n_587);
  not gc27 (wc27, n_582);
  or g764 (n_799, wc28, n_583);
  not gc28 (wc28, n_584);
  or g765 (n_801, wc29, n_593);
  not gc29 (wc29, n_588);
  or g766 (n_804, wc30, n_589);
  not gc30 (wc30, n_590);
  or g767 (n_807, wc31, n_599);
  not gc31 (wc31, n_594);
  or g768 (n_810, wc32, n_595);
  not gc32 (wc32, n_596);
  or g769 (n_812, wc33, n_605);
  not gc33 (wc33, n_600);
  or g770 (n_815, wc34, n_601);
  not gc34 (wc34, n_602);
  or g771 (n_816, wc35, n_611);
  not gc35 (wc35, n_606);
  or g772 (n_819, wc36, n_607);
  not gc36 (wc36, n_608);
  or g773 (n_821, wc37, n_617);
  not gc37 (wc37, n_612);
  or g774 (n_824, wc38, n_613);
  not gc38 (wc38, n_614);
  or g775 (n_827, wc39, n_623);
  not gc39 (wc39, n_618);
  or g776 (n_830, wc40, n_619);
  not gc40 (wc40, n_620);
  or g777 (n_832, wc41, n_629);
  not gc41 (wc41, n_624);
  or g778 (n_835, wc42, n_625);
  not gc42 (wc42, n_626);
  or g779 (n_837, wc43, n_633);
  not gc43 (wc43, n_630);
  and g780 (n_695, wc44, n_576);
  not gc44 (wc44, n_640);
  and g781 (n_647, wc45, n_644);
  not gc45 (wc45, n_639);
  and g782 (n_657, wc46, n_654);
  not gc46 (wc46, n_649);
  and g783 (n_667, wc47, n_664);
  not gc47 (wc47, n_659);
  and g784 (n_677, wc48, n_674);
  not gc48 (wc48, n_669);
  and g785 (n_687, wc49, n_684);
  not gc49 (wc49, n_679);
  or g786 (n_691, wc50, n_575);
  not gc50 (wc50, n_689);
  and g787 (n_744, wc51, n_662);
  not gc51 (wc51, n_704);
  and g788 (n_771, wc52, n_682);
  not gc52 (wc52, n_719);
  and g789 (n_699, wc53, n_646);
  not gc53 (wc53, n_647);
  and g790 (n_737, wc54, n_588);
  not gc54 (wc54, n_650);
  and g791 (n_701, wc55, n_656);
  not gc55 (wc55, n_657);
  and g792 (n_709, wc56, n_600);
  not gc56 (wc56, n_660);
  and g793 (n_713, wc57, n_666);
  not gc57 (wc57, n_667);
  and g794 (n_764, wc58, n_612);
  not gc58 (wc58, n_670);
  and g795 (n_716, wc59, n_676);
  not gc59 (wc59, n_677);
  and g796 (n_724, wc60, n_624);
  not gc60 (wc60, n_680);
  and g797 (n_728, wc61, n_686);
  not gc61 (wc61, n_687);
  or g798 (n_696, n_693, wc62);
  not gc62 (wc62, n_689);
  or g799 (n_700, n_697, wc63);
  not gc63 (wc63, n_689);
  or g800 (n_778, wc64, n_633);
  not gc64 (wc64, n_756);
  and g801 (n_706, wc65, n_662);
  not gc65 (wc65, n_701);
  and g802 (n_721, wc66, n_682);
  not gc66 (wc66, n_716);
  and g803 (n_742, wc67, n_594);
  not gc67 (wc67, n_702);
  and g804 (n_745, wc68, n_659);
  not gc68 (wc68, n_706);
  and g805 (n_748, n_709, wc69);
  not gc69 (wc69, n_710);
  and g806 (n_751, n_713, wc70);
  not gc70 (wc70, n_714);
  and g807 (n_769, wc71, n_618);
  not gc71 (wc71, n_717);
  and g808 (n_772, wc72, n_679);
  not gc72 (wc72, n_721);
  and g809 (n_775, n_724, wc73);
  not gc73 (wc73, n_725);
  and g810 (n_753, n_728, wc74);
  not gc74 (wc74, n_729);
  or g811 (n_733, wc75, n_587);
  not gc75 (wc75, n_731);
  or g812 (n_738, n_735, wc76);
  not gc76 (wc76, n_731);
  or g813 (n_740, wc77, n_704);
  not gc77 (wc77, n_731);
  and g814 (n_780, wc78, n_630);
  not gc78 (wc78, n_754);
  or g815 (n_760, wc79, n_611);
  not gc79 (wc79, n_758);
  or g816 (n_765, n_762, wc80);
  not gc80 (wc80, n_758);
  or g817 (n_767, wc81, n_719);
  not gc81 (wc81, n_758);
  or g818 (n_781, n_778, wc82);
  not gc82 (wc82, n_758);
  not g819 (out_0[25], n_839);
endmodule

module csa_tree_add_841_44_group_6807_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  csa_tree_add_841_44_group_6807_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module csa_tree_add_915_44_group_6805_GENERIC_REAL(in_0, in_1, in_2,
     in_3, in_4, out_0);
// synthesis_equation "assign out_0 = ( ( ( ( $signed(in_3) + $signed(in_4) )  + $signed(in_2) )  + $signed(in_1) )  + $signed(in_0) )  ;"
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  wire n_143, n_144, n_145, n_146, n_147, n_148, n_149, n_150;
  wire n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158;
  wire n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166;
  wire n_167, n_169, n_170, n_171, n_172, n_173, n_174, n_175;
  wire n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183;
  wire n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191;
  wire n_192, n_193, n_195, n_196, n_197, n_198, n_199, n_200;
  wire n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_213, n_214, n_215, n_216;
  wire n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224;
  wire n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232;
  wire n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240;
  wire n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248;
  wire n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256;
  wire n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264;
  wire n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_272;
  wire n_273, n_274, n_280, n_281, n_282, n_283, n_284, n_287;
  wire n_289, n_290, n_291, n_292, n_293, n_294, n_295, n_296;
  wire n_297, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_310, n_311, n_312;
  wire n_313, n_314, n_315, n_316, n_317, n_318, n_319, n_320;
  wire n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328;
  wire n_329, n_330, n_331, n_332, n_333, n_334, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352;
  wire n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_391, n_392;
  wire n_393, n_394, n_395, n_396, n_397, n_398, n_399, n_400;
  wire n_401, n_402, n_403, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448;
  wire n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504;
  wire n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512;
  wire n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520;
  wire n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528;
  wire n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_544, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_556, n_557;
  wire n_558, n_559, n_560, n_562, n_563, n_564, n_565, n_566;
  wire n_567, n_569, n_570, n_571, n_572, n_573, n_575, n_576;
  wire n_577, n_578, n_579, n_581, n_582, n_583, n_584, n_585;
  wire n_587, n_588, n_589, n_590, n_591, n_593, n_594, n_595;
  wire n_596, n_597, n_599, n_600, n_601, n_602, n_603, n_605;
  wire n_606, n_607, n_608, n_609, n_611, n_612, n_613, n_614;
  wire n_615, n_617, n_618, n_619, n_620, n_621, n_623, n_624;
  wire n_625, n_626, n_627, n_629, n_630, n_633, n_634, n_636;
  wire n_637, n_638, n_639, n_640, n_642, n_644, n_646, n_647;
  wire n_649, n_650, n_652, n_654, n_656, n_657, n_659, n_660;
  wire n_662, n_664, n_666, n_667, n_669, n_670, n_672, n_674;
  wire n_676, n_677, n_679, n_680, n_682, n_684, n_686, n_687;
  wire n_689, n_691, n_692, n_693, n_695, n_696, n_697, n_699;
  wire n_700, n_701, n_702, n_704, n_706, n_708, n_709, n_710;
  wire n_712, n_713, n_714, n_716, n_717, n_719, n_721, n_723;
  wire n_724, n_725, n_727, n_728, n_729, n_731, n_733, n_734;
  wire n_735, n_737, n_738, n_740, n_741, n_742, n_743, n_744;
  wire n_745, n_746, n_747, n_748, n_749, n_750, n_751, n_752;
  wire n_753, n_754, n_756, n_758, n_760, n_761, n_762, n_764;
  wire n_765, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_778, n_780, n_781, n_782;
  wire n_783, n_785, n_786, n_787, n_789, n_790, n_791, n_792;
  wire n_794, n_795, n_796, n_798, n_799, n_800, n_801, n_803;
  wire n_804, n_806, n_807, n_809, n_810, n_811, n_812, n_814;
  wire n_815, n_816, n_818, n_819, n_820, n_821, n_823, n_824;
  wire n_826, n_827, n_829, n_830, n_831, n_832, n_834, n_835;
  wire n_836, n_837, n_839, n_841;
  xor g75 (n_290, in_0[0], in_4[0]);
  xor g76 (n_193, n_290, in_3[0]);
  nand g77 (n_291, in_0[0], in_4[0]);
  nand g78 (n_292, in_3[0], in_4[0]);
  nand g79 (n_293, in_0[0], in_3[0]);
  nand g6 (n_195, n_291, n_292, n_293);
  xor g80 (n_294, in_0[1], in_1[1]);
  xor g81 (n_166, n_294, in_4[1]);
  nand g82 (n_295, in_0[1], in_1[1]);
  nand g83 (n_296, in_4[1], in_1[1]);
  nand g84 (n_297, in_0[1], in_4[1]);
  nand g85 (n_197, n_295, n_296, n_297);
  xor g86 (n_298, in_3[1], in_2[1]);
  xor g87 (n_192, n_298, n_195);
  nand g88 (n_299, in_3[1], in_2[1]);
  nand g89 (n_300, n_195, in_2[1]);
  nand g90 (n_301, in_3[1], n_195);
  nand g91 (n_165, n_299, n_300, n_301);
  xor g92 (n_196, in_0[2], in_1[2]);
  and g93 (n_199, in_0[2], in_1[2]);
  xor g94 (n_302, in_3[2], in_4[2]);
  xor g95 (n_198, n_302, in_2[2]);
  nand g96 (n_303, in_3[2], in_4[2]);
  nand g97 (n_304, in_2[2], in_4[2]);
  nand g98 (n_305, in_3[2], in_2[2]);
  nand g99 (n_200, n_303, n_304, n_305);
  xor g100 (n_306, n_196, n_197);
  xor g101 (n_191, n_306, n_198);
  nand g102 (n_307, n_196, n_197);
  nand g103 (n_308, n_198, n_197);
  nand g104 (n_309, n_196, n_198);
  nand g105 (n_164, n_307, n_308, n_309);
  xor g106 (n_310, in_0[3], in_1[3]);
  xor g107 (n_201, n_310, in_3[3]);
  nand g108 (n_311, in_0[3], in_1[3]);
  nand g109 (n_312, in_3[3], in_1[3]);
  nand g110 (n_313, in_0[3], in_3[3]);
  nand g111 (n_203, n_311, n_312, n_313);
  xor g112 (n_314, in_4[3], in_2[3]);
  xor g113 (n_202, n_314, n_199);
  nand g114 (n_315, in_4[3], in_2[3]);
  nand g115 (n_316, n_199, in_2[3]);
  nand g116 (n_317, in_4[3], n_199);
  nand g117 (n_205, n_315, n_316, n_317);
  xor g118 (n_318, n_200, n_201);
  xor g119 (n_190, n_318, n_202);
  nand g120 (n_319, n_200, n_201);
  nand g121 (n_320, n_202, n_201);
  nand g122 (n_321, n_200, n_202);
  nand g123 (n_163, n_319, n_320, n_321);
  xor g124 (n_322, in_0[4], in_1[4]);
  xor g125 (n_204, n_322, in_3[4]);
  nand g126 (n_323, in_0[4], in_1[4]);
  nand g127 (n_324, in_3[4], in_1[4]);
  nand g128 (n_325, in_0[4], in_3[4]);
  nand g129 (n_207, n_323, n_324, n_325);
  xor g130 (n_326, in_4[4], in_2[4]);
  xor g131 (n_206, n_326, n_203);
  nand g132 (n_327, in_4[4], in_2[4]);
  nand g133 (n_328, n_203, in_2[4]);
  nand g134 (n_329, in_4[4], n_203);
  nand g135 (n_210, n_327, n_328, n_329);
  xor g136 (n_330, n_204, n_205);
  xor g137 (n_189, n_330, n_206);
  nand g138 (n_331, n_204, n_205);
  nand g139 (n_332, n_206, n_205);
  nand g140 (n_333, n_204, n_206);
  nand g141 (n_162, n_331, n_332, n_333);
  xor g142 (n_334, in_0[5], in_1[5]);
  xor g143 (n_208, n_334, in_3[5]);
  nand g144 (n_335, in_0[5], in_1[5]);
  nand g145 (n_336, in_3[5], in_1[5]);
  nand g146 (n_337, in_0[5], in_3[5]);
  nand g147 (n_211, n_335, n_336, n_337);
  xor g148 (n_338, in_4[5], in_2[5]);
  xor g149 (n_209, n_338, n_207);
  nand g150 (n_339, in_4[5], in_2[5]);
  nand g151 (n_340, n_207, in_2[5]);
  nand g152 (n_341, in_4[5], n_207);
  nand g153 (n_214, n_339, n_340, n_341);
  xor g154 (n_342, n_208, n_209);
  xor g155 (n_188, n_342, n_210);
  nand g156 (n_343, n_208, n_209);
  nand g157 (n_344, n_210, n_209);
  nand g158 (n_345, n_208, n_210);
  nand g159 (n_161, n_343, n_344, n_345);
  xor g160 (n_346, in_0[6], in_1[6]);
  xor g161 (n_212, n_346, in_3[6]);
  nand g162 (n_347, in_0[6], in_1[6]);
  nand g163 (n_348, in_3[6], in_1[6]);
  nand g164 (n_349, in_0[6], in_3[6]);
  nand g165 (n_215, n_347, n_348, n_349);
  xor g166 (n_350, in_4[6], in_2[6]);
  xor g167 (n_213, n_350, n_211);
  nand g168 (n_351, in_4[6], in_2[6]);
  nand g169 (n_352, n_211, in_2[6]);
  nand g170 (n_353, in_4[6], n_211);
  nand g171 (n_218, n_351, n_352, n_353);
  xor g172 (n_354, n_212, n_213);
  xor g173 (n_187, n_354, n_214);
  nand g174 (n_355, n_212, n_213);
  nand g175 (n_356, n_214, n_213);
  nand g176 (n_357, n_212, n_214);
  nand g177 (n_160, n_355, n_356, n_357);
  xor g178 (n_358, in_0[7], in_1[7]);
  xor g179 (n_216, n_358, in_3[7]);
  nand g180 (n_359, in_0[7], in_1[7]);
  nand g181 (n_360, in_3[7], in_1[7]);
  nand g182 (n_361, in_0[7], in_3[7]);
  nand g183 (n_219, n_359, n_360, n_361);
  xor g184 (n_362, in_4[7], in_2[7]);
  xor g185 (n_217, n_362, n_215);
  nand g186 (n_363, in_4[7], in_2[7]);
  nand g187 (n_364, n_215, in_2[7]);
  nand g188 (n_365, in_4[7], n_215);
  nand g189 (n_222, n_363, n_364, n_365);
  xor g190 (n_366, n_216, n_217);
  xor g191 (n_186, n_366, n_218);
  nand g192 (n_367, n_216, n_217);
  nand g193 (n_368, n_218, n_217);
  nand g194 (n_369, n_216, n_218);
  nand g195 (n_159, n_367, n_368, n_369);
  xor g196 (n_370, in_0[8], in_1[8]);
  xor g197 (n_220, n_370, in_3[8]);
  nand g198 (n_371, in_0[8], in_1[8]);
  nand g199 (n_372, in_3[8], in_1[8]);
  nand g200 (n_373, in_0[8], in_3[8]);
  nand g201 (n_223, n_371, n_372, n_373);
  xor g202 (n_374, in_4[8], in_2[8]);
  xor g203 (n_221, n_374, n_219);
  nand g204 (n_375, in_4[8], in_2[8]);
  nand g205 (n_376, n_219, in_2[8]);
  nand g206 (n_377, in_4[8], n_219);
  nand g207 (n_226, n_375, n_376, n_377);
  xor g208 (n_378, n_220, n_221);
  xor g209 (n_185, n_378, n_222);
  nand g210 (n_379, n_220, n_221);
  nand g211 (n_380, n_222, n_221);
  nand g212 (n_381, n_220, n_222);
  nand g213 (n_158, n_379, n_380, n_381);
  xor g214 (n_382, in_0[9], in_1[9]);
  xor g215 (n_224, n_382, in_3[9]);
  nand g216 (n_383, in_0[9], in_1[9]);
  nand g217 (n_384, in_3[9], in_1[9]);
  nand g218 (n_385, in_0[9], in_3[9]);
  nand g219 (n_227, n_383, n_384, n_385);
  xor g220 (n_386, in_4[9], in_2[9]);
  xor g221 (n_225, n_386, n_223);
  nand g222 (n_387, in_4[9], in_2[9]);
  nand g223 (n_388, n_223, in_2[9]);
  nand g224 (n_389, in_4[9], n_223);
  nand g225 (n_230, n_387, n_388, n_389);
  xor g226 (n_390, n_224, n_225);
  xor g227 (n_184, n_390, n_226);
  nand g228 (n_391, n_224, n_225);
  nand g229 (n_392, n_226, n_225);
  nand g230 (n_393, n_224, n_226);
  nand g231 (n_157, n_391, n_392, n_393);
  xor g232 (n_394, in_0[10], in_1[10]);
  xor g233 (n_228, n_394, in_3[10]);
  nand g234 (n_395, in_0[10], in_1[10]);
  nand g235 (n_396, in_3[10], in_1[10]);
  nand g236 (n_397, in_0[10], in_3[10]);
  nand g237 (n_231, n_395, n_396, n_397);
  xor g238 (n_398, in_4[10], in_2[10]);
  xor g239 (n_229, n_398, n_227);
  nand g240 (n_399, in_4[10], in_2[10]);
  nand g241 (n_400, n_227, in_2[10]);
  nand g242 (n_401, in_4[10], n_227);
  nand g243 (n_234, n_399, n_400, n_401);
  xor g244 (n_402, n_228, n_229);
  xor g245 (n_183, n_402, n_230);
  nand g246 (n_403, n_228, n_229);
  nand g247 (n_404, n_230, n_229);
  nand g248 (n_405, n_228, n_230);
  nand g249 (n_156, n_403, n_404, n_405);
  xor g250 (n_406, in_0[11], in_1[11]);
  xor g251 (n_232, n_406, in_3[11]);
  nand g252 (n_407, in_0[11], in_1[11]);
  nand g253 (n_408, in_3[11], in_1[11]);
  nand g254 (n_409, in_0[11], in_3[11]);
  nand g255 (n_235, n_407, n_408, n_409);
  xor g256 (n_410, in_4[11], in_2[11]);
  xor g257 (n_233, n_410, n_231);
  nand g258 (n_411, in_4[11], in_2[11]);
  nand g259 (n_412, n_231, in_2[11]);
  nand g260 (n_413, in_4[11], n_231);
  nand g261 (n_238, n_411, n_412, n_413);
  xor g262 (n_414, n_232, n_233);
  xor g263 (n_182, n_414, n_234);
  nand g264 (n_415, n_232, n_233);
  nand g265 (n_416, n_234, n_233);
  nand g266 (n_417, n_232, n_234);
  nand g267 (n_155, n_415, n_416, n_417);
  xor g268 (n_418, in_0[12], in_1[12]);
  xor g269 (n_236, n_418, in_3[12]);
  nand g270 (n_419, in_0[12], in_1[12]);
  nand g271 (n_420, in_3[12], in_1[12]);
  nand g272 (n_421, in_0[12], in_3[12]);
  nand g273 (n_239, n_419, n_420, n_421);
  xor g274 (n_422, in_4[12], in_2[12]);
  xor g275 (n_237, n_422, n_235);
  nand g276 (n_423, in_4[12], in_2[12]);
  nand g277 (n_424, n_235, in_2[12]);
  nand g278 (n_425, in_4[12], n_235);
  nand g279 (n_242, n_423, n_424, n_425);
  xor g280 (n_426, n_236, n_237);
  xor g281 (n_181, n_426, n_238);
  nand g282 (n_427, n_236, n_237);
  nand g283 (n_428, n_238, n_237);
  nand g284 (n_429, n_236, n_238);
  nand g285 (n_154, n_427, n_428, n_429);
  xor g286 (n_430, in_0[13], in_1[13]);
  xor g287 (n_240, n_430, in_3[13]);
  nand g288 (n_431, in_0[13], in_1[13]);
  nand g289 (n_432, in_3[13], in_1[13]);
  nand g290 (n_433, in_0[13], in_3[13]);
  nand g291 (n_243, n_431, n_432, n_433);
  xor g292 (n_434, in_4[13], in_2[13]);
  xor g293 (n_241, n_434, n_239);
  nand g294 (n_435, in_4[13], in_2[13]);
  nand g295 (n_436, n_239, in_2[13]);
  nand g296 (n_437, in_4[13], n_239);
  nand g297 (n_246, n_435, n_436, n_437);
  xor g298 (n_438, n_240, n_241);
  xor g299 (n_180, n_438, n_242);
  nand g300 (n_439, n_240, n_241);
  nand g301 (n_440, n_242, n_241);
  nand g302 (n_441, n_240, n_242);
  nand g303 (n_153, n_439, n_440, n_441);
  xor g304 (n_442, in_0[14], in_1[14]);
  xor g305 (n_244, n_442, in_3[14]);
  nand g306 (n_443, in_0[14], in_1[14]);
  nand g307 (n_444, in_3[14], in_1[14]);
  nand g308 (n_445, in_0[14], in_3[14]);
  nand g309 (n_247, n_443, n_444, n_445);
  xor g310 (n_446, in_4[14], in_2[14]);
  xor g311 (n_245, n_446, n_243);
  nand g312 (n_447, in_4[14], in_2[14]);
  nand g313 (n_448, n_243, in_2[14]);
  nand g314 (n_449, in_4[14], n_243);
  nand g315 (n_250, n_447, n_448, n_449);
  xor g316 (n_450, n_244, n_245);
  xor g317 (n_179, n_450, n_246);
  nand g318 (n_451, n_244, n_245);
  nand g319 (n_452, n_246, n_245);
  nand g320 (n_453, n_244, n_246);
  nand g321 (n_152, n_451, n_452, n_453);
  xor g322 (n_454, in_0[15], in_1[15]);
  xor g323 (n_248, n_454, in_3[15]);
  nand g324 (n_455, in_0[15], in_1[15]);
  nand g325 (n_456, in_3[15], in_1[15]);
  nand g326 (n_457, in_0[15], in_3[15]);
  nand g327 (n_251, n_455, n_456, n_457);
  xor g328 (n_458, in_4[15], in_2[15]);
  xor g329 (n_249, n_458, n_247);
  nand g330 (n_459, in_4[15], in_2[15]);
  nand g331 (n_460, n_247, in_2[15]);
  nand g332 (n_461, in_4[15], n_247);
  nand g333 (n_254, n_459, n_460, n_461);
  xor g334 (n_462, n_248, n_249);
  xor g335 (n_178, n_462, n_250);
  nand g336 (n_463, n_248, n_249);
  nand g337 (n_464, n_250, n_249);
  nand g338 (n_465, n_248, n_250);
  nand g339 (n_151, n_463, n_464, n_465);
  xor g340 (n_466, in_0[16], in_1[16]);
  xor g341 (n_252, n_466, in_3[16]);
  nand g342 (n_467, in_0[16], in_1[16]);
  nand g343 (n_468, in_3[16], in_1[16]);
  nand g344 (n_469, in_0[16], in_3[16]);
  nand g345 (n_255, n_467, n_468, n_469);
  xor g346 (n_470, in_4[16], in_2[16]);
  xor g347 (n_253, n_470, n_251);
  nand g348 (n_471, in_4[16], in_2[16]);
  nand g349 (n_472, n_251, in_2[16]);
  nand g350 (n_473, in_4[16], n_251);
  nand g351 (n_258, n_471, n_472, n_473);
  xor g352 (n_474, n_252, n_253);
  xor g353 (n_177, n_474, n_254);
  nand g354 (n_475, n_252, n_253);
  nand g355 (n_476, n_254, n_253);
  nand g356 (n_477, n_252, n_254);
  nand g357 (n_150, n_475, n_476, n_477);
  xor g358 (n_478, in_0[17], in_1[17]);
  xor g359 (n_256, n_478, in_3[17]);
  nand g360 (n_479, in_0[17], in_1[17]);
  nand g361 (n_480, in_3[17], in_1[17]);
  nand g362 (n_481, in_0[17], in_3[17]);
  nand g363 (n_259, n_479, n_480, n_481);
  xor g364 (n_482, in_4[17], in_2[17]);
  xor g365 (n_257, n_482, n_255);
  nand g366 (n_483, in_4[17], in_2[17]);
  nand g367 (n_484, n_255, in_2[17]);
  nand g368 (n_485, in_4[17], n_255);
  nand g369 (n_262, n_483, n_484, n_485);
  xor g370 (n_486, n_256, n_257);
  xor g371 (n_176, n_486, n_258);
  nand g372 (n_487, n_256, n_257);
  nand g373 (n_488, n_258, n_257);
  nand g374 (n_489, n_256, n_258);
  nand g375 (n_149, n_487, n_488, n_489);
  xor g376 (n_490, in_0[18], in_1[18]);
  xor g377 (n_260, n_490, in_3[18]);
  nand g378 (n_491, in_0[18], in_1[18]);
  nand g379 (n_492, in_3[18], in_1[18]);
  nand g380 (n_493, in_0[18], in_3[18]);
  nand g381 (n_263, n_491, n_492, n_493);
  xor g382 (n_494, in_4[18], in_2[18]);
  xor g383 (n_261, n_494, n_259);
  nand g384 (n_495, in_4[18], in_2[18]);
  nand g385 (n_496, n_259, in_2[18]);
  nand g386 (n_497, in_4[18], n_259);
  nand g387 (n_266, n_495, n_496, n_497);
  xor g388 (n_498, n_260, n_261);
  xor g389 (n_175, n_498, n_262);
  nand g390 (n_499, n_260, n_261);
  nand g391 (n_500, n_262, n_261);
  nand g392 (n_501, n_260, n_262);
  nand g393 (n_148, n_499, n_500, n_501);
  xor g394 (n_502, in_0[19], in_1[19]);
  xor g395 (n_264, n_502, in_3[19]);
  nand g396 (n_503, in_0[19], in_1[19]);
  nand g397 (n_504, in_3[19], in_1[19]);
  nand g398 (n_505, in_0[19], in_3[19]);
  nand g399 (n_267, n_503, n_504, n_505);
  xor g400 (n_506, in_4[19], in_2[19]);
  xor g401 (n_265, n_506, n_263);
  nand g402 (n_507, in_4[19], in_2[19]);
  nand g403 (n_508, n_263, in_2[19]);
  nand g404 (n_509, in_4[19], n_263);
  nand g405 (n_270, n_507, n_508, n_509);
  xor g406 (n_510, n_264, n_265);
  xor g407 (n_174, n_510, n_266);
  nand g408 (n_511, n_264, n_265);
  nand g409 (n_512, n_266, n_265);
  nand g410 (n_513, n_264, n_266);
  nand g411 (n_147, n_511, n_512, n_513);
  xor g412 (n_514, in_0[20], in_1[20]);
  xor g413 (n_268, n_514, in_3[20]);
  nand g414 (n_515, in_0[20], in_1[20]);
  nand g415 (n_516, in_3[20], in_1[20]);
  nand g416 (n_517, in_0[20], in_3[20]);
  nand g417 (n_271, n_515, n_516, n_517);
  xor g418 (n_518, in_4[20], in_2[20]);
  xor g419 (n_269, n_518, n_267);
  nand g420 (n_519, in_4[20], in_2[20]);
  nand g421 (n_520, n_267, in_2[20]);
  nand g422 (n_521, in_4[20], n_267);
  nand g423 (n_274, n_519, n_520, n_521);
  xor g424 (n_522, n_268, n_269);
  xor g425 (n_173, n_522, n_270);
  nand g426 (n_523, n_268, n_269);
  nand g427 (n_524, n_270, n_269);
  nand g428 (n_525, n_268, n_270);
  nand g429 (n_146, n_523, n_524, n_525);
  xor g430 (n_526, in_0[21], in_1[21]);
  xor g431 (n_272, n_526, in_3[21]);
  nand g432 (n_527, in_0[21], in_1[21]);
  nand g433 (n_528, in_3[21], in_1[21]);
  nand g434 (n_529, in_0[21], in_3[21]);
  nand g435 (n_281, n_527, n_528, n_529);
  xor g436 (n_530, in_4[21], in_2[21]);
  xor g437 (n_273, n_530, n_271);
  nand g438 (n_531, in_4[21], in_2[21]);
  nand g439 (n_532, n_271, in_2[21]);
  nand g440 (n_533, in_4[21], n_271);
  nand g441 (n_284, n_531, n_532, n_533);
  xor g442 (n_534, n_272, n_273);
  xor g443 (n_172, n_534, n_274);
  nand g444 (n_535, n_272, n_273);
  nand g445 (n_536, n_274, n_273);
  nand g446 (n_537, n_272, n_274);
  nand g447 (n_145, n_535, n_536, n_537);
  nand g455 (n_287, n_539, n_540, n_541);
  nand g459 (n_544, n_281, n_280);
  xor g462 (n_546, n_282, n_283);
  xor g463 (n_171, n_546, n_284);
  nand g464 (n_547, n_282, n_283);
  nand g465 (n_548, n_284, n_283);
  nand g466 (n_549, n_282, n_284);
  nand g467 (n_144, n_547, n_548, n_549);
  xor g471 (n_170, n_550, n_289);
  nand g474 (n_553, n_287, n_289);
  nand g475 (n_169, n_551, n_552, n_553);
  xor g478 (n_841, in_1[0], n_193);
  nand g479 (n_556, in_1[0], n_193);
  nand g480 (n_557, in_1[0], in_2[0]);
  nand g7 (n_558, n_193, in_2[0]);
  nand g8 (n_560, n_556, n_557, n_558);
  nor g9 (n_559, n_166, n_192);
  nand g10 (n_562, n_166, n_192);
  nor g11 (n_569, n_165, n_191);
  nand g12 (n_564, n_165, n_191);
  nor g13 (n_565, n_164, n_190);
  nand g14 (n_566, n_164, n_190);
  nor g15 (n_575, n_163, n_189);
  nand g16 (n_570, n_163, n_189);
  nor g17 (n_571, n_162, n_188);
  nand g18 (n_572, n_162, n_188);
  nor g19 (n_581, n_161, n_187);
  nand g20 (n_576, n_161, n_187);
  nor g21 (n_577, n_160, n_186);
  nand g22 (n_578, n_160, n_186);
  nor g23 (n_587, n_159, n_185);
  nand g24 (n_582, n_159, n_185);
  nor g25 (n_583, n_158, n_184);
  nand g26 (n_584, n_158, n_184);
  nor g27 (n_593, n_157, n_183);
  nand g28 (n_588, n_157, n_183);
  nor g29 (n_589, n_156, n_182);
  nand g30 (n_590, n_156, n_182);
  nor g31 (n_599, n_155, n_181);
  nand g32 (n_594, n_155, n_181);
  nor g33 (n_595, n_154, n_180);
  nand g34 (n_596, n_154, n_180);
  nor g35 (n_605, n_153, n_179);
  nand g36 (n_600, n_153, n_179);
  nor g37 (n_601, n_152, n_178);
  nand g38 (n_602, n_152, n_178);
  nor g39 (n_611, n_151, n_177);
  nand g40 (n_606, n_151, n_177);
  nor g41 (n_607, n_150, n_176);
  nand g42 (n_608, n_150, n_176);
  nor g43 (n_617, n_149, n_175);
  nand g44 (n_612, n_149, n_175);
  nor g45 (n_613, n_148, n_174);
  nand g46 (n_614, n_148, n_174);
  nor g47 (n_623, n_147, n_173);
  nand g48 (n_618, n_147, n_173);
  nor g49 (n_619, n_146, n_172);
  nand g50 (n_620, n_146, n_172);
  nor g51 (n_629, n_145, n_171);
  nand g52 (n_624, n_145, n_171);
  nor g53 (n_625, n_144, n_170);
  nand g54 (n_626, n_144, n_170);
  nor g55 (n_633, n_143, n_169);
  nand g56 (n_630, n_143, n_169);
  nand g61 (n_634, n_562, n_563);
  nor g62 (n_567, n_564, n_565);
  nor g65 (n_167, n_569, n_565);
  nor g66 (n_573, n_570, n_571);
  nor g69 (n_642, n_575, n_571);
  nor g70 (n_579, n_576, n_577);
  nor g73 (n_644, n_581, n_577);
  nor g74 (n_585, n_582, n_583);
  nor g483 (n_652, n_587, n_583);
  nor g484 (n_591, n_588, n_589);
  nor g487 (n_654, n_593, n_589);
  nor g488 (n_597, n_594, n_595);
  nor g491 (n_662, n_599, n_595);
  nor g492 (n_603, n_600, n_601);
  nor g495 (n_664, n_605, n_601);
  nor g496 (n_609, n_606, n_607);
  nor g499 (n_672, n_611, n_607);
  nor g500 (n_615, n_612, n_613);
  nor g503 (n_674, n_617, n_613);
  nor g504 (n_621, n_618, n_619);
  nor g507 (n_682, n_623, n_619);
  nor g508 (n_627, n_624, n_625);
  nor g511 (n_684, n_629, n_625);
  nand g514 (n_785, n_564, n_636);
  nand g515 (n_638, n_167, n_634);
  nand g516 (n_689, n_637, n_638);
  nor g517 (n_640, n_581, n_639);
  nand g526 (n_697, n_642, n_644);
  nor g527 (n_650, n_593, n_649);
  nand g536 (n_704, n_652, n_654);
  nor g537 (n_660, n_605, n_659);
  nand g546 (n_712, n_662, n_664);
  nor g547 (n_670, n_617, n_669);
  nand g556 (n_719, n_672, n_674);
  nor g557 (n_680, n_629, n_679);
  nand g566 (n_727, n_682, n_684);
  nand g569 (n_789, n_570, n_691);
  nand g570 (n_692, n_642, n_689);
  nand g571 (n_791, n_639, n_692);
  nand g574 (n_794, n_695, n_696);
  nand g577 (n_731, n_699, n_700);
  nor g578 (n_702, n_599, n_701);
  nor g581 (n_741, n_599, n_704);
  nor g587 (n_710, n_708, n_701);
  nor g590 (n_747, n_704, n_708);
  nor g591 (n_714, n_712, n_701);
  nor g594 (n_750, n_704, n_712);
  nor g595 (n_717, n_623, n_716);
  nor g598 (n_768, n_623, n_719);
  nor g604 (n_725, n_723, n_716);
  nor g607 (n_774, n_719, n_723);
  nor g608 (n_729, n_727, n_716);
  nor g611 (n_756, n_719, n_727);
  nand g614 (n_798, n_582, n_733);
  nand g615 (n_734, n_652, n_731);
  nand g616 (n_800, n_649, n_734);
  nand g619 (n_803, n_737, n_738);
  nand g622 (n_806, n_701, n_740);
  nand g623 (n_743, n_741, n_731);
  nand g624 (n_809, n_742, n_743);
  nand g625 (n_746, n_744, n_731);
  nand g626 (n_811, n_745, n_746);
  nand g627 (n_749, n_747, n_731);
  nand g628 (n_814, n_748, n_749);
  nand g629 (n_752, n_750, n_731);
  nand g630 (n_758, n_751, n_752);
  nor g631 (n_754, n_633, n_753);
  nand g638 (n_818, n_606, n_760);
  nand g639 (n_761, n_672, n_758);
  nand g640 (n_820, n_669, n_761);
  nand g643 (n_823, n_764, n_765);
  nand g646 (n_826, n_716, n_767);
  nand g647 (n_770, n_768, n_758);
  nand g648 (n_829, n_769, n_770);
  nand g649 (n_773, n_771, n_758);
  nand g650 (n_831, n_772, n_773);
  nand g651 (n_776, n_774, n_758);
  nand g652 (n_834, n_775, n_776);
  nand g653 (n_777, n_756, n_758);
  nand g654 (n_836, n_753, n_777);
  nand g657 (n_839, n_780, n_781);
  xnor g659 (out_0[1], n_560, n_782);
  xnor g661 (out_0[2], n_634, n_783);
  xnor g664 (out_0[3], n_785, n_786);
  xnor g666 (out_0[4], n_689, n_787);
  xnor g669 (out_0[5], n_789, n_790);
  xnor g671 (out_0[6], n_791, n_792);
  xnor g674 (out_0[7], n_794, n_795);
  xnor g676 (out_0[8], n_731, n_796);
  xnor g679 (out_0[9], n_798, n_799);
  xnor g681 (out_0[10], n_800, n_801);
  xnor g684 (out_0[11], n_803, n_804);
  xnor g687 (out_0[12], n_806, n_807);
  xnor g690 (out_0[13], n_809, n_810);
  xnor g692 (out_0[14], n_811, n_812);
  xnor g695 (out_0[15], n_814, n_815);
  xnor g697 (out_0[16], n_758, n_816);
  xnor g700 (out_0[17], n_818, n_819);
  xnor g702 (out_0[18], n_820, n_821);
  xnor g705 (out_0[19], n_823, n_824);
  xnor g708 (out_0[20], n_826, n_827);
  xnor g711 (out_0[21], n_829, n_830);
  xnor g713 (out_0[22], n_831, n_832);
  xnor g716 (out_0[23], n_834, n_835);
  xnor g718 (out_0[24], n_836, n_837);
  xor g722 (out_0[0], in_2[0], n_841);
  xor g723 (n_280, in_0[22], in_1[22]);
  nor g724 (n_143, in_0[22], in_1[22]);
  xor g725 (n_538, in_3[22], in_4[22]);
  or g726 (n_539, in_3[22], in_4[22]);
  or g727 (n_540, in_2[22], in_4[22]);
  or g728 (n_541, in_2[22], in_3[22]);
  xnor g729 (n_282, n_538, in_2[22]);
  xnor g733 (n_283, n_281, n_280);
  or g734 (n_289, n_280, wc, n_281);
  not gc (wc, n_544);
  xnor g735 (n_550, n_287, n_143);
  or g736 (n_551, n_143, wc0);
  not gc0 (wc0, n_287);
  or g737 (n_552, wc1, n_143);
  not gc1 (wc1, n_289);
  or g738 (n_563, n_559, wc2);
  not gc2 (wc2, n_560);
  or g739 (n_782, wc3, n_559);
  not gc3 (wc3, n_562);
  and g740 (n_637, wc4, n_566);
  not gc4 (wc4, n_567);
  or g741 (n_783, wc5, n_569);
  not gc5 (wc5, n_564);
  or g742 (n_786, wc6, n_565);
  not gc6 (wc6, n_566);
  and g743 (n_639, wc7, n_572);
  not gc7 (wc7, n_573);
  or g744 (n_636, wc8, n_569);
  not gc8 (wc8, n_634);
  or g745 (n_787, wc9, n_575);
  not gc9 (wc9, n_570);
  or g746 (n_790, wc10, n_571);
  not gc10 (wc10, n_572);
  and g747 (n_646, wc11, n_578);
  not gc11 (wc11, n_579);
  and g748 (n_649, wc12, n_584);
  not gc12 (wc12, n_585);
  and g749 (n_656, wc13, n_590);
  not gc13 (wc13, n_591);
  and g750 (n_659, wc14, n_596);
  not gc14 (wc14, n_597);
  and g751 (n_666, wc15, n_602);
  not gc15 (wc15, n_603);
  and g752 (n_669, wc16, n_608);
  not gc16 (wc16, n_609);
  and g753 (n_676, wc17, n_614);
  not gc17 (wc17, n_615);
  and g754 (n_679, wc18, n_620);
  not gc18 (wc18, n_621);
  and g755 (n_686, wc19, n_626);
  not gc19 (wc19, n_627);
  or g756 (n_693, wc20, n_581);
  not gc20 (wc20, n_642);
  or g757 (n_735, wc21, n_593);
  not gc21 (wc21, n_652);
  or g758 (n_708, wc22, n_605);
  not gc22 (wc22, n_662);
  or g759 (n_762, wc23, n_617);
  not gc23 (wc23, n_672);
  or g760 (n_723, wc24, n_629);
  not gc24 (wc24, n_682);
  or g761 (n_792, wc25, n_581);
  not gc25 (wc25, n_576);
  or g762 (n_795, wc26, n_577);
  not gc26 (wc26, n_578);
  or g763 (n_796, wc27, n_587);
  not gc27 (wc27, n_582);
  or g764 (n_799, wc28, n_583);
  not gc28 (wc28, n_584);
  or g765 (n_801, wc29, n_593);
  not gc29 (wc29, n_588);
  or g766 (n_804, wc30, n_589);
  not gc30 (wc30, n_590);
  or g767 (n_807, wc31, n_599);
  not gc31 (wc31, n_594);
  or g768 (n_810, wc32, n_595);
  not gc32 (wc32, n_596);
  or g769 (n_812, wc33, n_605);
  not gc33 (wc33, n_600);
  or g770 (n_815, wc34, n_601);
  not gc34 (wc34, n_602);
  or g771 (n_816, wc35, n_611);
  not gc35 (wc35, n_606);
  or g772 (n_819, wc36, n_607);
  not gc36 (wc36, n_608);
  or g773 (n_821, wc37, n_617);
  not gc37 (wc37, n_612);
  or g774 (n_824, wc38, n_613);
  not gc38 (wc38, n_614);
  or g775 (n_827, wc39, n_623);
  not gc39 (wc39, n_618);
  or g776 (n_830, wc40, n_619);
  not gc40 (wc40, n_620);
  or g777 (n_832, wc41, n_629);
  not gc41 (wc41, n_624);
  or g778 (n_835, wc42, n_625);
  not gc42 (wc42, n_626);
  or g779 (n_837, wc43, n_633);
  not gc43 (wc43, n_630);
  and g780 (n_695, wc44, n_576);
  not gc44 (wc44, n_640);
  and g781 (n_647, wc45, n_644);
  not gc45 (wc45, n_639);
  and g782 (n_657, wc46, n_654);
  not gc46 (wc46, n_649);
  and g783 (n_667, wc47, n_664);
  not gc47 (wc47, n_659);
  and g784 (n_677, wc48, n_674);
  not gc48 (wc48, n_669);
  and g785 (n_687, wc49, n_684);
  not gc49 (wc49, n_679);
  or g786 (n_691, wc50, n_575);
  not gc50 (wc50, n_689);
  and g787 (n_744, wc51, n_662);
  not gc51 (wc51, n_704);
  and g788 (n_771, wc52, n_682);
  not gc52 (wc52, n_719);
  and g789 (n_699, wc53, n_646);
  not gc53 (wc53, n_647);
  and g790 (n_737, wc54, n_588);
  not gc54 (wc54, n_650);
  and g791 (n_701, wc55, n_656);
  not gc55 (wc55, n_657);
  and g792 (n_709, wc56, n_600);
  not gc56 (wc56, n_660);
  and g793 (n_713, wc57, n_666);
  not gc57 (wc57, n_667);
  and g794 (n_764, wc58, n_612);
  not gc58 (wc58, n_670);
  and g795 (n_716, wc59, n_676);
  not gc59 (wc59, n_677);
  and g796 (n_724, wc60, n_624);
  not gc60 (wc60, n_680);
  and g797 (n_728, wc61, n_686);
  not gc61 (wc61, n_687);
  or g798 (n_696, n_693, wc62);
  not gc62 (wc62, n_689);
  or g799 (n_700, n_697, wc63);
  not gc63 (wc63, n_689);
  or g800 (n_778, wc64, n_633);
  not gc64 (wc64, n_756);
  and g801 (n_706, wc65, n_662);
  not gc65 (wc65, n_701);
  and g802 (n_721, wc66, n_682);
  not gc66 (wc66, n_716);
  and g803 (n_742, wc67, n_594);
  not gc67 (wc67, n_702);
  and g804 (n_745, wc68, n_659);
  not gc68 (wc68, n_706);
  and g805 (n_748, n_709, wc69);
  not gc69 (wc69, n_710);
  and g806 (n_751, n_713, wc70);
  not gc70 (wc70, n_714);
  and g807 (n_769, wc71, n_618);
  not gc71 (wc71, n_717);
  and g808 (n_772, wc72, n_679);
  not gc72 (wc72, n_721);
  and g809 (n_775, n_724, wc73);
  not gc73 (wc73, n_725);
  and g810 (n_753, n_728, wc74);
  not gc74 (wc74, n_729);
  or g811 (n_733, wc75, n_587);
  not gc75 (wc75, n_731);
  or g812 (n_738, n_735, wc76);
  not gc76 (wc76, n_731);
  or g813 (n_740, wc77, n_704);
  not gc77 (wc77, n_731);
  and g814 (n_780, wc78, n_630);
  not gc78 (wc78, n_754);
  or g815 (n_760, wc79, n_611);
  not gc79 (wc79, n_758);
  or g816 (n_765, n_762, wc80);
  not gc80 (wc80, n_758);
  or g817 (n_767, wc81, n_719);
  not gc81 (wc81, n_758);
  or g818 (n_781, n_778, wc82);
  not gc82 (wc82, n_758);
  not g819 (out_0[25], n_839);
endmodule

module csa_tree_add_915_44_group_6805_GENERIC(in_0, in_1, in_2, in_3,
     in_4, out_0);
  input [22:0] in_0, in_1, in_2, in_3, in_4;
  output [25:0] out_0;
  wire [22:0] in_0, in_1, in_2, in_3, in_4;
  wire [25:0] out_0;
  csa_tree_add_915_44_group_6805_GENERIC_REAL g1(.in_0 (in_0), .in_1
       (in_1), .in_2 (in_2), .in_3 (in_3), .in_4 (in_4), .out_0
       (out_0));
endmodule

module mult_signed_const_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_119, n_171, n_172, n_173, n_174, n_181;
  wire n_182, n_184, n_185, n_186, n_190, n_191, n_196, n_197;
  wire n_198, n_204, n_205, n_206, n_210, n_211, n_212, n_213;
  wire n_214, n_218, n_220, n_221, n_226, n_227, n_228, n_229;
  wire n_235, n_237, n_238, n_239, n_240, n_241, n_246, n_247;
  wire n_248, n_249, n_250, n_251, n_252, n_253, n_259, n_260;
  wire n_261, n_262, n_263, n_264, n_267, n_269, n_271, n_272;
  wire n_273, n_274, n_275, n_276, n_277, n_278, n_279, n_283;
  wire n_284, n_285, n_286, n_287, n_288, n_289, n_290, n_291;
  wire n_292, n_293, n_294, n_295, n_298, n_300, n_301, n_302;
  wire n_303, n_304, n_305, n_306, n_307, n_308, n_309, n_310;
  wire n_311, n_317, n_319, n_320, n_321, n_322, n_323, n_324;
  wire n_325, n_326, n_327, n_328, n_338, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_346, n_347, n_355, n_357, n_359;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_368;
  wire n_369, n_373, n_374, n_375, n_376, n_377, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_390, n_391, n_392, n_394, n_395, n_396;
  wire n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404;
  wire n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412;
  wire n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420;
  wire n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_431, n_432, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_450, n_451, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_469, n_470, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_505, n_506, n_507, n_508;
  wire n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516;
  wire n_517, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_530, n_531, n_532, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_555, n_556, n_559, n_560, n_561, n_562;
  wire n_563, n_564, n_565, n_566, n_567, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_577, n_578, n_580, n_581, n_582;
  wire n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590;
  wire n_591, n_592, n_593, n_594, n_597, n_598, n_599, n_600;
  wire n_601, n_605, n_606, n_607, n_608, n_610, n_611, n_612;
  wire n_613, n_614, n_615, n_616, n_619, n_624, n_625, n_626;
  wire n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634;
  wire n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_642;
  wire n_643, n_648, n_649, n_650, n_651, n_652, n_653, n_654;
  wire n_655, n_656, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_666, n_667, n_672, n_673, n_674, n_675, n_676, n_677;
  wire n_678, n_679, n_684, n_688, n_689, n_690, n_691, n_692;
  wire n_693, n_694, n_695, n_706, n_707, n_708, n_709, n_710;
  wire n_711, n_712, n_713, n_714, n_715, n_720, n_721, n_723;
  wire n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_734, n_735, n_744, n_745, n_746, n_747;
  wire n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755;
  wire n_768, n_769, n_770, n_772, n_773, n_774, n_775, n_776;
  wire n_777, n_778, n_779, n_790, n_791, n_792, n_793, n_794;
  wire n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802;
  wire n_803, n_804, n_805, n_806, n_807, n_818, n_820, n_821;
  wire n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829;
  wire n_830, n_831, n_832, n_833, n_834, n_835, n_844, n_845;
  wire n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855;
  wire n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_863;
  wire n_864, n_868, n_869, n_870, n_874, n_875, n_878, n_879;
  wire n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887;
  wire n_888, n_889, n_890, n_891, n_892, n_893, n_894, n_895;
  wire n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909;
  wire n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917;
  wire n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925;
  wire n_926, n_927, n_928, n_929, n_930, n_931, n_940, n_941;
  wire n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950;
  wire n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958;
  wire n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966;
  wire n_967, n_980, n_981, n_982, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_996, n_997, n_998, n_999, n_1000, n_1001, n_1002, n_1003;
  wire n_1024, n_1025, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040;
  wire n_1041, n_1042, n_1043, n_1045, n_1046, n_1049, n_1051, n_1053;
  wire n_1054, n_1055, n_1058, n_1059, n_1062, n_1063, n_1066, n_1067;
  wire n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077;
  wire n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085;
  wire n_1086, n_1087, n_1088, n_1090, n_1092, n_1093, n_1094, n_1095;
  wire n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103;
  wire n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111;
  wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119;
  wire n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127;
  wire n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135;
  wire n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143;
  wire n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151;
  wire n_1152, n_1153, n_1154, n_1156, n_1157, n_1158, n_1159, n_1160;
  wire n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168;
  wire n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176;
  wire n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1184, n_1185;
  wire n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193;
  wire n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201;
  wire n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209;
  wire n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217;
  wire n_1218, n_1219, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227;
  wire n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235;
  wire n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243;
  wire n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251;
  wire n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1260;
  wire n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1268, n_1269;
  wire n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
  wire n_1278, n_1279, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287;
  wire n_1288, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298;
  wire n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306;
  wire n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314;
  wire n_1315, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1326;
  wire n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334;
  wire n_1335, n_1336, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343;
  wire n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351;
  wire n_1352, n_1353, n_1354, n_1355, n_1357, n_1358, n_1359, n_1360;
  wire n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368;
  wire n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1378;
  wire n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386;
  wire n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394;
  wire n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402;
  wire n_1403, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1414;
  wire n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422;
  wire n_1423, n_1424, n_1425, n_1426, n_1428, n_1429, n_1430, n_1431;
  wire n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1442, n_1443;
  wire n_1444, n_1445, n_1446, n_1448, n_1449, n_1450, n_1451, n_1452;
  wire n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460;
  wire n_1461, n_1462, n_1463, n_1465, n_1466, n_1467, n_1468, n_1470;
  wire n_1471, n_1472, n_1473, n_1474, n_1475, n_1478, n_1479, n_1480;
  wire n_1481, n_1482, n_1483, n_1486, n_1488, n_1489, n_1490, n_1491;
  wire n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1500;
  wire n_1501, n_1502, n_1503, n_1504, n_1506, n_1508, n_1509, n_1510;
  wire n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518;
  wire n_1519, n_1520, n_1521, n_1522, n_1523, n_1526, n_1527, n_1528;
  wire n_1529, n_1530, n_1531, n_1534, n_1535, n_1536, n_1537, n_1538;
  wire n_1539, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1548;
  wire n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556;
  wire n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564;
  wire n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575;
  wire n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583;
  wire n_1585, n_1586, n_1587, n_1588, n_1590, n_1591, n_1608, n_1613;
  wire n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621;
  wire n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629;
  wire n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637;
  wire n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645;
  wire n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653;
  wire n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661;
  wire n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669;
  wire n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677;
  wire n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685;
  wire n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693;
  wire n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701;
  wire n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709;
  wire n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717;
  wire n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725;
  wire n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733;
  wire n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741;
  wire n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749;
  wire n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757;
  wire n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765;
  wire n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773;
  wire n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781;
  wire n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789;
  wire n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797;
  wire n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805;
  wire n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813;
  wire n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821;
  wire n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829;
  wire n_1830, n_1831, n_1832, n_1833;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_70, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_624, A[1], n_171);
  xor g270 (n_69, n_624, A[2]);
  nand g3 (n_625, A[1], n_171);
  nand g271 (n_626, A[2], n_171);
  nand g272 (n_627, A[1], A[2]);
  nand g273 (n_172, n_625, n_626, n_627);
  xor g274 (n_628, A[2], n_172);
  xor g275 (n_116, n_628, A[3]);
  nand g276 (n_629, A[2], n_172);
  nand g4 (n_630, A[3], n_172);
  nand g277 (n_631, A[2], A[3]);
  nand g278 (n_174, n_629, n_630, n_631);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_71, A[0], A[3]);
  xor g281 (n_632, A[4], n_173);
  xor g282 (n_115, n_632, n_174);
  nand g283 (n_633, A[4], n_173);
  nand g284 (n_634, n_174, n_173);
  nand g5 (n_635, A[4], n_174);
  nand g6 (n_72, n_633, n_634, n_635);
  xor g287 (n_636, n_70, n_71);
  xor g288 (n_73, n_636, A[4]);
  nand g289 (n_637, n_70, n_71);
  nand g290 (n_638, A[4], n_71);
  nand g291 (n_639, n_70, A[4]);
  nand g292 (n_181, n_637, n_638, n_639);
  xor g293 (n_640, A[5], n_73);
  xor g294 (n_114, n_640, n_72);
  nand g295 (n_641, A[5], n_73);
  nand g296 (n_642, n_72, n_73);
  nand g297 (n_643, A[5], n_72);
  nand g298 (n_65, n_641, n_642, n_643);
  xor g305 (n_648, n_69, A[5]);
  xor g306 (n_182, n_648, n_181);
  nand g307 (n_649, n_69, A[5]);
  nand g308 (n_650, n_181, A[5]);
  nand g309 (n_651, n_69, n_181);
  nand g310 (n_185, n_649, n_650, n_651);
  xor g311 (n_652, A[6], n_182);
  xor g312 (n_113, n_652, A[8]);
  nand g313 (n_653, A[6], n_182);
  nand g314 (n_654, A[8], n_182);
  nand g315 (n_655, A[6], A[8]);
  nand g316 (n_64, n_653, n_654, n_655);
  xor g317 (n_656, A[2], A[3]);
  xor g318 (n_184, n_656, n_172);
  xor g323 (n_660, n_184, A[6]);
  xor g324 (n_186, n_660, A[7]);
  nand g325 (n_661, n_184, A[6]);
  nand g326 (n_662, A[7], A[6]);
  nand g327 (n_663, n_184, A[7]);
  nand g328 (n_190, n_661, n_662, n_663);
  xor g329 (n_664, n_185, n_186);
  xor g330 (n_112, n_664, A[9]);
  nand g331 (n_665, n_185, n_186);
  nand g332 (n_666, A[9], n_186);
  nand g333 (n_667, n_185, A[9]);
  nand g334 (n_63, n_665, n_666, n_667);
  xor g343 (n_672, A[7], n_115);
  xor g344 (n_191, n_672, A[8]);
  nand g345 (n_673, A[7], n_115);
  nand g346 (n_674, A[8], n_115);
  nand g347 (n_675, A[7], A[8]);
  nand g348 (n_197, n_673, n_674, n_675);
  xor g349 (n_676, n_190, A[10]);
  xor g350 (n_111, n_676, n_191);
  nand g351 (n_677, n_190, A[10]);
  nand g352 (n_678, n_191, A[10]);
  nand g353 (n_679, n_190, n_191);
  nand g354 (n_62, n_677, n_678, n_679);
  xor g363 (n_684, A[5], n_72);
  xor g364 (n_196, n_684, n_73);
  xor g369 (n_688, A[8], A[9]);
  xor g370 (n_198, n_688, n_196);
  nand g371 (n_689, A[8], A[9]);
  nand g372 (n_690, n_196, A[9]);
  nand g373 (n_691, A[8], n_196);
  nand g374 (n_205, n_689, n_690, n_691);
  xor g375 (n_692, A[11], n_197);
  xor g376 (n_110, n_692, n_198);
  nand g377 (n_693, A[11], n_197);
  nand g378 (n_694, n_198, n_197);
  nand g379 (n_695, A[11], n_198);
  nand g380 (n_61, n_693, n_694, n_695);
  xor g394 (n_204, n_652, A[9]);
  nand g396 (n_706, A[9], n_182);
  nand g397 (n_707, A[6], A[9]);
  nand g398 (n_211, n_653, n_706, n_707);
  xor g399 (n_708, n_65, A[10]);
  xor g400 (n_206, n_708, n_204);
  nand g401 (n_709, n_65, A[10]);
  nand g402 (n_710, n_204, A[10]);
  nand g403 (n_711, n_65, n_204);
  nand g404 (n_213, n_709, n_710, n_711);
  xor g405 (n_712, A[12], n_205);
  xor g406 (n_109, n_712, n_206);
  nand g407 (n_713, A[12], n_205);
  nand g408 (n_714, n_206, n_205);
  nand g409 (n_715, A[12], n_206);
  nand g410 (n_60, n_713, n_714, n_715);
  xor g417 (n_720, n_116, A[6]);
  xor g418 (n_210, n_720, A[7]);
  nand g419 (n_721, n_116, A[6]);
  nand g421 (n_723, n_116, A[7]);
  nand g422 (n_218, n_721, n_662, n_723);
  xor g423 (n_724, n_185, n_210);
  xor g424 (n_212, n_724, A[10]);
  nand g425 (n_725, n_185, n_210);
  nand g426 (n_726, A[10], n_210);
  nand g427 (n_727, n_185, A[10]);
  nand g428 (n_220, n_725, n_726, n_727);
  xor g429 (n_728, A[11], n_211);
  xor g430 (n_214, n_728, n_212);
  nand g431 (n_729, A[11], n_211);
  nand g432 (n_730, n_212, n_211);
  nand g433 (n_731, A[11], n_212);
  nand g434 (n_68, n_729, n_730, n_731);
  xor g435 (n_732, A[13], n_213);
  xor g436 (n_108, n_732, n_214);
  nand g437 (n_733, A[13], n_213);
  nand g438 (n_734, n_214, n_213);
  nand g439 (n_735, A[13], n_214);
  nand g440 (n_59, n_733, n_734, n_735);
  xor g455 (n_744, n_218, n_191);
  xor g456 (n_66, n_744, A[11]);
  nand g457 (n_745, n_218, n_191);
  nand g458 (n_746, A[11], n_191);
  nand g459 (n_747, n_218, A[11]);
  nand g460 (n_226, n_745, n_746, n_747);
  xor g461 (n_748, n_220, A[12]);
  xor g462 (n_221, n_748, n_66);
  nand g463 (n_749, n_220, A[12]);
  nand g464 (n_750, n_66, A[12]);
  nand g465 (n_751, n_220, n_66);
  nand g466 (n_228, n_749, n_750, n_751);
  xor g467 (n_752, A[14], n_68);
  xor g468 (n_107, n_752, n_221);
  nand g469 (n_753, A[14], n_68);
  nand g470 (n_754, n_221, n_68);
  nand g471 (n_755, A[14], n_221);
  nand g472 (n_58, n_753, n_754, n_755);
  xor g493 (n_768, n_197, A[12]);
  xor g494 (n_227, n_768, n_198);
  nand g495 (n_769, n_197, A[12]);
  nand g496 (n_770, n_198, A[12]);
  nand g498 (n_238, n_769, n_770, n_694);
  xor g499 (n_772, A[13], n_226);
  xor g500 (n_229, n_772, A[15]);
  nand g501 (n_773, A[13], n_226);
  nand g502 (n_774, A[15], n_226);
  nand g503 (n_775, A[13], A[15]);
  nand g504 (n_240, n_773, n_774, n_775);
  xor g505 (n_776, n_227, n_228);
  xor g506 (n_106, n_776, n_229);
  nand g507 (n_777, n_227, n_228);
  nand g508 (n_778, n_229, n_228);
  nand g509 (n_779, n_227, n_229);
  nand g510 (n_57, n_777, n_778, n_779);
  xor g524 (n_235, n_652, n_65);
  nand g526 (n_790, n_65, n_182);
  nand g527 (n_791, A[6], n_65);
  nand g528 (n_246, n_653, n_790, n_791);
  xor g529 (n_792, A[9], A[10]);
  xor g530 (n_237, n_792, n_235);
  nand g531 (n_793, A[9], A[10]);
  nand g532 (n_794, n_235, A[10]);
  nand g533 (n_795, A[9], n_235);
  nand g534 (n_248, n_793, n_794, n_795);
  xor g535 (n_796, n_205, A[13]);
  xor g536 (n_239, n_796, n_237);
  nand g537 (n_797, n_205, A[13]);
  nand g538 (n_798, n_237, A[13]);
  nand g539 (n_799, n_205, n_237);
  nand g540 (n_250, n_797, n_798, n_799);
  xor g541 (n_800, A[14], n_238);
  xor g542 (n_241, n_800, A[16]);
  nand g543 (n_801, A[14], n_238);
  nand g544 (n_802, A[16], n_238);
  nand g545 (n_803, A[14], A[16]);
  nand g546 (n_252, n_801, n_802, n_803);
  xor g547 (n_804, n_239, n_240);
  xor g548 (n_105, n_804, n_241);
  nand g549 (n_805, n_239, n_240);
  nand g550 (n_806, n_241, n_240);
  nand g551 (n_807, n_239, n_241);
  nand g552 (n_56, n_805, n_806, n_807);
  xor g566 (n_247, n_664, A[10]);
  nand g568 (n_818, A[10], n_186);
  nand g570 (n_259, n_665, n_818, n_727);
  xor g571 (n_820, A[11], n_246);
  xor g572 (n_249, n_820, n_247);
  nand g573 (n_821, A[11], n_246);
  nand g574 (n_822, n_247, n_246);
  nand g575 (n_823, A[11], n_247);
  nand g576 (n_261, n_821, n_822, n_823);
  xor g577 (n_824, n_248, A[14]);
  xor g578 (n_251, n_824, n_249);
  nand g579 (n_825, n_248, A[14]);
  nand g580 (n_826, n_249, A[14]);
  nand g581 (n_827, n_248, n_249);
  nand g582 (n_117, n_825, n_826, n_827);
  xor g583 (n_828, A[15], n_250);
  xor g584 (n_253, n_828, A[17]);
  nand g585 (n_829, A[15], n_250);
  nand g586 (n_830, A[17], n_250);
  nand g587 (n_831, A[15], A[17]);
  nand g588 (n_263, n_829, n_830, n_831);
  xor g589 (n_832, n_251, n_252);
  xor g590 (n_104, n_832, n_253);
  nand g591 (n_833, n_251, n_252);
  nand g592 (n_834, n_253, n_252);
  nand g593 (n_835, n_251, n_253);
  nand g594 (n_55, n_833, n_834, n_835);
  xor g609 (n_844, n_190, A[11]);
  xor g610 (n_260, n_844, n_191);
  nand g611 (n_845, n_190, A[11]);
  nand g614 (n_272, n_845, n_746, n_679);
  xor g615 (n_848, A[12], n_259);
  xor g616 (n_262, n_848, n_260);
  nand g617 (n_849, A[12], n_259);
  nand g618 (n_850, n_260, n_259);
  nand g619 (n_851, A[12], n_260);
  nand g620 (n_274, n_849, n_850, n_851);
  xor g621 (n_852, n_261, A[15]);
  xor g622 (n_119, n_852, n_262);
  nand g623 (n_853, n_261, A[15]);
  nand g624 (n_854, n_262, A[15]);
  nand g625 (n_855, n_261, n_262);
  nand g626 (n_276, n_853, n_854, n_855);
  xor g627 (n_856, A[16], n_117);
  xor g628 (n_264, n_856, A[18]);
  nand g629 (n_857, A[16], n_117);
  nand g630 (n_858, A[18], n_117);
  nand g631 (n_859, A[16], A[18]);
  nand g632 (n_278, n_857, n_858, n_859);
  xor g633 (n_860, n_119, n_263);
  xor g634 (n_103, n_860, n_264);
  nand g635 (n_861, n_119, n_263);
  nand g636 (n_862, n_264, n_263);
  nand g637 (n_863, n_119, n_264);
  nand g638 (n_54, n_861, n_862, n_863);
  xor g641 (n_864, n_70, A[4]);
  xor g642 (n_267, n_864, n_71);
  xor g647 (n_868, A[5], n_267);
  xor g648 (n_269, n_868, n_72);
  nand g649 (n_869, A[5], n_267);
  nand g650 (n_870, n_72, n_267);
  nand g652 (n_284, n_869, n_870, n_643);
  xor g654 (n_271, n_688, n_269);
  nand g656 (n_874, n_269, A[9]);
  nand g657 (n_875, A[8], n_269);
  nand g658 (n_286, n_689, n_874, n_875);
  xor g660 (n_273, n_768, n_271);
  nand g662 (n_878, n_271, A[12]);
  nand g663 (n_879, n_197, n_271);
  nand g664 (n_288, n_769, n_878, n_879);
  xor g665 (n_880, A[13], n_272);
  xor g666 (n_275, n_880, n_273);
  nand g667 (n_881, A[13], n_272);
  nand g668 (n_882, n_273, n_272);
  nand g669 (n_883, A[13], n_273);
  nand g670 (n_290, n_881, n_882, n_883);
  xor g671 (n_884, n_274, A[16]);
  xor g672 (n_277, n_884, A[17]);
  nand g673 (n_885, n_274, A[16]);
  nand g674 (n_886, A[17], A[16]);
  nand g675 (n_887, n_274, A[17]);
  nand g676 (n_292, n_885, n_886, n_887);
  xor g677 (n_888, n_275, n_276);
  xor g678 (n_279, n_888, A[19]);
  nand g679 (n_889, n_275, n_276);
  nand g680 (n_890, A[19], n_276);
  nand g681 (n_891, n_275, A[19]);
  nand g682 (n_294, n_889, n_890, n_891);
  xor g683 (n_892, n_277, n_278);
  xor g684 (n_102, n_892, n_279);
  nand g685 (n_893, n_277, n_278);
  nand g686 (n_894, n_279, n_278);
  nand g687 (n_895, n_277, n_279);
  nand g688 (n_53, n_893, n_894, n_895);
  xor g696 (n_283, n_648, A[6]);
  nand g698 (n_902, A[6], A[5]);
  nand g699 (n_903, n_69, A[6]);
  nand g700 (n_298, n_649, n_902, n_903);
  xor g701 (n_904, n_181, n_283);
  xor g702 (n_285, n_904, A[9]);
  nand g703 (n_905, n_181, n_283);
  nand g704 (n_906, A[9], n_283);
  nand g705 (n_907, n_181, A[9]);
  nand g706 (n_300, n_905, n_906, n_907);
  xor g707 (n_908, n_284, A[10]);
  xor g708 (n_287, n_908, n_285);
  nand g709 (n_909, n_284, A[10]);
  nand g710 (n_910, n_285, A[10]);
  nand g711 (n_911, n_284, n_285);
  nand g712 (n_302, n_909, n_910, n_911);
  xor g713 (n_912, n_286, A[13]);
  xor g714 (n_289, n_912, n_287);
  nand g715 (n_913, n_286, A[13]);
  nand g716 (n_914, n_287, A[13]);
  nand g717 (n_915, n_286, n_287);
  nand g718 (n_304, n_913, n_914, n_915);
  xor g719 (n_916, n_288, A[14]);
  xor g720 (n_291, n_916, n_289);
  nand g721 (n_917, n_288, A[14]);
  nand g722 (n_918, n_289, A[14]);
  nand g723 (n_919, n_288, n_289);
  nand g724 (n_306, n_917, n_918, n_919);
  xor g725 (n_920, n_290, A[17]);
  xor g726 (n_293, n_920, n_291);
  nand g727 (n_921, n_290, A[17]);
  nand g728 (n_922, n_291, A[17]);
  nand g729 (n_923, n_290, n_291);
  nand g730 (n_308, n_921, n_922, n_923);
  xor g731 (n_924, A[18], n_292);
  xor g732 (n_295, n_924, A[20]);
  nand g733 (n_925, A[18], n_292);
  nand g734 (n_926, A[20], n_292);
  nand g735 (n_927, A[18], A[20]);
  nand g736 (n_310, n_925, n_926, n_927);
  xor g737 (n_928, n_293, n_294);
  xor g738 (n_101, n_928, n_295);
  nand g739 (n_929, n_293, n_294);
  nand g740 (n_930, n_295, n_294);
  nand g741 (n_931, n_293, n_295);
  nand g742 (n_52, n_929, n_930, n_931);
  xor g755 (n_940, n_298, n_186);
  xor g756 (n_301, n_940, A[10]);
  nand g757 (n_941, n_298, n_186);
  nand g759 (n_943, n_298, A[10]);
  nand g760 (n_317, n_941, n_818, n_943);
  xor g761 (n_944, A[11], n_300);
  xor g762 (n_303, n_944, n_301);
  nand g763 (n_945, A[11], n_300);
  nand g764 (n_946, n_301, n_300);
  nand g765 (n_947, A[11], n_301);
  nand g766 (n_319, n_945, n_946, n_947);
  xor g767 (n_948, n_302, A[14]);
  xor g768 (n_305, n_948, n_303);
  nand g769 (n_949, n_302, A[14]);
  nand g770 (n_950, n_303, A[14]);
  nand g771 (n_951, n_302, n_303);
  nand g772 (n_321, n_949, n_950, n_951);
  xor g773 (n_952, A[15], n_304);
  xor g774 (n_307, n_952, n_305);
  nand g775 (n_953, A[15], n_304);
  nand g776 (n_954, n_305, n_304);
  nand g777 (n_955, A[15], n_305);
  nand g778 (n_323, n_953, n_954, n_955);
  xor g779 (n_956, n_306, A[18]);
  xor g780 (n_309, n_956, n_307);
  nand g781 (n_957, n_306, A[18]);
  nand g782 (n_958, n_307, A[18]);
  nand g783 (n_959, n_306, n_307);
  nand g784 (n_325, n_957, n_958, n_959);
  xor g785 (n_960, A[19], n_308);
  xor g786 (n_311, n_960, n_309);
  nand g787 (n_961, A[19], n_308);
  nand g788 (n_962, n_309, n_308);
  nand g789 (n_963, A[19], n_309);
  nand g790 (n_327, n_961, n_962, n_963);
  xor g791 (n_964, n_310, A[21]);
  xor g792 (n_100, n_964, n_311);
  nand g793 (n_965, n_310, A[21]);
  nand g794 (n_966, n_311, A[21]);
  nand g795 (n_967, n_310, n_311);
  nand g796 (n_51, n_965, n_966, n_967);
  xor g817 (n_980, A[12], n_317);
  xor g818 (n_320, n_980, n_260);
  nand g819 (n_981, A[12], n_317);
  nand g820 (n_982, n_260, n_317);
  nand g822 (n_338, n_981, n_982, n_851);
  xor g823 (n_984, n_319, A[15]);
  xor g824 (n_322, n_984, A[16]);
  nand g825 (n_985, n_319, A[15]);
  nand g826 (n_986, A[16], A[15]);
  nand g827 (n_987, n_319, A[16]);
  nand g828 (n_340, n_985, n_986, n_987);
  xor g829 (n_988, n_320, n_321);
  xor g830 (n_324, n_988, n_322);
  nand g831 (n_989, n_320, n_321);
  nand g832 (n_990, n_322, n_321);
  nand g833 (n_991, n_320, n_322);
  nand g834 (n_342, n_989, n_990, n_991);
  xor g835 (n_992, n_323, A[19]);
  xor g836 (n_326, n_992, n_324);
  nand g837 (n_993, n_323, A[19]);
  nand g838 (n_994, n_324, A[19]);
  nand g839 (n_995, n_323, n_324);
  nand g840 (n_344, n_993, n_994, n_995);
  xor g841 (n_996, A[20], n_325);
  xor g842 (n_328, n_996, n_326);
  nand g843 (n_997, A[20], n_325);
  nand g844 (n_998, n_326, n_325);
  nand g845 (n_999, A[20], n_326);
  nand g846 (n_346, n_997, n_998, n_999);
  xor g847 (n_1000, A[22], n_327);
  xor g848 (n_99, n_1000, n_328);
  nand g849 (n_1001, A[22], n_327);
  nand g850 (n_1002, n_328, n_327);
  nand g851 (n_1003, A[22], n_328);
  nand g852 (n_50, n_1001, n_1002, n_1003);
  xor g885 (n_1024, n_338, A[16]);
  xor g886 (n_341, n_1024, A[17]);
  nand g887 (n_1025, n_338, A[16]);
  nand g889 (n_1027, n_338, A[17]);
  nand g890 (n_362, n_1025, n_886, n_1027);
  xor g891 (n_1028, n_275, n_340);
  xor g892 (n_343, n_1028, n_341);
  nand g893 (n_1029, n_275, n_340);
  nand g894 (n_1030, n_341, n_340);
  nand g895 (n_1031, n_275, n_341);
  nand g896 (n_364, n_1029, n_1030, n_1031);
  xor g897 (n_1032, n_342, A[20]);
  xor g898 (n_345, n_1032, n_343);
  nand g899 (n_1033, n_342, A[20]);
  nand g900 (n_1034, n_343, A[20]);
  nand g901 (n_1035, n_342, n_343);
  nand g902 (n_366, n_1033, n_1034, n_1035);
  xor g903 (n_1036, n_344, A[21]);
  xor g904 (n_347, n_1036, A[23]);
  nand g905 (n_1037, n_344, A[21]);
  nand g906 (n_1038, A[23], A[21]);
  nand g907 (n_1039, n_344, A[23]);
  nand g908 (n_368, n_1037, n_1038, n_1039);
  xor g909 (n_1040, n_345, n_346);
  xor g910 (n_98, n_1040, n_347);
  nand g911 (n_1041, n_345, n_346);
  nand g912 (n_1042, n_347, n_346);
  nand g913 (n_1043, n_345, n_347);
  nand g914 (n_49, n_1041, n_1042, n_1043);
  nand g922 (n_373, n_1045, n_1046, n_626);
  nand g928 (n_375, n_1049, n_650, n_1051);
  nand g933 (n_1055, A[6], n_284);
  nand g934 (n_377, n_1053, n_1054, n_1055);
  xor g936 (n_357, n_792, n_355);
  nand g938 (n_1058, n_355, A[10]);
  nand g939 (n_1059, A[9], n_355);
  nand g940 (n_379, n_793, n_1058, n_1059);
  xor g942 (n_359, n_912, n_357);
  nand g944 (n_1062, n_357, A[13]);
  nand g945 (n_1063, n_286, n_357);
  nand g946 (n_381, n_913, n_1062, n_1063);
  xor g948 (n_361, n_916, n_359);
  nand g950 (n_1066, n_359, A[14]);
  nand g951 (n_1067, n_288, n_359);
  nand g952 (n_383, n_917, n_1066, n_1067);
  xor g954 (n_363, n_920, A[18]);
  nand g956 (n_1070, A[18], A[17]);
  nand g957 (n_1071, n_290, A[18]);
  nand g958 (n_385, n_921, n_1070, n_1071);
  xor g959 (n_1072, n_361, n_362);
  xor g960 (n_365, n_1072, n_363);
  nand g961 (n_1073, n_361, n_362);
  nand g962 (n_1074, n_363, n_362);
  nand g963 (n_1075, n_361, n_363);
  nand g964 (n_388, n_1073, n_1074, n_1075);
  xor g965 (n_1076, n_364, A[21]);
  xor g966 (n_367, n_1076, n_365);
  nand g967 (n_1077, n_364, A[21]);
  nand g968 (n_1078, n_365, A[21]);
  nand g969 (n_1079, n_364, n_365);
  nand g970 (n_389, n_1077, n_1078, n_1079);
  xor g971 (n_1080, A[22], n_366);
  nand g973 (n_1081, A[22], n_366);
  nand g976 (n_391, n_1081, n_1082, n_1083);
  xor g977 (n_1084, n_367, n_368);
  xor g978 (n_97, n_1084, n_369);
  nand g979 (n_1085, n_367, n_368);
  nand g980 (n_1086, n_369, n_368);
  nand g981 (n_1087, n_367, n_369);
  nand g982 (n_48, n_1085, n_1086, n_1087);
  xor g986 (n_374, n_1088, A[3]);
  nand g990 (n_394, n_1046, n_1090, n_631);
  xor g991 (n_1092, n_373, n_374);
  xor g992 (n_376, n_1092, A[6]);
  nand g993 (n_1093, n_373, n_374);
  nand g994 (n_1094, A[6], n_374);
  nand g995 (n_1095, n_373, A[6]);
  nand g996 (n_396, n_1093, n_1094, n_1095);
  xor g997 (n_1096, A[7], n_375);
  xor g998 (n_378, n_1096, n_376);
  nand g999 (n_1097, A[7], n_375);
  nand g1000 (n_1098, n_376, n_375);
  nand g1001 (n_1099, A[7], n_376);
  nand g1002 (n_398, n_1097, n_1098, n_1099);
  xor g1003 (n_1100, A[10], A[11]);
  xor g1004 (n_380, n_1100, n_377);
  nand g1005 (n_1101, A[10], A[11]);
  nand g1006 (n_1102, n_377, A[11]);
  nand g1007 (n_1103, A[10], n_377);
  nand g1008 (n_400, n_1101, n_1102, n_1103);
  xor g1009 (n_1104, n_378, n_379);
  xor g1010 (n_382, n_1104, n_380);
  nand g1011 (n_1105, n_378, n_379);
  nand g1012 (n_1106, n_380, n_379);
  nand g1013 (n_1107, n_378, n_380);
  nand g1014 (n_402, n_1105, n_1106, n_1107);
  xor g1015 (n_1108, A[14], A[15]);
  xor g1016 (n_384, n_1108, n_381);
  nand g1017 (n_1109, A[14], A[15]);
  nand g1018 (n_1110, n_381, A[15]);
  nand g1019 (n_1111, A[14], n_381);
  nand g1020 (n_404, n_1109, n_1110, n_1111);
  xor g1021 (n_1112, n_382, A[18]);
  xor g1022 (n_386, n_1112, n_383);
  nand g1023 (n_1113, n_382, A[18]);
  nand g1024 (n_1114, n_383, A[18]);
  nand g1025 (n_1115, n_382, n_383);
  nand g1026 (n_406, n_1113, n_1114, n_1115);
  xor g1027 (n_1116, n_384, A[19]);
  xor g1028 (n_387, n_1116, n_385);
  nand g1029 (n_1117, n_384, A[19]);
  nand g1030 (n_1118, n_385, A[19]);
  nand g1031 (n_1119, n_384, n_385);
  nand g1032 (n_408, n_1117, n_1118, n_1119);
  xor g1033 (n_1120, n_386, n_387);
  xor g1034 (n_390, n_1120, n_388);
  nand g1035 (n_1121, n_386, n_387);
  nand g1036 (n_1122, n_388, n_387);
  nand g1037 (n_1123, n_386, n_388);
  nand g1038 (n_410, n_1121, n_1122, n_1123);
  xor g1039 (n_1124, A[22], A[23]);
  xor g1040 (n_392, n_1124, n_389);
  nand g1041 (n_1125, A[22], A[23]);
  nand g1042 (n_1126, n_389, A[23]);
  nand g1043 (n_1127, A[22], n_389);
  nand g1044 (n_413, n_1125, n_1126, n_1127);
  xor g1045 (n_1128, n_390, n_391);
  xor g1046 (n_96, n_1128, n_392);
  nand g1047 (n_1129, n_390, n_391);
  nand g1048 (n_1130, n_392, n_391);
  nand g1049 (n_1131, n_390, n_392);
  nand g1050 (n_47, n_1129, n_1130, n_1131);
  xor g1051 (n_1132, A[1], A[3]);
  xor g1052 (n_395, n_1132, A[4]);
  nand g1053 (n_1133, A[1], A[3]);
  nand g1054 (n_1134, A[4], A[3]);
  nand g1055 (n_1135, A[1], A[4]);
  nand g1056 (n_414, n_1133, n_1134, n_1135);
  xor g1057 (n_1136, n_394, n_395);
  xor g1058 (n_397, n_1136, A[7]);
  nand g1059 (n_1137, n_394, n_395);
  nand g1060 (n_1138, A[7], n_395);
  nand g1061 (n_1139, n_394, A[7]);
  nand g1062 (n_416, n_1137, n_1138, n_1139);
  xor g1063 (n_1140, A[8], n_396);
  xor g1064 (n_399, n_1140, n_397);
  nand g1065 (n_1141, A[8], n_396);
  nand g1066 (n_1142, n_397, n_396);
  nand g1067 (n_1143, A[8], n_397);
  nand g1068 (n_418, n_1141, n_1142, n_1143);
  xor g1069 (n_1144, n_398, A[11]);
  xor g1070 (n_401, n_1144, n_399);
  nand g1071 (n_1145, n_398, A[11]);
  nand g1072 (n_1146, n_399, A[11]);
  nand g1073 (n_1147, n_398, n_399);
  nand g1074 (n_419, n_1145, n_1146, n_1147);
  xor g1075 (n_1148, A[12], n_400);
  xor g1076 (n_403, n_1148, n_401);
  nand g1077 (n_1149, A[12], n_400);
  nand g1078 (n_1150, n_401, n_400);
  nand g1079 (n_1151, A[12], n_401);
  nand g1080 (n_421, n_1149, n_1150, n_1151);
  xor g1081 (n_1152, A[15], n_402);
  xor g1082 (n_405, n_1152, A[16]);
  nand g1083 (n_1153, A[15], n_402);
  nand g1084 (n_1154, A[16], n_402);
  nand g1086 (n_423, n_1153, n_1154, n_986);
  xor g1087 (n_1156, n_403, n_404);
  xor g1088 (n_407, n_1156, n_405);
  nand g1089 (n_1157, n_403, n_404);
  nand g1090 (n_1158, n_405, n_404);
  nand g1091 (n_1159, n_403, n_405);
  nand g1092 (n_426, n_1157, n_1158, n_1159);
  xor g1093 (n_1160, A[19], n_406);
  xor g1094 (n_409, n_1160, A[20]);
  nand g1095 (n_1161, A[19], n_406);
  nand g1096 (n_1162, A[20], n_406);
  nand g1097 (n_1163, A[19], A[20]);
  nand g1098 (n_427, n_1161, n_1162, n_1163);
  xor g1099 (n_1164, n_407, n_408);
  xor g1100 (n_411, n_1164, n_409);
  nand g1101 (n_1165, n_407, n_408);
  nand g1102 (n_1166, n_409, n_408);
  nand g1103 (n_1167, n_407, n_409);
  nand g1104 (n_429, n_1165, n_1166, n_1167);
  xor g1106 (n_412, n_1168, n_410);
  nand g1109 (n_1171, A[23], n_410);
  nand g1110 (n_431, n_1169, n_1170, n_1171);
  xor g1111 (n_1172, n_411, n_412);
  xor g1112 (n_95, n_1172, n_413);
  nand g1113 (n_1173, n_411, n_412);
  nand g1114 (n_1174, n_413, n_412);
  nand g1115 (n_1175, n_411, n_413);
  nand g1116 (n_46, n_1173, n_1174, n_1175);
  xor g1117 (n_1176, A[4], A[5]);
  xor g1118 (n_415, n_1176, n_414);
  nand g1119 (n_1177, A[4], A[5]);
  nand g1120 (n_1178, n_414, A[5]);
  nand g1121 (n_1179, A[4], n_414);
  nand g1122 (n_435, n_1177, n_1178, n_1179);
  xor g1123 (n_1180, A[8], n_415);
  xor g1124 (n_417, n_1180, A[9]);
  nand g1125 (n_1181, A[8], n_415);
  nand g1126 (n_1182, A[9], n_415);
  nand g1128 (n_437, n_1181, n_1182, n_689);
  xor g1129 (n_1184, n_416, n_417);
  xor g1130 (n_420, n_1184, n_418);
  nand g1131 (n_1185, n_416, n_417);
  nand g1132 (n_1186, n_418, n_417);
  nand g1133 (n_1187, n_416, n_418);
  nand g1134 (n_439, n_1185, n_1186, n_1187);
  xor g1135 (n_1188, A[12], A[13]);
  xor g1136 (n_422, n_1188, n_419);
  nand g1137 (n_1189, A[12], A[13]);
  nand g1138 (n_1190, n_419, A[13]);
  nand g1139 (n_1191, A[12], n_419);
  nand g1140 (n_441, n_1189, n_1190, n_1191);
  xor g1141 (n_1192, n_420, n_421);
  xor g1142 (n_424, n_1192, A[16]);
  nand g1143 (n_1193, n_420, n_421);
  nand g1144 (n_1194, A[16], n_421);
  nand g1145 (n_1195, n_420, A[16]);
  nand g1146 (n_442, n_1193, n_1194, n_1195);
  xor g1147 (n_1196, n_422, A[17]);
  xor g1148 (n_425, n_1196, n_423);
  nand g1149 (n_1197, n_422, A[17]);
  nand g1150 (n_1198, n_423, A[17]);
  nand g1151 (n_1199, n_422, n_423);
  nand g1152 (n_444, n_1197, n_1198, n_1199);
  xor g1153 (n_1200, n_424, A[20]);
  xor g1154 (n_428, n_1200, n_425);
  nand g1155 (n_1201, n_424, A[20]);
  nand g1156 (n_1202, n_425, A[20]);
  nand g1157 (n_1203, n_424, n_425);
  nand g1158 (n_446, n_1201, n_1202, n_1203);
  xor g1159 (n_1204, n_426, n_427);
  xor g1160 (n_430, n_1204, A[21]);
  nand g1161 (n_1205, n_426, n_427);
  nand g1162 (n_1206, A[21], n_427);
  nand g1163 (n_1207, n_426, A[21]);
  nand g1164 (n_448, n_1205, n_1206, n_1207);
  xor g1166 (n_432, n_1208, n_429);
  nand g1169 (n_1211, n_428, n_429);
  nand g1170 (n_451, n_1209, n_1210, n_1211);
  xor g1171 (n_1212, n_430, n_431);
  xor g1172 (n_94, n_1212, n_432);
  nand g1173 (n_1213, n_430, n_431);
  nand g1174 (n_1214, n_432, n_431);
  nand g1175 (n_1215, n_430, n_432);
  nand g1176 (n_45, n_1213, n_1214, n_1215);
  xor g1180 (n_436, n_1216, n_435);
  nand g1183 (n_1219, A[6], n_435);
  nand g1184 (n_456, n_1217, n_1218, n_1219);
  xor g1186 (n_438, n_792, n_436);
  nand g1188 (n_1222, n_436, A[10]);
  nand g1189 (n_1223, A[9], n_436);
  nand g1190 (n_458, n_793, n_1222, n_1223);
  xor g1191 (n_1224, n_437, n_438);
  xor g1192 (n_440, n_1224, A[13]);
  nand g1193 (n_1225, n_437, n_438);
  nand g1194 (n_1226, A[13], n_438);
  nand g1195 (n_1227, n_437, A[13]);
  nand g1196 (n_459, n_1225, n_1226, n_1227);
  xor g1197 (n_1228, n_439, A[14]);
  xor g1198 (n_443, n_1228, n_440);
  nand g1199 (n_1229, n_439, A[14]);
  nand g1200 (n_1230, n_440, A[14]);
  nand g1201 (n_1231, n_439, n_440);
  nand g1202 (n_461, n_1229, n_1230, n_1231);
  xor g1203 (n_1232, n_441, A[17]);
  xor g1204 (n_445, n_1232, n_442);
  nand g1205 (n_1233, n_441, A[17]);
  nand g1206 (n_1234, n_442, A[17]);
  nand g1207 (n_1235, n_441, n_442);
  nand g1208 (n_463, n_1233, n_1234, n_1235);
  xor g1209 (n_1236, A[18], n_443);
  xor g1210 (n_447, n_1236, n_444);
  nand g1211 (n_1237, A[18], n_443);
  nand g1212 (n_1238, n_444, n_443);
  nand g1213 (n_1239, A[18], n_444);
  nand g1214 (n_465, n_1237, n_1238, n_1239);
  xor g1215 (n_1240, n_445, n_446);
  xor g1216 (n_449, n_1240, n_447);
  nand g1217 (n_1241, n_445, n_446);
  nand g1218 (n_1242, n_447, n_446);
  nand g1219 (n_1243, n_445, n_447);
  nand g1220 (n_467, n_1241, n_1242, n_1243);
  xor g1221 (n_1244, A[21], A[22]);
  xor g1222 (n_450, n_1244, n_448);
  nand g1223 (n_1245, A[21], A[22]);
  nand g1224 (n_1246, n_448, A[22]);
  nand g1225 (n_1247, A[21], n_448);
  nand g1226 (n_470, n_1245, n_1246, n_1247);
  xor g1227 (n_1248, n_449, n_450);
  xor g1228 (n_93, n_1248, n_451);
  nand g1229 (n_1249, n_449, n_450);
  nand g1230 (n_1250, n_451, n_450);
  nand g1231 (n_1251, n_449, n_451);
  nand g1232 (n_44, n_1249, n_1250, n_1251);
  xor g1235 (n_1252, A[5], A[7]);
  nand g1237 (n_1253, A[5], A[7]);
  nand g1240 (n_472, n_1253, n_1254, n_1255);
  xor g1241 (n_1256, A[10], n_455);
  xor g1242 (n_457, n_1256, A[11]);
  nand g1243 (n_1257, A[10], n_455);
  nand g1244 (n_1258, A[11], n_455);
  nand g1246 (n_474, n_1257, n_1258, n_1101);
  xor g1247 (n_1260, n_456, n_457);
  xor g1248 (n_460, n_1260, n_458);
  nand g1249 (n_1261, n_456, n_457);
  nand g1250 (n_1262, n_458, n_457);
  nand g1251 (n_1263, n_456, n_458);
  nand g1252 (n_476, n_1261, n_1262, n_1263);
  xor g1253 (n_1264, A[14], n_459);
  xor g1254 (n_462, n_1264, A[15]);
  nand g1255 (n_1265, A[14], n_459);
  nand g1256 (n_1266, A[15], n_459);
  nand g1258 (n_478, n_1265, n_1266, n_1109);
  xor g1259 (n_1268, n_460, A[18]);
  xor g1260 (n_464, n_1268, n_461);
  nand g1261 (n_1269, n_460, A[18]);
  nand g1262 (n_1270, n_461, A[18]);
  nand g1263 (n_1271, n_460, n_461);
  nand g1264 (n_481, n_1269, n_1270, n_1271);
  xor g1265 (n_1272, n_462, A[19]);
  xor g1266 (n_466, n_1272, n_463);
  nand g1267 (n_1273, n_462, A[19]);
  nand g1268 (n_1274, n_463, A[19]);
  nand g1269 (n_1275, n_462, n_463);
  nand g1270 (n_482, n_1273, n_1274, n_1275);
  xor g1271 (n_1276, n_464, n_465);
  xor g1272 (n_468, n_1276, n_466);
  nand g1273 (n_1277, n_464, n_465);
  nand g1274 (n_1278, n_466, n_465);
  nand g1275 (n_1279, n_464, n_466);
  nand g1276 (n_484, n_1277, n_1278, n_1279);
  xor g1278 (n_469, n_1124, n_467);
  nand g1280 (n_1282, n_467, A[23]);
  nand g1281 (n_1283, A[22], n_467);
  nand g1282 (n_487, n_1125, n_1282, n_1283);
  xor g1283 (n_1284, n_468, n_469);
  xor g1284 (n_92, n_1284, n_470);
  nand g1285 (n_1285, n_468, n_469);
  nand g1286 (n_1286, n_470, n_469);
  nand g1287 (n_1287, n_468, n_470);
  nand g1288 (n_43, n_1285, n_1286, n_1287);
  xor g1289 (n_1288, A[7], A[6]);
  xor g1290 (n_473, n_1288, A[8]);
  nand g1294 (n_488, n_662, n_655, n_675);
  xor g1295 (n_1292, n_472, A[11]);
  xor g1296 (n_475, n_1292, n_473);
  nand g1297 (n_1293, n_472, A[11]);
  nand g1298 (n_1294, n_473, A[11]);
  nand g1299 (n_1295, n_472, n_473);
  nand g1300 (n_489, n_1293, n_1294, n_1295);
  xor g1301 (n_1296, A[12], n_474);
  xor g1302 (n_477, n_1296, n_475);
  nand g1303 (n_1297, A[12], n_474);
  nand g1304 (n_1298, n_475, n_474);
  nand g1305 (n_1299, A[12], n_475);
  nand g1306 (n_492, n_1297, n_1298, n_1299);
  xor g1307 (n_1300, A[15], n_476);
  xor g1308 (n_479, n_1300, n_477);
  nand g1309 (n_1301, A[15], n_476);
  nand g1310 (n_1302, n_477, n_476);
  nand g1311 (n_1303, A[15], n_477);
  nand g1312 (n_493, n_1301, n_1302, n_1303);
  xor g1313 (n_1304, A[16], n_478);
  xor g1314 (n_480, n_1304, n_479);
  nand g1315 (n_1305, A[16], n_478);
  nand g1316 (n_1306, n_479, n_478);
  nand g1317 (n_1307, A[16], n_479);
  nand g1318 (n_496, n_1305, n_1306, n_1307);
  xor g1319 (n_1308, A[19], n_480);
  xor g1320 (n_483, n_1308, n_481);
  nand g1321 (n_1309, A[19], n_480);
  nand g1322 (n_1310, n_481, n_480);
  nand g1323 (n_1311, A[19], n_481);
  nand g1324 (n_497, n_1309, n_1310, n_1311);
  xor g1325 (n_1312, A[20], n_482);
  xor g1326 (n_485, n_1312, n_483);
  nand g1327 (n_1313, A[20], n_482);
  nand g1328 (n_1314, n_483, n_482);
  nand g1329 (n_1315, A[20], n_483);
  nand g1330 (n_500, n_1313, n_1314, n_1315);
  xor g1332 (n_486, n_1168, n_484);
  nand g1335 (n_1319, A[23], n_484);
  nand g1336 (n_501, n_1169, n_1318, n_1319);
  xor g1337 (n_1320, n_485, n_486);
  xor g1338 (n_91, n_1320, n_487);
  nand g1339 (n_1321, n_485, n_486);
  nand g1340 (n_1322, n_487, n_486);
  nand g1341 (n_1323, n_485, n_487);
  nand g1342 (n_42, n_1321, n_1322, n_1323);
  xor g1344 (n_490, n_688, n_488);
  nand g1346 (n_1326, n_488, A[9]);
  nand g1347 (n_1327, A[8], n_488);
  nand g1348 (n_505, n_689, n_1326, n_1327);
  xor g1349 (n_1328, A[12], n_489);
  xor g1350 (n_491, n_1328, n_490);
  nand g1351 (n_1329, A[12], n_489);
  nand g1352 (n_1330, n_490, n_489);
  nand g1353 (n_1331, A[12], n_490);
  nand g1354 (n_506, n_1329, n_1330, n_1331);
  xor g1355 (n_1332, A[13], n_491);
  xor g1356 (n_494, n_1332, n_492);
  nand g1357 (n_1333, A[13], n_491);
  nand g1358 (n_1334, n_492, n_491);
  nand g1359 (n_1335, A[13], n_492);
  nand g1360 (n_509, n_1333, n_1334, n_1335);
  xor g1361 (n_1336, A[16], A[17]);
  xor g1362 (n_495, n_1336, n_493);
  nand g1364 (n_1338, n_493, A[17]);
  nand g1365 (n_1339, A[16], n_493);
  nand g1366 (n_510, n_886, n_1338, n_1339);
  xor g1367 (n_1340, n_494, A[20]);
  xor g1368 (n_498, n_1340, n_495);
  nand g1369 (n_1341, n_494, A[20]);
  nand g1370 (n_1342, n_495, A[20]);
  nand g1371 (n_1343, n_494, n_495);
  nand g1372 (n_513, n_1341, n_1342, n_1343);
  xor g1373 (n_1344, n_496, n_497);
  xor g1374 (n_499, n_1344, A[21]);
  nand g1375 (n_1345, n_496, n_497);
  nand g1376 (n_1346, A[21], n_497);
  nand g1377 (n_1347, n_496, A[21]);
  nand g1378 (n_514, n_1345, n_1346, n_1347);
  xor g1380 (n_502, n_1348, n_499);
  nand g1383 (n_1351, n_498, n_499);
  nand g1384 (n_517, n_1349, n_1350, n_1351);
  xor g1385 (n_1352, n_500, n_501);
  xor g1386 (n_90, n_1352, n_502);
  nand g1387 (n_1353, n_500, n_501);
  nand g1388 (n_1354, n_502, n_501);
  nand g1389 (n_1355, n_500, n_502);
  nand g1390 (n_41, n_1353, n_1354, n_1355);
  nand g1397 (n_1359, A[10], n_505);
  nand g1398 (n_522, n_1357, n_1358, n_1359);
  xor g1399 (n_1360, A[13], A[14]);
  xor g1400 (n_508, n_1360, n_506);
  nand g1401 (n_1361, A[13], A[14]);
  nand g1402 (n_1362, n_506, A[14]);
  nand g1403 (n_1363, A[13], n_506);
  nand g1404 (n_523, n_1361, n_1362, n_1363);
  xor g1405 (n_1364, n_507, A[17]);
  xor g1406 (n_511, n_1364, n_508);
  nand g1407 (n_1365, n_507, A[17]);
  nand g1408 (n_1366, n_508, A[17]);
  nand g1409 (n_1367, n_507, n_508);
  nand g1410 (n_525, n_1365, n_1366, n_1367);
  xor g1411 (n_1368, A[18], n_509);
  xor g1412 (n_512, n_1368, n_510);
  nand g1413 (n_1369, A[18], n_509);
  nand g1414 (n_1370, n_510, n_509);
  nand g1415 (n_1371, A[18], n_510);
  nand g1416 (n_528, n_1369, n_1370, n_1371);
  xor g1417 (n_1372, n_511, n_512);
  xor g1418 (n_515, n_1372, n_513);
  nand g1419 (n_1373, n_511, n_512);
  nand g1420 (n_1374, n_513, n_512);
  nand g1421 (n_1375, n_511, n_513);
  nand g1422 (n_529, n_1373, n_1374, n_1375);
  xor g1424 (n_516, n_1244, n_514);
  nand g1426 (n_1378, n_514, A[22]);
  nand g1427 (n_1379, A[21], n_514);
  nand g1428 (n_532, n_1245, n_1378, n_1379);
  xor g1429 (n_1380, n_515, n_516);
  xor g1430 (n_89, n_1380, n_517);
  nand g1431 (n_1381, n_515, n_516);
  nand g1432 (n_1382, n_517, n_516);
  nand g1433 (n_1383, n_515, n_517);
  nand g1434 (n_40, n_1381, n_1382, n_1383);
  xor g1437 (n_1384, A[11], A[9]);
  nand g1439 (n_1385, A[11], A[9]);
  nand g1442 (n_534, n_1385, n_1386, n_1387);
  xor g1443 (n_1388, n_521, A[14]);
  xor g1444 (n_524, n_1388, n_522);
  nand g1445 (n_1389, n_521, A[14]);
  nand g1446 (n_1390, n_522, A[14]);
  nand g1447 (n_1391, n_521, n_522);
  nand g1448 (n_536, n_1389, n_1390, n_1391);
  xor g1449 (n_1392, A[15], n_523);
  xor g1450 (n_526, n_1392, n_524);
  nand g1451 (n_1393, A[15], n_523);
  nand g1452 (n_1394, n_524, n_523);
  nand g1453 (n_1395, A[15], n_524);
  nand g1454 (n_538, n_1393, n_1394, n_1395);
  xor g1455 (n_1396, A[18], n_525);
  xor g1456 (n_527, n_1396, A[19]);
  nand g1457 (n_1397, A[18], n_525);
  nand g1458 (n_1398, A[19], n_525);
  nand g1459 (n_1399, A[18], A[19]);
  nand g1460 (n_540, n_1397, n_1398, n_1399);
  xor g1461 (n_1400, n_526, n_527);
  xor g1462 (n_530, n_1400, n_528);
  nand g1463 (n_1401, n_526, n_527);
  nand g1464 (n_1402, n_528, n_527);
  nand g1465 (n_1403, n_526, n_528);
  nand g1466 (n_542, n_1401, n_1402, n_1403);
  xor g1468 (n_531, n_1124, n_529);
  nand g1470 (n_1406, n_529, A[23]);
  nand g1471 (n_1407, A[22], n_529);
  nand g1472 (n_545, n_1125, n_1406, n_1407);
  xor g1473 (n_1408, n_530, n_531);
  xor g1474 (n_88, n_1408, n_532);
  nand g1475 (n_1409, n_530, n_531);
  nand g1476 (n_1410, n_532, n_531);
  nand g1477 (n_1411, n_530, n_532);
  nand g1478 (n_39, n_1409, n_1410, n_1411);
  xor g1480 (n_535, n_1100, A[12]);
  nand g1482 (n_1414, A[12], A[10]);
  nand g1483 (n_1415, A[11], A[12]);
  nand g1484 (n_546, n_1101, n_1414, n_1415);
  xor g1485 (n_1416, n_534, n_535);
  xor g1486 (n_537, n_1416, A[15]);
  nand g1487 (n_1417, n_534, n_535);
  nand g1488 (n_1418, A[15], n_535);
  nand g1489 (n_1419, n_534, A[15]);
  nand g1490 (n_548, n_1417, n_1418, n_1419);
  xor g1491 (n_1420, A[16], n_536);
  xor g1492 (n_539, n_1420, n_537);
  nand g1493 (n_1421, A[16], n_536);
  nand g1494 (n_1422, n_537, n_536);
  nand g1495 (n_1423, A[16], n_537);
  nand g1496 (n_549, n_1421, n_1422, n_1423);
  xor g1497 (n_1424, A[19], n_538);
  xor g1498 (n_541, n_1424, A[20]);
  nand g1499 (n_1425, A[19], n_538);
  nand g1500 (n_1426, A[20], n_538);
  nand g1502 (n_551, n_1425, n_1426, n_1163);
  xor g1503 (n_1428, n_539, n_540);
  xor g1504 (n_543, n_1428, n_541);
  nand g1505 (n_1429, n_539, n_540);
  nand g1506 (n_1430, n_541, n_540);
  nand g1507 (n_1431, n_539, n_541);
  nand g1508 (n_553, n_1429, n_1430, n_1431);
  xor g1510 (n_544, n_1168, n_542);
  nand g1513 (n_1435, A[23], n_542);
  nand g1514 (n_556, n_1169, n_1434, n_1435);
  xor g1515 (n_1436, n_543, n_544);
  xor g1516 (n_87, n_1436, n_545);
  nand g1517 (n_1437, n_543, n_544);
  nand g1518 (n_1438, n_545, n_544);
  nand g1519 (n_1439, n_543, n_545);
  nand g1520 (n_38, n_1437, n_1438, n_1439);
  xor g1522 (n_547, n_1188, n_546);
  nand g1524 (n_1442, n_546, A[13]);
  nand g1525 (n_1443, A[12], n_546);
  nand g1526 (n_559, n_1189, n_1442, n_1443);
  xor g1527 (n_1444, A[16], n_547);
  xor g1528 (n_550, n_1444, A[17]);
  nand g1529 (n_1445, A[16], n_547);
  nand g1530 (n_1446, A[17], n_547);
  nand g1532 (n_561, n_1445, n_1446, n_886);
  xor g1533 (n_1448, n_548, n_549);
  xor g1534 (n_552, n_1448, n_550);
  nand g1535 (n_1449, n_548, n_549);
  nand g1536 (n_1450, n_550, n_549);
  nand g1537 (n_1451, n_548, n_550);
  nand g1538 (n_563, n_1449, n_1450, n_1451);
  xor g1539 (n_1452, A[20], n_551);
  xor g1540 (n_554, n_1452, n_552);
  nand g1541 (n_1453, A[20], n_551);
  nand g1542 (n_1454, n_552, n_551);
  nand g1543 (n_1455, A[20], n_552);
  nand g1544 (n_565, n_1453, n_1454, n_1455);
  xor g1546 (n_555, n_1456, n_553);
  nand g1549 (n_1459, A[21], n_553);
  nand g1550 (n_567, n_1457, n_1458, n_1459);
  xor g1551 (n_1460, n_554, n_555);
  xor g1552 (n_86, n_1460, n_556);
  nand g1553 (n_1461, n_554, n_555);
  nand g1554 (n_1462, n_556, n_555);
  nand g1555 (n_1463, n_554, n_556);
  nand g1556 (n_37, n_1461, n_1462, n_1463);
  nand g1563 (n_1467, A[14], n_559);
  nand g1564 (n_572, n_1465, n_1466, n_1467);
  xor g1565 (n_1468, A[17], A[18]);
  xor g1566 (n_562, n_1468, n_560);
  nand g1568 (n_1470, n_560, A[18]);
  nand g1569 (n_1471, A[17], n_560);
  nand g1570 (n_573, n_1070, n_1470, n_1471);
  xor g1571 (n_1472, n_561, n_562);
  xor g1572 (n_564, n_1472, n_563);
  nand g1573 (n_1473, n_561, n_562);
  nand g1574 (n_1474, n_563, n_562);
  nand g1575 (n_1475, n_561, n_563);
  nand g1576 (n_576, n_1473, n_1474, n_1475);
  xor g1578 (n_566, n_1244, n_564);
  nand g1580 (n_1478, n_564, A[22]);
  nand g1581 (n_1479, A[21], n_564);
  nand g1582 (n_577, n_1245, n_1478, n_1479);
  xor g1583 (n_1480, n_565, n_566);
  xor g1584 (n_85, n_1480, n_567);
  nand g1585 (n_1481, n_565, n_566);
  nand g1586 (n_1482, n_567, n_566);
  nand g1587 (n_1483, n_565, n_567);
  nand g1588 (n_36, n_1481, n_1482, n_1483);
  nand g1596 (n_580, n_1109, n_1486, n_1465);
  xor g1597 (n_1488, A[18], n_571);
  xor g1598 (n_574, n_1488, n_572);
  nand g1599 (n_1489, A[18], n_571);
  nand g1600 (n_1490, n_572, n_571);
  nand g1601 (n_1491, A[18], n_572);
  nand g1602 (n_582, n_1489, n_1490, n_1491);
  xor g1603 (n_1492, A[19], n_573);
  xor g1604 (n_575, n_1492, n_574);
  nand g1605 (n_1493, A[19], n_573);
  nand g1606 (n_1494, n_574, n_573);
  nand g1607 (n_1495, A[19], n_574);
  nand g1608 (n_584, n_1493, n_1494, n_1495);
  xor g1609 (n_1496, A[22], n_575);
  xor g1610 (n_578, n_1496, A[23]);
  nand g1611 (n_1497, A[22], n_575);
  nand g1612 (n_1498, A[23], n_575);
  nand g1614 (n_586, n_1497, n_1498, n_1125);
  xor g1615 (n_1500, n_576, n_577);
  xor g1616 (n_84, n_1500, n_578);
  nand g1617 (n_1501, n_576, n_577);
  nand g1618 (n_1502, n_578, n_577);
  nand g1619 (n_1503, n_576, n_578);
  nand g1620 (n_35, n_1501, n_1502, n_1503);
  xor g1621 (n_1504, A[15], A[16]);
  xor g1622 (n_581, n_1504, A[13]);
  nand g1624 (n_1506, A[13], A[16]);
  nand g1626 (n_588, n_986, n_1506, n_775);
  xor g1627 (n_1508, n_580, n_581);
  xor g1628 (n_583, n_1508, A[19]);
  nand g1629 (n_1509, n_580, n_581);
  nand g1630 (n_1510, A[19], n_581);
  nand g1631 (n_1511, n_580, A[19]);
  nand g1632 (n_590, n_1509, n_1510, n_1511);
  xor g1633 (n_1512, A[20], n_582);
  xor g1634 (n_585, n_1512, n_583);
  nand g1635 (n_1513, A[20], n_582);
  nand g1636 (n_1514, n_583, n_582);
  nand g1637 (n_1515, A[20], n_583);
  nand g1638 (n_591, n_1513, n_1514, n_1515);
  xor g1639 (n_1516, n_584, n_585);
  xor g1640 (n_587, n_1516, A[23]);
  nand g1641 (n_1517, n_584, n_585);
  nand g1642 (n_1518, A[23], n_585);
  nand g1643 (n_1519, n_584, A[23]);
  nand g1644 (n_593, n_1517, n_1518, n_1519);
  xor g1646 (n_83, n_1520, n_587);
  nand g1648 (n_1522, n_587, n_586);
  nand g1650 (n_34, n_1521, n_1522, n_1523);
  xor g1652 (n_589, n_1336, n_588);
  nand g1654 (n_1526, n_588, A[17]);
  nand g1655 (n_1527, A[16], n_588);
  nand g1656 (n_597, n_886, n_1526, n_1527);
  xor g1657 (n_1528, A[20], n_589);
  xor g1658 (n_592, n_1528, n_590);
  nand g1659 (n_1529, A[20], n_589);
  nand g1660 (n_1530, n_590, n_589);
  nand g1661 (n_1531, A[20], n_590);
  nand g1662 (n_599, n_1529, n_1530, n_1531);
  xor g1664 (n_594, n_1456, n_591);
  nand g1667 (n_1535, A[21], n_591);
  nand g1668 (n_601, n_1457, n_1534, n_1535);
  xor g1669 (n_1536, n_592, n_593);
  xor g1670 (n_82, n_1536, n_594);
  nand g1671 (n_1537, n_592, n_593);
  nand g1672 (n_1538, n_594, n_593);
  nand g1673 (n_1539, n_592, n_594);
  nand g1674 (n_81, n_1537, n_1538, n_1539);
  nand g1681 (n_1543, A[18], n_597);
  nand g1682 (n_605, n_1541, n_1542, n_1543);
  xor g1683 (n_1544, A[21], n_598);
  xor g1684 (n_600, n_1544, A[22]);
  nand g1685 (n_1545, A[21], n_598);
  nand g1686 (n_1546, A[22], n_598);
  nand g1688 (n_608, n_1545, n_1546, n_1245);
  xor g1689 (n_1548, n_599, n_600);
  xor g1690 (n_33, n_1548, n_601);
  nand g1691 (n_1549, n_599, n_600);
  nand g1692 (n_1550, n_601, n_600);
  nand g1693 (n_1551, n_599, n_601);
  nand g1694 (n_32, n_1549, n_1550, n_1551);
  xor g1697 (n_1552, A[17], A[19]);
  nand g1699 (n_1553, A[17], A[19]);
  nand g1702 (n_610, n_1553, n_1554, n_1555);
  xor g1703 (n_1556, n_605, n_606);
  xor g1704 (n_607, n_1556, A[22]);
  nand g1705 (n_1557, n_605, n_606);
  nand g1706 (n_1558, A[22], n_606);
  nand g1707 (n_1559, n_605, A[22]);
  nand g1708 (n_612, n_1557, n_1558, n_1559);
  xor g1709 (n_1560, A[23], n_607);
  xor g1710 (n_80, n_1560, n_608);
  nand g1711 (n_1561, A[23], n_607);
  nand g1712 (n_1562, n_608, n_607);
  nand g1713 (n_1563, A[23], n_608);
  nand g1714 (n_31, n_1561, n_1562, n_1563);
  xor g1715 (n_1564, A[19], A[18]);
  xor g1716 (n_611, n_1564, A[20]);
  nand g1720 (n_614, n_1399, n_927, n_1163);
  xor g1721 (n_1568, n_610, n_611);
  xor g1722 (n_613, n_1568, A[23]);
  nand g1723 (n_1569, n_610, n_611);
  nand g1724 (n_1570, A[23], n_611);
  nand g1725 (n_1571, n_610, A[23]);
  nand g1726 (n_616, n_1569, n_1570, n_1571);
  xor g1728 (n_79, n_1572, n_613);
  nand g1730 (n_1574, n_613, n_612);
  nand g1732 (n_30, n_1573, n_1574, n_1575);
  xor g1733 (n_1576, A[20], n_614);
  xor g1734 (n_615, n_1576, A[21]);
  nand g1735 (n_1577, A[20], n_614);
  nand g1736 (n_1578, A[21], n_614);
  nand g1737 (n_1579, A[20], A[21]);
  nand g1738 (n_619, n_1577, n_1578, n_1579);
  xor g1740 (n_78, n_1580, n_616);
  nand g1742 (n_1582, n_616, n_615);
  nand g1744 (n_77, n_1581, n_1582, n_1583);
  nand g1751 (n_1587, A[22], n_619);
  nand g1752 (n_28, n_1585, n_1586, n_1587);
  xor g1755 (n_1588, A[21], A[23]);
  nand g1760 (n_27, n_1038, n_1590, n_1591);
  xor g1762 (n_75, n_1168, A[22]);
  nand g1766 (n_74, n_1169, n_1125, n_1083);
  nand g16 (n_1608, A[0], A[2]);
  xor g20 (Z[2], A[0], A[2]);
  nand g22 (n_1613, n_70, A[3]);
  nand g25 (n_1617, n_1613, n_1614, n_1615);
  xor g26 (n_1616, n_70, A[3]);
  nand g28 (n_1618, n_69, A[4]);
  nand g29 (n_1619, n_69, n_1617);
  nand g30 (n_1620, A[4], n_1617);
  nand g31 (n_1622, n_1618, n_1619, n_1620);
  xor g32 (n_1621, n_69, A[4]);
  xor g33 (Z[4], n_1617, n_1621);
  nand g34 (n_1623, A[5], n_116);
  nand g35 (n_1624, A[5], n_1622);
  nand g36 (n_1625, n_116, n_1622);
  nand g37 (n_1627, n_1623, n_1624, n_1625);
  xor g38 (n_1626, A[5], n_116);
  xor g39 (Z[5], n_1622, n_1626);
  nand g40 (n_1628, A[6], n_115);
  nand g41 (n_1629, A[6], n_1627);
  nand g42 (n_1630, n_115, n_1627);
  nand g43 (n_1632, n_1628, n_1629, n_1630);
  xor g44 (n_1631, A[6], n_115);
  xor g45 (Z[6], n_1627, n_1631);
  nand g46 (n_1633, A[7], n_114);
  nand g47 (n_1634, A[7], n_1632);
  nand g48 (n_1635, n_114, n_1632);
  nand g49 (n_1637, n_1633, n_1634, n_1635);
  xor g50 (n_1636, A[7], n_114);
  xor g51 (Z[7], n_1632, n_1636);
  nand g52 (n_1638, n_65, n_113);
  nand g53 (n_1639, n_65, n_1637);
  nand g54 (n_1640, n_113, n_1637);
  nand g55 (n_1642, n_1638, n_1639, n_1640);
  xor g56 (n_1641, n_65, n_113);
  xor g57 (Z[8], n_1637, n_1641);
  nand g58 (n_1643, n_64, n_112);
  nand g59 (n_1644, n_64, n_1642);
  nand g60 (n_1645, n_112, n_1642);
  nand g61 (n_1647, n_1643, n_1644, n_1645);
  xor g62 (n_1646, n_64, n_112);
  xor g63 (Z[9], n_1642, n_1646);
  nand g64 (n_1648, n_63, n_111);
  nand g65 (n_1649, n_63, n_1647);
  nand g66 (n_1650, n_111, n_1647);
  nand g67 (n_1652, n_1648, n_1649, n_1650);
  xor g68 (n_1651, n_63, n_111);
  xor g69 (Z[10], n_1647, n_1651);
  nand g70 (n_1653, n_62, n_110);
  nand g71 (n_1654, n_62, n_1652);
  nand g72 (n_1655, n_110, n_1652);
  nand g73 (n_1657, n_1653, n_1654, n_1655);
  xor g74 (n_1656, n_62, n_110);
  xor g75 (Z[11], n_1652, n_1656);
  nand g76 (n_1658, n_61, n_109);
  nand g77 (n_1659, n_61, n_1657);
  nand g78 (n_1660, n_109, n_1657);
  nand g79 (n_1662, n_1658, n_1659, n_1660);
  xor g80 (n_1661, n_61, n_109);
  xor g81 (Z[12], n_1657, n_1661);
  nand g82 (n_1663, n_60, n_108);
  nand g83 (n_1664, n_60, n_1662);
  nand g84 (n_1665, n_108, n_1662);
  nand g85 (n_1667, n_1663, n_1664, n_1665);
  xor g86 (n_1666, n_60, n_108);
  xor g87 (Z[13], n_1662, n_1666);
  nand g88 (n_1668, n_59, n_107);
  nand g89 (n_1669, n_59, n_1667);
  nand g90 (n_1670, n_107, n_1667);
  nand g91 (n_1672, n_1668, n_1669, n_1670);
  xor g92 (n_1671, n_59, n_107);
  xor g93 (Z[14], n_1667, n_1671);
  nand g94 (n_1673, n_58, n_106);
  nand g95 (n_1674, n_58, n_1672);
  nand g96 (n_1675, n_106, n_1672);
  nand g97 (n_1677, n_1673, n_1674, n_1675);
  xor g98 (n_1676, n_58, n_106);
  xor g99 (Z[15], n_1672, n_1676);
  nand g100 (n_1678, n_57, n_105);
  nand g101 (n_1679, n_57, n_1677);
  nand g102 (n_1680, n_105, n_1677);
  nand g103 (n_1682, n_1678, n_1679, n_1680);
  xor g104 (n_1681, n_57, n_105);
  xor g105 (Z[16], n_1677, n_1681);
  nand g106 (n_1683, n_56, n_104);
  nand g107 (n_1684, n_56, n_1682);
  nand g108 (n_1685, n_104, n_1682);
  nand g109 (n_1687, n_1683, n_1684, n_1685);
  xor g110 (n_1686, n_56, n_104);
  xor g111 (Z[17], n_1682, n_1686);
  nand g112 (n_1688, n_55, n_103);
  nand g113 (n_1689, n_55, n_1687);
  nand g114 (n_1690, n_103, n_1687);
  nand g115 (n_1692, n_1688, n_1689, n_1690);
  xor g116 (n_1691, n_55, n_103);
  xor g117 (Z[18], n_1687, n_1691);
  nand g118 (n_1693, n_54, n_102);
  nand g119 (n_1694, n_54, n_1692);
  nand g120 (n_1695, n_102, n_1692);
  nand g121 (n_1697, n_1693, n_1694, n_1695);
  xor g122 (n_1696, n_54, n_102);
  xor g123 (Z[19], n_1692, n_1696);
  nand g124 (n_1698, n_53, n_101);
  nand g125 (n_1699, n_53, n_1697);
  nand g126 (n_1700, n_101, n_1697);
  nand g127 (n_1702, n_1698, n_1699, n_1700);
  xor g128 (n_1701, n_53, n_101);
  xor g129 (Z[20], n_1697, n_1701);
  nand g130 (n_1703, n_52, n_100);
  nand g131 (n_1704, n_52, n_1702);
  nand g132 (n_1705, n_100, n_1702);
  nand g133 (n_1707, n_1703, n_1704, n_1705);
  xor g134 (n_1706, n_52, n_100);
  xor g135 (Z[21], n_1702, n_1706);
  nand g136 (n_1708, n_51, n_99);
  nand g137 (n_1709, n_51, n_1707);
  nand g138 (n_1710, n_99, n_1707);
  nand g139 (n_1712, n_1708, n_1709, n_1710);
  xor g140 (n_1711, n_51, n_99);
  xor g141 (Z[22], n_1707, n_1711);
  nand g142 (n_1713, n_50, n_98);
  nand g143 (n_1714, n_50, n_1712);
  nand g144 (n_1715, n_98, n_1712);
  nand g145 (n_1717, n_1713, n_1714, n_1715);
  xor g146 (n_1716, n_50, n_98);
  xor g147 (Z[23], n_1712, n_1716);
  nand g148 (n_1718, n_49, n_97);
  nand g149 (n_1719, n_49, n_1717);
  nand g150 (n_1720, n_97, n_1717);
  nand g151 (n_1722, n_1718, n_1719, n_1720);
  xor g152 (n_1721, n_49, n_97);
  xor g153 (Z[24], n_1717, n_1721);
  nand g154 (n_1723, n_48, n_96);
  nand g155 (n_1724, n_48, n_1722);
  nand g156 (n_1725, n_96, n_1722);
  nand g157 (n_1727, n_1723, n_1724, n_1725);
  xor g158 (n_1726, n_48, n_96);
  xor g159 (Z[25], n_1722, n_1726);
  nand g160 (n_1728, n_47, n_95);
  nand g161 (n_1729, n_47, n_1727);
  nand g162 (n_1730, n_95, n_1727);
  nand g163 (n_1732, n_1728, n_1729, n_1730);
  xor g164 (n_1731, n_47, n_95);
  xor g165 (Z[26], n_1727, n_1731);
  nand g166 (n_1733, n_46, n_94);
  nand g167 (n_1734, n_46, n_1732);
  nand g168 (n_1735, n_94, n_1732);
  nand g169 (n_1737, n_1733, n_1734, n_1735);
  xor g170 (n_1736, n_46, n_94);
  xor g171 (Z[27], n_1732, n_1736);
  nand g172 (n_1738, n_45, n_93);
  nand g173 (n_1739, n_45, n_1737);
  nand g174 (n_1740, n_93, n_1737);
  nand g175 (n_1742, n_1738, n_1739, n_1740);
  xor g176 (n_1741, n_45, n_93);
  xor g177 (Z[28], n_1737, n_1741);
  nand g178 (n_1743, n_44, n_92);
  nand g179 (n_1744, n_44, n_1742);
  nand g180 (n_1745, n_92, n_1742);
  nand g181 (n_1747, n_1743, n_1744, n_1745);
  xor g182 (n_1746, n_44, n_92);
  xor g183 (Z[29], n_1742, n_1746);
  nand g184 (n_1748, n_43, n_91);
  nand g185 (n_1749, n_43, n_1747);
  nand g186 (n_1750, n_91, n_1747);
  nand g187 (n_1752, n_1748, n_1749, n_1750);
  xor g188 (n_1751, n_43, n_91);
  xor g189 (Z[30], n_1747, n_1751);
  nand g190 (n_1753, n_42, n_90);
  nand g191 (n_1754, n_42, n_1752);
  nand g192 (n_1755, n_90, n_1752);
  nand g193 (n_1757, n_1753, n_1754, n_1755);
  xor g194 (n_1756, n_42, n_90);
  xor g195 (Z[31], n_1752, n_1756);
  nand g196 (n_1758, n_41, n_89);
  nand g197 (n_1759, n_41, n_1757);
  nand g198 (n_1760, n_89, n_1757);
  nand g199 (n_1762, n_1758, n_1759, n_1760);
  xor g200 (n_1761, n_41, n_89);
  xor g201 (Z[32], n_1757, n_1761);
  nand g202 (n_1763, n_40, n_88);
  nand g203 (n_1764, n_40, n_1762);
  nand g204 (n_1765, n_88, n_1762);
  nand g205 (n_1767, n_1763, n_1764, n_1765);
  xor g206 (n_1766, n_40, n_88);
  xor g207 (Z[33], n_1762, n_1766);
  nand g208 (n_1768, n_39, n_87);
  nand g209 (n_1769, n_39, n_1767);
  nand g210 (n_1770, n_87, n_1767);
  nand g211 (n_1772, n_1768, n_1769, n_1770);
  xor g212 (n_1771, n_39, n_87);
  xor g213 (Z[34], n_1767, n_1771);
  nand g214 (n_1773, n_38, n_86);
  nand g215 (n_1774, n_38, n_1772);
  nand g216 (n_1775, n_86, n_1772);
  nand g217 (n_1777, n_1773, n_1774, n_1775);
  xor g218 (n_1776, n_38, n_86);
  xor g219 (Z[35], n_1772, n_1776);
  nand g220 (n_1778, n_37, n_85);
  nand g221 (n_1779, n_37, n_1777);
  nand g222 (n_1780, n_85, n_1777);
  nand g223 (n_1782, n_1778, n_1779, n_1780);
  xor g224 (n_1781, n_37, n_85);
  xor g225 (Z[36], n_1777, n_1781);
  nand g226 (n_1783, n_36, n_84);
  nand g227 (n_1784, n_36, n_1782);
  nand g228 (n_1785, n_84, n_1782);
  nand g229 (n_1787, n_1783, n_1784, n_1785);
  xor g230 (n_1786, n_36, n_84);
  xor g231 (Z[37], n_1782, n_1786);
  nand g232 (n_1788, n_35, n_83);
  nand g233 (n_1789, n_35, n_1787);
  nand g234 (n_1790, n_83, n_1787);
  nand g235 (n_1792, n_1788, n_1789, n_1790);
  xor g236 (n_1791, n_35, n_83);
  xor g237 (Z[38], n_1787, n_1791);
  nand g238 (n_1793, n_34, n_82);
  nand g239 (n_1794, n_34, n_1792);
  nand g240 (n_1795, n_82, n_1792);
  nand g241 (n_1797, n_1793, n_1794, n_1795);
  xor g242 (n_1796, n_34, n_82);
  xor g243 (Z[39], n_1792, n_1796);
  nand g244 (n_1798, n_33, n_81);
  nand g245 (n_1799, n_33, n_1797);
  nand g246 (n_1800, n_81, n_1797);
  nand g247 (n_1802, n_1798, n_1799, n_1800);
  xor g248 (n_1801, n_33, n_81);
  xor g249 (Z[40], n_1797, n_1801);
  nand g250 (n_1803, n_32, n_80);
  nand g251 (n_1804, n_32, n_1802);
  nand g252 (n_1805, n_80, n_1802);
  nand g253 (n_1807, n_1803, n_1804, n_1805);
  xor g254 (n_1806, n_32, n_80);
  xor g255 (Z[41], n_1802, n_1806);
  nand g256 (n_1808, n_31, n_79);
  nand g257 (n_1809, n_31, n_1807);
  nand g258 (n_1810, n_79, n_1807);
  nand g259 (n_1812, n_1808, n_1809, n_1810);
  xor g260 (n_1811, n_31, n_79);
  xor g261 (Z[42], n_1807, n_1811);
  nand g262 (n_1813, n_30, n_78);
  nand g263 (n_1814, n_30, n_1812);
  nand g264 (n_1815, n_78, n_1812);
  nand g265 (n_1817, n_1813, n_1814, n_1815);
  xor g266 (n_1816, n_30, n_78);
  xor g267 (Z[43], n_1812, n_1816);
  nand g1772 (n_1818, n_29, n_77);
  nand g1773 (n_1819, n_29, n_1817);
  nand g1774 (n_1820, n_77, n_1817);
  nand g1775 (n_1822, n_1818, n_1819, n_1820);
  xor g1776 (n_1821, n_29, n_77);
  xor g1777 (Z[44], n_1817, n_1821);
  nand g1778 (n_1823, n_28, n_76);
  nand g1779 (n_1824, n_28, n_1822);
  nand g1780 (n_1825, n_76, n_1822);
  nand g1781 (n_1827, n_1823, n_1824, n_1825);
  xor g1782 (n_1826, n_28, n_76);
  xor g1783 (Z[45], n_1822, n_1826);
  nand g1784 (n_1828, n_27, n_75);
  nand g1785 (n_1829, n_27, n_1827);
  nand g1786 (n_1830, n_75, n_1827);
  nand g1787 (n_1832, n_1828, n_1829, n_1830);
  xor g1788 (n_1831, n_27, n_75);
  xor g1789 (Z[46], n_1827, n_1831);
  xor g1791 (Z[47], n_1832, n_1833);
  or g1803 (n_1045, A[1], wc);
  not gc (wc, n_171);
  or g1804 (n_1046, A[1], wc0);
  not gc0 (wc0, A[2]);
  or g1805 (n_1083, wc1, A[24]);
  not gc1 (wc1, A[22]);
  xnor g1807 (n_1168, A[24], A[23]);
  or g1808 (n_1169, wc2, A[24]);
  not gc2 (wc2, A[23]);
  xnor g1809 (n_1216, A[6], A[5]);
  or g1810 (n_1217, A[5], wc3);
  not gc3 (wc3, A[6]);
  or g1811 (n_1254, A[6], wc4);
  not gc4 (wc4, A[7]);
  or g1812 (n_1255, wc5, A[6]);
  not gc5 (wc5, A[5]);
  or g1814 (n_1357, A[9], wc6);
  not gc6 (wc6, A[10]);
  or g1815 (n_1386, wc7, A[10]);
  not gc7 (wc7, A[9]);
  or g1816 (n_1387, A[10], wc8);
  not gc8 (wc8, A[11]);
  xnor g1817 (n_1456, A[24], A[21]);
  or g1818 (n_1457, wc9, A[24]);
  not gc9 (wc9, A[21]);
  or g1820 (n_1465, A[13], wc10);
  not gc10 (wc10, A[14]);
  or g1822 (n_1541, A[17], wc11);
  not gc11 (wc11, A[18]);
  or g1823 (n_1554, A[18], wc12);
  not gc12 (wc12, A[19]);
  or g1824 (n_1555, wc13, A[18]);
  not gc13 (wc13, A[17]);
  or g1826 (n_1585, A[21], wc14);
  not gc14 (wc14, A[22]);
  or g1827 (n_1590, A[22], wc15);
  not gc15 (wc15, A[23]);
  or g1828 (n_1591, wc16, A[22]);
  not gc16 (wc16, A[21]);
  xnor g1830 (n_1088, A[2], A[1]);
  or g1831 (n_1090, A[1], wc17);
  not gc17 (wc17, A[3]);
  xnor g1832 (n_455, n_1252, A[6]);
  xnor g1833 (n_521, n_1384, A[10]);
  xnor g1834 (n_571, n_1108, A[13]);
  or g1835 (n_1486, A[13], wc18);
  not gc18 (wc18, A[15]);
  xnor g1836 (n_606, n_1552, A[18]);
  xnor g1837 (n_76, n_1588, A[22]);
  or g1839 (n_1049, wc19, n_69);
  not gc19 (wc19, A[5]);
  or g1840 (n_1051, wc20, n_69);
  not gc20 (wc20, n_181);
  xnor g1842 (n_1833, n_74, A[24]);
  or g1844 (n_1053, wc21, n_182);
  not gc21 (wc21, A[6]);
  xnor g1845 (n_507, n_792, n_505);
  or g1846 (n_1358, A[9], wc22);
  not gc22 (wc22, n_505);
  xnor g1847 (n_560, n_1360, n_559);
  or g1848 (n_1466, A[13], wc23);
  not gc23 (wc23, n_559);
  or g1849 (n_1575, A[24], wc24);
  not gc24 (wc24, n_613);
  xnor g1850 (n_1580, n_615, A[24]);
  or g1851 (n_1581, A[24], wc25);
  not gc25 (wc25, n_615);
  or g1852 (n_1583, A[24], wc26);
  not gc26 (wc26, n_616);
  xnor g1853 (n_29, n_1244, n_619);
  or g1854 (n_1586, A[21], wc27);
  not gc27 (wc27, n_619);
  or g1856 (n_1218, A[5], wc28);
  not gc28 (wc28, n_435);
  xnor g1857 (n_598, n_1468, n_597);
  or g1858 (n_1542, A[17], wc29);
  not gc29 (wc29, n_597);
  or g1859 (n_1614, n_1608, wc30);
  not gc30 (wc30, n_70);
  or g1860 (n_1615, wc31, n_1608);
  not gc31 (wc31, A[3]);
  xnor g1861 (Z[3], n_1608, n_1616);
  xnor g1862 (n_355, n_652, n_284);
  or g1863 (n_1054, wc32, n_182);
  not gc32 (wc32, n_284);
  xnor g1864 (n_1572, n_612, A[24]);
  or g1865 (n_1573, A[24], wc33);
  not gc33 (wc33, n_612);
  or g1866 (n_1534, A[24], wc34);
  not gc34 (wc34, n_591);
  xnor g1867 (n_1520, n_586, A[24]);
  or g1868 (n_1521, A[24], wc35);
  not gc35 (wc35, n_586);
  or g1869 (n_1523, A[24], wc36);
  not gc36 (wc36, n_587);
  xnor g1870 (n_1348, n_498, A[24]);
  or g1871 (n_1349, A[24], wc37);
  not gc37 (wc37, n_498);
  or g1872 (n_1458, A[24], wc38);
  not gc38 (wc38, n_553);
  or g1873 (n_1082, A[24], wc39);
  not gc39 (wc39, n_366);
  xnor g1874 (n_369, n_1080, A[24]);
  or g1875 (n_1170, A[24], wc40);
  not gc40 (wc40, n_410);
  or g1876 (n_1350, A[24], wc41);
  not gc41 (wc41, n_499);
  xnor g1877 (n_1208, n_428, A[24]);
  or g1878 (n_1209, A[24], wc42);
  not gc42 (wc42, n_428);
  or g1879 (n_1434, A[24], wc43);
  not gc43 (wc43, n_542);
  or g1880 (n_1210, A[24], wc44);
  not gc44 (wc44, n_429);
  or g1881 (n_1318, A[24], wc45);
  not gc45 (wc45, n_484);
endmodule

module mult_signed_const_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_3885_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_176;
  wire n_179, n_180, n_183, n_184, n_187, n_188, n_189, n_195;
  wire n_196, n_201, n_202, n_203, n_204, n_209, n_210, n_211;
  wire n_212, n_217, n_218, n_219, n_220, n_221, n_223, n_224;
  wire n_225, n_226, n_227, n_233, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_246, n_248, n_249, n_250, n_251, n_260;
  wire n_261, n_262, n_265, n_267, n_269, n_271, n_272, n_273;
  wire n_274, n_275, n_276, n_277, n_282, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_300;
  wire n_302, n_303, n_304, n_305, n_306, n_307, n_308, n_309;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_332, n_333, n_335, n_337, n_338, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_349, n_351, n_352, n_353, n_354;
  wire n_355, n_356, n_357, n_358, n_359, n_361, n_362, n_363;
  wire n_364, n_365, n_366, n_367, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477;
  wire n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485;
  wire n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539;
  wire n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_595;
  wire n_596, n_597, n_598, n_599, n_603, n_604, n_605, n_606;
  wire n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_617;
  wire n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629;
  wire n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637;
  wire n_638, n_639, n_640, n_641, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_658, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_668, n_669, n_670, n_671;
  wire n_672, n_673, n_674, n_675, n_676, n_677, n_684, n_685;
  wire n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693;
  wire n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711;
  wire n_712, n_713, n_722, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_738, n_742, n_743;
  wire n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_751;
  wire n_752, n_753, n_760, n_761, n_762, n_763, n_764, n_765;
  wire n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_792, n_793, n_794, n_795;
  wire n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803;
  wire n_804, n_805, n_822, n_823, n_824, n_825, n_826, n_827;
  wire n_828, n_829, n_830, n_831, n_832, n_833, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_866, n_867, n_868;
  wire n_872, n_873, n_876, n_877, n_878, n_879, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_906, n_907, n_908, n_910;
  wire n_911, n_913, n_914, n_915, n_916, n_917, n_918, n_919;
  wire n_920, n_921, n_922, n_923, n_924, n_925, n_926, n_927;
  wire n_928, n_929, n_946, n_947, n_949, n_950, n_951, n_952;
  wire n_953, n_954, n_955, n_956, n_957, n_958, n_959, n_960;
  wire n_961, n_962, n_963, n_964, n_965, n_984, n_985, n_986;
  wire n_987, n_988, n_989, n_990, n_991, n_992, n_993, n_994;
  wire n_995, n_996, n_997, n_998, n_999, n_1000, n_1001, n_1008;
  wire n_1009, n_1010, n_1011, n_1012, n_1014, n_1015, n_1016, n_1017;
  wire n_1020, n_1021, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031;
  wire n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039;
  wire n_1040, n_1041, n_1042, n_1044, n_1045, n_1046, n_1047, n_1048;
  wire n_1050, n_1051, n_1052, n_1054, n_1055, n_1056, n_1057, n_1058;
  wire n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066;
  wire n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074;
  wire n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082;
  wire n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090;
  wire n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098;
  wire n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106;
  wire n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114;
  wire n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122;
  wire n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1132;
  wire n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140;
  wire n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148;
  wire n_1149, n_1150, n_1151, n_1152, n_1154, n_1155, n_1156, n_1157;
  wire n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165;
  wire n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173;
  wire n_1174, n_1175, n_1176, n_1177, n_1180, n_1181, n_1182, n_1183;
  wire n_1184, n_1185, n_1186, n_1188, n_1189, n_1190, n_1191, n_1192;
  wire n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200;
  wire n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208;
  wire n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216;
  wire n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224;
  wire n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1241;
  wire n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249;
  wire n_1250, n_1252, n_1253, n_1254, n_1255, n_1256, n_1258, n_1259;
  wire n_1260, n_1261, n_1262, n_1263, n_1264, n_1266, n_1267, n_1268;
  wire n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276;
  wire n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284;
  wire n_1285, n_1286, n_1288, n_1290, n_1291, n_1292, n_1293, n_1294;
  wire n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302;
  wire n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310;
  wire n_1311, n_1312, n_1313, n_1316, n_1317, n_1318, n_1319, n_1320;
  wire n_1321, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330;
  wire n_1331, n_1332, n_1333, n_1334, n_1336, n_1337, n_1338, n_1339;
  wire n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347;
  wire n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355;
  wire n_1356, n_1357, n_1358, n_1360, n_1361, n_1362, n_1363, n_1364;
  wire n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381;
  wire n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
  wire n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397;
  wire n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405;
  wire n_1406, n_1407, n_1408, n_1409, n_1412, n_1413, n_1414, n_1415;
  wire n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423;
  wire n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1432, n_1433;
  wire n_1434, n_1435, n_1436, n_1437, n_1440, n_1441, n_1444, n_1445;
  wire n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453;
  wire n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461;
  wire n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470;
  wire n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478;
  wire n_1479, n_1480, n_1481, n_1482, n_1484, n_1485, n_1486, n_1487;
  wire n_1488, n_1490, n_1491, n_1492, n_1493, n_1496, n_1497, n_1498;
  wire n_1499, n_1500, n_1501, n_1504, n_1506, n_1507, n_1508, n_1509;
  wire n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1518;
  wire n_1519, n_1520, n_1521, n_1524, n_1525, n_1526, n_1527, n_1528;
  wire n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536;
  wire n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1544, n_1545;
  wire n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553;
  wire n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561;
  wire n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573;
  wire n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1583, n_1584;
  wire n_1585, n_1587, n_1588, n_1589, n_1593, n_1606, n_1611, n_1612;
  wire n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620;
  wire n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628;
  wire n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636;
  wire n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644;
  wire n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652;
  wire n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660;
  wire n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668;
  wire n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676;
  wire n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684;
  wire n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692;
  wire n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700;
  wire n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708;
  wire n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716;
  wire n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724;
  wire n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732;
  wire n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740;
  wire n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748;
  wire n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756;
  wire n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764;
  wire n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772;
  wire n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780;
  wire n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788;
  wire n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796;
  wire n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804;
  wire n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812;
  wire n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820;
  wire n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828;
  wire n_1829, n_1830, n_1831;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], A[2]);
  xor g270 (n_117, n_622, n_171);
  nand g3 (n_623, A[1], A[2]);
  nand g271 (n_624, n_171, A[2]);
  nand g272 (n_625, A[1], n_171);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, n_69);
  xor g288 (n_176, n_634, A[4]);
  nand g289 (n_635, n_68, n_69);
  nand g290 (n_636, A[4], n_69);
  nand g291 (n_637, n_68, A[4]);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_176);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_176);
  nand g296 (n_640, A[7], n_176);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g305 (n_646, n_117, A[5]);
  xor g306 (n_180, n_646, A[6]);
  nand g307 (n_647, n_117, A[5]);
  nand g308 (n_648, A[6], A[5]);
  nand g309 (n_649, n_117, A[6]);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, n_179, n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, n_179, n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, n_179, A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_188, n_659, n_660, n_661);
  xor g329 (n_662, n_183, A[9]);
  xor g330 (n_112, n_662, n_184);
  nand g331 (n_663, n_183, A[9]);
  nand g332 (n_664, n_184, A[9]);
  nand g333 (n_665, n_183, n_184);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_187, n_630, n_67);
  nand g340 (n_668, n_67, n_173);
  nand g341 (n_669, A[4], n_67);
  nand g342 (n_71, n_631, n_668, n_669);
  xor g343 (n_670, A[7], n_187);
  xor g344 (n_189, n_670, A[8]);
  nand g345 (n_671, A[7], n_187);
  nand g346 (n_672, A[8], n_187);
  nand g347 (n_673, A[7], A[8]);
  nand g348 (n_73, n_671, n_672, n_673);
  xor g349 (n_674, n_188, A[10]);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, n_188, A[10]);
  nand g352 (n_676, n_189, A[10]);
  nand g353 (n_677, n_188, n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_195, n_638, n_71);
  nand g366 (n_684, n_71, n_176);
  nand g367 (n_685, A[5], n_71);
  nand g368 (n_202, n_639, n_684, n_685);
  xor g369 (n_686, A[9], A[8]);
  xor g370 (n_196, n_686, n_73);
  nand g371 (n_687, A[9], A[8]);
  nand g372 (n_688, n_73, A[8]);
  nand g373 (n_689, A[9], n_73);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, A[11], n_195);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, A[11], n_195);
  nand g378 (n_692, n_196, n_195);
  nand g379 (n_693, A[11], n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g394 (n_201, n_650, A[9]);
  nand g396 (n_704, A[9], n_180);
  nand g397 (n_705, n_179, A[9]);
  nand g398 (n_209, n_651, n_704, n_705);
  xor g399 (n_706, A[10], n_201);
  xor g400 (n_204, n_706, n_202);
  nand g401 (n_707, A[10], n_201);
  nand g402 (n_708, n_202, n_201);
  nand g403 (n_709, A[10], n_202);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, A[12], n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, A[12], n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, A[12], n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g423 (n_722, n_183, n_184);
  xor g424 (n_210, n_722, A[10]);
  nand g426 (n_724, A[10], n_184);
  nand g427 (n_725, n_183, A[10]);
  nand g428 (n_218, n_665, n_724, n_725);
  xor g429 (n_726, A[11], n_209);
  xor g430 (n_212, n_726, n_210);
  nand g431 (n_727, A[11], n_209);
  nand g432 (n_728, n_210, n_209);
  nand g433 (n_729, A[11], n_210);
  nand g434 (n_220, n_727, n_728, n_729);
  xor g435 (n_730, n_211, A[13]);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, n_211, A[13]);
  nand g438 (n_732, n_212, A[13]);
  nand g439 (n_733, n_211, n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_217, n_738, n_187);
  xor g455 (n_742, n_188, A[11]);
  xor g456 (n_219, n_742, n_217);
  nand g457 (n_743, n_188, A[11]);
  nand g458 (n_744, n_217, A[11]);
  nand g459 (n_745, n_188, n_217);
  nand g460 (n_224, n_743, n_744, n_745);
  xor g461 (n_746, n_218, A[12]);
  xor g462 (n_221, n_746, A[14]);
  nand g463 (n_747, n_218, A[12]);
  nand g464 (n_748, A[14], A[12]);
  nand g465 (n_749, n_218, A[14]);
  nand g466 (n_226, n_747, n_748, n_749);
  xor g467 (n_750, n_219, n_220);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, n_219, n_220);
  nand g470 (n_752, n_221, n_220);
  nand g471 (n_753, n_219, n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g482 (n_72, n_638, A[9]);
  nand g484 (n_760, A[9], n_176);
  nand g485 (n_761, A[5], A[9]);
  nand g486 (n_233, n_639, n_760, n_761);
  xor g487 (n_762, A[8], n_71);
  xor g488 (n_223, n_762, n_72);
  nand g489 (n_763, A[8], n_71);
  nand g490 (n_764, n_72, n_71);
  nand g491 (n_765, A[8], n_72);
  nand g492 (n_234, n_763, n_764, n_765);
  xor g493 (n_766, n_73, A[12]);
  xor g494 (n_225, n_766, n_223);
  nand g495 (n_767, n_73, A[12]);
  nand g496 (n_768, n_223, A[12]);
  nand g497 (n_769, n_73, n_223);
  nand g498 (n_236, n_767, n_768, n_769);
  xor g499 (n_770, A[13], n_224);
  xor g500 (n_227, n_770, A[15]);
  nand g501 (n_771, A[13], n_224);
  nand g502 (n_772, A[15], n_224);
  nand g503 (n_773, A[13], A[15]);
  nand g504 (n_238, n_771, n_772, n_773);
  xor g505 (n_774, n_225, n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, n_225, n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, n_225, n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g530 (n_235, n_706, n_233);
  nand g532 (n_792, n_233, n_201);
  nand g533 (n_793, A[10], n_233);
  nand g534 (n_246, n_707, n_792, n_793);
  xor g535 (n_794, A[13], n_234);
  xor g536 (n_237, n_794, A[14]);
  nand g537 (n_795, A[13], n_234);
  nand g538 (n_796, A[14], n_234);
  nand g539 (n_797, A[13], A[14]);
  nand g540 (n_248, n_795, n_796, n_797);
  xor g541 (n_798, n_235, n_236);
  xor g542 (n_239, n_798, n_237);
  nand g543 (n_799, n_235, n_236);
  nand g544 (n_800, n_237, n_236);
  nand g545 (n_801, n_235, n_237);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, A[16], n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, A[16], n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, A[16], n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g577 (n_822, n_246, A[14]);
  xor g578 (n_249, n_822, n_212);
  nand g579 (n_823, n_246, A[14]);
  nand g580 (n_824, n_212, A[14]);
  nand g581 (n_825, n_246, n_212);
  nand g582 (n_261, n_823, n_824, n_825);
  xor g583 (n_826, A[15], n_248);
  xor g584 (n_251, n_826, A[17]);
  nand g585 (n_827, A[15], n_248);
  nand g586 (n_828, A[17], n_248);
  nand g587 (n_829, A[15], A[17]);
  nand g588 (n_118, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g616 (n_260, n_746, n_219);
  nand g618 (n_848, n_219, n_218);
  nand g619 (n_849, A[12], n_219);
  nand g620 (n_272, n_747, n_848, n_849);
  xor g621 (n_850, n_220, A[15]);
  xor g622 (n_262, n_850, n_260);
  nand g623 (n_851, n_220, A[15]);
  nand g624 (n_852, n_260, A[15]);
  nand g625 (n_853, n_220, n_260);
  nand g626 (n_274, n_851, n_852, n_853);
  xor g627 (n_854, A[16], n_261);
  xor g628 (n_119, n_854, A[18]);
  nand g629 (n_855, A[16], n_261);
  nand g630 (n_856, A[18], n_261);
  nand g631 (n_857, A[16], A[18]);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_262, n_118);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_262, n_118);
  nand g636 (n_860, n_119, n_118);
  nand g637 (n_861, n_262, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g641 (n_862, n_68, A[4]);
  xor g642 (n_265, n_862, n_69);
  xor g647 (n_866, A[5], n_265);
  xor g648 (n_267, n_866, A[9]);
  nand g649 (n_867, A[5], n_265);
  nand g650 (n_868, A[9], n_265);
  nand g652 (n_282, n_867, n_868, n_761);
  xor g654 (n_269, n_762, n_267);
  nand g656 (n_872, n_267, n_71);
  nand g657 (n_873, A[8], n_267);
  nand g658 (n_284, n_763, n_872, n_873);
  xor g660 (n_271, n_766, A[13]);
  nand g662 (n_876, A[13], A[12]);
  nand g663 (n_877, n_73, A[13]);
  nand g664 (n_286, n_767, n_876, n_877);
  xor g665 (n_878, n_269, n_224);
  xor g666 (n_273, n_878, n_271);
  nand g667 (n_879, n_269, n_224);
  nand g668 (n_880, n_271, n_224);
  nand g669 (n_881, n_269, n_271);
  nand g670 (n_288, n_879, n_880, n_881);
  xor g671 (n_882, n_272, A[16]);
  xor g672 (n_275, n_882, A[17]);
  nand g673 (n_883, n_272, A[16]);
  nand g674 (n_884, A[17], A[16]);
  nand g675 (n_885, n_272, A[17]);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, n_273, n_274);
  xor g678 (n_277, n_886, A[19]);
  nand g679 (n_887, n_273, n_274);
  nand g680 (n_888, A[19], n_274);
  nand g681 (n_889, n_273, A[19]);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g707 (n_906, A[10], n_282);
  xor g708 (n_285, n_906, n_201);
  nand g709 (n_907, A[10], n_282);
  nand g710 (n_908, n_201, n_282);
  nand g712 (n_300, n_907, n_908, n_707);
  xor g713 (n_910, n_284, A[13]);
  xor g714 (n_287, n_910, A[14]);
  nand g715 (n_911, n_284, A[13]);
  nand g717 (n_913, n_284, A[14]);
  nand g718 (n_302, n_911, n_797, n_913);
  xor g719 (n_914, n_285, n_286);
  xor g720 (n_289, n_914, n_287);
  nand g721 (n_915, n_285, n_286);
  nand g722 (n_916, n_287, n_286);
  nand g723 (n_917, n_285, n_287);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, A[17], n_288);
  xor g726 (n_291, n_918, n_289);
  nand g727 (n_919, A[17], n_288);
  nand g728 (n_920, n_289, n_288);
  nand g729 (n_921, A[17], n_289);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, A[18], n_290);
  xor g732 (n_293, n_922, A[20]);
  nand g733 (n_923, A[18], n_290);
  nand g734 (n_924, A[20], n_290);
  nand g735 (n_925, A[18], A[20]);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g767 (n_946, n_300, A[14]);
  xor g768 (n_303, n_946, n_212);
  nand g769 (n_947, n_300, A[14]);
  nand g771 (n_949, n_300, n_212);
  nand g772 (n_319, n_947, n_824, n_949);
  xor g773 (n_950, A[15], n_302);
  xor g774 (n_305, n_950, n_303);
  nand g775 (n_951, A[15], n_302);
  nand g776 (n_952, n_303, n_302);
  nand g777 (n_953, A[15], n_303);
  nand g778 (n_321, n_951, n_952, n_953);
  xor g779 (n_954, n_304, A[18]);
  xor g780 (n_307, n_954, n_305);
  nand g781 (n_955, n_304, A[18]);
  nand g782 (n_956, n_305, A[18]);
  nand g783 (n_957, n_304, n_305);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, A[19], n_306);
  xor g786 (n_309, n_958, A[21]);
  nand g787 (n_959, A[19], n_306);
  nand g788 (n_960, A[21], n_306);
  nand g789 (n_961, A[19], A[21]);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g824 (n_320, n_850, A[16]);
  nand g826 (n_984, A[16], A[15]);
  nand g827 (n_985, n_220, A[16]);
  nand g828 (n_338, n_851, n_984, n_985);
  xor g829 (n_986, n_260, n_319);
  xor g830 (n_322, n_986, n_320);
  nand g831 (n_987, n_260, n_319);
  nand g832 (n_988, n_320, n_319);
  nand g833 (n_989, n_260, n_320);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, n_321, A[19]);
  xor g836 (n_324, n_990, n_322);
  nand g837 (n_991, n_321, A[19]);
  nand g838 (n_992, n_322, A[19]);
  nand g839 (n_993, n_321, n_322);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, A[20], n_323);
  xor g842 (n_326, n_994, A[22]);
  nand g843 (n_995, A[20], n_323);
  nand g844 (n_996, A[22], n_323);
  nand g845 (n_997, A[20], A[22]);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, n_324, n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, n_324, n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, n_324, n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g862 (n_332, n_866, A[8]);
  nand g864 (n_1008, A[8], n_265);
  nand g865 (n_1009, A[5], A[8]);
  nand g866 (n_352, n_867, n_1008, n_1009);
  xor g867 (n_1010, A[9], n_71);
  xor g868 (n_333, n_1010, n_73);
  nand g869 (n_1011, A[9], n_71);
  nand g870 (n_1012, n_73, n_71);
  nand g872 (n_354, n_1011, n_1012, n_689);
  xor g873 (n_1014, n_332, A[12]);
  xor g874 (n_335, n_1014, n_333);
  nand g875 (n_1015, n_332, A[12]);
  nand g876 (n_1016, n_333, A[12]);
  nand g877 (n_1017, n_332, n_333);
  nand g878 (n_356, n_1015, n_1016, n_1017);
  xor g880 (n_337, n_770, n_335);
  nand g882 (n_1020, n_335, n_224);
  nand g883 (n_1021, A[13], n_335);
  nand g884 (n_358, n_771, n_1020, n_1021);
  xor g891 (n_1026, n_337, n_338);
  xor g892 (n_341, n_1026, n_275);
  nand g893 (n_1027, n_337, n_338);
  nand g894 (n_1028, n_275, n_338);
  nand g895 (n_1029, n_337, n_275);
  nand g896 (n_362, n_1027, n_1028, n_1029);
  xor g897 (n_1030, n_340, A[20]);
  xor g898 (n_343, n_1030, n_341);
  nand g899 (n_1031, n_340, A[20]);
  nand g900 (n_1032, n_341, A[20]);
  nand g901 (n_1033, n_340, n_341);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, A[21], n_342);
  xor g904 (n_345, n_1034, n_343);
  nand g905 (n_1035, A[21], n_342);
  nand g906 (n_1036, n_343, n_342);
  nand g907 (n_1037, A[21], n_343);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, A[23], n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, A[23], n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, A[23], n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  xor g917 (n_1042, A[2], n_171);
  nand g922 (n_371, n_624, n_1044, n_1045);
  xor g923 (n_1046, A[5], n_349);
  xor g924 (n_351, n_1046, A[6]);
  nand g925 (n_1047, A[5], n_349);
  nand g926 (n_1048, A[6], n_349);
  nand g928 (n_373, n_1047, n_1048, n_648);
  xor g929 (n_1050, n_179, n_351);
  xor g930 (n_353, n_1050, A[9]);
  nand g931 (n_1051, n_179, n_351);
  nand g932 (n_1052, A[9], n_351);
  nand g934 (n_375, n_1051, n_1052, n_705);
  xor g935 (n_1054, A[10], n_352);
  xor g936 (n_355, n_1054, n_353);
  nand g937 (n_1055, A[10], n_352);
  nand g938 (n_1056, n_353, n_352);
  nand g939 (n_1057, A[10], n_353);
  nand g940 (n_377, n_1055, n_1056, n_1057);
  xor g941 (n_1058, n_354, A[13]);
  xor g942 (n_357, n_1058, n_355);
  nand g943 (n_1059, n_354, A[13]);
  nand g944 (n_1060, n_355, A[13]);
  nand g945 (n_1061, n_354, n_355);
  nand g946 (n_379, n_1059, n_1060, n_1061);
  xor g947 (n_1062, A[14], n_356);
  xor g948 (n_359, n_1062, n_357);
  nand g949 (n_1063, A[14], n_356);
  nand g950 (n_1064, n_357, n_356);
  nand g951 (n_1065, A[14], n_357);
  nand g952 (n_381, n_1063, n_1064, n_1065);
  xor g953 (n_1066, A[17], n_358);
  xor g954 (n_361, n_1066, A[18]);
  nand g955 (n_1067, A[17], n_358);
  nand g956 (n_1068, A[18], n_358);
  nand g957 (n_1069, A[17], A[18]);
  nand g958 (n_383, n_1067, n_1068, n_1069);
  xor g959 (n_1070, n_359, n_290);
  xor g960 (n_363, n_1070, n_361);
  nand g961 (n_1071, n_359, n_290);
  nand g962 (n_1072, n_361, n_290);
  nand g963 (n_1073, n_359, n_361);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, A[21], n_362);
  xor g966 (n_365, n_1074, A[22]);
  nand g967 (n_1075, A[21], n_362);
  nand g968 (n_1076, A[22], n_362);
  nand g969 (n_1077, A[21], A[22]);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g971 (n_1078, n_363, n_364);
  nand g973 (n_1079, n_363, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  xor g985 (n_1086, A[1], A[3]);
  nand g987 (n_1087, A[1], A[3]);
  nand g990 (n_392, n_1087, n_1088, n_1089);
  xor g991 (n_1090, n_371, A[6]);
  xor g992 (n_374, n_1090, n_372);
  nand g993 (n_1091, n_371, A[6]);
  nand g994 (n_1092, n_372, A[6]);
  nand g995 (n_1093, n_371, n_372);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, n_374);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, n_374, n_373);
  nand g1001 (n_1097, A[7], n_374);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, A[10], A[11]);
  xor g1004 (n_378, n_1098, n_375);
  nand g1005 (n_1099, A[10], A[11]);
  nand g1006 (n_1100, n_375, A[11]);
  nand g1007 (n_1101, A[10], n_375);
  nand g1008 (n_398, n_1099, n_1100, n_1101);
  xor g1009 (n_1102, n_376, n_377);
  xor g1010 (n_380, n_1102, n_378);
  nand g1011 (n_1103, n_376, n_377);
  nand g1012 (n_1104, n_378, n_377);
  nand g1013 (n_1105, n_376, n_378);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, A[14], A[15]);
  xor g1016 (n_382, n_1106, n_379);
  nand g1017 (n_1107, A[14], A[15]);
  nand g1018 (n_1108, n_379, A[15]);
  nand g1019 (n_1109, A[14], n_379);
  nand g1020 (n_402, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, n_380, A[18]);
  xor g1022 (n_384, n_1110, n_381);
  nand g1023 (n_1111, n_380, A[18]);
  nand g1024 (n_1112, n_381, A[18]);
  nand g1025 (n_1113, n_380, n_381);
  nand g1026 (n_404, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, n_382, A[19]);
  xor g1028 (n_386, n_1114, n_383);
  nand g1029 (n_1115, n_382, A[19]);
  nand g1030 (n_1116, n_383, A[19]);
  nand g1031 (n_1117, n_382, n_383);
  nand g1032 (n_406, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_384, A[22]);
  xor g1034 (n_388, n_1118, n_385);
  nand g1035 (n_1119, n_384, A[22]);
  nand g1036 (n_1120, n_385, A[22]);
  nand g1037 (n_1121, n_384, n_385);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, n_386, A[23]);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, n_386, A[23]);
  nand g1042 (n_1124, n_387, A[23]);
  nand g1043 (n_1125, n_386, n_387);
  nand g1044 (n_410, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1052 (n_393, n_626, A[4]);
  nand g1054 (n_1132, A[4], A[2]);
  nand g1055 (n_1133, A[3], A[4]);
  nand g1056 (n_412, n_627, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, n_394, A[8]);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, n_394, A[8]);
  nand g1066 (n_1140, n_395, A[8]);
  nand g1067 (n_1141, n_394, n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, n_396, A[11]);
  xor g1070 (n_399, n_1142, n_397);
  nand g1071 (n_1143, n_396, A[11]);
  nand g1072 (n_1144, n_397, A[11]);
  nand g1073 (n_1145, n_396, n_397);
  nand g1074 (n_417, n_1143, n_1144, n_1145);
  xor g1075 (n_1146, A[12], n_398);
  xor g1076 (n_401, n_1146, n_399);
  nand g1077 (n_1147, A[12], n_398);
  nand g1078 (n_1148, n_399, n_398);
  nand g1079 (n_1149, A[12], n_399);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, A[15], n_400);
  xor g1082 (n_403, n_1150, A[16]);
  nand g1083 (n_1151, A[15], n_400);
  nand g1084 (n_1152, A[16], n_400);
  nand g1086 (n_421, n_1151, n_1152, n_984);
  xor g1087 (n_1154, n_401, n_402);
  xor g1088 (n_405, n_1154, A[19]);
  nand g1089 (n_1155, n_401, n_402);
  nand g1090 (n_1156, A[19], n_402);
  nand g1091 (n_1157, n_401, A[19]);
  nand g1092 (n_424, n_1155, n_1156, n_1157);
  xor g1093 (n_1158, n_403, A[20]);
  xor g1094 (n_407, n_1158, n_404);
  nand g1095 (n_1159, n_403, A[20]);
  nand g1096 (n_1160, n_404, A[20]);
  nand g1097 (n_1161, n_403, n_404);
  nand g1098 (n_425, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_405, n_406);
  xor g1100 (n_409, n_1162, n_407);
  nand g1101 (n_1163, n_405, n_406);
  nand g1102 (n_1164, n_407, n_406);
  nand g1103 (n_1165, n_405, n_407);
  nand g1104 (n_428, n_1163, n_1164, n_1165);
  xor g1106 (n_411, n_1166, n_408);
  nand g1109 (n_1169, A[23], n_408);
  nand g1110 (n_430, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1124 (n_415, n_686, n_413);
  nand g1126 (n_1180, n_413, A[8]);
  nand g1127 (n_1181, A[9], n_413);
  nand g1128 (n_435, n_687, n_1180, n_1181);
  xor g1129 (n_1182, n_414, n_415);
  xor g1130 (n_418, n_1182, n_416);
  nand g1131 (n_1183, n_414, n_415);
  nand g1132 (n_1184, n_416, n_415);
  nand g1133 (n_1185, n_414, n_416);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, A[12], A[13]);
  xor g1136 (n_420, n_1186, n_417);
  nand g1138 (n_1188, n_417, A[13]);
  nand g1139 (n_1189, A[12], n_417);
  nand g1140 (n_439, n_876, n_1188, n_1189);
  xor g1141 (n_1190, n_418, n_419);
  xor g1142 (n_422, n_1190, A[16]);
  nand g1143 (n_1191, n_418, n_419);
  nand g1144 (n_1192, A[16], n_419);
  nand g1145 (n_1193, n_418, A[16]);
  nand g1146 (n_440, n_1191, n_1192, n_1193);
  xor g1147 (n_1194, n_420, A[17]);
  xor g1148 (n_423, n_1194, n_421);
  nand g1149 (n_1195, n_420, A[17]);
  nand g1150 (n_1196, n_421, A[17]);
  nand g1151 (n_1197, n_420, n_421);
  nand g1152 (n_442, n_1195, n_1196, n_1197);
  xor g1153 (n_1198, n_422, A[20]);
  xor g1154 (n_426, n_1198, n_423);
  nand g1155 (n_1199, n_422, A[20]);
  nand g1156 (n_1200, n_423, A[20]);
  nand g1157 (n_1201, n_422, n_423);
  nand g1158 (n_445, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_424, A[21]);
  xor g1160 (n_427, n_1202, n_425);
  nand g1161 (n_1203, n_424, A[21]);
  nand g1162 (n_1204, n_425, A[21]);
  nand g1163 (n_1205, n_424, n_425);
  nand g1164 (n_447, n_1203, n_1204, n_1205);
  xor g1166 (n_429, n_1206, n_427);
  nand g1168 (n_1208, n_427, n_426);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, A[9]);
  nand g1183 (n_1217, A[6], A[9]);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, n_433, A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, n_433, A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, n_433, n_434);
  nand g1190 (n_456, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, n_435, n_436);
  xor g1192 (n_438, n_1222, A[13]);
  nand g1193 (n_1223, n_435, n_436);
  nand g1194 (n_1224, A[13], n_436);
  nand g1195 (n_1225, n_435, A[13]);
  nand g1196 (n_457, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, A[14], n_437);
  xor g1198 (n_441, n_1226, n_438);
  nand g1199 (n_1227, A[14], n_437);
  nand g1200 (n_1228, n_438, n_437);
  nand g1201 (n_1229, A[14], n_438);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, n_439, A[17]);
  xor g1204 (n_443, n_1230, n_440);
  nand g1205 (n_1231, n_439, A[17]);
  nand g1206 (n_1232, n_440, A[17]);
  nand g1207 (n_1233, n_439, n_440);
  nand g1208 (n_461, n_1231, n_1232, n_1233);
  xor g1209 (n_1234, A[18], n_441);
  xor g1210 (n_444, n_1234, n_442);
  nand g1211 (n_1235, A[18], n_441);
  nand g1212 (n_1236, n_442, n_441);
  nand g1213 (n_1237, A[18], n_442);
  nand g1214 (n_463, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_443, A[21]);
  xor g1216 (n_446, n_1238, A[22]);
  nand g1217 (n_1239, n_443, A[21]);
  nand g1219 (n_1241, n_443, A[22]);
  nand g1220 (n_465, n_1239, n_1077, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[5], A[7]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], n_453);
  xor g1242 (n_455, n_1254, A[11]);
  nand g1243 (n_1255, A[10], n_453);
  nand g1244 (n_1256, A[11], n_453);
  nand g1246 (n_472, n_1255, n_1256, n_1099);
  xor g1247 (n_1258, n_454, n_455);
  xor g1248 (n_458, n_1258, n_456);
  nand g1249 (n_1259, n_454, n_455);
  nand g1250 (n_1260, n_456, n_455);
  nand g1251 (n_1261, n_454, n_456);
  nand g1252 (n_474, n_1259, n_1260, n_1261);
  xor g1253 (n_1262, A[14], n_457);
  xor g1254 (n_460, n_1262, A[15]);
  nand g1255 (n_1263, A[14], n_457);
  nand g1256 (n_1264, A[15], n_457);
  nand g1258 (n_476, n_1263, n_1264, n_1107);
  xor g1259 (n_1266, n_458, A[18]);
  xor g1260 (n_462, n_1266, n_459);
  nand g1261 (n_1267, n_458, A[18]);
  nand g1262 (n_1268, n_459, A[18]);
  nand g1263 (n_1269, n_458, n_459);
  nand g1264 (n_479, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, n_460, A[19]);
  xor g1266 (n_464, n_1270, n_461);
  nand g1267 (n_1271, n_460, A[19]);
  nand g1268 (n_1272, n_461, A[19]);
  nand g1269 (n_1273, n_460, n_461);
  nand g1270 (n_480, n_1271, n_1272, n_1273);
  xor g1271 (n_1274, n_462, A[22]);
  xor g1272 (n_466, n_1274, n_463);
  nand g1273 (n_1275, n_462, A[22]);
  nand g1274 (n_1276, n_463, A[22]);
  nand g1275 (n_1277, n_462, n_463);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1277 (n_1278, n_464, A[23]);
  xor g1278 (n_467, n_1278, n_465);
  nand g1279 (n_1279, n_464, A[23]);
  nand g1280 (n_1280, n_465, A[23]);
  nand g1281 (n_1281, n_464, n_465);
  nand g1282 (n_484, n_1279, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1289 (n_1286, A[7], A[6]);
  xor g1290 (n_471, n_1286, A[8]);
  nand g1292 (n_1288, A[8], A[6]);
  nand g1294 (n_486, n_661, n_1288, n_673);
  xor g1295 (n_1290, n_470, A[11]);
  xor g1296 (n_473, n_1290, n_471);
  nand g1297 (n_1291, n_470, A[11]);
  nand g1298 (n_1292, n_471, A[11]);
  nand g1299 (n_1293, n_470, n_471);
  nand g1300 (n_487, n_1291, n_1292, n_1293);
  xor g1301 (n_1294, A[12], n_472);
  xor g1302 (n_475, n_1294, n_473);
  nand g1303 (n_1295, A[12], n_472);
  nand g1304 (n_1296, n_473, n_472);
  nand g1305 (n_1297, A[12], n_473);
  nand g1306 (n_490, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, A[15], n_474);
  xor g1308 (n_477, n_1298, n_475);
  nand g1309 (n_1299, A[15], n_474);
  nand g1310 (n_1300, n_475, n_474);
  nand g1311 (n_1301, A[15], n_475);
  nand g1312 (n_491, n_1299, n_1300, n_1301);
  xor g1313 (n_1302, A[16], n_476);
  xor g1314 (n_478, n_1302, n_477);
  nand g1315 (n_1303, A[16], n_476);
  nand g1316 (n_1304, n_477, n_476);
  nand g1317 (n_1305, A[16], n_477);
  nand g1318 (n_494, n_1303, n_1304, n_1305);
  xor g1319 (n_1306, A[19], n_478);
  xor g1320 (n_481, n_1306, n_479);
  nand g1321 (n_1307, A[19], n_478);
  nand g1322 (n_1308, n_479, n_478);
  nand g1323 (n_1309, A[19], n_479);
  nand g1324 (n_495, n_1307, n_1308, n_1309);
  xor g1325 (n_1310, A[20], n_480);
  xor g1326 (n_483, n_1310, n_481);
  nand g1327 (n_1311, A[20], n_480);
  nand g1328 (n_1312, n_481, n_480);
  nand g1329 (n_1313, A[20], n_481);
  nand g1330 (n_498, n_1311, n_1312, n_1313);
  xor g1332 (n_485, n_1166, n_482);
  nand g1335 (n_1317, A[23], n_482);
  nand g1336 (n_500, n_1167, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1344 (n_488, n_686, n_486);
  nand g1346 (n_1324, n_486, A[8]);
  nand g1347 (n_1325, A[9], n_486);
  nand g1348 (n_503, n_687, n_1324, n_1325);
  xor g1349 (n_1326, A[12], n_487);
  xor g1350 (n_489, n_1326, n_488);
  nand g1351 (n_1327, A[12], n_487);
  nand g1352 (n_1328, n_488, n_487);
  nand g1353 (n_1329, A[12], n_488);
  nand g1354 (n_504, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, A[13], n_489);
  xor g1356 (n_492, n_1330, n_490);
  nand g1357 (n_1331, A[13], n_489);
  nand g1358 (n_1332, n_490, n_489);
  nand g1359 (n_1333, A[13], n_490);
  nand g1360 (n_507, n_1331, n_1332, n_1333);
  xor g1361 (n_1334, A[16], A[17]);
  xor g1362 (n_493, n_1334, n_491);
  nand g1364 (n_1336, n_491, A[17]);
  nand g1365 (n_1337, A[16], n_491);
  nand g1366 (n_509, n_884, n_1336, n_1337);
  xor g1367 (n_1338, n_492, A[20]);
  xor g1368 (n_496, n_1338, n_493);
  nand g1369 (n_1339, n_492, A[20]);
  nand g1370 (n_1340, n_493, A[20]);
  nand g1371 (n_1341, n_492, n_493);
  nand g1372 (n_511, n_1339, n_1340, n_1341);
  xor g1373 (n_1342, n_494, A[21]);
  xor g1374 (n_497, n_1342, n_495);
  nand g1375 (n_1343, n_494, A[21]);
  nand g1376 (n_1344, n_495, A[21]);
  nand g1377 (n_1345, n_494, n_495);
  nand g1378 (n_513, n_1343, n_1344, n_1345);
  xor g1380 (n_499, n_1346, n_497);
  nand g1383 (n_1349, n_496, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  xor g1394 (n_505, n_1354, n_503);
  nand g1397 (n_1357, A[10], n_503);
  nand g1398 (n_520, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], A[14]);
  xor g1400 (n_506, n_1358, n_504);
  nand g1402 (n_1360, n_504, A[14]);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_521, n_797, n_1360, n_1361);
  xor g1405 (n_1362, n_505, A[17]);
  xor g1406 (n_508, n_1362, n_506);
  nand g1407 (n_1363, n_505, A[17]);
  nand g1408 (n_1364, n_506, A[17]);
  nand g1409 (n_1365, n_505, n_506);
  nand g1410 (n_523, n_1363, n_1364, n_1365);
  xor g1411 (n_1366, A[18], n_507);
  xor g1412 (n_510, n_1366, n_508);
  nand g1413 (n_1367, A[18], n_507);
  nand g1414 (n_1368, n_508, n_507);
  nand g1415 (n_1369, A[18], n_508);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_509, A[21]);
  xor g1418 (n_512, n_1370, A[22]);
  nand g1419 (n_1371, n_509, A[21]);
  nand g1421 (n_1373, n_509, A[22]);
  nand g1422 (n_527, n_1371, n_1077, n_1373);
  xor g1423 (n_1374, n_510, n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, n_510, n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, n_510, n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1437 (n_1382, A[9], A[11]);
  nand g1439 (n_1383, A[9], A[11]);
  nand g1442 (n_532, n_1383, n_1384, n_1385);
  xor g1443 (n_1386, A[14], n_519);
  xor g1444 (n_522, n_1386, n_520);
  nand g1445 (n_1387, A[14], n_519);
  nand g1446 (n_1388, n_520, n_519);
  nand g1447 (n_1389, A[14], n_520);
  nand g1448 (n_534, n_1387, n_1388, n_1389);
  xor g1449 (n_1390, A[15], n_521);
  xor g1450 (n_524, n_1390, n_522);
  nand g1451 (n_1391, A[15], n_521);
  nand g1452 (n_1392, n_522, n_521);
  nand g1453 (n_1393, A[15], n_522);
  nand g1454 (n_536, n_1391, n_1392, n_1393);
  xor g1455 (n_1394, A[18], A[19]);
  xor g1456 (n_525, n_1394, n_523);
  nand g1457 (n_1395, A[18], A[19]);
  nand g1458 (n_1396, n_523, A[19]);
  nand g1459 (n_1397, A[18], n_523);
  nand g1460 (n_538, n_1395, n_1396, n_1397);
  xor g1461 (n_1398, n_524, n_525);
  xor g1462 (n_528, n_1398, n_526);
  nand g1463 (n_1399, n_524, n_525);
  nand g1464 (n_1400, n_526, n_525);
  nand g1465 (n_1401, n_524, n_526);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1467 (n_1402, A[22], A[23]);
  xor g1468 (n_529, n_1402, n_527);
  nand g1469 (n_1403, A[22], A[23]);
  nand g1470 (n_1404, n_527, A[23]);
  nand g1471 (n_1405, A[22], n_527);
  nand g1472 (n_543, n_1403, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1480 (n_533, n_1098, A[12]);
  nand g1482 (n_1412, A[12], A[10]);
  nand g1483 (n_1413, A[11], A[12]);
  nand g1484 (n_544, n_1099, n_1412, n_1413);
  xor g1485 (n_1414, n_532, n_533);
  xor g1486 (n_535, n_1414, A[15]);
  nand g1487 (n_1415, n_532, n_533);
  nand g1488 (n_1416, A[15], n_533);
  nand g1489 (n_1417, n_532, A[15]);
  nand g1490 (n_546, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, A[16], n_534);
  xor g1492 (n_537, n_1418, n_535);
  nand g1493 (n_1419, A[16], n_534);
  nand g1494 (n_1420, n_535, n_534);
  nand g1495 (n_1421, A[16], n_535);
  nand g1496 (n_547, n_1419, n_1420, n_1421);
  xor g1497 (n_1422, A[19], n_536);
  xor g1498 (n_539, n_1422, A[20]);
  nand g1499 (n_1423, A[19], n_536);
  nand g1500 (n_1424, A[20], n_536);
  nand g1501 (n_1425, A[19], A[20]);
  nand g1502 (n_550, n_1423, n_1424, n_1425);
  xor g1503 (n_1426, n_537, n_538);
  xor g1504 (n_541, n_1426, n_539);
  nand g1505 (n_1427, n_537, n_538);
  nand g1506 (n_1428, n_539, n_538);
  nand g1507 (n_1429, n_537, n_539);
  nand g1508 (n_552, n_1427, n_1428, n_1429);
  xor g1510 (n_542, n_1166, n_540);
  nand g1513 (n_1433, A[23], n_540);
  nand g1514 (n_553, n_1167, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1522 (n_545, n_1186, n_544);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_876, n_1440, n_1441);
  xor g1528 (n_548, n_1334, n_545);
  nand g1530 (n_1444, n_545, A[17]);
  nand g1531 (n_1445, A[16], n_545);
  nand g1532 (n_558, n_884, n_1444, n_1445);
  xor g1533 (n_1446, n_546, n_547);
  xor g1534 (n_549, n_1446, n_548);
  nand g1535 (n_1447, n_546, n_547);
  nand g1536 (n_1448, n_548, n_547);
  nand g1537 (n_1449, n_546, n_548);
  nand g1538 (n_561, n_1447, n_1448, n_1449);
  xor g1539 (n_1450, A[20], A[21]);
  xor g1540 (n_551, n_1450, n_549);
  nand g1541 (n_1451, A[20], A[21]);
  nand g1542 (n_1452, n_549, A[21]);
  nand g1543 (n_1453, A[20], n_549);
  nand g1544 (n_563, n_1451, n_1452, n_1453);
  xor g1546 (n_554, n_1454, n_551);
  nand g1549 (n_1457, n_550, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1563 (n_1465, A[14], A[17]);
  nand g1564 (n_570, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, n_557, A[18]);
  xor g1566 (n_560, n_1466, n_558);
  nand g1567 (n_1467, n_557, A[18]);
  nand g1568 (n_1468, n_558, A[18]);
  nand g1569 (n_1469, n_557, n_558);
  nand g1570 (n_571, n_1467, n_1468, n_1469);
  xor g1571 (n_1470, n_559, n_560);
  xor g1572 (n_562, n_1470, A[21]);
  nand g1573 (n_1471, n_559, n_560);
  nand g1574 (n_1472, A[21], n_560);
  nand g1575 (n_1473, n_559, A[21]);
  nand g1576 (n_573, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, n_561, A[22]);
  xor g1578 (n_564, n_1474, n_562);
  nand g1579 (n_1475, n_561, A[22]);
  nand g1580 (n_1476, n_562, A[22]);
  nand g1581 (n_1477, n_561, n_562);
  nand g1582 (n_576, n_1475, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  xor g1591 (n_1482, A[13], A[15]);
  nand g1596 (n_578, n_773, n_1484, n_1485);
  xor g1597 (n_1486, A[18], n_569);
  xor g1598 (n_572, n_1486, A[19]);
  nand g1599 (n_1487, A[18], n_569);
  nand g1600 (n_1488, A[19], n_569);
  nand g1602 (n_580, n_1487, n_1488, n_1395);
  xor g1603 (n_1490, n_570, n_571);
  xor g1604 (n_574, n_1490, n_572);
  nand g1605 (n_1491, n_570, n_571);
  nand g1606 (n_1492, n_572, n_571);
  nand g1607 (n_1493, n_570, n_572);
  nand g1608 (n_582, n_1491, n_1492, n_1493);
  xor g1610 (n_575, n_1402, n_573);
  nand g1612 (n_1496, n_573, A[23]);
  nand g1613 (n_1497, A[22], n_573);
  nand g1614 (n_584, n_1403, n_1496, n_1497);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1622 (n_579, n_1106, A[16]);
  nand g1624 (n_1504, A[16], A[14]);
  nand g1626 (n_586, n_1107, n_1504, n_984);
  xor g1627 (n_1506, n_578, n_579);
  xor g1628 (n_581, n_1506, A[19]);
  nand g1629 (n_1507, n_578, n_579);
  nand g1630 (n_1508, A[19], n_579);
  nand g1631 (n_1509, n_578, A[19]);
  nand g1632 (n_588, n_1507, n_1508, n_1509);
  xor g1633 (n_1510, A[20], n_580);
  xor g1634 (n_583, n_1510, n_581);
  nand g1635 (n_1511, A[20], n_580);
  nand g1636 (n_1512, n_581, n_580);
  nand g1637 (n_1513, A[20], n_581);
  nand g1638 (n_589, n_1511, n_1512, n_1513);
  xor g1639 (n_1514, A[23], n_582);
  nand g1641 (n_1515, A[23], n_582);
  nand g1644 (n_591, n_1515, n_1516, n_1167);
  xor g1645 (n_1518, n_583, n_584);
  xor g1646 (n_83, n_1518, n_585);
  nand g1647 (n_1519, n_583, n_584);
  nand g1648 (n_1520, n_585, n_584);
  nand g1649 (n_1521, n_583, n_585);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1652 (n_587, n_1334, n_586);
  nand g1654 (n_1524, n_586, A[17]);
  nand g1655 (n_1525, A[16], n_586);
  nand g1656 (n_595, n_884, n_1524, n_1525);
  xor g1657 (n_1526, A[20], n_587);
  xor g1658 (n_590, n_1526, n_588);
  nand g1659 (n_1527, A[20], n_587);
  nand g1660 (n_1528, n_588, n_587);
  nand g1661 (n_1529, A[20], n_588);
  nand g1662 (n_597, n_1527, n_1528, n_1529);
  xor g1664 (n_592, n_1530, n_589);
  nand g1667 (n_1533, A[21], n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_81, n_1535, n_1536, n_1537);
  xor g1678 (n_596, n_1538, n_595);
  nand g1681 (n_1541, A[18], n_595);
  nand g1682 (n_604, n_1539, n_1540, n_1541);
  xor g1683 (n_1542, A[21], A[22]);
  xor g1684 (n_598, n_1542, n_596);
  nand g1686 (n_1544, n_596, A[22]);
  nand g1687 (n_1545, A[21], n_596);
  nand g1688 (n_606, n_1077, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_33, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[17], A[19]);
  nand g1699 (n_1551, A[17], A[19]);
  nand g1702 (n_608, n_1551, n_1552, n_1553);
  xor g1703 (n_1554, A[22], n_603);
  xor g1704 (n_605, n_1554, n_604);
  nand g1705 (n_1555, A[22], n_603);
  nand g1706 (n_1556, n_604, n_603);
  nand g1707 (n_1557, A[22], n_604);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, A[23], n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, A[23], n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, A[23], n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1716 (n_609, n_1394, A[20]);
  nand g1720 (n_612, n_1395, n_925, n_1425);
  xor g1721 (n_1566, n_608, n_609);
  xor g1722 (n_611, n_1566, A[23]);
  nand g1723 (n_1567, n_608, n_609);
  nand g1724 (n_1568, A[23], n_609);
  nand g1725 (n_1569, n_608, A[23]);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1728 (n_79, n_1570, n_611);
  nand g1730 (n_1572, n_611, n_610);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1734 (n_613, n_1450, n_612);
  nand g1736 (n_1576, n_612, A[21]);
  nand g1737 (n_1577, A[20], n_612);
  nand g1738 (n_617, n_1451, n_1576, n_1577);
  xor g1740 (n_78, n_1578, n_614);
  nand g1742 (n_1580, n_614, n_613);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_617);
  nand g1752 (n_76, n_1583, n_1584, n_1585);
  nand g1759 (n_1589, A[21], A[23]);
  nand g1760 (n_27, n_1587, n_1588, n_1589);
  xor g1762 (n_75, n_1166, A[22]);
  nand g1766 (n_74, n_1167, n_1403, n_1593);
  nand g16 (n_1606, A[0], A[2]);
  xor g20 (Z[2], A[0], A[2]);
  nand g22 (n_1611, n_68, A[3]);
  nand g25 (n_1615, n_1611, n_1612, n_1613);
  xor g26 (n_1614, n_68, A[3]);
  nand g28 (n_1616, A[4], n_117);
  nand g29 (n_1617, A[4], n_1615);
  nand g30 (n_1618, n_117, n_1615);
  nand g31 (n_1620, n_1616, n_1617, n_1618);
  xor g32 (n_1619, A[4], n_117);
  xor g33 (Z[4], n_1615, n_1619);
  nand g34 (n_1621, A[5], n_116);
  nand g35 (n_1622, A[5], n_1620);
  nand g36 (n_1623, n_116, n_1620);
  nand g37 (n_1625, n_1621, n_1622, n_1623);
  xor g38 (n_1624, A[5], n_116);
  xor g39 (Z[5], n_1620, n_1624);
  nand g40 (n_1626, n_67, n_115);
  nand g41 (n_1627, n_67, n_1625);
  nand g42 (n_1628, n_115, n_1625);
  nand g43 (n_1630, n_1626, n_1627, n_1628);
  xor g44 (n_1629, n_67, n_115);
  xor g45 (Z[6], n_1625, n_1629);
  nand g46 (n_1631, n_66, n_114);
  nand g47 (n_1632, n_66, n_1630);
  nand g48 (n_1633, n_114, n_1630);
  nand g49 (n_1635, n_1631, n_1632, n_1633);
  xor g50 (n_1634, n_66, n_114);
  xor g51 (Z[7], n_1630, n_1634);
  nand g52 (n_1636, n_65, n_113);
  nand g53 (n_1637, n_65, n_1635);
  nand g54 (n_1638, n_113, n_1635);
  nand g55 (n_1640, n_1636, n_1637, n_1638);
  xor g56 (n_1639, n_65, n_113);
  xor g57 (Z[8], n_1635, n_1639);
  nand g58 (n_1641, n_64, n_112);
  nand g59 (n_1642, n_64, n_1640);
  nand g60 (n_1643, n_112, n_1640);
  nand g61 (n_1645, n_1641, n_1642, n_1643);
  xor g62 (n_1644, n_64, n_112);
  xor g63 (Z[9], n_1640, n_1644);
  nand g64 (n_1646, n_63, n_111);
  nand g65 (n_1647, n_63, n_1645);
  nand g66 (n_1648, n_111, n_1645);
  nand g67 (n_1650, n_1646, n_1647, n_1648);
  xor g68 (n_1649, n_63, n_111);
  xor g69 (Z[10], n_1645, n_1649);
  nand g70 (n_1651, n_62, n_110);
  nand g71 (n_1652, n_62, n_1650);
  nand g72 (n_1653, n_110, n_1650);
  nand g73 (n_1655, n_1651, n_1652, n_1653);
  xor g74 (n_1654, n_62, n_110);
  xor g75 (Z[11], n_1650, n_1654);
  nand g76 (n_1656, n_61, n_109);
  nand g77 (n_1657, n_61, n_1655);
  nand g78 (n_1658, n_109, n_1655);
  nand g79 (n_1660, n_1656, n_1657, n_1658);
  xor g80 (n_1659, n_61, n_109);
  xor g81 (Z[12], n_1655, n_1659);
  nand g82 (n_1661, n_60, n_108);
  nand g83 (n_1662, n_60, n_1660);
  nand g84 (n_1663, n_108, n_1660);
  nand g85 (n_1665, n_1661, n_1662, n_1663);
  xor g86 (n_1664, n_60, n_108);
  xor g87 (Z[13], n_1660, n_1664);
  nand g88 (n_1666, n_59, n_107);
  nand g89 (n_1667, n_59, n_1665);
  nand g90 (n_1668, n_107, n_1665);
  nand g91 (n_1670, n_1666, n_1667, n_1668);
  xor g92 (n_1669, n_59, n_107);
  xor g93 (Z[14], n_1665, n_1669);
  nand g94 (n_1671, n_58, n_106);
  nand g95 (n_1672, n_58, n_1670);
  nand g96 (n_1673, n_106, n_1670);
  nand g97 (n_1675, n_1671, n_1672, n_1673);
  xor g98 (n_1674, n_58, n_106);
  xor g99 (Z[15], n_1670, n_1674);
  nand g100 (n_1676, n_57, n_105);
  nand g101 (n_1677, n_57, n_1675);
  nand g102 (n_1678, n_105, n_1675);
  nand g103 (n_1680, n_1676, n_1677, n_1678);
  xor g104 (n_1679, n_57, n_105);
  xor g105 (Z[16], n_1675, n_1679);
  nand g106 (n_1681, n_56, n_104);
  nand g107 (n_1682, n_56, n_1680);
  nand g108 (n_1683, n_104, n_1680);
  nand g109 (n_1685, n_1681, n_1682, n_1683);
  xor g110 (n_1684, n_56, n_104);
  xor g111 (Z[17], n_1680, n_1684);
  nand g112 (n_1686, n_55, n_103);
  nand g113 (n_1687, n_55, n_1685);
  nand g114 (n_1688, n_103, n_1685);
  nand g115 (n_1690, n_1686, n_1687, n_1688);
  xor g116 (n_1689, n_55, n_103);
  xor g117 (Z[18], n_1685, n_1689);
  nand g118 (n_1691, n_54, n_102);
  nand g119 (n_1692, n_54, n_1690);
  nand g120 (n_1693, n_102, n_1690);
  nand g121 (n_1695, n_1691, n_1692, n_1693);
  xor g122 (n_1694, n_54, n_102);
  xor g123 (Z[19], n_1690, n_1694);
  nand g124 (n_1696, n_53, n_101);
  nand g125 (n_1697, n_53, n_1695);
  nand g126 (n_1698, n_101, n_1695);
  nand g127 (n_1700, n_1696, n_1697, n_1698);
  xor g128 (n_1699, n_53, n_101);
  xor g129 (Z[20], n_1695, n_1699);
  nand g130 (n_1701, n_52, n_100);
  nand g131 (n_1702, n_52, n_1700);
  nand g132 (n_1703, n_100, n_1700);
  nand g133 (n_1705, n_1701, n_1702, n_1703);
  xor g134 (n_1704, n_52, n_100);
  xor g135 (Z[21], n_1700, n_1704);
  nand g136 (n_1706, n_51, n_99);
  nand g137 (n_1707, n_51, n_1705);
  nand g138 (n_1708, n_99, n_1705);
  nand g139 (n_1710, n_1706, n_1707, n_1708);
  xor g140 (n_1709, n_51, n_99);
  xor g141 (Z[22], n_1705, n_1709);
  nand g142 (n_1711, n_50, n_98);
  nand g143 (n_1712, n_50, n_1710);
  nand g144 (n_1713, n_98, n_1710);
  nand g145 (n_1715, n_1711, n_1712, n_1713);
  xor g146 (n_1714, n_50, n_98);
  xor g147 (Z[23], n_1710, n_1714);
  nand g148 (n_1716, n_49, n_97);
  nand g149 (n_1717, n_49, n_1715);
  nand g150 (n_1718, n_97, n_1715);
  nand g151 (n_1720, n_1716, n_1717, n_1718);
  xor g152 (n_1719, n_49, n_97);
  xor g153 (Z[24], n_1715, n_1719);
  nand g154 (n_1721, n_48, n_96);
  nand g155 (n_1722, n_48, n_1720);
  nand g156 (n_1723, n_96, n_1720);
  nand g157 (n_1725, n_1721, n_1722, n_1723);
  xor g158 (n_1724, n_48, n_96);
  xor g159 (Z[25], n_1720, n_1724);
  nand g160 (n_1726, n_47, n_95);
  nand g161 (n_1727, n_47, n_1725);
  nand g162 (n_1728, n_95, n_1725);
  nand g163 (n_1730, n_1726, n_1727, n_1728);
  xor g164 (n_1729, n_47, n_95);
  xor g165 (Z[26], n_1725, n_1729);
  nand g166 (n_1731, n_46, n_94);
  nand g167 (n_1732, n_46, n_1730);
  nand g168 (n_1733, n_94, n_1730);
  nand g169 (n_1735, n_1731, n_1732, n_1733);
  xor g170 (n_1734, n_46, n_94);
  xor g171 (Z[27], n_1730, n_1734);
  nand g172 (n_1736, n_45, n_93);
  nand g173 (n_1737, n_45, n_1735);
  nand g174 (n_1738, n_93, n_1735);
  nand g175 (n_1740, n_1736, n_1737, n_1738);
  xor g176 (n_1739, n_45, n_93);
  xor g177 (Z[28], n_1735, n_1739);
  nand g178 (n_1741, n_44, n_92);
  nand g179 (n_1742, n_44, n_1740);
  nand g180 (n_1743, n_92, n_1740);
  nand g181 (n_1745, n_1741, n_1742, n_1743);
  xor g182 (n_1744, n_44, n_92);
  xor g183 (Z[29], n_1740, n_1744);
  nand g184 (n_1746, n_43, n_91);
  nand g185 (n_1747, n_43, n_1745);
  nand g186 (n_1748, n_91, n_1745);
  nand g187 (n_1750, n_1746, n_1747, n_1748);
  xor g188 (n_1749, n_43, n_91);
  xor g189 (Z[30], n_1745, n_1749);
  nand g190 (n_1751, n_42, n_90);
  nand g191 (n_1752, n_42, n_1750);
  nand g192 (n_1753, n_90, n_1750);
  nand g193 (n_1755, n_1751, n_1752, n_1753);
  xor g194 (n_1754, n_42, n_90);
  xor g195 (Z[31], n_1750, n_1754);
  nand g196 (n_1756, n_41, n_89);
  nand g197 (n_1757, n_41, n_1755);
  nand g198 (n_1758, n_89, n_1755);
  nand g199 (n_1760, n_1756, n_1757, n_1758);
  xor g200 (n_1759, n_41, n_89);
  xor g201 (Z[32], n_1755, n_1759);
  nand g202 (n_1761, n_40, n_88);
  nand g203 (n_1762, n_40, n_1760);
  nand g204 (n_1763, n_88, n_1760);
  nand g205 (n_1765, n_1761, n_1762, n_1763);
  xor g206 (n_1764, n_40, n_88);
  xor g207 (Z[33], n_1760, n_1764);
  nand g208 (n_1766, n_39, n_87);
  nand g209 (n_1767, n_39, n_1765);
  nand g210 (n_1768, n_87, n_1765);
  nand g211 (n_1770, n_1766, n_1767, n_1768);
  xor g212 (n_1769, n_39, n_87);
  xor g213 (Z[34], n_1765, n_1769);
  nand g214 (n_1771, n_38, n_86);
  nand g215 (n_1772, n_38, n_1770);
  nand g216 (n_1773, n_86, n_1770);
  nand g217 (n_1775, n_1771, n_1772, n_1773);
  xor g218 (n_1774, n_38, n_86);
  xor g219 (Z[35], n_1770, n_1774);
  nand g220 (n_1776, n_37, n_85);
  nand g221 (n_1777, n_37, n_1775);
  nand g222 (n_1778, n_85, n_1775);
  nand g223 (n_1780, n_1776, n_1777, n_1778);
  xor g224 (n_1779, n_37, n_85);
  xor g225 (Z[36], n_1775, n_1779);
  nand g226 (n_1781, n_36, n_84);
  nand g227 (n_1782, n_36, n_1780);
  nand g228 (n_1783, n_84, n_1780);
  nand g229 (n_1785, n_1781, n_1782, n_1783);
  xor g230 (n_1784, n_36, n_84);
  xor g231 (Z[37], n_1780, n_1784);
  nand g232 (n_1786, n_35, n_83);
  nand g233 (n_1787, n_35, n_1785);
  nand g234 (n_1788, n_83, n_1785);
  nand g235 (n_1790, n_1786, n_1787, n_1788);
  xor g236 (n_1789, n_35, n_83);
  xor g237 (Z[38], n_1785, n_1789);
  nand g238 (n_1791, n_34, n_82);
  nand g239 (n_1792, n_34, n_1790);
  nand g240 (n_1793, n_82, n_1790);
  nand g241 (n_1795, n_1791, n_1792, n_1793);
  xor g242 (n_1794, n_34, n_82);
  xor g243 (Z[39], n_1790, n_1794);
  nand g244 (n_1796, n_33, n_81);
  nand g245 (n_1797, n_33, n_1795);
  nand g246 (n_1798, n_81, n_1795);
  nand g247 (n_1800, n_1796, n_1797, n_1798);
  xor g248 (n_1799, n_33, n_81);
  xor g249 (Z[40], n_1795, n_1799);
  nand g250 (n_1801, n_32, n_80);
  nand g251 (n_1802, n_32, n_1800);
  nand g252 (n_1803, n_80, n_1800);
  nand g253 (n_1805, n_1801, n_1802, n_1803);
  xor g254 (n_1804, n_32, n_80);
  xor g255 (Z[41], n_1800, n_1804);
  nand g256 (n_1806, n_31, n_79);
  nand g257 (n_1807, n_31, n_1805);
  nand g258 (n_1808, n_79, n_1805);
  nand g259 (n_1810, n_1806, n_1807, n_1808);
  xor g260 (n_1809, n_31, n_79);
  xor g261 (Z[42], n_1805, n_1809);
  nand g262 (n_1811, n_30, n_78);
  nand g263 (n_1812, n_30, n_1810);
  nand g264 (n_1813, n_78, n_1810);
  nand g265 (n_1815, n_1811, n_1812, n_1813);
  xor g266 (n_1814, n_30, n_78);
  xor g267 (Z[43], n_1810, n_1814);
  nand g1772 (n_1816, n_29, n_77);
  nand g1773 (n_1817, n_29, n_1815);
  nand g1774 (n_1818, n_77, n_1815);
  nand g1775 (n_1820, n_1816, n_1817, n_1818);
  xor g1776 (n_1819, n_29, n_77);
  xor g1777 (Z[44], n_1815, n_1819);
  nand g1778 (n_1821, n_28, n_76);
  nand g1779 (n_1822, n_28, n_1820);
  nand g1780 (n_1823, n_76, n_1820);
  nand g1781 (n_1825, n_1821, n_1822, n_1823);
  xor g1782 (n_1824, n_28, n_76);
  xor g1783 (Z[45], n_1820, n_1824);
  nand g1784 (n_1826, n_27, n_75);
  nand g1785 (n_1827, n_27, n_1825);
  nand g1786 (n_1828, n_75, n_1825);
  nand g1787 (n_1830, n_1826, n_1827, n_1828);
  xor g1788 (n_1829, n_27, n_75);
  xor g1789 (Z[46], n_1825, n_1829);
  xor g1791 (Z[47], n_1830, n_1831);
  or g1804 (n_1044, A[1], wc);
  not gc (wc, n_171);
  or g1805 (n_1045, A[1], wc0);
  not gc0 (wc0, A[2]);
  or g1806 (n_1088, A[2], wc1);
  not gc1 (wc1, A[3]);
  or g1807 (n_1089, wc2, A[2]);
  not gc2 (wc2, A[1]);
  xnor g1808 (n_1166, A[24], A[23]);
  or g1809 (n_1167, wc3, A[24]);
  not gc3 (wc3, A[23]);
  xnor g1810 (n_1214, A[6], A[5]);
  or g1811 (n_1215, A[5], wc4);
  not gc4 (wc4, A[6]);
  or g1812 (n_1216, A[5], wc5);
  not gc5 (wc5, A[9]);
  or g1813 (n_1252, A[6], wc6);
  not gc6 (wc6, A[7]);
  or g1814 (n_1253, wc7, A[6]);
  not gc7 (wc7, A[5]);
  xnor g1815 (n_1354, A[10], A[9]);
  or g1816 (n_1355, A[9], wc8);
  not gc8 (wc8, A[10]);
  or g1817 (n_1384, A[10], wc9);
  not gc9 (wc9, A[11]);
  or g1818 (n_1385, wc10, A[10]);
  not gc10 (wc10, A[9]);
  or g1820 (n_1463, A[13], wc11);
  not gc11 (wc11, A[14]);
  or g1821 (n_1464, A[13], wc12);
  not gc12 (wc12, A[17]);
  or g1822 (n_1484, A[14], wc13);
  not gc13 (wc13, A[15]);
  or g1823 (n_1485, wc14, A[14]);
  not gc14 (wc14, A[13]);
  xnor g1824 (n_1530, A[24], A[21]);
  or g1825 (n_1531, wc15, A[24]);
  not gc15 (wc15, A[21]);
  xnor g1826 (n_1538, A[18], A[17]);
  or g1827 (n_1539, A[17], wc16);
  not gc16 (wc16, A[18]);
  or g1828 (n_1552, A[18], wc17);
  not gc17 (wc17, A[19]);
  or g1829 (n_1553, wc18, A[18]);
  not gc18 (wc18, A[17]);
  or g1831 (n_1583, A[21], wc19);
  not gc19 (wc19, A[22]);
  or g1832 (n_1587, wc20, A[22]);
  not gc20 (wc20, A[21]);
  or g1833 (n_1588, A[22], wc21);
  not gc21 (wc21, A[23]);
  or g1834 (n_1593, wc22, A[24]);
  not gc22 (wc22, A[22]);
  xnor g1835 (n_349, n_1042, A[1]);
  xnor g1836 (n_372, n_1086, A[2]);
  xnor g1837 (n_453, n_1250, A[6]);
  xnor g1838 (n_519, n_1382, A[10]);
  xnor g1839 (n_559, n_1358, A[17]);
  xnor g1840 (n_569, n_1482, A[14]);
  xnor g1841 (n_603, n_1550, A[18]);
  xnor g1842 (n_28, n_1542, A[23]);
  xnor g1843 (n_1578, n_613, A[24]);
  or g1844 (n_1579, A[24], wc23);
  not gc23 (wc23, n_613);
  xnor g1845 (n_1831, n_74, A[24]);
  or g1846 (n_1356, A[9], wc24);
  not gc24 (wc24, n_503);
  or g1847 (n_1540, A[17], wc25);
  not gc25 (wc25, n_595);
  or g1848 (n_1573, A[24], wc26);
  not gc26 (wc26, n_611);
  or g1849 (n_1581, A[24], wc27);
  not gc27 (wc27, n_614);
  xnor g1850 (n_29, n_1542, n_617);
  or g1851 (n_1584, A[21], wc28);
  not gc28 (wc28, n_617);
  or g1853 (n_1612, n_1606, wc29);
  not gc29 (wc29, n_68);
  or g1854 (n_1613, wc30, n_1606);
  not gc30 (wc30, A[3]);
  xnor g1855 (Z[3], n_1606, n_1614);
  or g1856 (n_1532, A[24], wc31);
  not gc31 (wc31, n_589);
  xnor g1857 (n_1570, n_610, A[24]);
  or g1858 (n_1571, A[24], wc32);
  not gc32 (wc32, n_610);
  or g1859 (n_1516, A[24], wc33);
  not gc33 (wc33, n_582);
  xnor g1860 (n_585, n_1514, A[24]);
  xnor g1861 (n_1346, n_496, A[24]);
  or g1862 (n_1347, A[24], wc34);
  not gc34 (wc34, n_496);
  or g1863 (n_1432, A[24], wc35);
  not gc35 (wc35, n_540);
  xnor g1864 (n_1454, n_550, A[24]);
  or g1865 (n_1455, A[24], wc36);
  not gc36 (wc36, n_550);
  or g1866 (n_1456, A[24], wc37);
  not gc37 (wc37, n_551);
  or g1867 (n_1081, A[24], wc38);
  not gc38 (wc38, n_363);
  xnor g1868 (n_1206, n_426, A[24]);
  or g1869 (n_1207, A[24], wc39);
  not gc39 (wc39, n_426);
  or g1870 (n_1080, A[24], wc40);
  not gc40 (wc40, n_364);
  or g1871 (n_1348, A[24], wc41);
  not gc41 (wc41, n_497);
  xnor g1872 (n_367, n_1078, A[24]);
  or g1873 (n_1168, A[24], wc42);
  not gc42 (wc42, n_408);
  or g1874 (n_1209, A[24], wc43);
  not gc43 (wc43, n_427);
  or g1875 (n_1316, A[24], wc44);
  not gc44 (wc44, n_482);
endmodule

module mult_signed_const_3885_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_3885_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_4152_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_171, n_172, n_173, n_174, n_176;
  wire n_180, n_181, n_184, n_185, n_189, n_190, n_195, n_197;
  wire n_202, n_203, n_204, n_205, n_210, n_211, n_212, n_213;
  wire n_218, n_219, n_220, n_223, n_224, n_225, n_226, n_227;
  wire n_234, n_235, n_236, n_237, n_238, n_239, n_246, n_248;
  wire n_249, n_250, n_251, n_258, n_260, n_261, n_262, n_267;
  wire n_269, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_281, n_282, n_283, n_284, n_285, n_286, n_287, n_288;
  wire n_289, n_290, n_291, n_292, n_293, n_296, n_298, n_299;
  wire n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307;
  wire n_308, n_309, n_315, n_317, n_318, n_319, n_320, n_321;
  wire n_322, n_323, n_324, n_325, n_326, n_333, n_335, n_336;
  wire n_337, n_338, n_339, n_340, n_341, n_342, n_343, n_344;
  wire n_345, n_354, n_355, n_356, n_357, n_358, n_359, n_360;
  wire n_361, n_362, n_363, n_364, n_365, n_366, n_367, n_371;
  wire n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379;
  wire n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387;
  wire n_388, n_389, n_390, n_392, n_393, n_394, n_395, n_396;
  wire n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404;
  wire n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412;
  wire n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420;
  wire n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428;
  wire n_429, n_430, n_433, n_434, n_435, n_436, n_437, n_438;
  wire n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446;
  wire n_447, n_448, n_449, n_453, n_454, n_455, n_456, n_457;
  wire n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465;
  wire n_466, n_467, n_468, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_503, n_504, n_505, n_506, n_507, n_508;
  wire n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_519;
  wire n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527;
  wire n_528, n_529, n_530, n_532, n_533, n_534, n_535, n_536;
  wire n_537, n_538, n_539, n_540, n_541, n_542, n_543, n_544;
  wire n_545, n_546, n_547, n_548, n_549, n_550, n_551, n_552;
  wire n_553, n_554, n_557, n_558, n_559, n_560, n_561, n_562;
  wire n_563, n_564, n_565, n_569, n_570, n_571, n_572, n_573;
  wire n_574, n_575, n_576, n_578, n_579, n_580, n_581, n_582;
  wire n_583, n_584, n_585, n_586, n_587, n_588, n_589, n_590;
  wire n_591, n_592, n_595, n_596, n_597, n_598, n_599, n_603;
  wire n_604, n_605, n_606, n_608, n_609, n_610, n_611, n_612;
  wire n_613, n_614, n_617, n_622, n_623, n_624, n_625, n_626;
  wire n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_634;
  wire n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_646;
  wire n_647, n_648, n_649, n_650, n_651, n_652, n_653, n_658;
  wire n_659, n_660, n_661, n_662, n_663, n_664, n_665, n_670;
  wire n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_684;
  wire n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692;
  wire n_693, n_702, n_703, n_704, n_706, n_707, n_708, n_709;
  wire n_710, n_711, n_712, n_713, n_722, n_724, n_725, n_726;
  wire n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_738;
  wire n_742, n_743, n_744, n_745, n_746, n_747, n_748, n_749;
  wire n_750, n_751, n_752, n_753, n_764, n_765, n_766, n_767;
  wire n_768, n_769, n_770, n_771, n_772, n_773, n_774, n_775;
  wire n_776, n_777, n_792, n_793, n_794, n_795, n_796, n_797;
  wire n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805;
  wire n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829;
  wire n_830, n_831, n_832, n_833, n_842, n_848, n_849, n_850;
  wire n_851, n_852, n_853, n_854, n_855, n_856, n_857, n_858;
  wire n_859, n_860, n_861, n_868, n_869, n_870, n_871, n_872;
  wire n_873, n_876, n_877, n_880, n_881, n_882, n_883, n_884;
  wire n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892;
  wire n_893, n_900, n_901, n_902, n_903, n_904, n_905, n_906;
  wire n_907, n_908, n_909, n_910, n_911, n_912, n_913, n_914;
  wire n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922;
  wire n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_938;
  wire n_939, n_941, n_942, n_943, n_944, n_945, n_946, n_947;
  wire n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955;
  wire n_956, n_957, n_958, n_959, n_960, n_961, n_962, n_963;
  wire n_964, n_965, n_978, n_979, n_980, n_982, n_983, n_984;
  wire n_985, n_986, n_987, n_988, n_989, n_990, n_991, n_992;
  wire n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000;
  wire n_1001, n_1013, n_1014, n_1015, n_1016, n_1017, n_1020, n_1021;
  wire n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029;
  wire n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037;
  wire n_1038, n_1039, n_1040, n_1041, n_1043, n_1044, n_1047, n_1049;
  wire n_1052, n_1053, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061;
  wire n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069;
  wire n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077;
  wire n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085;
  wire n_1086, n_1088, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095;
  wire n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103;
  wire n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111;
  wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119;
  wire n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127;
  wire n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135;
  wire n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143;
  wire n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151;
  wire n_1152, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160;
  wire n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168;
  wire n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176;
  wire n_1177, n_1178, n_1179, n_1180, n_1182, n_1183, n_1184, n_1185;
  wire n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193;
  wire n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201;
  wire n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209;
  wire n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217;
  wire n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225;
  wire n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233;
  wire n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1241, n_1242;
  wire n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250;
  wire n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259;
  wire n_1260, n_1261, n_1262, n_1263, n_1264, n_1266, n_1267, n_1268;
  wire n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276;
  wire n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284;
  wire n_1285, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304;
  wire n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312;
  wire n_1313, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1324;
  wire n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332;
  wire n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340;
  wire n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348;
  wire n_1349, n_1350, n_1351, n_1352, n_1353, n_1355, n_1356, n_1357;
  wire n_1358, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366;
  wire n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374;
  wire n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382;
  wire n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390;
  wire n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398;
  wire n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406;
  wire n_1407, n_1408, n_1409, n_1410, n_1414, n_1415, n_1416, n_1417;
  wire n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425;
  wire n_1426, n_1427, n_1428, n_1429, n_1432, n_1433, n_1434, n_1435;
  wire n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443;
  wire n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451;
  wire n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1460, n_1461, n_1463, n_1464, n_1465, n_1466, n_1468, n_1469;
  wire n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477;
  wire n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485;
  wire n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493;
  wire n_1494, n_1495, n_1496, n_1498, n_1499, n_1500, n_1501, n_1506;
  wire n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514;
  wire n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522;
  wire n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531;
  wire n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1539, n_1540;
  wire n_1541, n_1542, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558;
  wire n_1559, n_1560, n_1561, n_1562, n_1565, n_1566, n_1567, n_1568;
  wire n_1569, n_1570, n_1571, n_1572, n_1573, n_1576, n_1577, n_1578;
  wire n_1579, n_1580, n_1581, n_1583, n_1584, n_1585, n_1587, n_1588;
  wire n_1589, n_1593, n_1606, n_1611, n_1612, n_1613, n_1614, n_1615;
  wire n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623;
  wire n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631;
  wire n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639;
  wire n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647;
  wire n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655;
  wire n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663;
  wire n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671;
  wire n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679;
  wire n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687;
  wire n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695;
  wire n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703;
  wire n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711;
  wire n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719;
  wire n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727;
  wire n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735;
  wire n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743;
  wire n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751;
  wire n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759;
  wire n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767;
  wire n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775;
  wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
  wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
  wire n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815;
  wire n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823;
  wire n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_69, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], n_171);
  xor g270 (n_117, n_622, A[2]);
  nand g3 (n_623, A[1], n_171);
  nand g271 (n_624, A[2], n_171);
  nand g272 (n_625, A[1], A[2]);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_174, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_176, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, n_174);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, n_174, n_173);
  nand g5 (n_633, A[4], n_174);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_69, A[4]);
  xor g288 (n_71, n_634, n_176);
  nand g289 (n_635, n_69, A[4]);
  nand g290 (n_636, n_176, A[4]);
  nand g291 (n_637, n_69, n_176);
  nand g292 (n_180, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_71);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_71);
  nand g296 (n_640, A[7], n_71);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g305 (n_646, n_117, A[5]);
  xor g306 (n_181, n_646, n_180);
  nand g307 (n_647, n_117, A[5]);
  nand g308 (n_648, n_180, A[5]);
  nand g309 (n_649, n_117, n_180);
  nand g310 (n_184, n_647, n_648, n_649);
  xor g311 (n_650, A[6], A[8]);
  xor g312 (n_113, n_650, n_181);
  nand g313 (n_651, A[6], A[8]);
  nand g314 (n_652, n_181, A[8]);
  nand g315 (n_653, A[6], n_181);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, n_116, A[6]);
  xor g324 (n_185, n_658, A[7]);
  nand g325 (n_659, n_116, A[6]);
  nand g326 (n_660, A[7], A[6]);
  nand g327 (n_661, n_116, A[7]);
  nand g328 (n_189, n_659, n_660, n_661);
  xor g329 (n_662, A[9], n_184);
  xor g330 (n_112, n_662, n_185);
  nand g331 (n_663, A[9], n_184);
  nand g332 (n_664, n_185, n_184);
  nand g333 (n_665, A[9], n_185);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g343 (n_670, A[7], n_115);
  xor g344 (n_190, n_670, A[8]);
  nand g345 (n_671, A[7], n_115);
  nand g346 (n_672, A[8], n_115);
  nand g347 (n_673, A[7], A[8]);
  nand g348 (n_195, n_671, n_672, n_673);
  xor g349 (n_674, n_189, A[10]);
  xor g350 (n_111, n_674, n_190);
  nand g351 (n_675, n_189, A[10]);
  nand g352 (n_676, n_190, A[10]);
  nand g353 (n_677, n_189, n_190);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_73, n_638, n_66);
  nand g366 (n_684, n_66, n_71);
  nand g367 (n_685, A[5], n_66);
  nand g368 (n_202, n_639, n_684, n_685);
  xor g369 (n_686, A[8], A[9]);
  xor g370 (n_197, n_686, n_195);
  nand g371 (n_687, A[8], A[9]);
  nand g372 (n_688, n_195, A[9]);
  nand g373 (n_689, A[8], n_195);
  nand g374 (n_204, n_687, n_688, n_689);
  xor g375 (n_690, n_73, A[11]);
  xor g376 (n_110, n_690, n_197);
  nand g377 (n_691, n_73, A[11]);
  nand g378 (n_692, n_197, A[11]);
  nand g379 (n_693, n_73, n_197);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g393 (n_702, A[6], A[9]);
  xor g394 (n_203, n_702, n_181);
  nand g395 (n_703, A[6], A[9]);
  nand g396 (n_704, n_181, A[9]);
  nand g398 (n_210, n_703, n_704, n_653);
  xor g399 (n_706, A[10], n_202);
  xor g400 (n_205, n_706, A[12]);
  nand g401 (n_707, A[10], n_202);
  nand g402 (n_708, A[12], n_202);
  nand g403 (n_709, A[10], A[12]);
  nand g404 (n_212, n_707, n_708, n_709);
  xor g405 (n_710, n_203, n_204);
  xor g406 (n_109, n_710, n_205);
  nand g407 (n_711, n_203, n_204);
  nand g408 (n_712, n_205, n_204);
  nand g409 (n_713, n_203, n_205);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g423 (n_722, n_184, n_185);
  xor g424 (n_211, n_722, A[10]);
  nand g426 (n_724, A[10], n_185);
  nand g427 (n_725, n_184, A[10]);
  nand g428 (n_219, n_664, n_724, n_725);
  xor g429 (n_726, A[11], n_210);
  xor g430 (n_213, n_726, n_211);
  nand g431 (n_727, A[11], n_210);
  nand g432 (n_728, n_211, n_210);
  nand g433 (n_729, A[11], n_211);
  nand g434 (n_67, n_727, n_728, n_729);
  xor g435 (n_730, A[13], n_212);
  xor g436 (n_108, n_730, n_213);
  nand g437 (n_731, A[13], n_212);
  nand g438 (n_732, n_213, n_212);
  nand g439 (n_733, A[13], n_213);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_218, n_738, n_115);
  xor g455 (n_742, n_189, n_218);
  xor g456 (n_220, n_742, A[11]);
  nand g457 (n_743, n_189, n_218);
  nand g458 (n_744, A[11], n_218);
  nand g459 (n_745, n_189, A[11]);
  nand g460 (n_224, n_743, n_744, n_745);
  xor g461 (n_746, A[12], n_219);
  xor g462 (n_68, n_746, A[14]);
  nand g463 (n_747, A[12], n_219);
  nand g464 (n_748, A[14], n_219);
  nand g465 (n_749, A[12], A[14]);
  nand g466 (n_226, n_747, n_748, n_749);
  xor g467 (n_750, n_220, n_67);
  xor g468 (n_107, n_750, n_68);
  nand g469 (n_751, n_220, n_67);
  nand g470 (n_752, n_68, n_67);
  nand g471 (n_753, n_220, n_68);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g488 (n_223, n_686, n_73);
  nand g490 (n_764, n_73, A[9]);
  nand g491 (n_765, A[8], n_73);
  nand g492 (n_234, n_687, n_764, n_765);
  xor g493 (n_766, n_195, A[12]);
  xor g494 (n_225, n_766, n_223);
  nand g495 (n_767, n_195, A[12]);
  nand g496 (n_768, n_223, A[12]);
  nand g497 (n_769, n_195, n_223);
  nand g498 (n_236, n_767, n_768, n_769);
  xor g499 (n_770, A[13], n_224);
  xor g500 (n_227, n_770, n_225);
  nand g501 (n_771, A[13], n_224);
  nand g502 (n_772, n_225, n_224);
  nand g503 (n_773, A[13], n_225);
  nand g504 (n_238, n_771, n_772, n_773);
  xor g505 (n_774, A[15], n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, A[15], n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, A[15], n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g530 (n_235, n_706, n_203);
  nand g532 (n_792, n_203, n_202);
  nand g533 (n_793, A[10], n_203);
  nand g534 (n_246, n_707, n_792, n_793);
  xor g535 (n_794, n_234, A[13]);
  xor g536 (n_237, n_794, n_235);
  nand g537 (n_795, n_234, A[13]);
  nand g538 (n_796, n_235, A[13]);
  nand g539 (n_797, n_234, n_235);
  nand g540 (n_248, n_795, n_796, n_797);
  xor g541 (n_798, A[14], n_236);
  xor g542 (n_239, n_798, A[16]);
  nand g543 (n_799, A[14], n_236);
  nand g544 (n_800, A[16], n_236);
  nand g545 (n_801, A[14], A[16]);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, n_237, n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, n_237, n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, n_237, n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g577 (n_822, A[14], n_246);
  xor g578 (n_249, n_822, n_213);
  nand g579 (n_823, A[14], n_246);
  nand g580 (n_824, n_213, n_246);
  nand g581 (n_825, A[14], n_213);
  nand g582 (n_261, n_823, n_824, n_825);
  xor g583 (n_826, A[15], n_248);
  xor g584 (n_251, n_826, A[17]);
  nand g585 (n_827, A[15], n_248);
  nand g586 (n_828, A[17], n_248);
  nand g587 (n_829, A[15], A[17]);
  nand g588 (n_119, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g609 (n_842, n_189, A[11]);
  xor g610 (n_258, n_842, n_218);
  xor g616 (n_260, n_746, n_258);
  nand g618 (n_848, n_258, n_219);
  nand g619 (n_849, A[12], n_258);
  nand g620 (n_272, n_747, n_848, n_849);
  xor g621 (n_850, n_67, A[15]);
  xor g622 (n_118, n_850, n_260);
  nand g623 (n_851, n_67, A[15]);
  nand g624 (n_852, n_260, A[15]);
  nand g625 (n_853, n_67, n_260);
  nand g626 (n_274, n_851, n_852, n_853);
  xor g627 (n_854, A[16], n_261);
  xor g628 (n_262, n_854, A[18]);
  nand g629 (n_855, A[16], n_261);
  nand g630 (n_856, A[18], n_261);
  nand g631 (n_857, A[16], A[18]);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_118, n_119);
  xor g634 (n_103, n_858, n_262);
  nand g635 (n_859, n_118, n_119);
  nand g636 (n_860, n_262, n_119);
  nand g637 (n_861, n_118, n_262);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g648 (n_267, n_638, A[8]);
  nand g650 (n_868, A[8], n_71);
  nand g651 (n_869, A[5], A[8]);
  nand g652 (n_282, n_639, n_868, n_869);
  xor g653 (n_870, n_66, A[9]);
  xor g654 (n_269, n_870, n_267);
  nand g655 (n_871, n_66, A[9]);
  nand g656 (n_872, n_267, A[9]);
  nand g657 (n_873, n_66, n_267);
  nand g658 (n_284, n_871, n_872, n_873);
  xor g660 (n_271, n_766, n_269);
  nand g662 (n_876, n_269, A[12]);
  nand g663 (n_877, n_195, n_269);
  nand g664 (n_286, n_767, n_876, n_877);
  xor g666 (n_273, n_770, n_271);
  nand g668 (n_880, n_271, A[13]);
  nand g669 (n_881, n_224, n_271);
  nand g670 (n_288, n_771, n_880, n_881);
  xor g671 (n_882, n_272, A[16]);
  xor g672 (n_275, n_882, n_273);
  nand g673 (n_883, n_272, A[16]);
  nand g674 (n_884, n_273, A[16]);
  nand g675 (n_885, n_272, n_273);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, A[17], n_274);
  xor g678 (n_277, n_886, A[19]);
  nand g679 (n_887, A[17], n_274);
  nand g680 (n_888, A[19], n_274);
  nand g681 (n_889, A[17], A[19]);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g696 (n_281, n_646, A[6]);
  nand g698 (n_900, A[6], A[5]);
  nand g699 (n_901, n_117, A[6]);
  nand g700 (n_296, n_647, n_900, n_901);
  xor g701 (n_902, n_180, A[9]);
  xor g702 (n_283, n_902, n_281);
  nand g703 (n_903, n_180, A[9]);
  nand g704 (n_904, n_281, A[9]);
  nand g705 (n_905, n_180, n_281);
  nand g706 (n_298, n_903, n_904, n_905);
  xor g707 (n_906, A[10], n_282);
  xor g708 (n_285, n_906, n_283);
  nand g709 (n_907, A[10], n_282);
  nand g710 (n_908, n_283, n_282);
  nand g711 (n_909, A[10], n_283);
  nand g712 (n_300, n_907, n_908, n_909);
  xor g713 (n_910, n_284, A[13]);
  xor g714 (n_287, n_910, A[14]);
  nand g715 (n_911, n_284, A[13]);
  nand g716 (n_912, A[14], A[13]);
  nand g717 (n_913, n_284, A[14]);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, n_285, n_286);
  xor g720 (n_289, n_914, n_287);
  nand g721 (n_915, n_285, n_286);
  nand g722 (n_916, n_287, n_286);
  nand g723 (n_917, n_285, n_287);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, n_288, A[17]);
  xor g726 (n_291, n_918, n_289);
  nand g727 (n_919, n_288, A[17]);
  nand g728 (n_920, n_289, A[17]);
  nand g729 (n_921, n_288, n_289);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, A[18], n_290);
  xor g732 (n_293, n_922, A[20]);
  nand g733 (n_923, A[18], n_290);
  nand g734 (n_924, A[20], n_290);
  nand g735 (n_925, A[18], A[20]);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g755 (n_938, n_296, n_185);
  xor g756 (n_299, n_938, A[10]);
  nand g757 (n_939, n_296, n_185);
  nand g759 (n_941, n_296, A[10]);
  nand g760 (n_315, n_939, n_724, n_941);
  xor g761 (n_942, A[11], n_298);
  xor g762 (n_301, n_942, n_299);
  nand g763 (n_943, A[11], n_298);
  nand g764 (n_944, n_299, n_298);
  nand g765 (n_945, A[11], n_299);
  nand g766 (n_317, n_943, n_944, n_945);
  xor g767 (n_946, n_300, A[14]);
  xor g768 (n_303, n_946, n_301);
  nand g769 (n_947, n_300, A[14]);
  nand g770 (n_948, n_301, A[14]);
  nand g771 (n_949, n_300, n_301);
  nand g772 (n_319, n_947, n_948, n_949);
  xor g773 (n_950, A[15], n_302);
  xor g774 (n_305, n_950, n_303);
  nand g775 (n_951, A[15], n_302);
  nand g776 (n_952, n_303, n_302);
  nand g777 (n_953, A[15], n_303);
  nand g778 (n_321, n_951, n_952, n_953);
  xor g779 (n_954, n_304, A[18]);
  xor g780 (n_307, n_954, n_305);
  nand g781 (n_955, n_304, A[18]);
  nand g782 (n_956, n_305, A[18]);
  nand g783 (n_957, n_304, n_305);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, A[19], n_306);
  xor g786 (n_309, n_958, A[21]);
  nand g787 (n_959, A[19], n_306);
  nand g788 (n_960, A[21], n_306);
  nand g789 (n_961, A[19], A[21]);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g817 (n_978, A[12], n_315);
  xor g818 (n_318, n_978, n_258);
  nand g819 (n_979, A[12], n_315);
  nand g820 (n_980, n_258, n_315);
  nand g822 (n_336, n_979, n_980, n_849);
  xor g823 (n_982, n_317, A[15]);
  xor g824 (n_320, n_982, A[16]);
  nand g825 (n_983, n_317, A[15]);
  nand g826 (n_984, A[16], A[15]);
  nand g827 (n_985, n_317, A[16]);
  nand g828 (n_338, n_983, n_984, n_985);
  xor g829 (n_986, n_318, n_319);
  xor g830 (n_322, n_986, n_320);
  nand g831 (n_987, n_318, n_319);
  nand g832 (n_988, n_320, n_319);
  nand g833 (n_989, n_318, n_320);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, n_321, A[19]);
  xor g836 (n_324, n_990, n_322);
  nand g837 (n_991, n_321, A[19]);
  nand g838 (n_992, n_322, A[19]);
  nand g839 (n_993, n_321, n_322);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, A[20], n_323);
  xor g842 (n_326, n_994, A[22]);
  nand g843 (n_995, A[20], n_323);
  nand g844 (n_996, A[22], n_323);
  nand g845 (n_997, A[20], A[22]);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, n_324, n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, n_324, n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, n_324, n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g868 (n_333, n_870, n_195);
  nand g871 (n_1013, n_66, n_195);
  nand g872 (n_354, n_871, n_688, n_1013);
  xor g873 (n_1014, n_267, A[12]);
  xor g874 (n_335, n_1014, n_333);
  nand g875 (n_1015, n_267, A[12]);
  nand g876 (n_1016, n_333, A[12]);
  nand g877 (n_1017, n_267, n_333);
  nand g878 (n_356, n_1015, n_1016, n_1017);
  xor g880 (n_337, n_770, n_335);
  nand g882 (n_1020, n_335, A[13]);
  nand g883 (n_1021, n_224, n_335);
  nand g884 (n_358, n_771, n_1020, n_1021);
  xor g885 (n_1022, n_336, A[16]);
  xor g886 (n_339, n_1022, n_337);
  nand g887 (n_1023, n_336, A[16]);
  nand g888 (n_1024, n_337, A[16]);
  nand g889 (n_1025, n_336, n_337);
  nand g890 (n_360, n_1023, n_1024, n_1025);
  xor g891 (n_1026, A[17], n_338);
  xor g892 (n_341, n_1026, n_339);
  nand g893 (n_1027, A[17], n_338);
  nand g894 (n_1028, n_339, n_338);
  nand g895 (n_1029, A[17], n_339);
  nand g896 (n_362, n_1027, n_1028, n_1029);
  xor g897 (n_1030, A[20], n_340);
  xor g898 (n_343, n_1030, n_341);
  nand g899 (n_1031, A[20], n_340);
  nand g900 (n_1032, n_341, n_340);
  nand g901 (n_1033, A[20], n_341);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, A[21], n_342);
  xor g904 (n_345, n_1034, n_343);
  nand g905 (n_1035, A[21], n_342);
  nand g906 (n_1036, n_343, n_342);
  nand g907 (n_1037, A[21], n_343);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, A[23], n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, A[23], n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, A[23], n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  nand g922 (n_371, n_1043, n_1044, n_624);
  nand g928 (n_373, n_1047, n_648, n_1049);
  nand g934 (n_375, n_703, n_1052, n_1053);
  nand g940 (n_377, n_907, n_1056, n_1057);
  xor g941 (n_1058, n_354, A[13]);
  xor g942 (n_357, n_1058, n_355);
  nand g943 (n_1059, n_354, A[13]);
  nand g944 (n_1060, n_355, A[13]);
  nand g945 (n_1061, n_354, n_355);
  nand g946 (n_379, n_1059, n_1060, n_1061);
  xor g947 (n_1062, A[14], n_356);
  xor g948 (n_359, n_1062, n_357);
  nand g949 (n_1063, A[14], n_356);
  nand g950 (n_1064, n_357, n_356);
  nand g951 (n_1065, A[14], n_357);
  nand g952 (n_381, n_1063, n_1064, n_1065);
  xor g953 (n_1066, n_358, A[17]);
  xor g954 (n_361, n_1066, A[18]);
  nand g955 (n_1067, n_358, A[17]);
  nand g956 (n_1068, A[18], A[17]);
  nand g957 (n_1069, n_358, A[18]);
  nand g958 (n_383, n_1067, n_1068, n_1069);
  xor g959 (n_1070, n_359, n_360);
  xor g960 (n_363, n_1070, n_361);
  nand g961 (n_1071, n_359, n_360);
  nand g962 (n_1072, n_361, n_360);
  nand g963 (n_1073, n_359, n_361);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, A[21], n_362);
  xor g966 (n_365, n_1074, A[22]);
  nand g967 (n_1075, A[21], n_362);
  nand g968 (n_1076, A[22], n_362);
  nand g969 (n_1077, A[21], A[22]);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g971 (n_1078, n_363, n_364);
  nand g973 (n_1079, n_363, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  xor g986 (n_372, n_1086, A[3]);
  nand g990 (n_392, n_1044, n_1088, n_627);
  xor g991 (n_1090, n_371, n_372);
  xor g992 (n_374, n_1090, A[6]);
  nand g993 (n_1091, n_371, n_372);
  nand g994 (n_1092, A[6], n_372);
  nand g995 (n_1093, n_371, A[6]);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, n_374);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, n_374, n_373);
  nand g1001 (n_1097, A[7], n_374);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, A[10], A[11]);
  xor g1004 (n_378, n_1098, n_375);
  nand g1005 (n_1099, A[10], A[11]);
  nand g1006 (n_1100, n_375, A[11]);
  nand g1007 (n_1101, A[10], n_375);
  nand g1008 (n_398, n_1099, n_1100, n_1101);
  xor g1009 (n_1102, n_376, n_377);
  xor g1010 (n_380, n_1102, n_378);
  nand g1011 (n_1103, n_376, n_377);
  nand g1012 (n_1104, n_378, n_377);
  nand g1013 (n_1105, n_376, n_378);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, A[14], A[15]);
  xor g1016 (n_382, n_1106, n_379);
  nand g1017 (n_1107, A[14], A[15]);
  nand g1018 (n_1108, n_379, A[15]);
  nand g1019 (n_1109, A[14], n_379);
  nand g1020 (n_402, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, n_380, A[18]);
  xor g1022 (n_384, n_1110, n_381);
  nand g1023 (n_1111, n_380, A[18]);
  nand g1024 (n_1112, n_381, A[18]);
  nand g1025 (n_1113, n_380, n_381);
  nand g1026 (n_404, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, n_382, A[19]);
  xor g1028 (n_386, n_1114, n_383);
  nand g1029 (n_1115, n_382, A[19]);
  nand g1030 (n_1116, n_383, A[19]);
  nand g1031 (n_1117, n_382, n_383);
  nand g1032 (n_406, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_384, A[22]);
  xor g1034 (n_388, n_1118, n_385);
  nand g1035 (n_1119, n_384, A[22]);
  nand g1036 (n_1120, n_385, A[22]);
  nand g1037 (n_1121, n_384, n_385);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, n_386, A[23]);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, n_386, A[23]);
  nand g1042 (n_1124, n_387, A[23]);
  nand g1043 (n_1125, n_386, n_387);
  nand g1044 (n_410, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1051 (n_1130, A[1], A[3]);
  xor g1052 (n_393, n_1130, A[4]);
  nand g1053 (n_1131, A[1], A[3]);
  nand g1054 (n_1132, A[4], A[3]);
  nand g1055 (n_1133, A[1], A[4]);
  nand g1056 (n_412, n_1131, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, n_396, A[11]);
  xor g1070 (n_399, n_1142, A[12]);
  nand g1071 (n_1143, n_396, A[11]);
  nand g1072 (n_1144, A[12], A[11]);
  nand g1073 (n_1145, n_396, A[12]);
  nand g1074 (n_418, n_1143, n_1144, n_1145);
  xor g1075 (n_1146, n_397, n_398);
  xor g1076 (n_401, n_1146, n_399);
  nand g1077 (n_1147, n_397, n_398);
  nand g1078 (n_1148, n_399, n_398);
  nand g1079 (n_1149, n_397, n_399);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, A[15], n_400);
  xor g1082 (n_403, n_1150, A[16]);
  nand g1083 (n_1151, A[15], n_400);
  nand g1084 (n_1152, A[16], n_400);
  nand g1086 (n_421, n_1151, n_1152, n_984);
  xor g1087 (n_1154, n_401, n_402);
  xor g1088 (n_405, n_1154, A[19]);
  nand g1089 (n_1155, n_401, n_402);
  nand g1090 (n_1156, A[19], n_402);
  nand g1091 (n_1157, n_401, A[19]);
  nand g1092 (n_424, n_1155, n_1156, n_1157);
  xor g1093 (n_1158, n_403, n_404);
  xor g1094 (n_407, n_1158, A[20]);
  nand g1095 (n_1159, n_403, n_404);
  nand g1096 (n_1160, A[20], n_404);
  nand g1097 (n_1161, n_403, A[20]);
  nand g1098 (n_425, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_405, n_406);
  xor g1100 (n_409, n_1162, n_407);
  nand g1101 (n_1163, n_405, n_406);
  nand g1102 (n_1164, n_407, n_406);
  nand g1103 (n_1165, n_405, n_407);
  nand g1104 (n_428, n_1163, n_1164, n_1165);
  xor g1106 (n_411, n_1166, n_408);
  nand g1108 (n_1168, n_408, A[23]);
  nand g1110 (n_430, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1123 (n_1178, A[8], n_413);
  xor g1124 (n_415, n_1178, A[9]);
  nand g1125 (n_1179, A[8], n_413);
  nand g1126 (n_1180, A[9], n_413);
  nand g1128 (n_435, n_1179, n_1180, n_687);
  xor g1129 (n_1182, n_414, n_415);
  xor g1130 (n_417, n_1182, A[12]);
  nand g1131 (n_1183, n_414, n_415);
  nand g1132 (n_1184, A[12], n_415);
  nand g1133 (n_1185, n_414, A[12]);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, n_416, A[13]);
  xor g1136 (n_420, n_1186, n_417);
  nand g1137 (n_1187, n_416, A[13]);
  nand g1138 (n_1188, n_417, A[13]);
  nand g1139 (n_1189, n_416, n_417);
  nand g1140 (n_439, n_1187, n_1188, n_1189);
  xor g1141 (n_1190, n_418, n_419);
  xor g1142 (n_422, n_1190, A[16]);
  nand g1143 (n_1191, n_418, n_419);
  nand g1144 (n_1192, A[16], n_419);
  nand g1145 (n_1193, n_418, A[16]);
  nand g1146 (n_440, n_1191, n_1192, n_1193);
  xor g1147 (n_1194, n_420, A[17]);
  xor g1148 (n_423, n_1194, n_421);
  nand g1149 (n_1195, n_420, A[17]);
  nand g1150 (n_1196, n_421, A[17]);
  nand g1151 (n_1197, n_420, n_421);
  nand g1152 (n_442, n_1195, n_1196, n_1197);
  xor g1153 (n_1198, n_422, A[20]);
  xor g1154 (n_426, n_1198, n_423);
  nand g1155 (n_1199, n_422, A[20]);
  nand g1156 (n_1200, n_423, A[20]);
  nand g1157 (n_1201, n_422, n_423);
  nand g1158 (n_445, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_424, A[21]);
  xor g1160 (n_427, n_1202, n_425);
  nand g1161 (n_1203, n_424, A[21]);
  nand g1162 (n_1204, n_425, A[21]);
  nand g1163 (n_1205, n_424, n_425);
  nand g1164 (n_447, n_1203, n_1204, n_1205);
  xor g1166 (n_429, n_1206, n_427);
  nand g1168 (n_1208, n_427, n_426);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, n_433);
  nand g1183 (n_1217, A[6], n_433);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, A[9], A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, A[9], A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, A[9], n_434);
  nand g1190 (n_455, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, n_435, n_436);
  xor g1192 (n_438, n_1222, A[13]);
  nand g1193 (n_1223, n_435, n_436);
  nand g1194 (n_1224, A[13], n_436);
  nand g1195 (n_1225, n_435, A[13]);
  nand g1196 (n_457, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, A[14], n_437);
  xor g1198 (n_441, n_1226, n_438);
  nand g1199 (n_1227, A[14], n_437);
  nand g1200 (n_1228, n_438, n_437);
  nand g1201 (n_1229, A[14], n_438);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, n_439, A[17]);
  xor g1204 (n_443, n_1230, n_440);
  nand g1205 (n_1231, n_439, A[17]);
  nand g1206 (n_1232, n_440, A[17]);
  nand g1207 (n_1233, n_439, n_440);
  nand g1208 (n_461, n_1231, n_1232, n_1233);
  xor g1209 (n_1234, A[18], n_441);
  xor g1210 (n_444, n_1234, n_442);
  nand g1211 (n_1235, A[18], n_441);
  nand g1212 (n_1236, n_442, n_441);
  nand g1213 (n_1237, A[18], n_442);
  nand g1214 (n_464, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_443, A[21]);
  xor g1216 (n_446, n_1238, A[22]);
  nand g1217 (n_1239, n_443, A[21]);
  nand g1219 (n_1241, n_443, A[22]);
  nand g1220 (n_465, n_1239, n_1077, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[5], A[7]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], n_453);
  xor g1242 (n_456, n_1254, n_454);
  nand g1243 (n_1255, A[10], n_453);
  nand g1244 (n_1256, n_454, n_453);
  nand g1245 (n_1257, A[10], n_454);
  nand g1246 (n_472, n_1255, n_1256, n_1257);
  xor g1247 (n_1258, A[11], n_455);
  xor g1248 (n_458, n_1258, n_456);
  nand g1249 (n_1259, A[11], n_455);
  nand g1250 (n_1260, n_456, n_455);
  nand g1251 (n_1261, A[11], n_456);
  nand g1252 (n_474, n_1259, n_1260, n_1261);
  xor g1253 (n_1262, A[14], n_457);
  xor g1254 (n_460, n_1262, A[15]);
  nand g1255 (n_1263, A[14], n_457);
  nand g1256 (n_1264, A[15], n_457);
  nand g1258 (n_476, n_1263, n_1264, n_1107);
  xor g1259 (n_1266, n_458, A[18]);
  xor g1260 (n_462, n_1266, n_459);
  nand g1261 (n_1267, n_458, A[18]);
  nand g1262 (n_1268, n_459, A[18]);
  nand g1263 (n_1269, n_458, n_459);
  nand g1264 (n_479, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, n_460, A[19]);
  xor g1266 (n_463, n_1270, n_461);
  nand g1267 (n_1271, n_460, A[19]);
  nand g1268 (n_1272, n_461, A[19]);
  nand g1269 (n_1273, n_460, n_461);
  nand g1270 (n_480, n_1271, n_1272, n_1273);
  xor g1271 (n_1274, n_462, A[22]);
  xor g1272 (n_466, n_1274, n_463);
  nand g1273 (n_1275, n_462, A[22]);
  nand g1274 (n_1276, n_463, A[22]);
  nand g1275 (n_1277, n_462, n_463);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1277 (n_1278, n_464, A[23]);
  xor g1278 (n_467, n_1278, n_465);
  nand g1279 (n_1279, n_464, A[23]);
  nand g1280 (n_1280, n_465, A[23]);
  nand g1281 (n_1281, n_464, n_465);
  nand g1282 (n_484, n_1279, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1290 (n_471, n_738, A[6]);
  nand g1294 (n_486, n_673, n_651, n_660);
  xor g1295 (n_1290, n_470, A[11]);
  xor g1296 (n_473, n_1290, n_471);
  nand g1297 (n_1291, n_470, A[11]);
  nand g1298 (n_1292, n_471, A[11]);
  nand g1299 (n_1293, n_470, n_471);
  nand g1300 (n_488, n_1291, n_1292, n_1293);
  xor g1301 (n_1294, A[12], n_472);
  xor g1302 (n_475, n_1294, n_473);
  nand g1303 (n_1295, A[12], n_472);
  nand g1304 (n_1296, n_473, n_472);
  nand g1305 (n_1297, A[12], n_473);
  nand g1306 (n_490, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, A[15], n_474);
  xor g1308 (n_477, n_1298, n_475);
  nand g1309 (n_1299, A[15], n_474);
  nand g1310 (n_1300, n_475, n_474);
  nand g1311 (n_1301, A[15], n_475);
  nand g1312 (n_491, n_1299, n_1300, n_1301);
  xor g1313 (n_1302, A[16], n_476);
  xor g1314 (n_478, n_1302, n_477);
  nand g1315 (n_1303, A[16], n_476);
  nand g1316 (n_1304, n_477, n_476);
  nand g1317 (n_1305, A[16], n_477);
  nand g1318 (n_494, n_1303, n_1304, n_1305);
  xor g1319 (n_1306, A[19], n_478);
  xor g1320 (n_481, n_1306, n_479);
  nand g1321 (n_1307, A[19], n_478);
  nand g1322 (n_1308, n_479, n_478);
  nand g1323 (n_1309, A[19], n_479);
  nand g1324 (n_495, n_1307, n_1308, n_1309);
  xor g1325 (n_1310, A[20], n_480);
  xor g1326 (n_483, n_1310, n_481);
  nand g1327 (n_1311, A[20], n_480);
  nand g1328 (n_1312, n_481, n_480);
  nand g1329 (n_1313, A[20], n_481);
  nand g1330 (n_498, n_1311, n_1312, n_1313);
  xor g1332 (n_485, n_1166, n_482);
  nand g1335 (n_1317, A[23], n_482);
  nand g1336 (n_500, n_1167, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1344 (n_487, n_686, n_486);
  nand g1346 (n_1324, n_486, A[9]);
  nand g1347 (n_1325, A[8], n_486);
  nand g1348 (n_503, n_687, n_1324, n_1325);
  xor g1349 (n_1326, A[12], n_487);
  xor g1350 (n_489, n_1326, n_488);
  nand g1351 (n_1327, A[12], n_487);
  nand g1352 (n_1328, n_488, n_487);
  nand g1353 (n_1329, A[12], n_488);
  nand g1354 (n_505, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, A[13], n_489);
  xor g1356 (n_492, n_1330, A[16]);
  nand g1357 (n_1331, A[13], n_489);
  nand g1358 (n_1332, A[16], n_489);
  nand g1359 (n_1333, A[13], A[16]);
  nand g1360 (n_507, n_1331, n_1332, n_1333);
  xor g1361 (n_1334, n_490, A[17]);
  xor g1362 (n_493, n_1334, n_491);
  nand g1363 (n_1335, n_490, A[17]);
  nand g1364 (n_1336, n_491, A[17]);
  nand g1365 (n_1337, n_490, n_491);
  nand g1366 (n_509, n_1335, n_1336, n_1337);
  xor g1367 (n_1338, n_492, A[20]);
  xor g1368 (n_496, n_1338, n_493);
  nand g1369 (n_1339, n_492, A[20]);
  nand g1370 (n_1340, n_493, A[20]);
  nand g1371 (n_1341, n_492, n_493);
  nand g1372 (n_511, n_1339, n_1340, n_1341);
  xor g1373 (n_1342, n_494, A[21]);
  xor g1374 (n_497, n_1342, n_495);
  nand g1375 (n_1343, n_494, A[21]);
  nand g1376 (n_1344, n_495, A[21]);
  nand g1377 (n_1345, n_494, n_495);
  nand g1378 (n_513, n_1343, n_1344, n_1345);
  xor g1380 (n_499, n_1346, n_497);
  nand g1383 (n_1349, n_496, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  nand g1397 (n_1357, A[10], n_503);
  nand g1398 (n_520, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], A[14]);
  xor g1400 (n_506, n_1358, n_504);
  nand g1402 (n_1360, n_504, A[14]);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_521, n_912, n_1360, n_1361);
  xor g1405 (n_1362, n_505, A[17]);
  xor g1406 (n_508, n_1362, n_506);
  nand g1407 (n_1363, n_505, A[17]);
  nand g1408 (n_1364, n_506, A[17]);
  nand g1409 (n_1365, n_505, n_506);
  nand g1410 (n_523, n_1363, n_1364, n_1365);
  xor g1411 (n_1366, A[18], n_507);
  xor g1412 (n_510, n_1366, n_508);
  nand g1413 (n_1367, A[18], n_507);
  nand g1414 (n_1368, n_508, n_507);
  nand g1415 (n_1369, A[18], n_508);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_509, A[21]);
  xor g1418 (n_512, n_1370, n_510);
  nand g1419 (n_1371, n_509, A[21]);
  nand g1420 (n_1372, n_510, A[21]);
  nand g1421 (n_1373, n_509, n_510);
  nand g1422 (n_527, n_1371, n_1372, n_1373);
  xor g1423 (n_1374, A[22], n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, A[22], n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, A[22], n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1437 (n_1382, A[9], A[11]);
  nand g1439 (n_1383, A[9], A[11]);
  nand g1442 (n_532, n_1383, n_1384, n_1385);
  xor g1443 (n_1386, A[14], n_519);
  xor g1444 (n_522, n_1386, n_520);
  nand g1445 (n_1387, A[14], n_519);
  nand g1446 (n_1388, n_520, n_519);
  nand g1447 (n_1389, A[14], n_520);
  nand g1448 (n_534, n_1387, n_1388, n_1389);
  xor g1449 (n_1390, A[15], n_521);
  xor g1450 (n_524, n_1390, n_522);
  nand g1451 (n_1391, A[15], n_521);
  nand g1452 (n_1392, n_522, n_521);
  nand g1453 (n_1393, A[15], n_522);
  nand g1454 (n_536, n_1391, n_1392, n_1393);
  xor g1455 (n_1394, A[18], n_523);
  xor g1456 (n_525, n_1394, A[19]);
  nand g1457 (n_1395, A[18], n_523);
  nand g1458 (n_1396, A[19], n_523);
  nand g1459 (n_1397, A[18], A[19]);
  nand g1460 (n_538, n_1395, n_1396, n_1397);
  xor g1461 (n_1398, n_524, n_525);
  xor g1462 (n_528, n_1398, n_526);
  nand g1463 (n_1399, n_524, n_525);
  nand g1464 (n_1400, n_526, n_525);
  nand g1465 (n_1401, n_524, n_526);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1467 (n_1402, A[22], A[23]);
  xor g1468 (n_529, n_1402, n_527);
  nand g1469 (n_1403, A[22], A[23]);
  nand g1470 (n_1404, n_527, A[23]);
  nand g1471 (n_1405, A[22], n_527);
  nand g1472 (n_543, n_1403, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1479 (n_1410, A[11], A[12]);
  xor g1480 (n_533, n_1410, A[10]);
  nand g1484 (n_544, n_1144, n_709, n_1099);
  xor g1485 (n_1414, n_532, n_533);
  xor g1486 (n_535, n_1414, A[15]);
  nand g1487 (n_1415, n_532, n_533);
  nand g1488 (n_1416, A[15], n_533);
  nand g1489 (n_1417, n_532, A[15]);
  nand g1490 (n_546, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, A[16], n_534);
  xor g1492 (n_537, n_1418, n_535);
  nand g1493 (n_1419, A[16], n_534);
  nand g1494 (n_1420, n_535, n_534);
  nand g1495 (n_1421, A[16], n_535);
  nand g1496 (n_548, n_1419, n_1420, n_1421);
  xor g1497 (n_1422, A[19], n_536);
  xor g1498 (n_539, n_1422, n_537);
  nand g1499 (n_1423, A[19], n_536);
  nand g1500 (n_1424, n_537, n_536);
  nand g1501 (n_1425, A[19], n_537);
  nand g1502 (n_549, n_1423, n_1424, n_1425);
  xor g1503 (n_1426, A[20], n_538);
  xor g1504 (n_541, n_1426, n_539);
  nand g1505 (n_1427, A[20], n_538);
  nand g1506 (n_1428, n_539, n_538);
  nand g1507 (n_1429, A[20], n_539);
  nand g1508 (n_551, n_1427, n_1428, n_1429);
  xor g1510 (n_542, n_1166, n_540);
  nand g1513 (n_1433, A[23], n_540);
  nand g1514 (n_554, n_1167, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1521 (n_1438, A[12], A[13]);
  xor g1522 (n_545, n_1438, n_544);
  nand g1523 (n_1439, A[12], A[13]);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_1439, n_1440, n_1441);
  xor g1527 (n_1442, A[16], n_545);
  xor g1528 (n_547, n_1442, A[17]);
  nand g1529 (n_1443, A[16], n_545);
  nand g1530 (n_1444, A[17], n_545);
  nand g1531 (n_1445, A[16], A[17]);
  nand g1532 (n_559, n_1443, n_1444, n_1445);
  xor g1533 (n_1446, n_546, n_547);
  xor g1534 (n_550, n_1446, n_548);
  nand g1535 (n_1447, n_546, n_547);
  nand g1536 (n_1448, n_548, n_547);
  nand g1537 (n_1449, n_546, n_548);
  nand g1538 (n_561, n_1447, n_1448, n_1449);
  xor g1539 (n_1450, A[20], A[21]);
  xor g1540 (n_552, n_1450, n_549);
  nand g1541 (n_1451, A[20], A[21]);
  nand g1542 (n_1452, n_549, A[21]);
  nand g1543 (n_1453, A[20], n_549);
  nand g1544 (n_562, n_1451, n_1452, n_1453);
  xor g1546 (n_553, n_1454, n_551);
  nand g1549 (n_1457, n_550, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1563 (n_1465, A[14], n_557);
  nand g1564 (n_569, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, A[17], A[18]);
  xor g1566 (n_560, n_1466, n_558);
  nand g1568 (n_1468, n_558, A[18]);
  nand g1569 (n_1469, A[17], n_558);
  nand g1570 (n_571, n_1068, n_1468, n_1469);
  xor g1571 (n_1470, n_559, n_560);
  xor g1572 (n_563, n_1470, A[21]);
  nand g1573 (n_1471, n_559, n_560);
  nand g1574 (n_1472, A[21], n_560);
  nand g1575 (n_1473, n_559, A[21]);
  nand g1576 (n_574, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, A[22], n_561);
  xor g1578 (n_564, n_1474, n_562);
  nand g1579 (n_1475, A[22], n_561);
  nand g1580 (n_1476, n_562, n_561);
  nand g1581 (n_1477, A[22], n_562);
  nand g1582 (n_576, n_1475, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  xor g1591 (n_1482, A[13], A[15]);
  nand g1593 (n_1483, A[13], A[15]);
  nand g1596 (n_578, n_1483, n_1484, n_1485);
  xor g1597 (n_1486, A[18], n_569);
  xor g1598 (n_572, n_1486, n_570);
  nand g1599 (n_1487, A[18], n_569);
  nand g1600 (n_1488, n_570, n_569);
  nand g1601 (n_1489, A[18], n_570);
  nand g1602 (n_580, n_1487, n_1488, n_1489);
  xor g1603 (n_1490, A[19], n_571);
  xor g1604 (n_573, n_1490, n_572);
  nand g1605 (n_1491, A[19], n_571);
  nand g1606 (n_1492, n_572, n_571);
  nand g1607 (n_1493, A[19], n_572);
  nand g1608 (n_582, n_1491, n_1492, n_1493);
  xor g1609 (n_1494, A[22], n_573);
  xor g1610 (n_575, n_1494, A[23]);
  nand g1611 (n_1495, A[22], n_573);
  nand g1612 (n_1496, A[23], n_573);
  nand g1614 (n_584, n_1495, n_1496, n_1403);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1622 (n_579, n_1106, A[16]);
  nand g1626 (n_586, n_1107, n_801, n_984);
  xor g1627 (n_1506, n_578, n_579);
  xor g1628 (n_581, n_1506, A[19]);
  nand g1629 (n_1507, n_578, n_579);
  nand g1630 (n_1508, A[19], n_579);
  nand g1631 (n_1509, n_578, A[19]);
  nand g1632 (n_588, n_1507, n_1508, n_1509);
  xor g1633 (n_1510, n_580, A[20]);
  xor g1634 (n_583, n_1510, n_581);
  nand g1635 (n_1511, n_580, A[20]);
  nand g1636 (n_1512, n_581, A[20]);
  nand g1637 (n_1513, n_580, n_581);
  nand g1638 (n_589, n_1511, n_1512, n_1513);
  xor g1639 (n_1514, n_582, n_583);
  xor g1640 (n_585, n_1514, A[23]);
  nand g1641 (n_1515, n_582, n_583);
  nand g1642 (n_1516, A[23], n_583);
  nand g1643 (n_1517, n_582, A[23]);
  nand g1644 (n_591, n_1515, n_1516, n_1517);
  xor g1646 (n_83, n_1518, n_585);
  nand g1648 (n_1520, n_585, n_584);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1651 (n_1522, A[16], A[17]);
  xor g1652 (n_587, n_1522, n_586);
  nand g1654 (n_1524, n_586, A[17]);
  nand g1655 (n_1525, A[16], n_586);
  nand g1656 (n_595, n_1445, n_1524, n_1525);
  xor g1657 (n_1526, A[20], n_587);
  xor g1658 (n_590, n_1526, n_588);
  nand g1659 (n_1527, A[20], n_587);
  nand g1660 (n_1528, n_588, n_587);
  nand g1661 (n_1529, A[20], n_588);
  nand g1662 (n_597, n_1527, n_1528, n_1529);
  xor g1664 (n_592, n_1530, n_589);
  nand g1667 (n_1533, A[21], n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_81, n_1535, n_1536, n_1537);
  nand g1681 (n_1541, A[18], n_595);
  nand g1682 (n_604, n_1539, n_1540, n_1541);
  xor g1683 (n_1542, A[21], A[22]);
  xor g1684 (n_598, n_1542, n_596);
  nand g1686 (n_1544, n_596, A[22]);
  nand g1687 (n_1545, A[21], n_596);
  nand g1688 (n_606, n_1077, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_33, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[17], A[19]);
  nand g1702 (n_608, n_889, n_1552, n_1553);
  xor g1703 (n_1554, A[22], n_603);
  xor g1704 (n_605, n_1554, n_604);
  nand g1705 (n_1555, A[22], n_603);
  nand g1706 (n_1556, n_604, n_603);
  nand g1707 (n_1557, A[22], n_604);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, A[23], n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, A[23], n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, A[23], n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1715 (n_1562, A[19], A[18]);
  xor g1716 (n_609, n_1562, A[20]);
  nand g1719 (n_1565, A[19], A[20]);
  nand g1720 (n_612, n_1397, n_925, n_1565);
  xor g1721 (n_1566, n_608, n_609);
  xor g1722 (n_611, n_1566, A[23]);
  nand g1723 (n_1567, n_608, n_609);
  nand g1724 (n_1568, A[23], n_609);
  nand g1725 (n_1569, n_608, A[23]);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1728 (n_79, n_1570, n_611);
  nand g1730 (n_1572, n_611, n_610);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1734 (n_613, n_1450, n_612);
  nand g1736 (n_1576, n_612, A[21]);
  nand g1737 (n_1577, A[20], n_612);
  nand g1738 (n_617, n_1451, n_1576, n_1577);
  xor g1740 (n_78, n_1578, n_614);
  nand g1742 (n_1580, n_614, n_613);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_617);
  nand g1752 (n_76, n_1583, n_1584, n_1585);
  nand g1759 (n_1589, A[21], A[23]);
  nand g1760 (n_27, n_1587, n_1588, n_1589);
  xor g1762 (n_75, n_1166, A[22]);
  nand g1766 (n_74, n_1167, n_1403, n_1593);
  nand g16 (n_1606, A[0], A[2]);
  xor g20 (Z[2], A[0], A[2]);
  nand g22 (n_1611, n_69, A[3]);
  nand g25 (n_1615, n_1611, n_1612, n_1613);
  xor g26 (n_1614, n_69, A[3]);
  nand g28 (n_1616, A[4], n_117);
  nand g29 (n_1617, A[4], n_1615);
  nand g30 (n_1618, n_117, n_1615);
  nand g31 (n_1620, n_1616, n_1617, n_1618);
  xor g32 (n_1619, A[4], n_117);
  xor g33 (Z[4], n_1615, n_1619);
  nand g34 (n_1621, A[5], n_116);
  nand g35 (n_1622, A[5], n_1620);
  nand g36 (n_1623, n_116, n_1620);
  nand g37 (n_1625, n_1621, n_1622, n_1623);
  xor g38 (n_1624, A[5], n_116);
  xor g39 (Z[5], n_1620, n_1624);
  nand g40 (n_1626, A[6], n_115);
  nand g41 (n_1627, A[6], n_1625);
  nand g42 (n_1628, n_115, n_1625);
  nand g43 (n_1630, n_1626, n_1627, n_1628);
  xor g44 (n_1629, A[6], n_115);
  xor g45 (Z[6], n_1625, n_1629);
  nand g46 (n_1631, n_66, n_114);
  nand g47 (n_1632, n_66, n_1630);
  nand g48 (n_1633, n_114, n_1630);
  nand g49 (n_1635, n_1631, n_1632, n_1633);
  xor g50 (n_1634, n_66, n_114);
  xor g51 (Z[7], n_1630, n_1634);
  nand g52 (n_1636, n_65, n_113);
  nand g53 (n_1637, n_65, n_1635);
  nand g54 (n_1638, n_113, n_1635);
  nand g55 (n_1640, n_1636, n_1637, n_1638);
  xor g56 (n_1639, n_65, n_113);
  xor g57 (Z[8], n_1635, n_1639);
  nand g58 (n_1641, n_64, n_112);
  nand g59 (n_1642, n_64, n_1640);
  nand g60 (n_1643, n_112, n_1640);
  nand g61 (n_1645, n_1641, n_1642, n_1643);
  xor g62 (n_1644, n_64, n_112);
  xor g63 (Z[9], n_1640, n_1644);
  nand g64 (n_1646, n_63, n_111);
  nand g65 (n_1647, n_63, n_1645);
  nand g66 (n_1648, n_111, n_1645);
  nand g67 (n_1650, n_1646, n_1647, n_1648);
  xor g68 (n_1649, n_63, n_111);
  xor g69 (Z[10], n_1645, n_1649);
  nand g70 (n_1651, n_62, n_110);
  nand g71 (n_1652, n_62, n_1650);
  nand g72 (n_1653, n_110, n_1650);
  nand g73 (n_1655, n_1651, n_1652, n_1653);
  xor g74 (n_1654, n_62, n_110);
  xor g75 (Z[11], n_1650, n_1654);
  nand g76 (n_1656, n_61, n_109);
  nand g77 (n_1657, n_61, n_1655);
  nand g78 (n_1658, n_109, n_1655);
  nand g79 (n_1660, n_1656, n_1657, n_1658);
  xor g80 (n_1659, n_61, n_109);
  xor g81 (Z[12], n_1655, n_1659);
  nand g82 (n_1661, n_60, n_108);
  nand g83 (n_1662, n_60, n_1660);
  nand g84 (n_1663, n_108, n_1660);
  nand g85 (n_1665, n_1661, n_1662, n_1663);
  xor g86 (n_1664, n_60, n_108);
  xor g87 (Z[13], n_1660, n_1664);
  nand g88 (n_1666, n_59, n_107);
  nand g89 (n_1667, n_59, n_1665);
  nand g90 (n_1668, n_107, n_1665);
  nand g91 (n_1670, n_1666, n_1667, n_1668);
  xor g92 (n_1669, n_59, n_107);
  xor g93 (Z[14], n_1665, n_1669);
  nand g94 (n_1671, n_58, n_106);
  nand g95 (n_1672, n_58, n_1670);
  nand g96 (n_1673, n_106, n_1670);
  nand g97 (n_1675, n_1671, n_1672, n_1673);
  xor g98 (n_1674, n_58, n_106);
  xor g99 (Z[15], n_1670, n_1674);
  nand g100 (n_1676, n_57, n_105);
  nand g101 (n_1677, n_57, n_1675);
  nand g102 (n_1678, n_105, n_1675);
  nand g103 (n_1680, n_1676, n_1677, n_1678);
  xor g104 (n_1679, n_57, n_105);
  xor g105 (Z[16], n_1675, n_1679);
  nand g106 (n_1681, n_56, n_104);
  nand g107 (n_1682, n_56, n_1680);
  nand g108 (n_1683, n_104, n_1680);
  nand g109 (n_1685, n_1681, n_1682, n_1683);
  xor g110 (n_1684, n_56, n_104);
  xor g111 (Z[17], n_1680, n_1684);
  nand g112 (n_1686, n_55, n_103);
  nand g113 (n_1687, n_55, n_1685);
  nand g114 (n_1688, n_103, n_1685);
  nand g115 (n_1690, n_1686, n_1687, n_1688);
  xor g116 (n_1689, n_55, n_103);
  xor g117 (Z[18], n_1685, n_1689);
  nand g118 (n_1691, n_54, n_102);
  nand g119 (n_1692, n_54, n_1690);
  nand g120 (n_1693, n_102, n_1690);
  nand g121 (n_1695, n_1691, n_1692, n_1693);
  xor g122 (n_1694, n_54, n_102);
  xor g123 (Z[19], n_1690, n_1694);
  nand g124 (n_1696, n_53, n_101);
  nand g125 (n_1697, n_53, n_1695);
  nand g126 (n_1698, n_101, n_1695);
  nand g127 (n_1700, n_1696, n_1697, n_1698);
  xor g128 (n_1699, n_53, n_101);
  xor g129 (Z[20], n_1695, n_1699);
  nand g130 (n_1701, n_52, n_100);
  nand g131 (n_1702, n_52, n_1700);
  nand g132 (n_1703, n_100, n_1700);
  nand g133 (n_1705, n_1701, n_1702, n_1703);
  xor g134 (n_1704, n_52, n_100);
  xor g135 (Z[21], n_1700, n_1704);
  nand g136 (n_1706, n_51, n_99);
  nand g137 (n_1707, n_51, n_1705);
  nand g138 (n_1708, n_99, n_1705);
  nand g139 (n_1710, n_1706, n_1707, n_1708);
  xor g140 (n_1709, n_51, n_99);
  xor g141 (Z[22], n_1705, n_1709);
  nand g142 (n_1711, n_50, n_98);
  nand g143 (n_1712, n_50, n_1710);
  nand g144 (n_1713, n_98, n_1710);
  nand g145 (n_1715, n_1711, n_1712, n_1713);
  xor g146 (n_1714, n_50, n_98);
  xor g147 (Z[23], n_1710, n_1714);
  nand g148 (n_1716, n_49, n_97);
  nand g149 (n_1717, n_49, n_1715);
  nand g150 (n_1718, n_97, n_1715);
  nand g151 (n_1720, n_1716, n_1717, n_1718);
  xor g152 (n_1719, n_49, n_97);
  xor g153 (Z[24], n_1715, n_1719);
  nand g154 (n_1721, n_48, n_96);
  nand g155 (n_1722, n_48, n_1720);
  nand g156 (n_1723, n_96, n_1720);
  nand g157 (n_1725, n_1721, n_1722, n_1723);
  xor g158 (n_1724, n_48, n_96);
  xor g159 (Z[25], n_1720, n_1724);
  nand g160 (n_1726, n_47, n_95);
  nand g161 (n_1727, n_47, n_1725);
  nand g162 (n_1728, n_95, n_1725);
  nand g163 (n_1730, n_1726, n_1727, n_1728);
  xor g164 (n_1729, n_47, n_95);
  xor g165 (Z[26], n_1725, n_1729);
  nand g166 (n_1731, n_46, n_94);
  nand g167 (n_1732, n_46, n_1730);
  nand g168 (n_1733, n_94, n_1730);
  nand g169 (n_1735, n_1731, n_1732, n_1733);
  xor g170 (n_1734, n_46, n_94);
  xor g171 (Z[27], n_1730, n_1734);
  nand g172 (n_1736, n_45, n_93);
  nand g173 (n_1737, n_45, n_1735);
  nand g174 (n_1738, n_93, n_1735);
  nand g175 (n_1740, n_1736, n_1737, n_1738);
  xor g176 (n_1739, n_45, n_93);
  xor g177 (Z[28], n_1735, n_1739);
  nand g178 (n_1741, n_44, n_92);
  nand g179 (n_1742, n_44, n_1740);
  nand g180 (n_1743, n_92, n_1740);
  nand g181 (n_1745, n_1741, n_1742, n_1743);
  xor g182 (n_1744, n_44, n_92);
  xor g183 (Z[29], n_1740, n_1744);
  nand g184 (n_1746, n_43, n_91);
  nand g185 (n_1747, n_43, n_1745);
  nand g186 (n_1748, n_91, n_1745);
  nand g187 (n_1750, n_1746, n_1747, n_1748);
  xor g188 (n_1749, n_43, n_91);
  xor g189 (Z[30], n_1745, n_1749);
  nand g190 (n_1751, n_42, n_90);
  nand g191 (n_1752, n_42, n_1750);
  nand g192 (n_1753, n_90, n_1750);
  nand g193 (n_1755, n_1751, n_1752, n_1753);
  xor g194 (n_1754, n_42, n_90);
  xor g195 (Z[31], n_1750, n_1754);
  nand g196 (n_1756, n_41, n_89);
  nand g197 (n_1757, n_41, n_1755);
  nand g198 (n_1758, n_89, n_1755);
  nand g199 (n_1760, n_1756, n_1757, n_1758);
  xor g200 (n_1759, n_41, n_89);
  xor g201 (Z[32], n_1755, n_1759);
  nand g202 (n_1761, n_40, n_88);
  nand g203 (n_1762, n_40, n_1760);
  nand g204 (n_1763, n_88, n_1760);
  nand g205 (n_1765, n_1761, n_1762, n_1763);
  xor g206 (n_1764, n_40, n_88);
  xor g207 (Z[33], n_1760, n_1764);
  nand g208 (n_1766, n_39, n_87);
  nand g209 (n_1767, n_39, n_1765);
  nand g210 (n_1768, n_87, n_1765);
  nand g211 (n_1770, n_1766, n_1767, n_1768);
  xor g212 (n_1769, n_39, n_87);
  xor g213 (Z[34], n_1765, n_1769);
  nand g214 (n_1771, n_38, n_86);
  nand g215 (n_1772, n_38, n_1770);
  nand g216 (n_1773, n_86, n_1770);
  nand g217 (n_1775, n_1771, n_1772, n_1773);
  xor g218 (n_1774, n_38, n_86);
  xor g219 (Z[35], n_1770, n_1774);
  nand g220 (n_1776, n_37, n_85);
  nand g221 (n_1777, n_37, n_1775);
  nand g222 (n_1778, n_85, n_1775);
  nand g223 (n_1780, n_1776, n_1777, n_1778);
  xor g224 (n_1779, n_37, n_85);
  xor g225 (Z[36], n_1775, n_1779);
  nand g226 (n_1781, n_36, n_84);
  nand g227 (n_1782, n_36, n_1780);
  nand g228 (n_1783, n_84, n_1780);
  nand g229 (n_1785, n_1781, n_1782, n_1783);
  xor g230 (n_1784, n_36, n_84);
  xor g231 (Z[37], n_1780, n_1784);
  nand g232 (n_1786, n_35, n_83);
  nand g233 (n_1787, n_35, n_1785);
  nand g234 (n_1788, n_83, n_1785);
  nand g235 (n_1790, n_1786, n_1787, n_1788);
  xor g236 (n_1789, n_35, n_83);
  xor g237 (Z[38], n_1785, n_1789);
  nand g238 (n_1791, n_34, n_82);
  nand g239 (n_1792, n_34, n_1790);
  nand g240 (n_1793, n_82, n_1790);
  nand g241 (n_1795, n_1791, n_1792, n_1793);
  xor g242 (n_1794, n_34, n_82);
  xor g243 (Z[39], n_1790, n_1794);
  nand g244 (n_1796, n_33, n_81);
  nand g245 (n_1797, n_33, n_1795);
  nand g246 (n_1798, n_81, n_1795);
  nand g247 (n_1800, n_1796, n_1797, n_1798);
  xor g248 (n_1799, n_33, n_81);
  xor g249 (Z[40], n_1795, n_1799);
  nand g250 (n_1801, n_32, n_80);
  nand g251 (n_1802, n_32, n_1800);
  nand g252 (n_1803, n_80, n_1800);
  nand g253 (n_1805, n_1801, n_1802, n_1803);
  xor g254 (n_1804, n_32, n_80);
  xor g255 (Z[41], n_1800, n_1804);
  nand g256 (n_1806, n_31, n_79);
  nand g257 (n_1807, n_31, n_1805);
  nand g258 (n_1808, n_79, n_1805);
  nand g259 (n_1810, n_1806, n_1807, n_1808);
  xor g260 (n_1809, n_31, n_79);
  xor g261 (Z[42], n_1805, n_1809);
  nand g262 (n_1811, n_30, n_78);
  nand g263 (n_1812, n_30, n_1810);
  nand g264 (n_1813, n_78, n_1810);
  nand g265 (n_1815, n_1811, n_1812, n_1813);
  xor g266 (n_1814, n_30, n_78);
  xor g267 (Z[43], n_1810, n_1814);
  nand g1772 (n_1816, n_29, n_77);
  nand g1773 (n_1817, n_29, n_1815);
  nand g1774 (n_1818, n_77, n_1815);
  nand g1775 (n_1820, n_1816, n_1817, n_1818);
  xor g1776 (n_1819, n_29, n_77);
  xor g1777 (Z[44], n_1815, n_1819);
  nand g1778 (n_1821, n_28, n_76);
  nand g1779 (n_1822, n_28, n_1820);
  nand g1780 (n_1823, n_76, n_1820);
  nand g1781 (n_1825, n_1821, n_1822, n_1823);
  xor g1782 (n_1824, n_28, n_76);
  xor g1783 (Z[45], n_1820, n_1824);
  nand g1784 (n_1826, n_27, n_75);
  nand g1785 (n_1827, n_27, n_1825);
  nand g1786 (n_1828, n_75, n_1825);
  nand g1787 (n_1830, n_1826, n_1827, n_1828);
  xor g1788 (n_1829, n_27, n_75);
  xor g1789 (Z[46], n_1825, n_1829);
  xor g1791 (Z[47], n_1830, n_1831);
  or g1804 (n_1043, A[1], wc);
  not gc (wc, n_171);
  or g1805 (n_1044, A[1], wc0);
  not gc0 (wc0, A[2]);
  xnor g1807 (n_1166, A[24], A[23]);
  or g1808 (n_1167, wc1, A[24]);
  not gc1 (wc1, A[23]);
  xnor g1809 (n_1214, A[6], A[5]);
  or g1810 (n_1215, A[5], wc2);
  not gc2 (wc2, A[6]);
  or g1811 (n_1252, A[6], wc3);
  not gc3 (wc3, A[7]);
  or g1812 (n_1253, wc4, A[6]);
  not gc4 (wc4, A[5]);
  or g1814 (n_1355, A[9], wc5);
  not gc5 (wc5, A[10]);
  or g1815 (n_1384, A[10], wc6);
  not gc6 (wc6, A[11]);
  or g1816 (n_1385, wc7, A[10]);
  not gc7 (wc7, A[9]);
  or g1818 (n_1463, A[13], wc8);
  not gc8 (wc8, A[14]);
  or g1819 (n_1484, A[14], wc9);
  not gc9 (wc9, A[15]);
  or g1820 (n_1485, wc10, A[14]);
  not gc10 (wc10, A[13]);
  xnor g1821 (n_1530, A[24], A[21]);
  or g1822 (n_1531, wc11, A[24]);
  not gc11 (wc11, A[21]);
  or g1824 (n_1539, A[17], wc12);
  not gc12 (wc12, A[18]);
  or g1825 (n_1552, A[18], wc13);
  not gc13 (wc13, A[19]);
  or g1826 (n_1553, wc14, A[18]);
  not gc14 (wc14, A[17]);
  or g1828 (n_1583, A[21], wc15);
  not gc15 (wc15, A[22]);
  or g1829 (n_1587, wc16, A[22]);
  not gc16 (wc16, A[21]);
  or g1830 (n_1588, A[22], wc17);
  not gc17 (wc17, A[23]);
  or g1831 (n_1593, wc18, A[24]);
  not gc18 (wc18, A[22]);
  xnor g1833 (n_1086, A[2], A[1]);
  or g1834 (n_1088, A[1], wc19);
  not gc19 (wc19, A[3]);
  xnor g1835 (n_453, n_1250, A[6]);
  xnor g1836 (n_519, n_1382, A[10]);
  xnor g1837 (n_570, n_1482, A[14]);
  xnor g1838 (n_603, n_1550, A[18]);
  xnor g1839 (n_28, n_1542, A[23]);
  or g1841 (n_1047, wc20, n_117);
  not gc20 (wc20, A[5]);
  or g1842 (n_1049, wc21, n_117);
  not gc21 (wc21, n_180);
  xnor g1844 (n_1578, n_613, A[24]);
  or g1845 (n_1579, A[24], wc22);
  not gc22 (wc22, n_613);
  xnor g1846 (n_1831, n_74, A[24]);
  or g1848 (n_1052, wc23, n_181);
  not gc23 (wc23, A[9]);
  or g1849 (n_1053, wc24, n_181);
  not gc24 (wc24, A[6]);
  xnor g1850 (n_504, n_1218, n_503);
  or g1851 (n_1356, A[9], wc25);
  not gc25 (wc25, n_503);
  xnor g1852 (n_558, n_1358, n_557);
  or g1853 (n_1464, A[13], wc26);
  not gc26 (wc26, n_557);
  xnor g1854 (n_596, n_1466, n_595);
  or g1855 (n_1540, A[17], wc27);
  not gc27 (wc27, n_595);
  or g1856 (n_1573, A[24], wc28);
  not gc28 (wc28, n_611);
  or g1857 (n_1581, A[24], wc29);
  not gc29 (wc29, n_614);
  xnor g1858 (n_29, n_1542, n_617);
  or g1859 (n_1584, A[21], wc30);
  not gc30 (wc30, n_617);
  xnor g1861 (n_355, n_203, n_906);
  or g1862 (n_1056, wc31, n_203);
  not gc31 (wc31, n_282);
  or g1863 (n_1057, wc32, n_203);
  not gc32 (wc32, A[10]);
  or g1864 (n_1216, A[5], wc33);
  not gc33 (wc33, n_433);
  or g1865 (n_1612, n_1606, wc34);
  not gc34 (wc34, n_69);
  or g1866 (n_1613, wc35, n_1606);
  not gc35 (wc35, A[3]);
  xnor g1867 (Z[3], n_1606, n_1614);
  xnor g1868 (n_1570, n_610, A[24]);
  or g1869 (n_1571, A[24], wc36);
  not gc36 (wc36, n_610);
  or g1870 (n_1532, A[24], wc37);
  not gc37 (wc37, n_589);
  xnor g1871 (n_1454, n_550, A[24]);
  or g1872 (n_1455, A[24], wc38);
  not gc38 (wc38, n_550);
  xnor g1873 (n_1518, n_584, A[24]);
  or g1874 (n_1519, A[24], wc39);
  not gc39 (wc39, n_584);
  or g1875 (n_1432, A[24], wc40);
  not gc40 (wc40, n_540);
  or g1876 (n_1521, A[24], wc41);
  not gc41 (wc41, n_585);
  or g1877 (n_1456, A[24], wc42);
  not gc42 (wc42, n_551);
  or g1878 (n_1081, A[24], wc43);
  not gc43 (wc43, n_363);
  or g1879 (n_1080, A[24], wc44);
  not gc44 (wc44, n_364);
  xnor g1880 (n_1206, n_426, A[24]);
  or g1881 (n_1207, A[24], wc45);
  not gc45 (wc45, n_426);
  xnor g1882 (n_1346, n_496, A[24]);
  or g1883 (n_1347, A[24], wc46);
  not gc46 (wc46, n_496);
  xnor g1884 (n_367, n_1078, A[24]);
  or g1885 (n_1348, A[24], wc47);
  not gc47 (wc47, n_497);
  or g1886 (n_1169, A[24], wc48);
  not gc48 (wc48, n_408);
  or g1887 (n_1209, A[24], wc49);
  not gc49 (wc49, n_427);
  or g1888 (n_1316, A[24], wc50);
  not gc50 (wc50, n_482);
endmodule

module mult_signed_const_4152_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_4152_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_4419_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_176;
  wire n_179, n_180, n_183, n_184, n_187, n_188, n_189, n_196;
  wire n_201, n_202, n_203, n_204, n_209, n_210, n_211, n_212;
  wire n_218, n_219, n_220, n_221, n_224, n_225, n_226, n_227;
  wire n_236, n_237, n_238, n_239, n_248, n_249, n_250, n_251;
  wire n_258, n_260, n_261, n_262, n_265, n_267, n_269, n_271;
  wire n_272, n_273, n_274, n_275, n_276, n_277, n_282, n_284;
  wire n_285, n_286, n_287, n_288, n_289, n_290, n_291, n_292;
  wire n_293, n_300, n_302, n_303, n_304, n_305, n_306, n_307;
  wire n_308, n_309, n_319, n_320, n_321, n_322, n_323, n_324;
  wire n_325, n_326, n_338, n_339, n_340, n_341, n_342, n_343;
  wire n_344, n_345, n_349, n_351, n_353, n_355, n_357, n_359;
  wire n_360, n_361, n_362, n_363, n_364, n_365, n_366, n_367;
  wire n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378;
  wire n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386;
  wire n_387, n_388, n_389, n_390, n_392, n_393, n_394, n_395;
  wire n_396, n_397, n_398, n_399, n_400, n_401, n_402, n_403;
  wire n_404, n_405, n_406, n_407, n_408, n_409, n_410, n_411;
  wire n_412, n_413, n_414, n_415, n_416, n_417, n_418, n_419;
  wire n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427;
  wire n_428, n_429, n_430, n_433, n_434, n_435, n_436, n_437;
  wire n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445;
  wire n_446, n_447, n_448, n_449, n_453, n_454, n_455, n_456;
  wire n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464;
  wire n_465, n_466, n_467, n_468, n_470, n_471, n_472, n_473;
  wire n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481;
  wire n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489;
  wire n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497;
  wire n_498, n_499, n_500, n_503, n_504, n_505, n_506, n_507;
  wire n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515;
  wire n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526;
  wire n_527, n_528, n_529, n_530, n_532, n_533, n_534, n_535;
  wire n_536, n_537, n_538, n_539, n_540, n_541, n_542, n_543;
  wire n_544, n_545, n_546, n_547, n_548, n_549, n_550, n_551;
  wire n_552, n_553, n_554, n_557, n_558, n_559, n_560, n_561;
  wire n_562, n_563, n_564, n_565, n_569, n_570, n_571, n_572;
  wire n_573, n_574, n_575, n_576, n_578, n_579, n_580, n_581;
  wire n_582, n_583, n_584, n_585, n_586, n_587, n_588, n_589;
  wire n_590, n_591, n_592, n_595, n_596, n_597, n_598, n_599;
  wire n_603, n_604, n_605, n_606, n_608, n_609, n_610, n_611;
  wire n_612, n_613, n_614, n_617, n_622, n_623, n_624, n_625;
  wire n_626, n_627, n_628, n_629, n_630, n_631, n_632, n_633;
  wire n_634, n_635, n_636, n_637, n_638, n_639, n_640, n_641;
  wire n_646, n_647, n_648, n_649, n_650, n_651, n_652, n_653;
  wire n_658, n_659, n_660, n_661, n_662, n_663, n_664, n_665;
  wire n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675;
  wire n_676, n_677, n_684, n_685, n_686, n_687, n_688, n_689;
  wire n_690, n_691, n_692, n_693, n_704, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_711, n_712, n_713, n_722, n_724;
  wire n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732;
  wire n_733, n_742, n_744, n_745, n_746, n_747, n_748, n_749;
  wire n_750, n_751, n_752, n_753, n_766, n_767, n_768, n_770;
  wire n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_794;
  wire n_795, n_796, n_798, n_799, n_800, n_801, n_802, n_803;
  wire n_804, n_805, n_822, n_823, n_824, n_826, n_827, n_828;
  wire n_829, n_830, n_831, n_832, n_833, n_842, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_866, n_867, n_868;
  wire n_872, n_873, n_876, n_877, n_880, n_881, n_882, n_883;
  wire n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891;
  wire n_892, n_893, n_906, n_907, n_908, n_910, n_911, n_912;
  wire n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920;
  wire n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928;
  wire n_929, n_946, n_947, n_949, n_950, n_951, n_952, n_953;
  wire n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961;
  wire n_962, n_963, n_964, n_965, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_996, n_997, n_998, n_999, n_1000, n_1001, n_1024, n_1025;
  wire n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033;
  wire n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041;
  wire n_1042, n_1044, n_1045, n_1046, n_1047, n_1048, n_1050, n_1051;
  wire n_1052, n_1056, n_1057, n_1060, n_1061, n_1064, n_1065, n_1068;
  wire n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
  wire n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084;
  wire n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092;
  wire n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100;
  wire n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108;
  wire n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116;
  wire n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124;
  wire n_1125, n_1126, n_1127, n_1128, n_1129, n_1132, n_1133, n_1134;
  wire n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142;
  wire n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150;
  wire n_1151, n_1152, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159;
  wire n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167;
  wire n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175;
  wire n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183;
  wire n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191;
  wire n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199;
  wire n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207;
  wire n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215;
  wire n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223;
  wire n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231;
  wire n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239;
  wire n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248;
  wire n_1249, n_1250, n_1252, n_1253, n_1254, n_1255, n_1256, n_1258;
  wire n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1266, n_1267;
  wire n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275;
  wire n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283;
  wire n_1284, n_1285, n_1286, n_1288, n_1290, n_1291, n_1292, n_1293;
  wire n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301;
  wire n_1302, n_1303, n_1304, n_1305, n_1306, n_1308, n_1309, n_1310;
  wire n_1311, n_1312, n_1313, n_1316, n_1317, n_1318, n_1319, n_1320;
  wire n_1321, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330;
  wire n_1331, n_1332, n_1333, n_1334, n_1336, n_1337, n_1338, n_1339;
  wire n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347;
  wire n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355;
  wire n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363;
  wire n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371;
  wire n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379;
  wire n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387;
  wire n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395;
  wire n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403;
  wire n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1412;
  wire n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421;
  wire n_1422, n_1423, n_1424, n_1426, n_1427, n_1428, n_1429, n_1432;
  wire n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440;
  wire n_1441, n_1442, n_1443, n_1444, n_1446, n_1447, n_1448, n_1449;
  wire n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457;
  wire n_1458, n_1459, n_1460, n_1461, n_1463, n_1464, n_1465, n_1466;
  wire n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475;
  wire n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483;
  wire n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491;
  wire n_1492, n_1493, n_1494, n_1495, n_1496, n_1498, n_1499, n_1500;
  wire n_1501, n_1502, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511;
  wire n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519;
  wire n_1520, n_1521, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529;
  wire n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537;
  wire n_1539, n_1540, n_1541, n_1542, n_1544, n_1545, n_1546, n_1547;
  wire n_1548, n_1549, n_1550, n_1552, n_1553, n_1554, n_1555, n_1556;
  wire n_1557, n_1558, n_1559, n_1560, n_1561, n_1566, n_1567, n_1568;
  wire n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576;
  wire n_1577, n_1578, n_1579, n_1580, n_1581, n_1583, n_1584, n_1585;
  wire n_1587, n_1588, n_1589, n_1593, n_1606, n_1611, n_1612, n_1613;
  wire n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621;
  wire n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629;
  wire n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637;
  wire n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645;
  wire n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653;
  wire n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661;
  wire n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669;
  wire n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677;
  wire n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685;
  wire n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693;
  wire n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701;
  wire n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709;
  wire n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717;
  wire n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725;
  wire n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733;
  wire n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741;
  wire n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749;
  wire n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757;
  wire n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765;
  wire n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773;
  wire n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781;
  wire n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789;
  wire n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797;
  wire n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805;
  wire n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813;
  wire n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821;
  wire n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829;
  wire n_1830, n_1831;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], A[2]);
  xor g270 (n_117, n_622, n_171);
  nand g3 (n_623, A[1], A[2]);
  nand g271 (n_624, n_171, A[2]);
  nand g272 (n_625, A[1], n_171);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, n_69);
  xor g288 (n_176, n_634, A[4]);
  nand g289 (n_635, n_68, n_69);
  nand g290 (n_636, A[4], n_69);
  nand g291 (n_637, n_68, A[4]);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_176);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_176);
  nand g296 (n_640, A[7], n_176);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g305 (n_646, n_117, A[5]);
  xor g306 (n_180, n_646, A[6]);
  nand g307 (n_647, n_117, A[5]);
  nand g308 (n_648, A[6], A[5]);
  nand g309 (n_649, n_117, A[6]);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, n_179, n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, n_179, n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, n_179, A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_188, n_659, n_660, n_661);
  xor g329 (n_662, n_183, A[9]);
  xor g330 (n_112, n_662, n_184);
  nand g331 (n_663, n_183, A[9]);
  nand g332 (n_664, n_184, A[9]);
  nand g333 (n_665, n_183, n_184);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_187, n_630, n_67);
  nand g340 (n_668, n_67, n_173);
  nand g341 (n_669, A[4], n_67);
  nand g342 (n_71, n_631, n_668, n_669);
  xor g343 (n_670, A[7], A[8]);
  xor g344 (n_189, n_670, n_187);
  nand g345 (n_671, A[7], A[8]);
  nand g346 (n_672, n_187, A[8]);
  nand g347 (n_673, A[7], n_187);
  nand g348 (n_73, n_671, n_672, n_673);
  xor g349 (n_674, n_188, A[10]);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, n_188, A[10]);
  nand g352 (n_676, n_189, A[10]);
  nand g353 (n_677, n_188, n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_72, n_638, A[8]);
  nand g366 (n_684, A[8], n_176);
  nand g367 (n_685, A[5], A[8]);
  nand g368 (n_201, n_639, n_684, n_685);
  xor g369 (n_686, n_71, A[9]);
  xor g370 (n_196, n_686, n_72);
  nand g371 (n_687, n_71, A[9]);
  nand g372 (n_688, n_72, A[9]);
  nand g373 (n_689, n_71, n_72);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, n_73, A[11]);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, n_73, A[11]);
  nand g378 (n_692, n_196, A[11]);
  nand g379 (n_693, n_73, n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g394 (n_202, n_650, A[9]);
  nand g396 (n_704, A[9], n_180);
  nand g397 (n_705, n_179, A[9]);
  nand g398 (n_209, n_651, n_704, n_705);
  xor g399 (n_706, A[10], n_201);
  xor g400 (n_204, n_706, n_202);
  nand g401 (n_707, A[10], n_201);
  nand g402 (n_708, n_202, n_201);
  nand g403 (n_709, A[10], n_202);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, A[12], n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, A[12], n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, A[12], n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g423 (n_722, n_183, n_184);
  xor g424 (n_210, n_722, A[10]);
  nand g426 (n_724, A[10], n_184);
  nand g427 (n_725, n_183, A[10]);
  nand g428 (n_218, n_665, n_724, n_725);
  xor g429 (n_726, A[11], n_209);
  xor g430 (n_212, n_726, n_210);
  nand g431 (n_727, A[11], n_209);
  nand g432 (n_728, n_210, n_209);
  nand g433 (n_729, A[11], n_210);
  nand g434 (n_220, n_727, n_728, n_729);
  xor g435 (n_730, n_211, A[13]);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, n_211, A[13]);
  nand g438 (n_732, n_212, A[13]);
  nand g439 (n_733, n_211, n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g455 (n_742, n_188, n_189);
  xor g456 (n_219, n_742, A[11]);
  nand g458 (n_744, A[11], n_189);
  nand g459 (n_745, n_188, A[11]);
  nand g460 (n_224, n_677, n_744, n_745);
  xor g461 (n_746, A[12], n_218);
  xor g462 (n_221, n_746, A[14]);
  nand g463 (n_747, A[12], n_218);
  nand g464 (n_748, A[14], n_218);
  nand g465 (n_749, A[12], A[14]);
  nand g466 (n_226, n_747, n_748, n_749);
  xor g467 (n_750, n_219, n_220);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, n_219, n_220);
  nand g470 (n_752, n_221, n_220);
  nand g471 (n_753, n_219, n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g493 (n_766, n_73, A[12]);
  xor g494 (n_225, n_766, n_196);
  nand g495 (n_767, n_73, A[12]);
  nand g496 (n_768, n_196, A[12]);
  nand g498 (n_236, n_767, n_768, n_693);
  xor g499 (n_770, n_224, A[13]);
  xor g500 (n_227, n_770, n_225);
  nand g501 (n_771, n_224, A[13]);
  nand g502 (n_772, n_225, A[13]);
  nand g503 (n_773, n_224, n_225);
  nand g504 (n_238, n_771, n_772, n_773);
  xor g505 (n_774, A[15], n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, A[15], n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, A[15], n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g535 (n_794, n_203, A[13]);
  xor g536 (n_237, n_794, n_204);
  nand g537 (n_795, n_203, A[13]);
  nand g538 (n_796, n_204, A[13]);
  nand g540 (n_248, n_795, n_796, n_712);
  xor g541 (n_798, A[14], n_236);
  xor g542 (n_239, n_798, A[16]);
  nand g543 (n_799, A[14], n_236);
  nand g544 (n_800, A[16], n_236);
  nand g545 (n_801, A[14], A[16]);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, n_237, n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, n_237, n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, n_237, n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g577 (n_822, n_211, A[14]);
  xor g578 (n_249, n_822, n_212);
  nand g579 (n_823, n_211, A[14]);
  nand g580 (n_824, n_212, A[14]);
  nand g582 (n_261, n_823, n_824, n_733);
  xor g583 (n_826, A[15], n_248);
  xor g584 (n_251, n_826, A[17]);
  nand g585 (n_827, A[15], n_248);
  nand g586 (n_828, A[17], n_248);
  nand g587 (n_829, A[15], A[17]);
  nand g588 (n_118, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g609 (n_842, n_188, A[11]);
  xor g610 (n_258, n_842, n_189);
  xor g616 (n_260, n_746, n_258);
  nand g618 (n_848, n_258, n_218);
  nand g619 (n_849, A[12], n_258);
  nand g620 (n_272, n_747, n_848, n_849);
  xor g621 (n_850, n_220, A[15]);
  xor g622 (n_262, n_850, n_260);
  nand g623 (n_851, n_220, A[15]);
  nand g624 (n_852, n_260, A[15]);
  nand g625 (n_853, n_220, n_260);
  nand g626 (n_274, n_851, n_852, n_853);
  xor g627 (n_854, A[16], n_261);
  xor g628 (n_119, n_854, A[18]);
  nand g629 (n_855, A[16], n_261);
  nand g630 (n_856, A[18], n_261);
  nand g631 (n_857, A[16], A[18]);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_262, n_118);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_262, n_118);
  nand g636 (n_860, n_119, n_118);
  nand g637 (n_861, n_262, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g641 (n_862, n_68, A[4]);
  xor g642 (n_265, n_862, n_69);
  xor g647 (n_866, A[5], n_265);
  xor g648 (n_267, n_866, A[8]);
  nand g649 (n_867, A[5], n_265);
  nand g650 (n_868, A[8], n_265);
  nand g652 (n_282, n_867, n_868, n_685);
  xor g654 (n_269, n_686, n_267);
  nand g656 (n_872, n_267, n_71);
  nand g657 (n_873, A[9], n_267);
  nand g658 (n_284, n_687, n_872, n_873);
  xor g660 (n_271, n_766, n_269);
  nand g662 (n_876, n_269, A[12]);
  nand g663 (n_877, n_73, n_269);
  nand g664 (n_286, n_767, n_876, n_877);
  xor g666 (n_273, n_770, n_271);
  nand g668 (n_880, n_271, A[13]);
  nand g669 (n_881, n_224, n_271);
  nand g670 (n_288, n_771, n_880, n_881);
  xor g671 (n_882, n_272, A[16]);
  xor g672 (n_275, n_882, n_273);
  nand g673 (n_883, n_272, A[16]);
  nand g674 (n_884, n_273, A[16]);
  nand g675 (n_885, n_272, n_273);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, A[17], n_274);
  xor g678 (n_277, n_886, A[19]);
  nand g679 (n_887, A[17], n_274);
  nand g680 (n_888, A[19], n_274);
  nand g681 (n_889, A[17], A[19]);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g707 (n_906, A[10], n_282);
  xor g708 (n_285, n_906, n_202);
  nand g709 (n_907, A[10], n_282);
  nand g710 (n_908, n_202, n_282);
  nand g712 (n_300, n_907, n_908, n_709);
  xor g713 (n_910, n_284, A[13]);
  xor g714 (n_287, n_910, n_285);
  nand g715 (n_911, n_284, A[13]);
  nand g716 (n_912, n_285, A[13]);
  nand g717 (n_913, n_284, n_285);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, A[14], n_286);
  xor g720 (n_289, n_914, n_287);
  nand g721 (n_915, A[14], n_286);
  nand g722 (n_916, n_287, n_286);
  nand g723 (n_917, A[14], n_287);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, n_288, A[17]);
  xor g726 (n_291, n_918, n_289);
  nand g727 (n_919, n_288, A[17]);
  nand g728 (n_920, n_289, A[17]);
  nand g729 (n_921, n_288, n_289);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, A[18], n_290);
  xor g732 (n_293, n_922, A[20]);
  nand g733 (n_923, A[18], n_290);
  nand g734 (n_924, A[20], n_290);
  nand g735 (n_925, A[18], A[20]);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g767 (n_946, n_300, A[14]);
  xor g768 (n_303, n_946, n_212);
  nand g769 (n_947, n_300, A[14]);
  nand g771 (n_949, n_300, n_212);
  nand g772 (n_319, n_947, n_824, n_949);
  xor g773 (n_950, n_302, A[15]);
  xor g774 (n_305, n_950, n_303);
  nand g775 (n_951, n_302, A[15]);
  nand g776 (n_952, n_303, A[15]);
  nand g777 (n_953, n_302, n_303);
  nand g778 (n_321, n_951, n_952, n_953);
  xor g779 (n_954, n_304, A[18]);
  xor g780 (n_307, n_954, n_305);
  nand g781 (n_955, n_304, A[18]);
  nand g782 (n_956, n_305, A[18]);
  nand g783 (n_957, n_304, n_305);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, A[19], n_306);
  xor g786 (n_309, n_958, A[21]);
  nand g787 (n_959, A[19], n_306);
  nand g788 (n_960, A[21], n_306);
  nand g789 (n_961, A[19], A[21]);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g824 (n_320, n_850, A[16]);
  nand g826 (n_984, A[16], A[15]);
  nand g827 (n_985, n_220, A[16]);
  nand g828 (n_338, n_851, n_984, n_985);
  xor g829 (n_986, n_260, n_319);
  xor g830 (n_322, n_986, n_320);
  nand g831 (n_987, n_260, n_319);
  nand g832 (n_988, n_320, n_319);
  nand g833 (n_989, n_260, n_320);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, n_321, A[19]);
  xor g836 (n_324, n_990, A[20]);
  nand g837 (n_991, n_321, A[19]);
  nand g838 (n_992, A[20], A[19]);
  nand g839 (n_993, n_321, A[20]);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, n_322, n_323);
  xor g842 (n_326, n_994, n_324);
  nand g843 (n_995, n_322, n_323);
  nand g844 (n_996, n_324, n_323);
  nand g845 (n_997, n_322, n_324);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, A[22], n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, A[22], n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, A[22], n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g886 (n_339, n_882, A[17]);
  nand g888 (n_1024, A[17], A[16]);
  nand g889 (n_1025, n_272, A[17]);
  nand g890 (n_360, n_883, n_1024, n_1025);
  xor g891 (n_1026, n_273, n_338);
  xor g892 (n_341, n_1026, n_339);
  nand g893 (n_1027, n_273, n_338);
  nand g894 (n_1028, n_339, n_338);
  nand g895 (n_1029, n_273, n_339);
  nand g896 (n_362, n_1027, n_1028, n_1029);
  xor g897 (n_1030, A[20], n_340);
  xor g898 (n_343, n_1030, n_341);
  nand g899 (n_1031, A[20], n_340);
  nand g900 (n_1032, n_341, n_340);
  nand g901 (n_1033, A[20], n_341);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, A[21], n_342);
  xor g904 (n_345, n_1034, n_343);
  nand g905 (n_1035, A[21], n_342);
  nand g906 (n_1036, n_343, n_342);
  nand g907 (n_1037, A[21], n_343);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, A[23], n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, A[23], n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, A[23], n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  xor g917 (n_1042, A[2], n_171);
  nand g922 (n_371, n_624, n_1044, n_1045);
  xor g923 (n_1046, A[5], n_349);
  xor g924 (n_351, n_1046, A[6]);
  nand g925 (n_1047, A[5], n_349);
  nand g926 (n_1048, A[6], n_349);
  nand g928 (n_373, n_1047, n_1048, n_648);
  xor g929 (n_1050, n_179, n_351);
  xor g930 (n_353, n_1050, A[9]);
  nand g931 (n_1051, n_179, n_351);
  nand g932 (n_1052, A[9], n_351);
  nand g934 (n_375, n_1051, n_1052, n_705);
  xor g936 (n_355, n_906, n_353);
  nand g938 (n_1056, n_353, A[10]);
  nand g939 (n_1057, n_282, n_353);
  nand g940 (n_377, n_907, n_1056, n_1057);
  xor g942 (n_357, n_910, n_355);
  nand g944 (n_1060, n_355, A[13]);
  nand g945 (n_1061, n_284, n_355);
  nand g946 (n_379, n_911, n_1060, n_1061);
  xor g948 (n_359, n_914, n_357);
  nand g950 (n_1064, n_357, n_286);
  nand g951 (n_1065, A[14], n_357);
  nand g952 (n_381, n_915, n_1064, n_1065);
  xor g954 (n_361, n_918, A[18]);
  nand g956 (n_1068, A[18], A[17]);
  nand g957 (n_1069, n_288, A[18]);
  nand g958 (n_383, n_919, n_1068, n_1069);
  xor g959 (n_1070, n_359, n_360);
  xor g960 (n_363, n_1070, n_361);
  nand g961 (n_1071, n_359, n_360);
  nand g962 (n_1072, n_361, n_360);
  nand g963 (n_1073, n_359, n_361);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, A[21], n_362);
  xor g966 (n_365, n_1074, A[22]);
  nand g967 (n_1075, A[21], n_362);
  nand g968 (n_1076, A[22], n_362);
  nand g969 (n_1077, A[21], A[22]);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g972 (n_367, n_1078, n_364);
  nand g975 (n_1081, n_363, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  xor g985 (n_1086, A[1], A[3]);
  nand g987 (n_1087, A[1], A[3]);
  nand g990 (n_392, n_1087, n_1088, n_1089);
  xor g991 (n_1090, n_371, A[6]);
  xor g992 (n_374, n_1090, n_372);
  nand g993 (n_1091, n_371, A[6]);
  nand g994 (n_1092, n_372, A[6]);
  nand g995 (n_1093, n_371, n_372);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, n_374);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, n_374, n_373);
  nand g1001 (n_1097, A[7], n_374);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, A[10], A[11]);
  xor g1004 (n_378, n_1098, n_375);
  nand g1005 (n_1099, A[10], A[11]);
  nand g1006 (n_1100, n_375, A[11]);
  nand g1007 (n_1101, A[10], n_375);
  nand g1008 (n_398, n_1099, n_1100, n_1101);
  xor g1009 (n_1102, n_376, n_377);
  xor g1010 (n_380, n_1102, n_378);
  nand g1011 (n_1103, n_376, n_377);
  nand g1012 (n_1104, n_378, n_377);
  nand g1013 (n_1105, n_376, n_378);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, A[14], n_379);
  xor g1016 (n_382, n_1106, A[15]);
  nand g1017 (n_1107, A[14], n_379);
  nand g1018 (n_1108, A[15], n_379);
  nand g1019 (n_1109, A[14], A[15]);
  nand g1020 (n_402, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, n_380, A[18]);
  xor g1022 (n_384, n_1110, n_381);
  nand g1023 (n_1111, n_380, A[18]);
  nand g1024 (n_1112, n_381, A[18]);
  nand g1025 (n_1113, n_380, n_381);
  nand g1026 (n_404, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, n_382, A[19]);
  xor g1028 (n_386, n_1114, n_383);
  nand g1029 (n_1115, n_382, A[19]);
  nand g1030 (n_1116, n_383, A[19]);
  nand g1031 (n_1117, n_382, n_383);
  nand g1032 (n_407, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_384, A[22]);
  xor g1034 (n_388, n_1118, n_385);
  nand g1035 (n_1119, n_384, A[22]);
  nand g1036 (n_1120, n_385, A[22]);
  nand g1037 (n_1121, n_384, n_385);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, n_386, A[23]);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, n_386, A[23]);
  nand g1042 (n_1124, n_387, A[23]);
  nand g1043 (n_1125, n_386, n_387);
  nand g1044 (n_410, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1052 (n_393, n_626, A[4]);
  nand g1054 (n_1132, A[4], A[2]);
  nand g1055 (n_1133, A[3], A[4]);
  nand g1056 (n_412, n_627, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, n_396, A[11]);
  xor g1070 (n_399, n_1142, A[12]);
  nand g1071 (n_1143, n_396, A[11]);
  nand g1072 (n_1144, A[12], A[11]);
  nand g1073 (n_1145, n_396, A[12]);
  nand g1074 (n_417, n_1143, n_1144, n_1145);
  xor g1075 (n_1146, n_397, n_398);
  xor g1076 (n_401, n_1146, n_399);
  nand g1077 (n_1147, n_397, n_398);
  nand g1078 (n_1148, n_399, n_398);
  nand g1079 (n_1149, n_397, n_399);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, A[15], n_400);
  xor g1082 (n_403, n_1150, A[16]);
  nand g1083 (n_1151, A[15], n_400);
  nand g1084 (n_1152, A[16], n_400);
  nand g1086 (n_421, n_1151, n_1152, n_984);
  xor g1087 (n_1154, n_401, n_402);
  xor g1088 (n_405, n_1154, A[19]);
  nand g1089 (n_1155, n_401, n_402);
  nand g1090 (n_1156, A[19], n_402);
  nand g1091 (n_1157, n_401, A[19]);
  nand g1092 (n_424, n_1155, n_1156, n_1157);
  xor g1093 (n_1158, n_403, A[20]);
  xor g1094 (n_406, n_1158, n_404);
  nand g1095 (n_1159, n_403, A[20]);
  nand g1096 (n_1160, n_404, A[20]);
  nand g1097 (n_1161, n_403, n_404);
  nand g1098 (n_425, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_405, n_406);
  xor g1100 (n_409, n_1162, n_407);
  nand g1101 (n_1163, n_405, n_406);
  nand g1102 (n_1164, n_407, n_406);
  nand g1103 (n_1165, n_405, n_407);
  nand g1104 (n_427, n_1163, n_1164, n_1165);
  xor g1106 (n_411, n_1166, n_408);
  nand g1108 (n_1168, n_408, A[23]);
  nand g1110 (n_430, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1123 (n_1178, A[8], A[9]);
  xor g1124 (n_415, n_1178, n_413);
  nand g1125 (n_1179, A[8], A[9]);
  nand g1126 (n_1180, n_413, A[9]);
  nand g1127 (n_1181, A[8], n_413);
  nand g1128 (n_435, n_1179, n_1180, n_1181);
  xor g1129 (n_1182, n_414, A[12]);
  xor g1130 (n_418, n_1182, n_415);
  nand g1131 (n_1183, n_414, A[12]);
  nand g1132 (n_1184, n_415, A[12]);
  nand g1133 (n_1185, n_414, n_415);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, n_416, A[13]);
  xor g1136 (n_420, n_1186, n_417);
  nand g1137 (n_1187, n_416, A[13]);
  nand g1138 (n_1188, n_417, A[13]);
  nand g1139 (n_1189, n_416, n_417);
  nand g1140 (n_439, n_1187, n_1188, n_1189);
  xor g1141 (n_1190, n_418, n_419);
  xor g1142 (n_422, n_1190, A[16]);
  nand g1143 (n_1191, n_418, n_419);
  nand g1144 (n_1192, A[16], n_419);
  nand g1145 (n_1193, n_418, A[16]);
  nand g1146 (n_440, n_1191, n_1192, n_1193);
  xor g1147 (n_1194, n_420, A[17]);
  xor g1148 (n_423, n_1194, n_421);
  nand g1149 (n_1195, n_420, A[17]);
  nand g1150 (n_1196, n_421, A[17]);
  nand g1151 (n_1197, n_420, n_421);
  nand g1152 (n_442, n_1195, n_1196, n_1197);
  xor g1153 (n_1198, n_422, A[20]);
  xor g1154 (n_426, n_1198, n_423);
  nand g1155 (n_1199, n_422, A[20]);
  nand g1156 (n_1200, n_423, A[20]);
  nand g1157 (n_1201, n_422, n_423);
  nand g1158 (n_445, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_424, A[21]);
  xor g1160 (n_428, n_1202, n_425);
  nand g1161 (n_1203, n_424, A[21]);
  nand g1162 (n_1204, n_425, A[21]);
  nand g1163 (n_1205, n_424, n_425);
  nand g1164 (n_447, n_1203, n_1204, n_1205);
  xor g1166 (n_429, n_1206, n_427);
  nand g1169 (n_1209, n_426, n_427);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, A[9]);
  nand g1183 (n_1217, A[6], A[9]);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, n_433, A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, n_433, A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, n_433, n_434);
  nand g1190 (n_456, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, n_435, n_436);
  xor g1192 (n_438, n_1222, A[13]);
  nand g1193 (n_1223, n_435, n_436);
  nand g1194 (n_1224, A[13], n_436);
  nand g1195 (n_1225, n_435, A[13]);
  nand g1196 (n_457, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, A[14], n_437);
  xor g1198 (n_441, n_1226, n_438);
  nand g1199 (n_1227, A[14], n_437);
  nand g1200 (n_1228, n_438, n_437);
  nand g1201 (n_1229, A[14], n_438);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, n_439, A[17]);
  xor g1204 (n_443, n_1230, n_440);
  nand g1205 (n_1231, n_439, A[17]);
  nand g1206 (n_1232, n_440, A[17]);
  nand g1207 (n_1233, n_439, n_440);
  nand g1208 (n_461, n_1231, n_1232, n_1233);
  xor g1209 (n_1234, A[18], n_441);
  xor g1210 (n_444, n_1234, n_442);
  nand g1211 (n_1235, A[18], n_441);
  nand g1212 (n_1236, n_442, n_441);
  nand g1213 (n_1237, A[18], n_442);
  nand g1214 (n_463, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_443, A[21]);
  xor g1216 (n_446, n_1238, A[22]);
  nand g1217 (n_1239, n_443, A[21]);
  nand g1219 (n_1241, n_443, A[22]);
  nand g1220 (n_465, n_1239, n_1077, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[5], A[7]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], n_453);
  xor g1242 (n_455, n_1254, A[11]);
  nand g1243 (n_1255, A[10], n_453);
  nand g1244 (n_1256, A[11], n_453);
  nand g1246 (n_473, n_1255, n_1256, n_1099);
  xor g1247 (n_1258, n_454, n_455);
  xor g1248 (n_458, n_1258, n_456);
  nand g1249 (n_1259, n_454, n_455);
  nand g1250 (n_1260, n_456, n_455);
  nand g1251 (n_1261, n_454, n_456);
  nand g1252 (n_474, n_1259, n_1260, n_1261);
  xor g1253 (n_1262, A[14], n_457);
  xor g1254 (n_460, n_1262, A[15]);
  nand g1255 (n_1263, A[14], n_457);
  nand g1256 (n_1264, A[15], n_457);
  nand g1258 (n_476, n_1263, n_1264, n_1109);
  xor g1259 (n_1266, n_458, A[18]);
  xor g1260 (n_462, n_1266, n_459);
  nand g1261 (n_1267, n_458, A[18]);
  nand g1262 (n_1268, n_459, A[18]);
  nand g1263 (n_1269, n_458, n_459);
  nand g1264 (n_478, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, n_460, A[19]);
  xor g1266 (n_464, n_1270, n_461);
  nand g1267 (n_1271, n_460, A[19]);
  nand g1268 (n_1272, n_461, A[19]);
  nand g1269 (n_1273, n_460, n_461);
  nand g1270 (n_480, n_1271, n_1272, n_1273);
  xor g1271 (n_1274, n_462, A[22]);
  xor g1272 (n_466, n_1274, n_463);
  nand g1273 (n_1275, n_462, A[22]);
  nand g1274 (n_1276, n_463, A[22]);
  nand g1275 (n_1277, n_462, n_463);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1277 (n_1278, n_464, A[23]);
  xor g1278 (n_467, n_1278, n_465);
  nand g1279 (n_1279, n_464, A[23]);
  nand g1280 (n_1280, n_465, A[23]);
  nand g1281 (n_1281, n_464, n_465);
  nand g1282 (n_484, n_1279, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1289 (n_1286, A[7], A[6]);
  xor g1290 (n_471, n_1286, A[8]);
  nand g1292 (n_1288, A[8], A[6]);
  nand g1294 (n_486, n_661, n_1288, n_671);
  xor g1295 (n_1290, n_470, n_471);
  xor g1296 (n_472, n_1290, A[11]);
  nand g1297 (n_1291, n_470, n_471);
  nand g1298 (n_1292, A[11], n_471);
  nand g1299 (n_1293, n_470, A[11]);
  nand g1300 (n_488, n_1291, n_1292, n_1293);
  xor g1301 (n_1294, A[12], n_472);
  xor g1302 (n_475, n_1294, n_473);
  nand g1303 (n_1295, A[12], n_472);
  nand g1304 (n_1296, n_473, n_472);
  nand g1305 (n_1297, A[12], n_473);
  nand g1306 (n_489, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, A[15], n_474);
  xor g1308 (n_477, n_1298, n_475);
  nand g1309 (n_1299, A[15], n_474);
  nand g1310 (n_1300, n_475, n_474);
  nand g1311 (n_1301, A[15], n_475);
  nand g1312 (n_491, n_1299, n_1300, n_1301);
  xor g1313 (n_1302, A[16], n_476);
  xor g1314 (n_479, n_1302, n_477);
  nand g1315 (n_1303, A[16], n_476);
  nand g1316 (n_1304, n_477, n_476);
  nand g1317 (n_1305, A[16], n_477);
  nand g1318 (n_494, n_1303, n_1304, n_1305);
  xor g1319 (n_1306, A[19], A[20]);
  xor g1320 (n_481, n_1306, n_478);
  nand g1322 (n_1308, n_478, A[20]);
  nand g1323 (n_1309, A[19], n_478);
  nand g1324 (n_496, n_992, n_1308, n_1309);
  xor g1325 (n_1310, n_479, n_480);
  xor g1326 (n_483, n_1310, n_481);
  nand g1327 (n_1311, n_479, n_480);
  nand g1328 (n_1312, n_481, n_480);
  nand g1329 (n_1313, n_479, n_481);
  nand g1330 (n_497, n_1311, n_1312, n_1313);
  xor g1332 (n_485, n_1166, n_482);
  nand g1335 (n_1317, A[23], n_482);
  nand g1336 (n_500, n_1167, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1344 (n_487, n_1178, n_486);
  nand g1346 (n_1324, n_486, A[9]);
  nand g1347 (n_1325, A[8], n_486);
  nand g1348 (n_503, n_1179, n_1324, n_1325);
  xor g1349 (n_1326, A[12], n_487);
  xor g1350 (n_490, n_1326, n_488);
  nand g1351 (n_1327, A[12], n_487);
  nand g1352 (n_1328, n_488, n_487);
  nand g1353 (n_1329, A[12], n_488);
  nand g1354 (n_505, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, A[13], n_489);
  xor g1356 (n_492, n_1330, n_490);
  nand g1357 (n_1331, A[13], n_489);
  nand g1358 (n_1332, n_490, n_489);
  nand g1359 (n_1333, A[13], n_490);
  nand g1360 (n_507, n_1331, n_1332, n_1333);
  xor g1361 (n_1334, A[16], A[17]);
  xor g1362 (n_493, n_1334, n_491);
  nand g1364 (n_1336, n_491, A[17]);
  nand g1365 (n_1337, A[16], n_491);
  nand g1366 (n_509, n_1024, n_1336, n_1337);
  xor g1367 (n_1338, n_492, A[20]);
  xor g1368 (n_495, n_1338, n_493);
  nand g1369 (n_1339, n_492, A[20]);
  nand g1370 (n_1340, n_493, A[20]);
  nand g1371 (n_1341, n_492, n_493);
  nand g1372 (n_511, n_1339, n_1340, n_1341);
  xor g1373 (n_1342, n_494, A[21]);
  xor g1374 (n_498, n_1342, n_495);
  nand g1375 (n_1343, n_494, A[21]);
  nand g1376 (n_1344, n_495, A[21]);
  nand g1377 (n_1345, n_494, n_495);
  nand g1378 (n_513, n_1343, n_1344, n_1345);
  xor g1380 (n_499, n_1346, n_497);
  nand g1383 (n_1349, n_496, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  xor g1394 (n_504, n_1354, n_503);
  nand g1397 (n_1357, A[10], n_503);
  nand g1398 (n_520, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], A[14]);
  xor g1400 (n_506, n_1358, n_504);
  nand g1401 (n_1359, A[13], A[14]);
  nand g1402 (n_1360, n_504, A[14]);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_521, n_1359, n_1360, n_1361);
  xor g1405 (n_1362, n_505, A[17]);
  xor g1406 (n_508, n_1362, n_506);
  nand g1407 (n_1363, n_505, A[17]);
  nand g1408 (n_1364, n_506, A[17]);
  nand g1409 (n_1365, n_505, n_506);
  nand g1410 (n_523, n_1363, n_1364, n_1365);
  xor g1411 (n_1366, n_507, A[18]);
  xor g1412 (n_510, n_1366, n_508);
  nand g1413 (n_1367, n_507, A[18]);
  nand g1414 (n_1368, n_508, A[18]);
  nand g1415 (n_1369, n_507, n_508);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_509, A[21]);
  xor g1418 (n_512, n_1370, n_510);
  nand g1419 (n_1371, n_509, A[21]);
  nand g1420 (n_1372, n_510, A[21]);
  nand g1421 (n_1373, n_509, n_510);
  nand g1422 (n_527, n_1371, n_1372, n_1373);
  xor g1423 (n_1374, A[22], n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, A[22], n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, A[22], n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1437 (n_1382, A[9], A[11]);
  nand g1439 (n_1383, A[9], A[11]);
  nand g1442 (n_532, n_1383, n_1384, n_1385);
  xor g1443 (n_1386, A[14], n_519);
  xor g1444 (n_522, n_1386, n_520);
  nand g1445 (n_1387, A[14], n_519);
  nand g1446 (n_1388, n_520, n_519);
  nand g1447 (n_1389, A[14], n_520);
  nand g1448 (n_534, n_1387, n_1388, n_1389);
  xor g1449 (n_1390, A[15], n_521);
  xor g1450 (n_524, n_1390, n_522);
  nand g1451 (n_1391, A[15], n_521);
  nand g1452 (n_1392, n_522, n_521);
  nand g1453 (n_1393, A[15], n_522);
  nand g1454 (n_536, n_1391, n_1392, n_1393);
  xor g1455 (n_1394, A[18], n_523);
  xor g1456 (n_525, n_1394, A[19]);
  nand g1457 (n_1395, A[18], n_523);
  nand g1458 (n_1396, A[19], n_523);
  nand g1459 (n_1397, A[18], A[19]);
  nand g1460 (n_538, n_1395, n_1396, n_1397);
  xor g1461 (n_1398, n_524, n_525);
  xor g1462 (n_528, n_1398, n_526);
  nand g1463 (n_1399, n_524, n_525);
  nand g1464 (n_1400, n_526, n_525);
  nand g1465 (n_1401, n_524, n_526);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1467 (n_1402, A[22], A[23]);
  xor g1468 (n_529, n_1402, n_527);
  nand g1469 (n_1403, A[22], A[23]);
  nand g1470 (n_1404, n_527, A[23]);
  nand g1471 (n_1405, A[22], n_527);
  nand g1472 (n_543, n_1403, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1479 (n_1410, A[11], A[12]);
  xor g1480 (n_533, n_1410, A[10]);
  nand g1482 (n_1412, A[10], A[12]);
  nand g1484 (n_544, n_1144, n_1412, n_1099);
  xor g1485 (n_1414, n_532, n_533);
  xor g1486 (n_535, n_1414, A[15]);
  nand g1487 (n_1415, n_532, n_533);
  nand g1488 (n_1416, A[15], n_533);
  nand g1489 (n_1417, n_532, A[15]);
  nand g1490 (n_546, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, A[16], n_534);
  xor g1492 (n_537, n_1418, n_535);
  nand g1493 (n_1419, A[16], n_534);
  nand g1494 (n_1420, n_535, n_534);
  nand g1495 (n_1421, A[16], n_535);
  nand g1496 (n_548, n_1419, n_1420, n_1421);
  xor g1497 (n_1422, A[19], n_536);
  xor g1498 (n_539, n_1422, A[20]);
  nand g1499 (n_1423, A[19], n_536);
  nand g1500 (n_1424, A[20], n_536);
  nand g1502 (n_549, n_1423, n_1424, n_992);
  xor g1503 (n_1426, n_537, n_538);
  xor g1504 (n_541, n_1426, n_539);
  nand g1505 (n_1427, n_537, n_538);
  nand g1506 (n_1428, n_539, n_538);
  nand g1507 (n_1429, n_537, n_539);
  nand g1508 (n_551, n_1427, n_1428, n_1429);
  xor g1510 (n_542, n_1166, n_540);
  nand g1513 (n_1433, A[23], n_540);
  nand g1514 (n_554, n_1167, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1521 (n_1438, A[12], A[13]);
  xor g1522 (n_545, n_1438, n_544);
  nand g1523 (n_1439, A[12], A[13]);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_1439, n_1440, n_1441);
  xor g1527 (n_1442, A[16], n_545);
  xor g1528 (n_547, n_1442, A[17]);
  nand g1529 (n_1443, A[16], n_545);
  nand g1530 (n_1444, A[17], n_545);
  nand g1532 (n_559, n_1443, n_1444, n_1024);
  xor g1533 (n_1446, n_546, n_547);
  xor g1534 (n_550, n_1446, A[20]);
  nand g1535 (n_1447, n_546, n_547);
  nand g1536 (n_1448, A[20], n_547);
  nand g1537 (n_1449, n_546, A[20]);
  nand g1538 (n_561, n_1447, n_1448, n_1449);
  xor g1539 (n_1450, n_548, A[21]);
  xor g1540 (n_552, n_1450, n_549);
  nand g1541 (n_1451, n_548, A[21]);
  nand g1542 (n_1452, n_549, A[21]);
  nand g1543 (n_1453, n_548, n_549);
  nand g1544 (n_562, n_1451, n_1452, n_1453);
  xor g1546 (n_553, n_1454, n_551);
  nand g1549 (n_1457, n_550, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1563 (n_1465, A[14], n_557);
  nand g1564 (n_569, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, A[17], A[18]);
  xor g1566 (n_560, n_1466, n_558);
  nand g1568 (n_1468, n_558, A[18]);
  nand g1569 (n_1469, A[17], n_558);
  nand g1570 (n_571, n_1068, n_1468, n_1469);
  xor g1571 (n_1470, n_559, n_560);
  xor g1572 (n_563, n_1470, A[21]);
  nand g1573 (n_1471, n_559, n_560);
  nand g1574 (n_1472, A[21], n_560);
  nand g1575 (n_1473, n_559, A[21]);
  nand g1576 (n_574, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, A[22], n_561);
  xor g1578 (n_564, n_1474, n_562);
  nand g1579 (n_1475, A[22], n_561);
  nand g1580 (n_1476, n_562, n_561);
  nand g1581 (n_1477, A[22], n_562);
  nand g1582 (n_576, n_1475, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  xor g1591 (n_1482, A[13], A[15]);
  nand g1593 (n_1483, A[13], A[15]);
  nand g1596 (n_578, n_1483, n_1484, n_1485);
  xor g1597 (n_1486, A[18], n_569);
  xor g1598 (n_572, n_1486, n_570);
  nand g1599 (n_1487, A[18], n_569);
  nand g1600 (n_1488, n_570, n_569);
  nand g1601 (n_1489, A[18], n_570);
  nand g1602 (n_580, n_1487, n_1488, n_1489);
  xor g1603 (n_1490, A[19], n_571);
  xor g1604 (n_573, n_1490, n_572);
  nand g1605 (n_1491, A[19], n_571);
  nand g1606 (n_1492, n_572, n_571);
  nand g1607 (n_1493, A[19], n_572);
  nand g1608 (n_583, n_1491, n_1492, n_1493);
  xor g1609 (n_1494, A[22], n_573);
  xor g1610 (n_575, n_1494, A[23]);
  nand g1611 (n_1495, A[22], n_573);
  nand g1612 (n_1496, A[23], n_573);
  nand g1614 (n_584, n_1495, n_1496, n_1403);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1621 (n_1502, A[15], A[14]);
  xor g1622 (n_579, n_1502, A[16]);
  nand g1626 (n_586, n_1109, n_801, n_984);
  xor g1627 (n_1506, n_578, n_579);
  xor g1628 (n_581, n_1506, A[19]);
  nand g1629 (n_1507, n_578, n_579);
  nand g1630 (n_1508, A[19], n_579);
  nand g1631 (n_1509, n_578, A[19]);
  nand g1632 (n_588, n_1507, n_1508, n_1509);
  xor g1633 (n_1510, A[20], n_580);
  xor g1634 (n_582, n_1510, n_581);
  nand g1635 (n_1511, A[20], n_580);
  nand g1636 (n_1512, n_581, n_580);
  nand g1637 (n_1513, A[20], n_581);
  nand g1638 (n_589, n_1511, n_1512, n_1513);
  xor g1639 (n_1514, A[23], n_582);
  xor g1640 (n_585, n_1514, n_583);
  nand g1641 (n_1515, A[23], n_582);
  nand g1642 (n_1516, n_583, n_582);
  nand g1643 (n_1517, A[23], n_583);
  nand g1644 (n_591, n_1515, n_1516, n_1517);
  xor g1646 (n_83, n_1518, n_585);
  nand g1648 (n_1520, n_585, n_584);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1652 (n_587, n_1334, n_586);
  nand g1654 (n_1524, n_586, A[17]);
  nand g1655 (n_1525, A[16], n_586);
  nand g1656 (n_595, n_1024, n_1524, n_1525);
  xor g1657 (n_1526, A[20], n_587);
  xor g1658 (n_590, n_1526, n_588);
  nand g1659 (n_1527, A[20], n_587);
  nand g1660 (n_1528, n_588, n_587);
  nand g1661 (n_1529, A[20], n_588);
  nand g1662 (n_597, n_1527, n_1528, n_1529);
  xor g1664 (n_592, n_1530, n_589);
  nand g1667 (n_1533, A[21], n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_81, n_1535, n_1536, n_1537);
  nand g1681 (n_1541, A[18], n_595);
  nand g1682 (n_604, n_1539, n_1540, n_1541);
  xor g1683 (n_1542, A[21], A[22]);
  xor g1684 (n_598, n_1542, n_596);
  nand g1686 (n_1544, n_596, A[22]);
  nand g1687 (n_1545, A[21], n_596);
  nand g1688 (n_606, n_1077, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_33, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[17], A[19]);
  nand g1702 (n_608, n_889, n_1552, n_1553);
  xor g1703 (n_1554, A[22], n_603);
  xor g1704 (n_605, n_1554, n_604);
  nand g1705 (n_1555, A[22], n_603);
  nand g1706 (n_1556, n_604, n_603);
  nand g1707 (n_1557, A[22], n_604);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, A[23], n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, A[23], n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, A[23], n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1716 (n_609, n_1306, A[18]);
  nand g1720 (n_612, n_992, n_925, n_1397);
  xor g1721 (n_1566, n_608, n_609);
  xor g1722 (n_611, n_1566, A[23]);
  nand g1723 (n_1567, n_608, n_609);
  nand g1724 (n_1568, A[23], n_609);
  nand g1725 (n_1569, n_608, A[23]);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1728 (n_79, n_1570, n_611);
  nand g1730 (n_1572, n_611, n_610);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1733 (n_1574, A[20], A[21]);
  xor g1734 (n_613, n_1574, n_612);
  nand g1735 (n_1575, A[20], A[21]);
  nand g1736 (n_1576, n_612, A[21]);
  nand g1737 (n_1577, A[20], n_612);
  nand g1738 (n_617, n_1575, n_1576, n_1577);
  xor g1740 (n_78, n_1578, n_614);
  nand g1742 (n_1580, n_614, n_613);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_617);
  nand g1752 (n_28, n_1583, n_1584, n_1585);
  nand g1759 (n_1589, A[21], A[23]);
  nand g1760 (n_27, n_1587, n_1588, n_1589);
  xor g1762 (n_75, n_1166, A[22]);
  nand g1766 (n_74, n_1167, n_1403, n_1593);
  nand g16 (n_1606, A[0], A[2]);
  xor g20 (Z[2], A[0], A[2]);
  nand g22 (n_1611, n_68, A[3]);
  nand g25 (n_1615, n_1611, n_1612, n_1613);
  xor g26 (n_1614, n_68, A[3]);
  nand g28 (n_1616, A[4], n_117);
  nand g29 (n_1617, A[4], n_1615);
  nand g30 (n_1618, n_117, n_1615);
  nand g31 (n_1620, n_1616, n_1617, n_1618);
  xor g32 (n_1619, A[4], n_117);
  xor g33 (Z[4], n_1615, n_1619);
  nand g34 (n_1621, A[5], n_116);
  nand g35 (n_1622, A[5], n_1620);
  nand g36 (n_1623, n_116, n_1620);
  nand g37 (n_1625, n_1621, n_1622, n_1623);
  xor g38 (n_1624, A[5], n_116);
  xor g39 (Z[5], n_1620, n_1624);
  nand g40 (n_1626, n_67, n_115);
  nand g41 (n_1627, n_67, n_1625);
  nand g42 (n_1628, n_115, n_1625);
  nand g43 (n_1630, n_1626, n_1627, n_1628);
  xor g44 (n_1629, n_67, n_115);
  xor g45 (Z[6], n_1625, n_1629);
  nand g46 (n_1631, n_66, n_114);
  nand g47 (n_1632, n_66, n_1630);
  nand g48 (n_1633, n_114, n_1630);
  nand g49 (n_1635, n_1631, n_1632, n_1633);
  xor g50 (n_1634, n_66, n_114);
  xor g51 (Z[7], n_1630, n_1634);
  nand g52 (n_1636, n_65, n_113);
  nand g53 (n_1637, n_65, n_1635);
  nand g54 (n_1638, n_113, n_1635);
  nand g55 (n_1640, n_1636, n_1637, n_1638);
  xor g56 (n_1639, n_65, n_113);
  xor g57 (Z[8], n_1635, n_1639);
  nand g58 (n_1641, n_64, n_112);
  nand g59 (n_1642, n_64, n_1640);
  nand g60 (n_1643, n_112, n_1640);
  nand g61 (n_1645, n_1641, n_1642, n_1643);
  xor g62 (n_1644, n_64, n_112);
  xor g63 (Z[9], n_1640, n_1644);
  nand g64 (n_1646, n_63, n_111);
  nand g65 (n_1647, n_63, n_1645);
  nand g66 (n_1648, n_111, n_1645);
  nand g67 (n_1650, n_1646, n_1647, n_1648);
  xor g68 (n_1649, n_63, n_111);
  xor g69 (Z[10], n_1645, n_1649);
  nand g70 (n_1651, n_62, n_110);
  nand g71 (n_1652, n_62, n_1650);
  nand g72 (n_1653, n_110, n_1650);
  nand g73 (n_1655, n_1651, n_1652, n_1653);
  xor g74 (n_1654, n_62, n_110);
  xor g75 (Z[11], n_1650, n_1654);
  nand g76 (n_1656, n_61, n_109);
  nand g77 (n_1657, n_61, n_1655);
  nand g78 (n_1658, n_109, n_1655);
  nand g79 (n_1660, n_1656, n_1657, n_1658);
  xor g80 (n_1659, n_61, n_109);
  xor g81 (Z[12], n_1655, n_1659);
  nand g82 (n_1661, n_60, n_108);
  nand g83 (n_1662, n_60, n_1660);
  nand g84 (n_1663, n_108, n_1660);
  nand g85 (n_1665, n_1661, n_1662, n_1663);
  xor g86 (n_1664, n_60, n_108);
  xor g87 (Z[13], n_1660, n_1664);
  nand g88 (n_1666, n_59, n_107);
  nand g89 (n_1667, n_59, n_1665);
  nand g90 (n_1668, n_107, n_1665);
  nand g91 (n_1670, n_1666, n_1667, n_1668);
  xor g92 (n_1669, n_59, n_107);
  xor g93 (Z[14], n_1665, n_1669);
  nand g94 (n_1671, n_58, n_106);
  nand g95 (n_1672, n_58, n_1670);
  nand g96 (n_1673, n_106, n_1670);
  nand g97 (n_1675, n_1671, n_1672, n_1673);
  xor g98 (n_1674, n_58, n_106);
  xor g99 (Z[15], n_1670, n_1674);
  nand g100 (n_1676, n_57, n_105);
  nand g101 (n_1677, n_57, n_1675);
  nand g102 (n_1678, n_105, n_1675);
  nand g103 (n_1680, n_1676, n_1677, n_1678);
  xor g104 (n_1679, n_57, n_105);
  xor g105 (Z[16], n_1675, n_1679);
  nand g106 (n_1681, n_56, n_104);
  nand g107 (n_1682, n_56, n_1680);
  nand g108 (n_1683, n_104, n_1680);
  nand g109 (n_1685, n_1681, n_1682, n_1683);
  xor g110 (n_1684, n_56, n_104);
  xor g111 (Z[17], n_1680, n_1684);
  nand g112 (n_1686, n_55, n_103);
  nand g113 (n_1687, n_55, n_1685);
  nand g114 (n_1688, n_103, n_1685);
  nand g115 (n_1690, n_1686, n_1687, n_1688);
  xor g116 (n_1689, n_55, n_103);
  xor g117 (Z[18], n_1685, n_1689);
  nand g118 (n_1691, n_54, n_102);
  nand g119 (n_1692, n_54, n_1690);
  nand g120 (n_1693, n_102, n_1690);
  nand g121 (n_1695, n_1691, n_1692, n_1693);
  xor g122 (n_1694, n_54, n_102);
  xor g123 (Z[19], n_1690, n_1694);
  nand g124 (n_1696, n_53, n_101);
  nand g125 (n_1697, n_53, n_1695);
  nand g126 (n_1698, n_101, n_1695);
  nand g127 (n_1700, n_1696, n_1697, n_1698);
  xor g128 (n_1699, n_53, n_101);
  xor g129 (Z[20], n_1695, n_1699);
  nand g130 (n_1701, n_52, n_100);
  nand g131 (n_1702, n_52, n_1700);
  nand g132 (n_1703, n_100, n_1700);
  nand g133 (n_1705, n_1701, n_1702, n_1703);
  xor g134 (n_1704, n_52, n_100);
  xor g135 (Z[21], n_1700, n_1704);
  nand g136 (n_1706, n_51, n_99);
  nand g137 (n_1707, n_51, n_1705);
  nand g138 (n_1708, n_99, n_1705);
  nand g139 (n_1710, n_1706, n_1707, n_1708);
  xor g140 (n_1709, n_51, n_99);
  xor g141 (Z[22], n_1705, n_1709);
  nand g142 (n_1711, n_50, n_98);
  nand g143 (n_1712, n_50, n_1710);
  nand g144 (n_1713, n_98, n_1710);
  nand g145 (n_1715, n_1711, n_1712, n_1713);
  xor g146 (n_1714, n_50, n_98);
  xor g147 (Z[23], n_1710, n_1714);
  nand g148 (n_1716, n_49, n_97);
  nand g149 (n_1717, n_49, n_1715);
  nand g150 (n_1718, n_97, n_1715);
  nand g151 (n_1720, n_1716, n_1717, n_1718);
  xor g152 (n_1719, n_49, n_97);
  xor g153 (Z[24], n_1715, n_1719);
  nand g154 (n_1721, n_48, n_96);
  nand g155 (n_1722, n_48, n_1720);
  nand g156 (n_1723, n_96, n_1720);
  nand g157 (n_1725, n_1721, n_1722, n_1723);
  xor g158 (n_1724, n_48, n_96);
  xor g159 (Z[25], n_1720, n_1724);
  nand g160 (n_1726, n_47, n_95);
  nand g161 (n_1727, n_47, n_1725);
  nand g162 (n_1728, n_95, n_1725);
  nand g163 (n_1730, n_1726, n_1727, n_1728);
  xor g164 (n_1729, n_47, n_95);
  xor g165 (Z[26], n_1725, n_1729);
  nand g166 (n_1731, n_46, n_94);
  nand g167 (n_1732, n_46, n_1730);
  nand g168 (n_1733, n_94, n_1730);
  nand g169 (n_1735, n_1731, n_1732, n_1733);
  xor g170 (n_1734, n_46, n_94);
  xor g171 (Z[27], n_1730, n_1734);
  nand g172 (n_1736, n_45, n_93);
  nand g173 (n_1737, n_45, n_1735);
  nand g174 (n_1738, n_93, n_1735);
  nand g175 (n_1740, n_1736, n_1737, n_1738);
  xor g176 (n_1739, n_45, n_93);
  xor g177 (Z[28], n_1735, n_1739);
  nand g178 (n_1741, n_44, n_92);
  nand g179 (n_1742, n_44, n_1740);
  nand g180 (n_1743, n_92, n_1740);
  nand g181 (n_1745, n_1741, n_1742, n_1743);
  xor g182 (n_1744, n_44, n_92);
  xor g183 (Z[29], n_1740, n_1744);
  nand g184 (n_1746, n_43, n_91);
  nand g185 (n_1747, n_43, n_1745);
  nand g186 (n_1748, n_91, n_1745);
  nand g187 (n_1750, n_1746, n_1747, n_1748);
  xor g188 (n_1749, n_43, n_91);
  xor g189 (Z[30], n_1745, n_1749);
  nand g190 (n_1751, n_42, n_90);
  nand g191 (n_1752, n_42, n_1750);
  nand g192 (n_1753, n_90, n_1750);
  nand g193 (n_1755, n_1751, n_1752, n_1753);
  xor g194 (n_1754, n_42, n_90);
  xor g195 (Z[31], n_1750, n_1754);
  nand g196 (n_1756, n_41, n_89);
  nand g197 (n_1757, n_41, n_1755);
  nand g198 (n_1758, n_89, n_1755);
  nand g199 (n_1760, n_1756, n_1757, n_1758);
  xor g200 (n_1759, n_41, n_89);
  xor g201 (Z[32], n_1755, n_1759);
  nand g202 (n_1761, n_40, n_88);
  nand g203 (n_1762, n_40, n_1760);
  nand g204 (n_1763, n_88, n_1760);
  nand g205 (n_1765, n_1761, n_1762, n_1763);
  xor g206 (n_1764, n_40, n_88);
  xor g207 (Z[33], n_1760, n_1764);
  nand g208 (n_1766, n_39, n_87);
  nand g209 (n_1767, n_39, n_1765);
  nand g210 (n_1768, n_87, n_1765);
  nand g211 (n_1770, n_1766, n_1767, n_1768);
  xor g212 (n_1769, n_39, n_87);
  xor g213 (Z[34], n_1765, n_1769);
  nand g214 (n_1771, n_38, n_86);
  nand g215 (n_1772, n_38, n_1770);
  nand g216 (n_1773, n_86, n_1770);
  nand g217 (n_1775, n_1771, n_1772, n_1773);
  xor g218 (n_1774, n_38, n_86);
  xor g219 (Z[35], n_1770, n_1774);
  nand g220 (n_1776, n_37, n_85);
  nand g221 (n_1777, n_37, n_1775);
  nand g222 (n_1778, n_85, n_1775);
  nand g223 (n_1780, n_1776, n_1777, n_1778);
  xor g224 (n_1779, n_37, n_85);
  xor g225 (Z[36], n_1775, n_1779);
  nand g226 (n_1781, n_36, n_84);
  nand g227 (n_1782, n_36, n_1780);
  nand g228 (n_1783, n_84, n_1780);
  nand g229 (n_1785, n_1781, n_1782, n_1783);
  xor g230 (n_1784, n_36, n_84);
  xor g231 (Z[37], n_1780, n_1784);
  nand g232 (n_1786, n_35, n_83);
  nand g233 (n_1787, n_35, n_1785);
  nand g234 (n_1788, n_83, n_1785);
  nand g235 (n_1790, n_1786, n_1787, n_1788);
  xor g236 (n_1789, n_35, n_83);
  xor g237 (Z[38], n_1785, n_1789);
  nand g238 (n_1791, n_34, n_82);
  nand g239 (n_1792, n_34, n_1790);
  nand g240 (n_1793, n_82, n_1790);
  nand g241 (n_1795, n_1791, n_1792, n_1793);
  xor g242 (n_1794, n_34, n_82);
  xor g243 (Z[39], n_1790, n_1794);
  nand g244 (n_1796, n_33, n_81);
  nand g245 (n_1797, n_33, n_1795);
  nand g246 (n_1798, n_81, n_1795);
  nand g247 (n_1800, n_1796, n_1797, n_1798);
  xor g248 (n_1799, n_33, n_81);
  xor g249 (Z[40], n_1795, n_1799);
  nand g250 (n_1801, n_32, n_80);
  nand g251 (n_1802, n_32, n_1800);
  nand g252 (n_1803, n_80, n_1800);
  nand g253 (n_1805, n_1801, n_1802, n_1803);
  xor g254 (n_1804, n_32, n_80);
  xor g255 (Z[41], n_1800, n_1804);
  nand g256 (n_1806, n_31, n_79);
  nand g257 (n_1807, n_31, n_1805);
  nand g258 (n_1808, n_79, n_1805);
  nand g259 (n_1810, n_1806, n_1807, n_1808);
  xor g260 (n_1809, n_31, n_79);
  xor g261 (Z[42], n_1805, n_1809);
  nand g262 (n_1811, n_30, n_78);
  nand g263 (n_1812, n_30, n_1810);
  nand g264 (n_1813, n_78, n_1810);
  nand g265 (n_1815, n_1811, n_1812, n_1813);
  xor g266 (n_1814, n_30, n_78);
  xor g267 (Z[43], n_1810, n_1814);
  nand g1772 (n_1816, n_29, n_77);
  nand g1773 (n_1817, n_29, n_1815);
  nand g1774 (n_1818, n_77, n_1815);
  nand g1775 (n_1820, n_1816, n_1817, n_1818);
  xor g1776 (n_1819, n_29, n_77);
  xor g1777 (Z[44], n_1815, n_1819);
  nand g1778 (n_1821, n_28, n_76);
  nand g1779 (n_1822, n_28, n_1820);
  nand g1780 (n_1823, n_76, n_1820);
  nand g1781 (n_1825, n_1821, n_1822, n_1823);
  xor g1782 (n_1824, n_28, n_76);
  xor g1783 (Z[45], n_1820, n_1824);
  nand g1784 (n_1826, n_27, n_75);
  nand g1785 (n_1827, n_27, n_1825);
  nand g1786 (n_1828, n_75, n_1825);
  nand g1787 (n_1830, n_1826, n_1827, n_1828);
  xor g1788 (n_1829, n_27, n_75);
  xor g1789 (Z[46], n_1825, n_1829);
  xor g1791 (Z[47], n_1830, n_1831);
  or g1804 (n_1044, A[1], wc);
  not gc (wc, n_171);
  or g1805 (n_1045, A[1], wc0);
  not gc0 (wc0, A[2]);
  or g1806 (n_1088, A[2], wc1);
  not gc1 (wc1, A[3]);
  or g1807 (n_1089, wc2, A[2]);
  not gc2 (wc2, A[1]);
  xnor g1808 (n_1166, A[24], A[23]);
  or g1809 (n_1167, wc3, A[24]);
  not gc3 (wc3, A[23]);
  xnor g1810 (n_1214, A[6], A[5]);
  or g1811 (n_1215, A[5], wc4);
  not gc4 (wc4, A[6]);
  or g1812 (n_1216, A[5], wc5);
  not gc5 (wc5, A[9]);
  or g1813 (n_1252, A[6], wc6);
  not gc6 (wc6, A[7]);
  or g1814 (n_1253, wc7, A[6]);
  not gc7 (wc7, A[5]);
  xnor g1815 (n_1354, A[10], A[9]);
  or g1816 (n_1355, A[9], wc8);
  not gc8 (wc8, A[10]);
  or g1817 (n_1384, A[10], wc9);
  not gc9 (wc9, A[11]);
  or g1818 (n_1385, wc10, A[10]);
  not gc10 (wc10, A[9]);
  or g1820 (n_1463, A[13], wc11);
  not gc11 (wc11, A[14]);
  or g1821 (n_1484, A[14], wc12);
  not gc12 (wc12, A[15]);
  or g1822 (n_1485, wc13, A[14]);
  not gc13 (wc13, A[13]);
  xnor g1823 (n_1530, A[24], A[21]);
  or g1824 (n_1531, wc14, A[24]);
  not gc14 (wc14, A[21]);
  or g1826 (n_1539, A[17], wc15);
  not gc15 (wc15, A[18]);
  or g1827 (n_1552, A[18], wc16);
  not gc16 (wc16, A[19]);
  or g1828 (n_1553, wc17, A[18]);
  not gc17 (wc17, A[17]);
  or g1830 (n_1583, A[21], wc18);
  not gc18 (wc18, A[22]);
  or g1831 (n_1587, wc19, A[22]);
  not gc19 (wc19, A[21]);
  or g1832 (n_1588, A[22], wc20);
  not gc20 (wc20, A[23]);
  or g1833 (n_1593, wc21, A[24]);
  not gc21 (wc21, A[22]);
  xnor g1834 (n_349, n_1042, A[1]);
  xnor g1835 (n_372, n_1086, A[2]);
  xnor g1836 (n_453, n_1250, A[6]);
  xnor g1837 (n_519, n_1382, A[10]);
  xnor g1838 (n_570, n_1482, A[14]);
  xnor g1839 (n_603, n_1550, A[18]);
  xnor g1840 (n_76, n_1542, A[23]);
  xnor g1841 (n_1578, n_613, A[24]);
  or g1842 (n_1579, A[24], wc22);
  not gc22 (wc22, n_613);
  xnor g1843 (n_1831, n_74, A[24]);
  or g1844 (n_1356, A[9], wc23);
  not gc23 (wc23, n_503);
  xnor g1845 (n_558, n_1358, n_557);
  or g1846 (n_1464, A[13], wc24);
  not gc24 (wc24, n_557);
  xnor g1847 (n_596, n_1466, n_595);
  or g1848 (n_1540, A[17], wc25);
  not gc25 (wc25, n_595);
  or g1849 (n_1573, A[24], wc26);
  not gc26 (wc26, n_611);
  or g1850 (n_1581, A[24], wc27);
  not gc27 (wc27, n_614);
  xnor g1851 (n_29, n_1542, n_617);
  or g1852 (n_1584, A[21], wc28);
  not gc28 (wc28, n_617);
  or g1854 (n_1612, n_1606, wc29);
  not gc29 (wc29, n_68);
  or g1855 (n_1613, wc30, n_1606);
  not gc30 (wc30, A[3]);
  xnor g1856 (Z[3], n_1606, n_1614);
  xnor g1857 (n_1454, n_550, A[24]);
  or g1858 (n_1455, A[24], wc31);
  not gc31 (wc31, n_550);
  xnor g1859 (n_1570, n_610, A[24]);
  or g1860 (n_1571, A[24], wc32);
  not gc32 (wc32, n_610);
  or g1861 (n_1532, A[24], wc33);
  not gc33 (wc33, n_589);
  xnor g1862 (n_1518, n_584, A[24]);
  or g1863 (n_1519, A[24], wc34);
  not gc34 (wc34, n_584);
  or g1864 (n_1432, A[24], wc35);
  not gc35 (wc35, n_540);
  or g1865 (n_1521, A[24], wc36);
  not gc36 (wc36, n_585);
  or g1866 (n_1456, A[24], wc37);
  not gc37 (wc37, n_551);
  xnor g1867 (n_1078, n_363, A[24]);
  or g1868 (n_1079, A[24], wc38);
  not gc38 (wc38, n_363);
  xnor g1869 (n_1206, n_426, A[24]);
  or g1870 (n_1207, A[24], wc39);
  not gc39 (wc39, n_426);
  xnor g1871 (n_1346, n_496, A[24]);
  or g1872 (n_1347, A[24], wc40);
  not gc40 (wc40, n_496);
  or g1873 (n_1080, A[24], wc41);
  not gc41 (wc41, n_364);
  or g1874 (n_1169, A[24], wc42);
  not gc42 (wc42, n_408);
  or g1875 (n_1208, A[24], wc43);
  not gc43 (wc43, n_427);
  or g1876 (n_1316, A[24], wc44);
  not gc44 (wc44, n_482);
  or g1877 (n_1348, A[24], wc45);
  not gc45 (wc45, n_497);
endmodule

module mult_signed_const_4419_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_4419_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_4686_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_176;
  wire n_179, n_180, n_183, n_184, n_187, n_188, n_189, n_196;
  wire n_201, n_202, n_203, n_204, n_209, n_210, n_211, n_212;
  wire n_217, n_218, n_219, n_220, n_221, n_223, n_224, n_225;
  wire n_226, n_227, n_234, n_236, n_237, n_238, n_239, n_248;
  wire n_249, n_250, n_251, n_258, n_260, n_261, n_262, n_267;
  wire n_269, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_282, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_300, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_333, n_335, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_354;
  wire n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_366, n_367, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477;
  wire n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485;
  wire n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539;
  wire n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_595;
  wire n_596, n_597, n_598, n_599, n_603, n_604, n_605, n_606;
  wire n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_617;
  wire n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629;
  wire n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637;
  wire n_638, n_639, n_640, n_641, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_658, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_668, n_669, n_670, n_671;
  wire n_672, n_673, n_674, n_675, n_676, n_677, n_684, n_685;
  wire n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693;
  wire n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711;
  wire n_712, n_713, n_722, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_738, n_742, n_743;
  wire n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_751;
  wire n_752, n_753, n_764, n_765, n_766, n_767, n_768, n_769;
  wire n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777;
  wire n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801;
  wire n_802, n_803, n_804, n_805, n_822, n_823, n_824, n_826;
  wire n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_842;
  wire n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855;
  wire n_856, n_857, n_858, n_859, n_860, n_861, n_868, n_869;
  wire n_870, n_871, n_872, n_873, n_876, n_877, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_906, n_907, n_908, n_910;
  wire n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918;
  wire n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926;
  wire n_927, n_928, n_929, n_946, n_947, n_949, n_950, n_951;
  wire n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959;
  wire n_960, n_961, n_962, n_963, n_964, n_965, n_984, n_985;
  wire n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993;
  wire n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001;
  wire n_1013, n_1014, n_1015, n_1016, n_1017, n_1020, n_1021, n_1024;
  wire n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040;
  wire n_1041, n_1043, n_1044, n_1047, n_1049, n_1051, n_1052, n_1056;
  wire n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064;
  wire n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072;
  wire n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080;
  wire n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1088, n_1090;
  wire n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098;
  wire n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106;
  wire n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114;
  wire n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122;
  wire n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130;
  wire n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138;
  wire n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146;
  wire n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1154, n_1155;
  wire n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163;
  wire n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171;
  wire n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179;
  wire n_1180, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188;
  wire n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196;
  wire n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204;
  wire n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212;
  wire n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220;
  wire n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228;
  wire n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236;
  wire n_1237, n_1238, n_1239, n_1241, n_1242, n_1243, n_1244, n_1245;
  wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1252, n_1253, n_1254;
  wire n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262;
  wire n_1263, n_1264, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271;
  wire n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279;
  wire n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1288;
  wire n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297;
  wire n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305;
  wire n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313;
  wire n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1324, n_1325;
  wire n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333;
  wire n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341;
  wire n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349;
  wire n_1350, n_1351, n_1352, n_1353, n_1355, n_1356, n_1357, n_1358;
  wire n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366;
  wire n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374;
  wire n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382;
  wire n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390;
  wire n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398;
  wire n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406;
  wire n_1407, n_1408, n_1409, n_1410, n_1412, n_1414, n_1415, n_1416;
  wire n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424;
  wire n_1425, n_1426, n_1427, n_1428, n_1429, n_1432, n_1433, n_1434;
  wire n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442;
  wire n_1443, n_1444, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451;
  wire n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1460, n_1461, n_1463, n_1464, n_1465, n_1466, n_1468, n_1469;
  wire n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477;
  wire n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485;
  wire n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493;
  wire n_1494, n_1495, n_1496, n_1498, n_1499, n_1500, n_1501, n_1502;
  wire n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513;
  wire n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521;
  wire n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531;
  wire n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1539, n_1540;
  wire n_1541, n_1542, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558;
  wire n_1559, n_1560, n_1561, n_1562, n_1565, n_1566, n_1567, n_1568;
  wire n_1569, n_1570, n_1571, n_1572, n_1573, n_1576, n_1577, n_1578;
  wire n_1579, n_1580, n_1581, n_1583, n_1584, n_1585, n_1587, n_1588;
  wire n_1589, n_1593, n_1606, n_1611, n_1612, n_1613, n_1614, n_1615;
  wire n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623;
  wire n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631;
  wire n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639;
  wire n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647;
  wire n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655;
  wire n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663;
  wire n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671;
  wire n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679;
  wire n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687;
  wire n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695;
  wire n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703;
  wire n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711;
  wire n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719;
  wire n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727;
  wire n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735;
  wire n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743;
  wire n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751;
  wire n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759;
  wire n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767;
  wire n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775;
  wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
  wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
  wire n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815;
  wire n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823;
  wire n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], n_171);
  xor g270 (n_117, n_622, A[2]);
  nand g3 (n_623, A[1], n_171);
  nand g271 (n_624, A[2], n_171);
  nand g272 (n_625, A[1], A[2]);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, A[4]);
  xor g288 (n_176, n_634, n_69);
  nand g289 (n_635, n_68, A[4]);
  nand g290 (n_636, n_69, A[4]);
  nand g291 (n_637, n_68, n_69);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_176);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_176);
  nand g296 (n_640, A[7], n_176);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g305 (n_646, n_117, A[5]);
  xor g306 (n_180, n_646, A[6]);
  nand g307 (n_647, n_117, A[5]);
  nand g308 (n_648, A[6], A[5]);
  nand g309 (n_649, n_117, A[6]);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, n_179, n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, n_179, n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, n_179, A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_188, n_659, n_660, n_661);
  xor g329 (n_662, n_183, A[9]);
  xor g330 (n_112, n_662, n_184);
  nand g331 (n_663, n_183, A[9]);
  nand g332 (n_664, n_184, A[9]);
  nand g333 (n_665, n_183, n_184);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_187, n_630, n_67);
  nand g340 (n_668, n_67, n_173);
  nand g341 (n_669, A[4], n_67);
  nand g342 (n_71, n_631, n_668, n_669);
  xor g343 (n_670, A[7], n_187);
  xor g344 (n_189, n_670, A[8]);
  nand g345 (n_671, A[7], n_187);
  nand g346 (n_672, A[8], n_187);
  nand g347 (n_673, A[7], A[8]);
  nand g348 (n_73, n_671, n_672, n_673);
  xor g349 (n_674, n_188, A[10]);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, n_188, A[10]);
  nand g352 (n_676, n_189, A[10]);
  nand g353 (n_677, n_188, n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_72, n_638, n_71);
  nand g366 (n_684, n_71, n_176);
  nand g367 (n_685, A[5], n_71);
  nand g368 (n_201, n_639, n_684, n_685);
  xor g369 (n_686, A[8], A[9]);
  xor g370 (n_196, n_686, n_73);
  nand g371 (n_687, A[8], A[9]);
  nand g372 (n_688, n_73, A[9]);
  nand g373 (n_689, A[8], n_73);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, n_72, A[11]);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, n_72, A[11]);
  nand g378 (n_692, n_196, A[11]);
  nand g379 (n_693, n_72, n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g394 (n_202, n_650, A[9]);
  nand g396 (n_704, A[9], n_180);
  nand g397 (n_705, n_179, A[9]);
  nand g398 (n_209, n_651, n_704, n_705);
  xor g399 (n_706, A[10], n_201);
  xor g400 (n_204, n_706, n_202);
  nand g401 (n_707, A[10], n_201);
  nand g402 (n_708, n_202, n_201);
  nand g403 (n_709, A[10], n_202);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, A[12], n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, A[12], n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, A[12], n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g423 (n_722, n_183, n_184);
  xor g424 (n_210, n_722, A[10]);
  nand g426 (n_724, A[10], n_184);
  nand g427 (n_725, n_183, A[10]);
  nand g428 (n_218, n_665, n_724, n_725);
  xor g429 (n_726, A[11], n_209);
  xor g430 (n_212, n_726, n_210);
  nand g431 (n_727, A[11], n_209);
  nand g432 (n_728, n_210, n_209);
  nand g433 (n_729, A[11], n_210);
  nand g434 (n_220, n_727, n_728, n_729);
  xor g435 (n_730, n_211, A[13]);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, n_211, A[13]);
  nand g438 (n_732, n_212, A[13]);
  nand g439 (n_733, n_211, n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_217, n_738, n_187);
  xor g455 (n_742, n_188, n_217);
  xor g456 (n_219, n_742, A[11]);
  nand g457 (n_743, n_188, n_217);
  nand g458 (n_744, A[11], n_217);
  nand g459 (n_745, n_188, A[11]);
  nand g460 (n_224, n_743, n_744, n_745);
  xor g461 (n_746, A[12], n_218);
  xor g462 (n_221, n_746, A[14]);
  nand g463 (n_747, A[12], n_218);
  nand g464 (n_748, A[14], n_218);
  nand g465 (n_749, A[12], A[14]);
  nand g466 (n_226, n_747, n_748, n_749);
  xor g467 (n_750, n_219, n_220);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, n_219, n_220);
  nand g470 (n_752, n_221, n_220);
  nand g471 (n_753, n_219, n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g488 (n_223, n_686, n_72);
  nand g490 (n_764, n_72, A[9]);
  nand g491 (n_765, A[8], n_72);
  nand g492 (n_234, n_687, n_764, n_765);
  xor g493 (n_766, n_73, A[12]);
  xor g494 (n_225, n_766, n_223);
  nand g495 (n_767, n_73, A[12]);
  nand g496 (n_768, n_223, A[12]);
  nand g497 (n_769, n_73, n_223);
  nand g498 (n_236, n_767, n_768, n_769);
  xor g499 (n_770, A[13], n_224);
  xor g500 (n_227, n_770, n_225);
  nand g501 (n_771, A[13], n_224);
  nand g502 (n_772, n_225, n_224);
  nand g503 (n_773, A[13], n_225);
  nand g504 (n_238, n_771, n_772, n_773);
  xor g505 (n_774, A[15], n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, A[15], n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, A[15], n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g535 (n_794, n_234, A[13]);
  xor g536 (n_237, n_794, n_204);
  nand g537 (n_795, n_234, A[13]);
  nand g538 (n_796, n_204, A[13]);
  nand g539 (n_797, n_234, n_204);
  nand g540 (n_248, n_795, n_796, n_797);
  xor g541 (n_798, A[14], n_236);
  xor g542 (n_239, n_798, A[16]);
  nand g543 (n_799, A[14], n_236);
  nand g544 (n_800, A[16], n_236);
  nand g545 (n_801, A[14], A[16]);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, n_237, n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, n_237, n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, n_237, n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g577 (n_822, n_211, A[14]);
  xor g578 (n_249, n_822, n_212);
  nand g579 (n_823, n_211, A[14]);
  nand g580 (n_824, n_212, A[14]);
  nand g582 (n_261, n_823, n_824, n_733);
  xor g583 (n_826, A[15], n_248);
  xor g584 (n_251, n_826, A[17]);
  nand g585 (n_827, A[15], n_248);
  nand g586 (n_828, A[17], n_248);
  nand g587 (n_829, A[15], A[17]);
  nand g588 (n_118, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g609 (n_842, n_188, A[11]);
  xor g610 (n_258, n_842, n_217);
  xor g616 (n_260, n_746, n_258);
  nand g618 (n_848, n_258, n_218);
  nand g619 (n_849, A[12], n_258);
  nand g620 (n_272, n_747, n_848, n_849);
  xor g621 (n_850, n_220, A[15]);
  xor g622 (n_262, n_850, n_260);
  nand g623 (n_851, n_220, A[15]);
  nand g624 (n_852, n_260, A[15]);
  nand g625 (n_853, n_220, n_260);
  nand g626 (n_274, n_851, n_852, n_853);
  xor g627 (n_854, A[16], n_261);
  xor g628 (n_119, n_854, A[18]);
  nand g629 (n_855, A[16], n_261);
  nand g630 (n_856, A[18], n_261);
  nand g631 (n_857, A[16], A[18]);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_262, n_118);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_262, n_118);
  nand g636 (n_860, n_119, n_118);
  nand g637 (n_861, n_262, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g648 (n_267, n_638, A[8]);
  nand g650 (n_868, A[8], n_176);
  nand g651 (n_869, A[5], A[8]);
  nand g652 (n_282, n_639, n_868, n_869);
  xor g653 (n_870, n_71, A[9]);
  xor g654 (n_269, n_870, n_267);
  nand g655 (n_871, n_71, A[9]);
  nand g656 (n_872, n_267, A[9]);
  nand g657 (n_873, n_71, n_267);
  nand g658 (n_284, n_871, n_872, n_873);
  xor g660 (n_271, n_766, n_269);
  nand g662 (n_876, n_269, A[12]);
  nand g663 (n_877, n_73, n_269);
  nand g664 (n_286, n_767, n_876, n_877);
  xor g666 (n_273, n_770, n_271);
  nand g668 (n_880, n_271, A[13]);
  nand g669 (n_881, n_224, n_271);
  nand g670 (n_288, n_771, n_880, n_881);
  xor g671 (n_882, n_272, A[16]);
  xor g672 (n_275, n_882, n_273);
  nand g673 (n_883, n_272, A[16]);
  nand g674 (n_884, n_273, A[16]);
  nand g675 (n_885, n_272, n_273);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, A[17], n_274);
  xor g678 (n_277, n_886, A[19]);
  nand g679 (n_887, A[17], n_274);
  nand g680 (n_888, A[19], n_274);
  nand g681 (n_889, A[17], A[19]);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g707 (n_906, A[10], n_282);
  xor g708 (n_285, n_906, n_202);
  nand g709 (n_907, A[10], n_282);
  nand g710 (n_908, n_202, n_282);
  nand g712 (n_300, n_907, n_908, n_709);
  xor g713 (n_910, n_284, A[13]);
  xor g714 (n_287, n_910, n_285);
  nand g715 (n_911, n_284, A[13]);
  nand g716 (n_912, n_285, A[13]);
  nand g717 (n_913, n_284, n_285);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, A[14], n_286);
  xor g720 (n_289, n_914, n_287);
  nand g721 (n_915, A[14], n_286);
  nand g722 (n_916, n_287, n_286);
  nand g723 (n_917, A[14], n_287);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, n_288, A[17]);
  xor g726 (n_291, n_918, n_289);
  nand g727 (n_919, n_288, A[17]);
  nand g728 (n_920, n_289, A[17]);
  nand g729 (n_921, n_288, n_289);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, A[18], n_290);
  xor g732 (n_293, n_922, A[20]);
  nand g733 (n_923, A[18], n_290);
  nand g734 (n_924, A[20], n_290);
  nand g735 (n_925, A[18], A[20]);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g767 (n_946, n_300, A[14]);
  xor g768 (n_303, n_946, n_212);
  nand g769 (n_947, n_300, A[14]);
  nand g771 (n_949, n_300, n_212);
  nand g772 (n_319, n_947, n_824, n_949);
  xor g773 (n_950, n_302, A[15]);
  xor g774 (n_305, n_950, n_303);
  nand g775 (n_951, n_302, A[15]);
  nand g776 (n_952, n_303, A[15]);
  nand g777 (n_953, n_302, n_303);
  nand g778 (n_321, n_951, n_952, n_953);
  xor g779 (n_954, n_304, A[18]);
  xor g780 (n_307, n_954, n_305);
  nand g781 (n_955, n_304, A[18]);
  nand g782 (n_956, n_305, A[18]);
  nand g783 (n_957, n_304, n_305);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, A[19], n_306);
  xor g786 (n_309, n_958, A[21]);
  nand g787 (n_959, A[19], n_306);
  nand g788 (n_960, A[21], n_306);
  nand g789 (n_961, A[19], A[21]);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g824 (n_320, n_850, A[16]);
  nand g826 (n_984, A[16], A[15]);
  nand g827 (n_985, n_220, A[16]);
  nand g828 (n_338, n_851, n_984, n_985);
  xor g829 (n_986, n_260, n_319);
  xor g830 (n_322, n_986, n_320);
  nand g831 (n_987, n_260, n_319);
  nand g832 (n_988, n_320, n_319);
  nand g833 (n_989, n_260, n_320);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, n_321, A[19]);
  xor g836 (n_324, n_990, n_322);
  nand g837 (n_991, n_321, A[19]);
  nand g838 (n_992, n_322, A[19]);
  nand g839 (n_993, n_321, n_322);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, A[20], n_323);
  xor g842 (n_326, n_994, A[22]);
  nand g843 (n_995, A[20], n_323);
  nand g844 (n_996, A[22], n_323);
  nand g845 (n_997, A[20], A[22]);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, n_324, n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, n_324, n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, n_324, n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g868 (n_333, n_870, n_73);
  nand g871 (n_1013, n_71, n_73);
  nand g872 (n_354, n_871, n_688, n_1013);
  xor g873 (n_1014, n_267, A[12]);
  xor g874 (n_335, n_1014, n_333);
  nand g875 (n_1015, n_267, A[12]);
  nand g876 (n_1016, n_333, A[12]);
  nand g877 (n_1017, n_267, n_333);
  nand g878 (n_356, n_1015, n_1016, n_1017);
  xor g880 (n_337, n_770, n_335);
  nand g882 (n_1020, n_335, A[13]);
  nand g883 (n_1021, n_224, n_335);
  nand g884 (n_358, n_771, n_1020, n_1021);
  xor g886 (n_339, n_882, n_337);
  nand g888 (n_1024, n_337, A[16]);
  nand g889 (n_1025, n_272, n_337);
  nand g890 (n_360, n_883, n_1024, n_1025);
  xor g891 (n_1026, A[17], n_338);
  xor g892 (n_341, n_1026, n_339);
  nand g893 (n_1027, A[17], n_338);
  nand g894 (n_1028, n_339, n_338);
  nand g895 (n_1029, A[17], n_339);
  nand g896 (n_362, n_1027, n_1028, n_1029);
  xor g897 (n_1030, A[20], n_340);
  xor g898 (n_343, n_1030, n_341);
  nand g899 (n_1031, A[20], n_340);
  nand g900 (n_1032, n_341, n_340);
  nand g901 (n_1033, A[20], n_341);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, A[21], n_342);
  xor g904 (n_345, n_1034, n_343);
  nand g905 (n_1035, A[21], n_342);
  nand g906 (n_1036, n_343, n_342);
  nand g907 (n_1037, A[21], n_343);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, A[23], n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, A[23], n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, A[23], n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  nand g922 (n_371, n_1043, n_1044, n_624);
  nand g928 (n_373, n_1047, n_648, n_1049);
  nand g934 (n_375, n_1051, n_1052, n_705);
  nand g940 (n_377, n_907, n_1056, n_1057);
  xor g941 (n_1058, n_354, A[13]);
  nand g943 (n_1059, n_354, A[13]);
  nand g946 (n_379, n_1059, n_1060, n_1061);
  xor g947 (n_1062, A[14], n_356);
  xor g948 (n_359, n_1062, n_357);
  nand g949 (n_1063, A[14], n_356);
  nand g950 (n_1064, n_357, n_356);
  nand g951 (n_1065, A[14], n_357);
  nand g952 (n_381, n_1063, n_1064, n_1065);
  xor g953 (n_1066, n_358, A[17]);
  xor g954 (n_361, n_1066, A[18]);
  nand g955 (n_1067, n_358, A[17]);
  nand g956 (n_1068, A[18], A[17]);
  nand g957 (n_1069, n_358, A[18]);
  nand g958 (n_383, n_1067, n_1068, n_1069);
  xor g959 (n_1070, n_359, n_360);
  xor g960 (n_363, n_1070, n_361);
  nand g961 (n_1071, n_359, n_360);
  nand g962 (n_1072, n_361, n_360);
  nand g963 (n_1073, n_359, n_361);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, A[21], n_362);
  xor g966 (n_365, n_1074, A[22]);
  nand g967 (n_1075, A[21], n_362);
  nand g968 (n_1076, A[22], n_362);
  nand g969 (n_1077, A[21], A[22]);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g972 (n_367, n_1078, n_364);
  nand g975 (n_1081, n_363, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  xor g986 (n_372, n_1086, A[3]);
  nand g990 (n_392, n_1044, n_1088, n_627);
  xor g991 (n_1090, n_371, n_372);
  xor g992 (n_374, n_1090, A[6]);
  nand g993 (n_1091, n_371, n_372);
  nand g994 (n_1092, A[6], n_372);
  nand g995 (n_1093, n_371, A[6]);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, n_374);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, n_374, n_373);
  nand g1001 (n_1097, A[7], n_374);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, A[10], A[11]);
  xor g1004 (n_378, n_1098, n_375);
  nand g1005 (n_1099, A[10], A[11]);
  nand g1006 (n_1100, n_375, A[11]);
  nand g1007 (n_1101, A[10], n_375);
  nand g1008 (n_398, n_1099, n_1100, n_1101);
  xor g1009 (n_1102, n_376, n_377);
  xor g1010 (n_380, n_1102, n_378);
  nand g1011 (n_1103, n_376, n_377);
  nand g1012 (n_1104, n_378, n_377);
  nand g1013 (n_1105, n_376, n_378);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, A[14], n_379);
  xor g1016 (n_382, n_1106, A[15]);
  nand g1017 (n_1107, A[14], n_379);
  nand g1018 (n_1108, A[15], n_379);
  nand g1019 (n_1109, A[14], A[15]);
  nand g1020 (n_402, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, n_380, A[18]);
  xor g1022 (n_384, n_1110, n_381);
  nand g1023 (n_1111, n_380, A[18]);
  nand g1024 (n_1112, n_381, A[18]);
  nand g1025 (n_1113, n_380, n_381);
  nand g1026 (n_404, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, n_382, A[19]);
  xor g1028 (n_386, n_1114, n_383);
  nand g1029 (n_1115, n_382, A[19]);
  nand g1030 (n_1116, n_383, A[19]);
  nand g1031 (n_1117, n_382, n_383);
  nand g1032 (n_406, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_384, A[22]);
  xor g1034 (n_388, n_1118, n_385);
  nand g1035 (n_1119, n_384, A[22]);
  nand g1036 (n_1120, n_385, A[22]);
  nand g1037 (n_1121, n_384, n_385);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, n_386, A[23]);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, n_386, A[23]);
  nand g1042 (n_1124, n_387, A[23]);
  nand g1043 (n_1125, n_386, n_387);
  nand g1044 (n_410, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1051 (n_1130, A[1], A[3]);
  xor g1052 (n_393, n_1130, A[4]);
  nand g1053 (n_1131, A[1], A[3]);
  nand g1054 (n_1132, A[4], A[3]);
  nand g1055 (n_1133, A[1], A[4]);
  nand g1056 (n_412, n_1131, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, n_396, A[11]);
  xor g1070 (n_399, n_1142, A[12]);
  nand g1071 (n_1143, n_396, A[11]);
  nand g1072 (n_1144, A[12], A[11]);
  nand g1073 (n_1145, n_396, A[12]);
  nand g1074 (n_418, n_1143, n_1144, n_1145);
  xor g1075 (n_1146, n_397, n_398);
  xor g1076 (n_401, n_1146, n_399);
  nand g1077 (n_1147, n_397, n_398);
  nand g1078 (n_1148, n_399, n_398);
  nand g1079 (n_1149, n_397, n_399);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, A[15], n_400);
  xor g1082 (n_403, n_1150, A[16]);
  nand g1083 (n_1151, A[15], n_400);
  nand g1084 (n_1152, A[16], n_400);
  nand g1086 (n_421, n_1151, n_1152, n_984);
  xor g1087 (n_1154, n_401, n_402);
  xor g1088 (n_405, n_1154, A[19]);
  nand g1089 (n_1155, n_401, n_402);
  nand g1090 (n_1156, A[19], n_402);
  nand g1091 (n_1157, n_401, A[19]);
  nand g1092 (n_424, n_1155, n_1156, n_1157);
  xor g1093 (n_1158, n_403, n_404);
  xor g1094 (n_407, n_1158, A[20]);
  nand g1095 (n_1159, n_403, n_404);
  nand g1096 (n_1160, A[20], n_404);
  nand g1097 (n_1161, n_403, A[20]);
  nand g1098 (n_425, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_405, n_406);
  xor g1100 (n_409, n_1162, n_407);
  nand g1101 (n_1163, n_405, n_406);
  nand g1102 (n_1164, n_407, n_406);
  nand g1103 (n_1165, n_405, n_407);
  nand g1104 (n_428, n_1163, n_1164, n_1165);
  xor g1106 (n_411, n_1166, n_408);
  nand g1108 (n_1168, n_408, A[23]);
  nand g1110 (n_430, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1123 (n_1178, A[8], n_413);
  xor g1124 (n_415, n_1178, A[9]);
  nand g1125 (n_1179, A[8], n_413);
  nand g1126 (n_1180, A[9], n_413);
  nand g1128 (n_435, n_1179, n_1180, n_687);
  xor g1129 (n_1182, n_414, n_415);
  xor g1130 (n_417, n_1182, A[12]);
  nand g1131 (n_1183, n_414, n_415);
  nand g1132 (n_1184, A[12], n_415);
  nand g1133 (n_1185, n_414, A[12]);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, n_416, A[13]);
  xor g1136 (n_420, n_1186, n_417);
  nand g1137 (n_1187, n_416, A[13]);
  nand g1138 (n_1188, n_417, A[13]);
  nand g1139 (n_1189, n_416, n_417);
  nand g1140 (n_439, n_1187, n_1188, n_1189);
  xor g1141 (n_1190, n_418, n_419);
  xor g1142 (n_422, n_1190, A[16]);
  nand g1143 (n_1191, n_418, n_419);
  nand g1144 (n_1192, A[16], n_419);
  nand g1145 (n_1193, n_418, A[16]);
  nand g1146 (n_440, n_1191, n_1192, n_1193);
  xor g1147 (n_1194, n_420, A[17]);
  xor g1148 (n_423, n_1194, n_421);
  nand g1149 (n_1195, n_420, A[17]);
  nand g1150 (n_1196, n_421, A[17]);
  nand g1151 (n_1197, n_420, n_421);
  nand g1152 (n_442, n_1195, n_1196, n_1197);
  xor g1153 (n_1198, n_422, A[20]);
  xor g1154 (n_426, n_1198, n_423);
  nand g1155 (n_1199, n_422, A[20]);
  nand g1156 (n_1200, n_423, A[20]);
  nand g1157 (n_1201, n_422, n_423);
  nand g1158 (n_445, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_424, A[21]);
  xor g1160 (n_427, n_1202, n_425);
  nand g1161 (n_1203, n_424, A[21]);
  nand g1162 (n_1204, n_425, A[21]);
  nand g1163 (n_1205, n_424, n_425);
  nand g1164 (n_447, n_1203, n_1204, n_1205);
  xor g1166 (n_429, n_1206, n_427);
  nand g1168 (n_1208, n_427, n_426);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, n_433);
  nand g1183 (n_1217, A[6], n_433);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, A[9], A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, A[9], A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, A[9], n_434);
  nand g1190 (n_455, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, n_435, n_436);
  xor g1192 (n_438, n_1222, A[13]);
  nand g1193 (n_1223, n_435, n_436);
  nand g1194 (n_1224, A[13], n_436);
  nand g1195 (n_1225, n_435, A[13]);
  nand g1196 (n_457, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, A[14], n_437);
  xor g1198 (n_441, n_1226, n_438);
  nand g1199 (n_1227, A[14], n_437);
  nand g1200 (n_1228, n_438, n_437);
  nand g1201 (n_1229, A[14], n_438);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, n_439, A[17]);
  xor g1204 (n_443, n_1230, n_440);
  nand g1205 (n_1231, n_439, A[17]);
  nand g1206 (n_1232, n_440, A[17]);
  nand g1207 (n_1233, n_439, n_440);
  nand g1208 (n_461, n_1231, n_1232, n_1233);
  xor g1209 (n_1234, A[18], n_441);
  xor g1210 (n_444, n_1234, n_442);
  nand g1211 (n_1235, A[18], n_441);
  nand g1212 (n_1236, n_442, n_441);
  nand g1213 (n_1237, A[18], n_442);
  nand g1214 (n_464, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_443, A[21]);
  xor g1216 (n_446, n_1238, A[22]);
  nand g1217 (n_1239, n_443, A[21]);
  nand g1219 (n_1241, n_443, A[22]);
  nand g1220 (n_465, n_1239, n_1077, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[5], A[7]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], n_453);
  xor g1242 (n_456, n_1254, n_454);
  nand g1243 (n_1255, A[10], n_453);
  nand g1244 (n_1256, n_454, n_453);
  nand g1245 (n_1257, A[10], n_454);
  nand g1246 (n_472, n_1255, n_1256, n_1257);
  xor g1247 (n_1258, A[11], n_455);
  xor g1248 (n_458, n_1258, n_456);
  nand g1249 (n_1259, A[11], n_455);
  nand g1250 (n_1260, n_456, n_455);
  nand g1251 (n_1261, A[11], n_456);
  nand g1252 (n_474, n_1259, n_1260, n_1261);
  xor g1253 (n_1262, A[14], n_457);
  xor g1254 (n_460, n_1262, A[15]);
  nand g1255 (n_1263, A[14], n_457);
  nand g1256 (n_1264, A[15], n_457);
  nand g1258 (n_476, n_1263, n_1264, n_1109);
  xor g1259 (n_1266, n_458, A[18]);
  xor g1260 (n_462, n_1266, n_459);
  nand g1261 (n_1267, n_458, A[18]);
  nand g1262 (n_1268, n_459, A[18]);
  nand g1263 (n_1269, n_458, n_459);
  nand g1264 (n_479, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, n_460, A[19]);
  xor g1266 (n_463, n_1270, n_461);
  nand g1267 (n_1271, n_460, A[19]);
  nand g1268 (n_1272, n_461, A[19]);
  nand g1269 (n_1273, n_460, n_461);
  nand g1270 (n_480, n_1271, n_1272, n_1273);
  xor g1271 (n_1274, n_462, A[22]);
  xor g1272 (n_466, n_1274, n_463);
  nand g1273 (n_1275, n_462, A[22]);
  nand g1274 (n_1276, n_463, A[22]);
  nand g1275 (n_1277, n_462, n_463);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1277 (n_1278, n_464, A[23]);
  xor g1278 (n_467, n_1278, n_465);
  nand g1279 (n_1279, n_464, A[23]);
  nand g1280 (n_1280, n_465, A[23]);
  nand g1281 (n_1281, n_464, n_465);
  nand g1282 (n_484, n_1279, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1289 (n_1286, A[7], A[6]);
  xor g1290 (n_471, n_1286, A[8]);
  nand g1292 (n_1288, A[8], A[6]);
  nand g1294 (n_486, n_661, n_1288, n_673);
  xor g1295 (n_1290, n_470, n_471);
  xor g1296 (n_473, n_1290, A[11]);
  nand g1297 (n_1291, n_470, n_471);
  nand g1298 (n_1292, A[11], n_471);
  nand g1299 (n_1293, n_470, A[11]);
  nand g1300 (n_488, n_1291, n_1292, n_1293);
  xor g1301 (n_1294, A[12], n_472);
  xor g1302 (n_475, n_1294, n_473);
  nand g1303 (n_1295, A[12], n_472);
  nand g1304 (n_1296, n_473, n_472);
  nand g1305 (n_1297, A[12], n_473);
  nand g1306 (n_489, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, A[15], n_474);
  xor g1308 (n_477, n_1298, n_475);
  nand g1309 (n_1299, A[15], n_474);
  nand g1310 (n_1300, n_475, n_474);
  nand g1311 (n_1301, A[15], n_475);
  nand g1312 (n_491, n_1299, n_1300, n_1301);
  xor g1313 (n_1302, A[16], n_476);
  xor g1314 (n_478, n_1302, n_477);
  nand g1315 (n_1303, A[16], n_476);
  nand g1316 (n_1304, n_477, n_476);
  nand g1317 (n_1305, A[16], n_477);
  nand g1318 (n_494, n_1303, n_1304, n_1305);
  xor g1319 (n_1306, A[19], n_478);
  xor g1320 (n_481, n_1306, n_479);
  nand g1321 (n_1307, A[19], n_478);
  nand g1322 (n_1308, n_479, n_478);
  nand g1323 (n_1309, A[19], n_479);
  nand g1324 (n_496, n_1307, n_1308, n_1309);
  xor g1325 (n_1310, A[20], n_480);
  xor g1326 (n_483, n_1310, n_481);
  nand g1327 (n_1311, A[20], n_480);
  nand g1328 (n_1312, n_481, n_480);
  nand g1329 (n_1313, A[20], n_481);
  nand g1330 (n_498, n_1311, n_1312, n_1313);
  xor g1332 (n_485, n_1166, n_482);
  nand g1335 (n_1317, A[23], n_482);
  nand g1336 (n_500, n_1167, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1344 (n_487, n_686, n_486);
  nand g1346 (n_1324, n_486, A[9]);
  nand g1347 (n_1325, A[8], n_486);
  nand g1348 (n_503, n_687, n_1324, n_1325);
  xor g1349 (n_1326, A[12], n_487);
  xor g1350 (n_490, n_1326, n_488);
  nand g1351 (n_1327, A[12], n_487);
  nand g1352 (n_1328, n_488, n_487);
  nand g1353 (n_1329, A[12], n_488);
  nand g1354 (n_505, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, A[13], n_489);
  xor g1356 (n_492, n_1330, n_490);
  nand g1357 (n_1331, A[13], n_489);
  nand g1358 (n_1332, n_490, n_489);
  nand g1359 (n_1333, A[13], n_490);
  nand g1360 (n_507, n_1331, n_1332, n_1333);
  xor g1361 (n_1334, A[16], A[17]);
  xor g1362 (n_493, n_1334, n_491);
  nand g1363 (n_1335, A[16], A[17]);
  nand g1364 (n_1336, n_491, A[17]);
  nand g1365 (n_1337, A[16], n_491);
  nand g1366 (n_509, n_1335, n_1336, n_1337);
  xor g1367 (n_1338, n_492, n_493);
  xor g1368 (n_495, n_1338, A[20]);
  nand g1369 (n_1339, n_492, n_493);
  nand g1370 (n_1340, A[20], n_493);
  nand g1371 (n_1341, n_492, A[20]);
  nand g1372 (n_511, n_1339, n_1340, n_1341);
  xor g1373 (n_1342, n_494, A[21]);
  xor g1374 (n_497, n_1342, n_495);
  nand g1375 (n_1343, n_494, A[21]);
  nand g1376 (n_1344, n_495, A[21]);
  nand g1377 (n_1345, n_494, n_495);
  nand g1378 (n_513, n_1343, n_1344, n_1345);
  xor g1380 (n_499, n_1346, n_497);
  nand g1383 (n_1349, n_496, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  nand g1397 (n_1357, A[10], n_503);
  nand g1398 (n_520, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], A[14]);
  xor g1400 (n_506, n_1358, n_504);
  nand g1401 (n_1359, A[13], A[14]);
  nand g1402 (n_1360, n_504, A[14]);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_521, n_1359, n_1360, n_1361);
  xor g1405 (n_1362, n_505, A[17]);
  xor g1406 (n_508, n_1362, n_506);
  nand g1407 (n_1363, n_505, A[17]);
  nand g1408 (n_1364, n_506, A[17]);
  nand g1409 (n_1365, n_505, n_506);
  nand g1410 (n_523, n_1363, n_1364, n_1365);
  xor g1411 (n_1366, n_507, A[18]);
  xor g1412 (n_510, n_1366, n_508);
  nand g1413 (n_1367, n_507, A[18]);
  nand g1414 (n_1368, n_508, A[18]);
  nand g1415 (n_1369, n_507, n_508);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_509, A[21]);
  xor g1418 (n_512, n_1370, n_510);
  nand g1419 (n_1371, n_509, A[21]);
  nand g1420 (n_1372, n_510, A[21]);
  nand g1421 (n_1373, n_509, n_510);
  nand g1422 (n_527, n_1371, n_1372, n_1373);
  xor g1423 (n_1374, A[22], n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, A[22], n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, A[22], n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1437 (n_1382, A[9], A[11]);
  nand g1439 (n_1383, A[9], A[11]);
  nand g1442 (n_532, n_1383, n_1384, n_1385);
  xor g1443 (n_1386, A[14], n_519);
  xor g1444 (n_522, n_1386, n_520);
  nand g1445 (n_1387, A[14], n_519);
  nand g1446 (n_1388, n_520, n_519);
  nand g1447 (n_1389, A[14], n_520);
  nand g1448 (n_534, n_1387, n_1388, n_1389);
  xor g1449 (n_1390, A[15], n_521);
  xor g1450 (n_524, n_1390, n_522);
  nand g1451 (n_1391, A[15], n_521);
  nand g1452 (n_1392, n_522, n_521);
  nand g1453 (n_1393, A[15], n_522);
  nand g1454 (n_536, n_1391, n_1392, n_1393);
  xor g1455 (n_1394, A[18], n_523);
  xor g1456 (n_525, n_1394, A[19]);
  nand g1457 (n_1395, A[18], n_523);
  nand g1458 (n_1396, A[19], n_523);
  nand g1459 (n_1397, A[18], A[19]);
  nand g1460 (n_538, n_1395, n_1396, n_1397);
  xor g1461 (n_1398, n_524, n_525);
  xor g1462 (n_528, n_1398, n_526);
  nand g1463 (n_1399, n_524, n_525);
  nand g1464 (n_1400, n_526, n_525);
  nand g1465 (n_1401, n_524, n_526);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1467 (n_1402, A[22], A[23]);
  xor g1468 (n_529, n_1402, n_527);
  nand g1469 (n_1403, A[22], A[23]);
  nand g1470 (n_1404, n_527, A[23]);
  nand g1471 (n_1405, A[22], n_527);
  nand g1472 (n_543, n_1403, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1479 (n_1410, A[11], A[12]);
  xor g1480 (n_533, n_1410, A[10]);
  nand g1482 (n_1412, A[10], A[12]);
  nand g1484 (n_544, n_1144, n_1412, n_1099);
  xor g1485 (n_1414, n_532, n_533);
  xor g1486 (n_535, n_1414, A[15]);
  nand g1487 (n_1415, n_532, n_533);
  nand g1488 (n_1416, A[15], n_533);
  nand g1489 (n_1417, n_532, A[15]);
  nand g1490 (n_546, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, A[16], n_534);
  xor g1492 (n_537, n_1418, n_535);
  nand g1493 (n_1419, A[16], n_534);
  nand g1494 (n_1420, n_535, n_534);
  nand g1495 (n_1421, A[16], n_535);
  nand g1496 (n_548, n_1419, n_1420, n_1421);
  xor g1497 (n_1422, A[19], n_536);
  xor g1498 (n_539, n_1422, n_537);
  nand g1499 (n_1423, A[19], n_536);
  nand g1500 (n_1424, n_537, n_536);
  nand g1501 (n_1425, A[19], n_537);
  nand g1502 (n_549, n_1423, n_1424, n_1425);
  xor g1503 (n_1426, A[20], n_538);
  xor g1504 (n_541, n_1426, n_539);
  nand g1505 (n_1427, A[20], n_538);
  nand g1506 (n_1428, n_539, n_538);
  nand g1507 (n_1429, A[20], n_539);
  nand g1508 (n_551, n_1427, n_1428, n_1429);
  xor g1510 (n_542, n_1166, n_540);
  nand g1513 (n_1433, A[23], n_540);
  nand g1514 (n_554, n_1167, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1521 (n_1438, A[12], A[13]);
  xor g1522 (n_545, n_1438, n_544);
  nand g1523 (n_1439, A[12], A[13]);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_1439, n_1440, n_1441);
  xor g1527 (n_1442, A[16], n_545);
  xor g1528 (n_547, n_1442, A[17]);
  nand g1529 (n_1443, A[16], n_545);
  nand g1530 (n_1444, A[17], n_545);
  nand g1532 (n_559, n_1443, n_1444, n_1335);
  xor g1533 (n_1446, n_546, n_547);
  xor g1534 (n_550, n_1446, n_548);
  nand g1535 (n_1447, n_546, n_547);
  nand g1536 (n_1448, n_548, n_547);
  nand g1537 (n_1449, n_546, n_548);
  nand g1538 (n_561, n_1447, n_1448, n_1449);
  xor g1539 (n_1450, A[20], A[21]);
  xor g1540 (n_552, n_1450, n_549);
  nand g1541 (n_1451, A[20], A[21]);
  nand g1542 (n_1452, n_549, A[21]);
  nand g1543 (n_1453, A[20], n_549);
  nand g1544 (n_562, n_1451, n_1452, n_1453);
  xor g1546 (n_553, n_1454, n_551);
  nand g1549 (n_1457, n_550, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1563 (n_1465, A[14], n_557);
  nand g1564 (n_569, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, A[17], A[18]);
  xor g1566 (n_560, n_1466, n_558);
  nand g1568 (n_1468, n_558, A[18]);
  nand g1569 (n_1469, A[17], n_558);
  nand g1570 (n_571, n_1068, n_1468, n_1469);
  xor g1571 (n_1470, n_559, n_560);
  xor g1572 (n_563, n_1470, A[21]);
  nand g1573 (n_1471, n_559, n_560);
  nand g1574 (n_1472, A[21], n_560);
  nand g1575 (n_1473, n_559, A[21]);
  nand g1576 (n_574, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, A[22], n_561);
  xor g1578 (n_564, n_1474, n_562);
  nand g1579 (n_1475, A[22], n_561);
  nand g1580 (n_1476, n_562, n_561);
  nand g1581 (n_1477, A[22], n_562);
  nand g1582 (n_576, n_1475, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  xor g1591 (n_1482, A[13], A[15]);
  nand g1593 (n_1483, A[13], A[15]);
  nand g1596 (n_578, n_1483, n_1484, n_1485);
  xor g1597 (n_1486, A[18], n_569);
  xor g1598 (n_572, n_1486, n_570);
  nand g1599 (n_1487, A[18], n_569);
  nand g1600 (n_1488, n_570, n_569);
  nand g1601 (n_1489, A[18], n_570);
  nand g1602 (n_580, n_1487, n_1488, n_1489);
  xor g1603 (n_1490, A[19], n_571);
  xor g1604 (n_573, n_1490, n_572);
  nand g1605 (n_1491, A[19], n_571);
  nand g1606 (n_1492, n_572, n_571);
  nand g1607 (n_1493, A[19], n_572);
  nand g1608 (n_582, n_1491, n_1492, n_1493);
  xor g1609 (n_1494, A[22], n_573);
  xor g1610 (n_575, n_1494, A[23]);
  nand g1611 (n_1495, A[22], n_573);
  nand g1612 (n_1496, A[23], n_573);
  nand g1614 (n_584, n_1495, n_1496, n_1403);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1621 (n_1502, A[15], A[14]);
  xor g1622 (n_579, n_1502, A[16]);
  nand g1626 (n_586, n_1109, n_801, n_984);
  xor g1627 (n_1506, n_578, n_579);
  xor g1628 (n_581, n_1506, A[19]);
  nand g1629 (n_1507, n_578, n_579);
  nand g1630 (n_1508, A[19], n_579);
  nand g1631 (n_1509, n_578, A[19]);
  nand g1632 (n_588, n_1507, n_1508, n_1509);
  xor g1633 (n_1510, n_580, A[20]);
  xor g1634 (n_583, n_1510, n_581);
  nand g1635 (n_1511, n_580, A[20]);
  nand g1636 (n_1512, n_581, A[20]);
  nand g1637 (n_1513, n_580, n_581);
  nand g1638 (n_589, n_1511, n_1512, n_1513);
  xor g1639 (n_1514, n_582, n_583);
  xor g1640 (n_585, n_1514, A[23]);
  nand g1641 (n_1515, n_582, n_583);
  nand g1642 (n_1516, A[23], n_583);
  nand g1643 (n_1517, n_582, A[23]);
  nand g1644 (n_591, n_1515, n_1516, n_1517);
  xor g1646 (n_83, n_1518, n_585);
  nand g1648 (n_1520, n_585, n_584);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1652 (n_587, n_1334, n_586);
  nand g1654 (n_1524, n_586, A[17]);
  nand g1655 (n_1525, A[16], n_586);
  nand g1656 (n_595, n_1335, n_1524, n_1525);
  xor g1657 (n_1526, A[20], n_587);
  xor g1658 (n_590, n_1526, n_588);
  nand g1659 (n_1527, A[20], n_587);
  nand g1660 (n_1528, n_588, n_587);
  nand g1661 (n_1529, A[20], n_588);
  nand g1662 (n_597, n_1527, n_1528, n_1529);
  xor g1664 (n_592, n_1530, n_589);
  nand g1667 (n_1533, A[21], n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_81, n_1535, n_1536, n_1537);
  nand g1681 (n_1541, A[18], n_595);
  nand g1682 (n_604, n_1539, n_1540, n_1541);
  xor g1683 (n_1542, A[21], A[22]);
  xor g1684 (n_598, n_1542, n_596);
  nand g1686 (n_1544, n_596, A[22]);
  nand g1687 (n_1545, A[21], n_596);
  nand g1688 (n_606, n_1077, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_33, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[17], A[19]);
  nand g1702 (n_608, n_889, n_1552, n_1553);
  xor g1703 (n_1554, A[22], n_603);
  xor g1704 (n_605, n_1554, n_604);
  nand g1705 (n_1555, A[22], n_603);
  nand g1706 (n_1556, n_604, n_603);
  nand g1707 (n_1557, A[22], n_604);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, A[23], n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, A[23], n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, A[23], n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1715 (n_1562, A[19], A[18]);
  xor g1716 (n_609, n_1562, A[20]);
  nand g1719 (n_1565, A[19], A[20]);
  nand g1720 (n_612, n_1397, n_925, n_1565);
  xor g1721 (n_1566, n_608, n_609);
  xor g1722 (n_611, n_1566, A[23]);
  nand g1723 (n_1567, n_608, n_609);
  nand g1724 (n_1568, A[23], n_609);
  nand g1725 (n_1569, n_608, A[23]);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1728 (n_79, n_1570, n_611);
  nand g1730 (n_1572, n_611, n_610);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1734 (n_613, n_1450, n_612);
  nand g1736 (n_1576, n_612, A[21]);
  nand g1737 (n_1577, A[20], n_612);
  nand g1738 (n_617, n_1451, n_1576, n_1577);
  xor g1740 (n_78, n_1578, n_614);
  nand g1742 (n_1580, n_614, n_613);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_617);
  nand g1752 (n_76, n_1583, n_1584, n_1585);
  nand g1759 (n_1589, A[21], A[23]);
  nand g1760 (n_27, n_1587, n_1588, n_1589);
  xor g1762 (n_75, n_1166, A[22]);
  nand g1766 (n_74, n_1167, n_1403, n_1593);
  nand g16 (n_1606, A[0], A[2]);
  xor g20 (Z[2], A[0], A[2]);
  nand g22 (n_1611, n_68, A[3]);
  nand g25 (n_1615, n_1611, n_1612, n_1613);
  xor g26 (n_1614, n_68, A[3]);
  nand g28 (n_1616, A[4], n_117);
  nand g29 (n_1617, A[4], n_1615);
  nand g30 (n_1618, n_117, n_1615);
  nand g31 (n_1620, n_1616, n_1617, n_1618);
  xor g32 (n_1619, A[4], n_117);
  xor g33 (Z[4], n_1615, n_1619);
  nand g34 (n_1621, A[5], n_116);
  nand g35 (n_1622, A[5], n_1620);
  nand g36 (n_1623, n_116, n_1620);
  nand g37 (n_1625, n_1621, n_1622, n_1623);
  xor g38 (n_1624, A[5], n_116);
  xor g39 (Z[5], n_1620, n_1624);
  nand g40 (n_1626, n_67, n_115);
  nand g41 (n_1627, n_67, n_1625);
  nand g42 (n_1628, n_115, n_1625);
  nand g43 (n_1630, n_1626, n_1627, n_1628);
  xor g44 (n_1629, n_67, n_115);
  xor g45 (Z[6], n_1625, n_1629);
  nand g46 (n_1631, n_66, n_114);
  nand g47 (n_1632, n_66, n_1630);
  nand g48 (n_1633, n_114, n_1630);
  nand g49 (n_1635, n_1631, n_1632, n_1633);
  xor g50 (n_1634, n_66, n_114);
  xor g51 (Z[7], n_1630, n_1634);
  nand g52 (n_1636, n_65, n_113);
  nand g53 (n_1637, n_65, n_1635);
  nand g54 (n_1638, n_113, n_1635);
  nand g55 (n_1640, n_1636, n_1637, n_1638);
  xor g56 (n_1639, n_65, n_113);
  xor g57 (Z[8], n_1635, n_1639);
  nand g58 (n_1641, n_64, n_112);
  nand g59 (n_1642, n_64, n_1640);
  nand g60 (n_1643, n_112, n_1640);
  nand g61 (n_1645, n_1641, n_1642, n_1643);
  xor g62 (n_1644, n_64, n_112);
  xor g63 (Z[9], n_1640, n_1644);
  nand g64 (n_1646, n_63, n_111);
  nand g65 (n_1647, n_63, n_1645);
  nand g66 (n_1648, n_111, n_1645);
  nand g67 (n_1650, n_1646, n_1647, n_1648);
  xor g68 (n_1649, n_63, n_111);
  xor g69 (Z[10], n_1645, n_1649);
  nand g70 (n_1651, n_62, n_110);
  nand g71 (n_1652, n_62, n_1650);
  nand g72 (n_1653, n_110, n_1650);
  nand g73 (n_1655, n_1651, n_1652, n_1653);
  xor g74 (n_1654, n_62, n_110);
  xor g75 (Z[11], n_1650, n_1654);
  nand g76 (n_1656, n_61, n_109);
  nand g77 (n_1657, n_61, n_1655);
  nand g78 (n_1658, n_109, n_1655);
  nand g79 (n_1660, n_1656, n_1657, n_1658);
  xor g80 (n_1659, n_61, n_109);
  xor g81 (Z[12], n_1655, n_1659);
  nand g82 (n_1661, n_60, n_108);
  nand g83 (n_1662, n_60, n_1660);
  nand g84 (n_1663, n_108, n_1660);
  nand g85 (n_1665, n_1661, n_1662, n_1663);
  xor g86 (n_1664, n_60, n_108);
  xor g87 (Z[13], n_1660, n_1664);
  nand g88 (n_1666, n_59, n_107);
  nand g89 (n_1667, n_59, n_1665);
  nand g90 (n_1668, n_107, n_1665);
  nand g91 (n_1670, n_1666, n_1667, n_1668);
  xor g92 (n_1669, n_59, n_107);
  xor g93 (Z[14], n_1665, n_1669);
  nand g94 (n_1671, n_58, n_106);
  nand g95 (n_1672, n_58, n_1670);
  nand g96 (n_1673, n_106, n_1670);
  nand g97 (n_1675, n_1671, n_1672, n_1673);
  xor g98 (n_1674, n_58, n_106);
  xor g99 (Z[15], n_1670, n_1674);
  nand g100 (n_1676, n_57, n_105);
  nand g101 (n_1677, n_57, n_1675);
  nand g102 (n_1678, n_105, n_1675);
  nand g103 (n_1680, n_1676, n_1677, n_1678);
  xor g104 (n_1679, n_57, n_105);
  xor g105 (Z[16], n_1675, n_1679);
  nand g106 (n_1681, n_56, n_104);
  nand g107 (n_1682, n_56, n_1680);
  nand g108 (n_1683, n_104, n_1680);
  nand g109 (n_1685, n_1681, n_1682, n_1683);
  xor g110 (n_1684, n_56, n_104);
  xor g111 (Z[17], n_1680, n_1684);
  nand g112 (n_1686, n_55, n_103);
  nand g113 (n_1687, n_55, n_1685);
  nand g114 (n_1688, n_103, n_1685);
  nand g115 (n_1690, n_1686, n_1687, n_1688);
  xor g116 (n_1689, n_55, n_103);
  xor g117 (Z[18], n_1685, n_1689);
  nand g118 (n_1691, n_54, n_102);
  nand g119 (n_1692, n_54, n_1690);
  nand g120 (n_1693, n_102, n_1690);
  nand g121 (n_1695, n_1691, n_1692, n_1693);
  xor g122 (n_1694, n_54, n_102);
  xor g123 (Z[19], n_1690, n_1694);
  nand g124 (n_1696, n_53, n_101);
  nand g125 (n_1697, n_53, n_1695);
  nand g126 (n_1698, n_101, n_1695);
  nand g127 (n_1700, n_1696, n_1697, n_1698);
  xor g128 (n_1699, n_53, n_101);
  xor g129 (Z[20], n_1695, n_1699);
  nand g130 (n_1701, n_52, n_100);
  nand g131 (n_1702, n_52, n_1700);
  nand g132 (n_1703, n_100, n_1700);
  nand g133 (n_1705, n_1701, n_1702, n_1703);
  xor g134 (n_1704, n_52, n_100);
  xor g135 (Z[21], n_1700, n_1704);
  nand g136 (n_1706, n_51, n_99);
  nand g137 (n_1707, n_51, n_1705);
  nand g138 (n_1708, n_99, n_1705);
  nand g139 (n_1710, n_1706, n_1707, n_1708);
  xor g140 (n_1709, n_51, n_99);
  xor g141 (Z[22], n_1705, n_1709);
  nand g142 (n_1711, n_50, n_98);
  nand g143 (n_1712, n_50, n_1710);
  nand g144 (n_1713, n_98, n_1710);
  nand g145 (n_1715, n_1711, n_1712, n_1713);
  xor g146 (n_1714, n_50, n_98);
  xor g147 (Z[23], n_1710, n_1714);
  nand g148 (n_1716, n_49, n_97);
  nand g149 (n_1717, n_49, n_1715);
  nand g150 (n_1718, n_97, n_1715);
  nand g151 (n_1720, n_1716, n_1717, n_1718);
  xor g152 (n_1719, n_49, n_97);
  xor g153 (Z[24], n_1715, n_1719);
  nand g154 (n_1721, n_48, n_96);
  nand g155 (n_1722, n_48, n_1720);
  nand g156 (n_1723, n_96, n_1720);
  nand g157 (n_1725, n_1721, n_1722, n_1723);
  xor g158 (n_1724, n_48, n_96);
  xor g159 (Z[25], n_1720, n_1724);
  nand g160 (n_1726, n_47, n_95);
  nand g161 (n_1727, n_47, n_1725);
  nand g162 (n_1728, n_95, n_1725);
  nand g163 (n_1730, n_1726, n_1727, n_1728);
  xor g164 (n_1729, n_47, n_95);
  xor g165 (Z[26], n_1725, n_1729);
  nand g166 (n_1731, n_46, n_94);
  nand g167 (n_1732, n_46, n_1730);
  nand g168 (n_1733, n_94, n_1730);
  nand g169 (n_1735, n_1731, n_1732, n_1733);
  xor g170 (n_1734, n_46, n_94);
  xor g171 (Z[27], n_1730, n_1734);
  nand g172 (n_1736, n_45, n_93);
  nand g173 (n_1737, n_45, n_1735);
  nand g174 (n_1738, n_93, n_1735);
  nand g175 (n_1740, n_1736, n_1737, n_1738);
  xor g176 (n_1739, n_45, n_93);
  xor g177 (Z[28], n_1735, n_1739);
  nand g178 (n_1741, n_44, n_92);
  nand g179 (n_1742, n_44, n_1740);
  nand g180 (n_1743, n_92, n_1740);
  nand g181 (n_1745, n_1741, n_1742, n_1743);
  xor g182 (n_1744, n_44, n_92);
  xor g183 (Z[29], n_1740, n_1744);
  nand g184 (n_1746, n_43, n_91);
  nand g185 (n_1747, n_43, n_1745);
  nand g186 (n_1748, n_91, n_1745);
  nand g187 (n_1750, n_1746, n_1747, n_1748);
  xor g188 (n_1749, n_43, n_91);
  xor g189 (Z[30], n_1745, n_1749);
  nand g190 (n_1751, n_42, n_90);
  nand g191 (n_1752, n_42, n_1750);
  nand g192 (n_1753, n_90, n_1750);
  nand g193 (n_1755, n_1751, n_1752, n_1753);
  xor g194 (n_1754, n_42, n_90);
  xor g195 (Z[31], n_1750, n_1754);
  nand g196 (n_1756, n_41, n_89);
  nand g197 (n_1757, n_41, n_1755);
  nand g198 (n_1758, n_89, n_1755);
  nand g199 (n_1760, n_1756, n_1757, n_1758);
  xor g200 (n_1759, n_41, n_89);
  xor g201 (Z[32], n_1755, n_1759);
  nand g202 (n_1761, n_40, n_88);
  nand g203 (n_1762, n_40, n_1760);
  nand g204 (n_1763, n_88, n_1760);
  nand g205 (n_1765, n_1761, n_1762, n_1763);
  xor g206 (n_1764, n_40, n_88);
  xor g207 (Z[33], n_1760, n_1764);
  nand g208 (n_1766, n_39, n_87);
  nand g209 (n_1767, n_39, n_1765);
  nand g210 (n_1768, n_87, n_1765);
  nand g211 (n_1770, n_1766, n_1767, n_1768);
  xor g212 (n_1769, n_39, n_87);
  xor g213 (Z[34], n_1765, n_1769);
  nand g214 (n_1771, n_38, n_86);
  nand g215 (n_1772, n_38, n_1770);
  nand g216 (n_1773, n_86, n_1770);
  nand g217 (n_1775, n_1771, n_1772, n_1773);
  xor g218 (n_1774, n_38, n_86);
  xor g219 (Z[35], n_1770, n_1774);
  nand g220 (n_1776, n_37, n_85);
  nand g221 (n_1777, n_37, n_1775);
  nand g222 (n_1778, n_85, n_1775);
  nand g223 (n_1780, n_1776, n_1777, n_1778);
  xor g224 (n_1779, n_37, n_85);
  xor g225 (Z[36], n_1775, n_1779);
  nand g226 (n_1781, n_36, n_84);
  nand g227 (n_1782, n_36, n_1780);
  nand g228 (n_1783, n_84, n_1780);
  nand g229 (n_1785, n_1781, n_1782, n_1783);
  xor g230 (n_1784, n_36, n_84);
  xor g231 (Z[37], n_1780, n_1784);
  nand g232 (n_1786, n_35, n_83);
  nand g233 (n_1787, n_35, n_1785);
  nand g234 (n_1788, n_83, n_1785);
  nand g235 (n_1790, n_1786, n_1787, n_1788);
  xor g236 (n_1789, n_35, n_83);
  xor g237 (Z[38], n_1785, n_1789);
  nand g238 (n_1791, n_34, n_82);
  nand g239 (n_1792, n_34, n_1790);
  nand g240 (n_1793, n_82, n_1790);
  nand g241 (n_1795, n_1791, n_1792, n_1793);
  xor g242 (n_1794, n_34, n_82);
  xor g243 (Z[39], n_1790, n_1794);
  nand g244 (n_1796, n_33, n_81);
  nand g245 (n_1797, n_33, n_1795);
  nand g246 (n_1798, n_81, n_1795);
  nand g247 (n_1800, n_1796, n_1797, n_1798);
  xor g248 (n_1799, n_33, n_81);
  xor g249 (Z[40], n_1795, n_1799);
  nand g250 (n_1801, n_32, n_80);
  nand g251 (n_1802, n_32, n_1800);
  nand g252 (n_1803, n_80, n_1800);
  nand g253 (n_1805, n_1801, n_1802, n_1803);
  xor g254 (n_1804, n_32, n_80);
  xor g255 (Z[41], n_1800, n_1804);
  nand g256 (n_1806, n_31, n_79);
  nand g257 (n_1807, n_31, n_1805);
  nand g258 (n_1808, n_79, n_1805);
  nand g259 (n_1810, n_1806, n_1807, n_1808);
  xor g260 (n_1809, n_31, n_79);
  xor g261 (Z[42], n_1805, n_1809);
  nand g262 (n_1811, n_30, n_78);
  nand g263 (n_1812, n_30, n_1810);
  nand g264 (n_1813, n_78, n_1810);
  nand g265 (n_1815, n_1811, n_1812, n_1813);
  xor g266 (n_1814, n_30, n_78);
  xor g267 (Z[43], n_1810, n_1814);
  nand g1772 (n_1816, n_29, n_77);
  nand g1773 (n_1817, n_29, n_1815);
  nand g1774 (n_1818, n_77, n_1815);
  nand g1775 (n_1820, n_1816, n_1817, n_1818);
  xor g1776 (n_1819, n_29, n_77);
  xor g1777 (Z[44], n_1815, n_1819);
  nand g1778 (n_1821, n_28, n_76);
  nand g1779 (n_1822, n_28, n_1820);
  nand g1780 (n_1823, n_76, n_1820);
  nand g1781 (n_1825, n_1821, n_1822, n_1823);
  xor g1782 (n_1824, n_28, n_76);
  xor g1783 (Z[45], n_1820, n_1824);
  nand g1784 (n_1826, n_27, n_75);
  nand g1785 (n_1827, n_27, n_1825);
  nand g1786 (n_1828, n_75, n_1825);
  nand g1787 (n_1830, n_1826, n_1827, n_1828);
  xor g1788 (n_1829, n_27, n_75);
  xor g1789 (Z[46], n_1825, n_1829);
  xor g1791 (Z[47], n_1830, n_1831);
  or g1804 (n_1043, A[1], wc);
  not gc (wc, n_171);
  or g1805 (n_1044, A[1], wc0);
  not gc0 (wc0, A[2]);
  xnor g1807 (n_1166, A[24], A[23]);
  or g1808 (n_1167, wc1, A[24]);
  not gc1 (wc1, A[23]);
  xnor g1809 (n_1214, A[6], A[5]);
  or g1810 (n_1215, A[5], wc2);
  not gc2 (wc2, A[6]);
  or g1811 (n_1252, A[6], wc3);
  not gc3 (wc3, A[7]);
  or g1812 (n_1253, wc4, A[6]);
  not gc4 (wc4, A[5]);
  or g1814 (n_1355, A[9], wc5);
  not gc5 (wc5, A[10]);
  or g1815 (n_1384, A[10], wc6);
  not gc6 (wc6, A[11]);
  or g1816 (n_1385, wc7, A[10]);
  not gc7 (wc7, A[9]);
  or g1818 (n_1463, A[13], wc8);
  not gc8 (wc8, A[14]);
  or g1819 (n_1484, A[14], wc9);
  not gc9 (wc9, A[15]);
  or g1820 (n_1485, wc10, A[14]);
  not gc10 (wc10, A[13]);
  xnor g1821 (n_1530, A[24], A[21]);
  or g1822 (n_1531, wc11, A[24]);
  not gc11 (wc11, A[21]);
  or g1824 (n_1539, A[17], wc12);
  not gc12 (wc12, A[18]);
  or g1825 (n_1552, A[18], wc13);
  not gc13 (wc13, A[19]);
  or g1826 (n_1553, wc14, A[18]);
  not gc14 (wc14, A[17]);
  or g1828 (n_1583, A[21], wc15);
  not gc15 (wc15, A[22]);
  or g1829 (n_1587, wc16, A[22]);
  not gc16 (wc16, A[21]);
  or g1830 (n_1588, A[22], wc17);
  not gc17 (wc17, A[23]);
  or g1831 (n_1593, wc18, A[24]);
  not gc18 (wc18, A[22]);
  xnor g1833 (n_1086, A[2], A[1]);
  or g1834 (n_1088, A[1], wc19);
  not gc19 (wc19, A[3]);
  xnor g1835 (n_453, n_1250, A[6]);
  xnor g1836 (n_519, n_1382, A[10]);
  xnor g1837 (n_570, n_1482, A[14]);
  xnor g1838 (n_603, n_1550, A[18]);
  xnor g1839 (n_28, n_1542, A[23]);
  or g1841 (n_1047, wc20, n_117);
  not gc20 (wc20, A[5]);
  or g1842 (n_1049, wc21, n_117);
  not gc21 (wc21, A[6]);
  xnor g1844 (n_1578, n_613, A[24]);
  or g1845 (n_1579, A[24], wc22);
  not gc22 (wc22, n_613);
  xnor g1846 (n_1831, n_74, A[24]);
  or g1848 (n_1051, n_180, wc23);
  not gc23 (wc23, n_179);
  or g1849 (n_1052, wc24, n_180);
  not gc24 (wc24, A[9]);
  xnor g1850 (n_504, n_1218, n_503);
  or g1851 (n_1356, A[9], wc25);
  not gc25 (wc25, n_503);
  xnor g1852 (n_558, n_1358, n_557);
  or g1853 (n_1464, A[13], wc26);
  not gc26 (wc26, n_557);
  xnor g1854 (n_596, n_1466, n_595);
  or g1855 (n_1540, A[17], wc27);
  not gc27 (wc27, n_595);
  or g1856 (n_1573, A[24], wc28);
  not gc28 (wc28, n_611);
  or g1857 (n_1581, A[24], wc29);
  not gc29 (wc29, n_614);
  xnor g1858 (n_29, n_1542, n_617);
  or g1859 (n_1584, A[21], wc30);
  not gc30 (wc30, n_617);
  or g1862 (n_1216, A[5], wc31);
  not gc31 (wc31, n_433);
  or g1863 (n_1612, n_1606, wc32);
  not gc32 (wc32, n_68);
  or g1864 (n_1613, wc33, n_1606);
  not gc33 (wc33, A[3]);
  xnor g1865 (Z[3], n_1606, n_1614);
  or g1867 (n_1056, wc34, n_202);
  not gc34 (wc34, A[10]);
  or g1868 (n_1057, wc35, n_202);
  not gc35 (wc35, n_282);
  or g1869 (n_1060, wc36, n_285);
  not gc36 (wc36, A[13]);
  xnor g1870 (n_1570, n_610, A[24]);
  or g1871 (n_1571, A[24], wc37);
  not gc37 (wc37, n_610);
  or g1872 (n_1061, wc38, n_285);
  not gc38 (wc38, n_354);
  xnor g1873 (n_357, n_285, n_1058);
  or g1874 (n_1532, A[24], wc39);
  not gc39 (wc39, n_589);
  xnor g1875 (n_1454, n_550, A[24]);
  or g1876 (n_1455, A[24], wc40);
  not gc40 (wc40, n_550);
  xnor g1877 (n_1518, n_584, A[24]);
  or g1878 (n_1519, A[24], wc41);
  not gc41 (wc41, n_584);
  or g1879 (n_1521, A[24], wc42);
  not gc42 (wc42, n_585);
  or g1880 (n_1456, A[24], wc43);
  not gc43 (wc43, n_551);
  xnor g1881 (n_1078, n_363, A[24]);
  or g1882 (n_1079, A[24], wc44);
  not gc44 (wc44, n_363);
  or g1883 (n_1080, A[24], wc45);
  not gc45 (wc45, n_364);
  xnor g1884 (n_1206, n_426, A[24]);
  or g1885 (n_1207, A[24], wc46);
  not gc46 (wc46, n_426);
  xnor g1886 (n_1346, n_496, A[24]);
  or g1887 (n_1347, A[24], wc47);
  not gc47 (wc47, n_496);
  or g1888 (n_1169, A[24], wc48);
  not gc48 (wc48, n_408);
  or g1889 (n_1348, A[24], wc49);
  not gc49 (wc49, n_497);
  or g1890 (n_1432, A[24], wc50);
  not gc50 (wc50, n_540);
  or g1891 (n_1209, A[24], wc51);
  not gc51 (wc51, n_427);
  or g1892 (n_1316, A[24], wc52);
  not gc52 (wc52, n_482);
endmodule

module mult_signed_const_4686_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_4686_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_4953_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74;
  wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_82;
  wire n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90;
  wire n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_119, n_171, n_172, n_173, n_179;
  wire n_180, n_183, n_184, n_187, n_188, n_189, n_193, n_195;
  wire n_196, n_200, n_201, n_202, n_203, n_204, n_207, n_208;
  wire n_209, n_210, n_211, n_212, n_215, n_217, n_218, n_219;
  wire n_220, n_221, n_222, n_223, n_224, n_225, n_226, n_233;
  wire n_235, n_236, n_237, n_238, n_246, n_247, n_248, n_249;
  wire n_250, n_257, n_258, n_259, n_260, n_261, n_262, n_265;
  wire n_267, n_269, n_270, n_271, n_272, n_273, n_274, n_275;
  wire n_276, n_277, n_282, n_283, n_284, n_285, n_286, n_287;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_298, n_299;
  wire n_300, n_301, n_302, n_303, n_304, n_305, n_306, n_307;
  wire n_308, n_309, n_314, n_315, n_316, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_332;
  wire n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_349, n_351, n_353, n_355;
  wire n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_366, n_367, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477;
  wire n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485;
  wire n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539;
  wire n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_595;
  wire n_596, n_597, n_598, n_599, n_603, n_604, n_605, n_606;
  wire n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_617;
  wire n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629;
  wire n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637;
  wire n_638, n_639, n_640, n_641, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_658, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_668, n_669, n_670, n_671;
  wire n_672, n_673, n_674, n_675, n_676, n_677, n_684, n_685;
  wire n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693;
  wire n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_711, n_712, n_713, n_718, n_722;
  wire n_723, n_724, n_725, n_726, n_727, n_728, n_729, n_730;
  wire n_731, n_732, n_733, n_736, n_737, n_738, n_739, n_740;
  wire n_741, n_742, n_743, n_744, n_745, n_746, n_747, n_748;
  wire n_749, n_750, n_751, n_752, n_753, n_762, n_763, n_764;
  wire n_766, n_767, n_768, n_769, n_770, n_771, n_772, n_773;
  wire n_774, n_775, n_776, n_777, n_794, n_795, n_796, n_797;
  wire n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805;
  wire n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827;
  wire n_828, n_829, n_830, n_831, n_832, n_833, n_842, n_843;
  wire n_844, n_848, n_849, n_850, n_851, n_852, n_853, n_854;
  wire n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862;
  wire n_866, n_867, n_868, n_872, n_873, n_874, n_875, n_876;
  wire n_877, n_878, n_879, n_880, n_881, n_882, n_883, n_884;
  wire n_885, n_886, n_887, n_888, n_889, n_890, n_891, n_892;
  wire n_893, n_904, n_905, n_906, n_907, n_908, n_909, n_910;
  wire n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918;
  wire n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926;
  wire n_927, n_928, n_929, n_938, n_939, n_941, n_942, n_943;
  wire n_944, n_945, n_946, n_947, n_948, n_949, n_950, n_951;
  wire n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959;
  wire n_960, n_961, n_962, n_963, n_964, n_965, n_972, n_973;
  wire n_974, n_976, n_977, n_978, n_979, n_980, n_981, n_982;
  wire n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990;
  wire n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998;
  wire n_999, n_1000, n_1001, n_1014, n_1015, n_1016, n_1017, n_1018;
  wire n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026;
  wire n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034;
  wire n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042;
  wire n_1044, n_1045, n_1046, n_1047, n_1048, n_1050, n_1051, n_1052;
  wire n_1056, n_1057, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065;
  wire n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073;
  wire n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081;
  wire n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089;
  wire n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097;
  wire n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105;
  wire n_1106, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114;
  wire n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122;
  wire n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1132;
  wire n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140;
  wire n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148;
  wire n_1149, n_1150, n_1151, n_1152, n_1154, n_1155, n_1156, n_1157;
  wire n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165;
  wire n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173;
  wire n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181;
  wire n_1182, n_1183, n_1184, n_1185, n_1186, n_1188, n_1189, n_1190;
  wire n_1191, n_1192, n_1193, n_1194, n_1196, n_1197, n_1198, n_1199;
  wire n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207;
  wire n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215;
  wire n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223;
  wire n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1241;
  wire n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249;
  wire n_1250, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258;
  wire n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1266, n_1267;
  wire n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275;
  wire n_1276, n_1277, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285;
  wire n_1288, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296;
  wire n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304;
  wire n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312;
  wire n_1313, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322;
  wire n_1324, n_1325, n_1326, n_1327, n_1328, n_1330, n_1331, n_1332;
  wire n_1333, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342;
  wire n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350;
  wire n_1351, n_1352, n_1353, n_1355, n_1356, n_1357, n_1358, n_1359;
  wire n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367;
  wire n_1368, n_1369, n_1370, n_1371, n_1373, n_1374, n_1375, n_1376;
  wire n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384;
  wire n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392;
  wire n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400;
  wire n_1401, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1412;
  wire n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420;
  wire n_1421, n_1422, n_1423, n_1424, n_1426, n_1427, n_1428, n_1429;
  wire n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1440, n_1441;
  wire n_1442, n_1443, n_1444, n_1446, n_1447, n_1448, n_1449, n_1452;
  wire n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460;
  wire n_1461, n_1463, n_1464, n_1465, n_1466, n_1468, n_1469, n_1470;
  wire n_1471, n_1472, n_1473, n_1474, n_1476, n_1477, n_1478, n_1479;
  wire n_1480, n_1481, n_1484, n_1486, n_1487, n_1488, n_1489, n_1490;
  wire n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1498, n_1499;
  wire n_1500, n_1501, n_1502, n_1504, n_1506, n_1507, n_1508, n_1509;
  wire n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517;
  wire n_1518, n_1519, n_1520, n_1521, n_1524, n_1525, n_1526, n_1527;
  wire n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535;
  wire n_1536, n_1537, n_1539, n_1540, n_1541, n_1544, n_1545, n_1546;
  wire n_1547, n_1548, n_1549, n_1550, n_1552, n_1553, n_1554, n_1555;
  wire n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1566;
  wire n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1576;
  wire n_1577, n_1578, n_1579, n_1580, n_1581, n_1583, n_1584, n_1585;
  wire n_1587, n_1588, n_1589, n_1593, n_1606, n_1611, n_1612, n_1613;
  wire n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621;
  wire n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629;
  wire n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637;
  wire n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645;
  wire n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653;
  wire n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661;
  wire n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669;
  wire n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677;
  wire n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685;
  wire n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693;
  wire n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701;
  wire n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709;
  wire n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717;
  wire n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725;
  wire n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733;
  wire n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741;
  wire n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749;
  wire n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757;
  wire n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765;
  wire n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773;
  wire n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781;
  wire n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789;
  wire n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797;
  wire n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805;
  wire n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813;
  wire n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821;
  wire n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829;
  wire n_1830, n_1831;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], A[2]);
  xor g270 (n_117, n_622, n_171);
  nand g3 (n_623, A[1], A[2]);
  nand g271 (n_624, n_171, A[2]);
  nand g272 (n_625, A[1], n_171);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, n_69);
  xor g288 (n_70, n_634, A[4]);
  nand g289 (n_635, n_68, n_69);
  nand g290 (n_636, A[4], n_69);
  nand g291 (n_637, n_68, A[4]);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_70);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_70);
  nand g296 (n_640, A[7], n_70);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g305 (n_646, A[5], n_117);
  xor g306 (n_180, n_646, A[6]);
  nand g307 (n_647, A[5], n_117);
  nand g308 (n_648, A[6], n_117);
  nand g309 (n_649, A[5], A[6]);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, n_179, n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, n_179, n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, n_179, A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_187, n_659, n_660, n_661);
  xor g329 (n_662, n_183, A[9]);
  xor g330 (n_112, n_662, n_184);
  nand g331 (n_663, n_183, A[9]);
  nand g332 (n_664, n_184, A[9]);
  nand g333 (n_665, n_183, n_184);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_188, n_630, A[7]);
  nand g340 (n_668, A[7], n_173);
  nand g341 (n_669, A[4], A[7]);
  nand g342 (n_193, n_631, n_668, n_669);
  xor g343 (n_670, n_67, A[8]);
  xor g344 (n_189, n_670, n_187);
  nand g345 (n_671, n_67, A[8]);
  nand g346 (n_672, n_187, A[8]);
  nand g347 (n_673, n_67, n_187);
  nand g348 (n_195, n_671, n_672, n_673);
  xor g349 (n_674, n_188, A[10]);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, n_188, A[10]);
  nand g352 (n_676, n_189, A[10]);
  nand g353 (n_677, n_188, n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_72, n_638, A[8]);
  nand g366 (n_684, A[8], n_70);
  nand g367 (n_685, A[5], A[8]);
  nand g368 (n_201, n_639, n_684, n_685);
  xor g369 (n_686, n_193, A[9]);
  xor g370 (n_196, n_686, n_72);
  nand g371 (n_687, n_193, A[9]);
  nand g372 (n_688, n_72, A[9]);
  nand g373 (n_689, n_193, n_72);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, n_195, A[11]);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, n_195, A[11]);
  nand g378 (n_692, n_196, A[11]);
  nand g379 (n_693, n_195, n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g388 (n_200, n_646, n_179);
  nand g390 (n_700, n_179, n_117);
  nand g391 (n_701, A[5], n_179);
  nand g392 (n_207, n_647, n_700, n_701);
  xor g393 (n_702, A[6], n_200);
  xor g394 (n_202, n_702, A[9]);
  nand g395 (n_703, A[6], n_200);
  nand g396 (n_704, A[9], n_200);
  nand g397 (n_705, A[6], A[9]);
  nand g398 (n_209, n_703, n_704, n_705);
  xor g399 (n_706, A[10], n_201);
  xor g400 (n_204, n_706, n_202);
  nand g401 (n_707, A[10], n_201);
  nand g402 (n_708, n_202, n_201);
  nand g403 (n_709, A[10], n_202);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, A[12], n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, A[12], n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, A[12], n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g417 (n_718, A[6], A[7]);
  xor g418 (n_208, n_718, n_116);
  xor g423 (n_722, n_207, A[10]);
  xor g424 (n_210, n_722, n_208);
  nand g425 (n_723, n_207, A[10]);
  nand g426 (n_724, n_208, A[10]);
  nand g427 (n_725, n_207, n_208);
  nand g428 (n_218, n_723, n_724, n_725);
  xor g429 (n_726, A[11], n_209);
  xor g430 (n_212, n_726, A[13]);
  nand g431 (n_727, A[11], n_209);
  nand g432 (n_728, A[13], n_209);
  nand g433 (n_729, A[11], A[13]);
  nand g434 (n_220, n_727, n_728, n_729);
  xor g435 (n_730, n_210, n_211);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, n_210, n_211);
  nand g438 (n_732, n_212, n_211);
  nand g439 (n_733, n_210, n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g444 (n_215, n_630, n_67);
  nand g446 (n_736, n_67, n_173);
  nand g447 (n_737, A[4], n_67);
  nand g448 (n_71, n_631, n_736, n_737);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_217, n_738, n_215);
  nand g451 (n_739, A[7], A[8]);
  nand g452 (n_740, n_215, A[8]);
  nand g453 (n_741, A[7], n_215);
  nand g454 (n_73, n_739, n_740, n_741);
  xor g455 (n_742, n_187, n_217);
  xor g456 (n_219, n_742, A[11]);
  nand g457 (n_743, n_187, n_217);
  nand g458 (n_744, A[11], n_217);
  nand g459 (n_745, n_187, A[11]);
  nand g460 (n_223, n_743, n_744, n_745);
  xor g461 (n_746, n_218, A[12]);
  xor g462 (n_221, n_746, A[14]);
  nand g463 (n_747, n_218, A[12]);
  nand g464 (n_748, A[14], A[12]);
  nand g465 (n_749, n_218, A[14]);
  nand g466 (n_225, n_747, n_748, n_749);
  xor g467 (n_750, n_219, n_220);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, n_219, n_220);
  nand g470 (n_752, n_221, n_220);
  nand g471 (n_753, n_219, n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g487 (n_762, A[9], n_71);
  xor g488 (n_222, n_762, n_72);
  nand g489 (n_763, A[9], n_71);
  nand g490 (n_764, n_72, n_71);
  nand g492 (n_233, n_763, n_764, n_688);
  xor g493 (n_766, n_73, A[12]);
  xor g494 (n_224, n_766, n_222);
  nand g495 (n_767, n_73, A[12]);
  nand g496 (n_768, n_222, A[12]);
  nand g497 (n_769, n_73, n_222);
  nand g498 (n_235, n_767, n_768, n_769);
  xor g499 (n_770, A[13], n_223);
  xor g500 (n_226, n_770, A[15]);
  nand g501 (n_771, A[13], n_223);
  nand g502 (n_772, A[15], n_223);
  nand g503 (n_773, A[13], A[15]);
  nand g504 (n_237, n_771, n_772, n_773);
  xor g505 (n_774, n_224, n_225);
  xor g506 (n_106, n_774, n_226);
  nand g507 (n_775, n_224, n_225);
  nand g508 (n_776, n_226, n_225);
  nand g509 (n_777, n_224, n_226);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g535 (n_794, n_233, A[13]);
  xor g536 (n_236, n_794, n_204);
  nand g537 (n_795, n_233, A[13]);
  nand g538 (n_796, n_204, A[13]);
  nand g539 (n_797, n_233, n_204);
  nand g540 (n_247, n_795, n_796, n_797);
  xor g541 (n_798, A[14], n_235);
  xor g542 (n_238, n_798, n_236);
  nand g543 (n_799, A[14], n_235);
  nand g544 (n_800, n_236, n_235);
  nand g545 (n_801, A[14], n_236);
  nand g546 (n_249, n_799, n_800, n_801);
  xor g547 (n_802, A[16], n_237);
  xor g548 (n_105, n_802, n_238);
  nand g549 (n_803, A[16], n_237);
  nand g550 (n_804, n_238, n_237);
  nand g551 (n_805, A[16], n_238);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g572 (n_246, n_726, n_210);
  nand g574 (n_820, n_210, n_209);
  nand g575 (n_821, A[11], n_210);
  nand g576 (n_258, n_727, n_820, n_821);
  xor g577 (n_822, n_211, A[14]);
  xor g578 (n_248, n_822, n_246);
  nand g579 (n_823, n_211, A[14]);
  nand g580 (n_824, n_246, A[14]);
  nand g581 (n_825, n_211, n_246);
  nand g582 (n_260, n_823, n_824, n_825);
  xor g583 (n_826, A[15], n_247);
  xor g584 (n_250, n_826, A[17]);
  nand g585 (n_827, A[15], n_247);
  nand g586 (n_828, A[17], n_247);
  nand g587 (n_829, A[15], A[17]);
  nand g588 (n_262, n_827, n_828, n_829);
  xor g589 (n_830, n_248, n_249);
  xor g590 (n_104, n_830, n_250);
  nand g591 (n_831, n_248, n_249);
  nand g592 (n_832, n_250, n_249);
  nand g593 (n_833, n_248, n_250);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g609 (n_842, n_188, A[11]);
  xor g610 (n_257, n_842, n_189);
  nand g611 (n_843, n_188, A[11]);
  nand g612 (n_844, n_189, A[11]);
  nand g614 (n_270, n_843, n_844, n_677);
  xor g616 (n_259, n_746, n_257);
  nand g618 (n_848, n_257, n_218);
  nand g619 (n_849, A[12], n_257);
  nand g620 (n_272, n_747, n_848, n_849);
  xor g621 (n_850, n_258, A[15]);
  xor g622 (n_261, n_850, n_259);
  nand g623 (n_851, n_258, A[15]);
  nand g624 (n_852, n_259, A[15]);
  nand g625 (n_853, n_258, n_259);
  nand g626 (n_274, n_851, n_852, n_853);
  xor g627 (n_854, A[16], n_260);
  xor g628 (n_119, n_854, A[18]);
  nand g629 (n_855, A[16], n_260);
  nand g630 (n_856, A[18], n_260);
  nand g631 (n_857, A[16], A[18]);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_261, n_262);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_261, n_262);
  nand g636 (n_860, n_119, n_262);
  nand g637 (n_861, n_261, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g641 (n_862, n_68, A[4]);
  xor g642 (n_265, n_862, n_69);
  xor g647 (n_866, A[5], n_265);
  xor g648 (n_267, n_866, A[8]);
  nand g649 (n_867, A[5], n_265);
  nand g650 (n_868, A[8], n_265);
  nand g652 (n_282, n_867, n_868, n_685);
  xor g654 (n_269, n_686, n_267);
  nand g656 (n_872, n_267, n_193);
  nand g657 (n_873, A[9], n_267);
  nand g658 (n_284, n_687, n_872, n_873);
  xor g659 (n_874, n_195, A[12]);
  xor g660 (n_271, n_874, A[13]);
  nand g661 (n_875, n_195, A[12]);
  nand g662 (n_876, A[13], A[12]);
  nand g663 (n_877, n_195, A[13]);
  nand g664 (n_286, n_875, n_876, n_877);
  xor g665 (n_878, n_269, n_270);
  xor g666 (n_273, n_878, n_271);
  nand g667 (n_879, n_269, n_270);
  nand g668 (n_880, n_271, n_270);
  nand g669 (n_881, n_269, n_271);
  nand g670 (n_288, n_879, n_880, n_881);
  xor g671 (n_882, n_272, A[16]);
  xor g672 (n_275, n_882, n_273);
  nand g673 (n_883, n_272, A[16]);
  nand g674 (n_884, n_273, A[16]);
  nand g675 (n_885, n_272, n_273);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, A[17], n_274);
  xor g678 (n_277, n_886, A[19]);
  nand g679 (n_887, A[17], n_274);
  nand g680 (n_888, A[19], n_274);
  nand g681 (n_889, A[17], A[19]);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g702 (n_283, n_650, A[9]);
  nand g704 (n_904, A[9], n_180);
  nand g705 (n_905, n_179, A[9]);
  nand g706 (n_298, n_651, n_904, n_905);
  xor g707 (n_906, A[10], n_282);
  xor g708 (n_285, n_906, n_283);
  nand g709 (n_907, A[10], n_282);
  nand g710 (n_908, n_283, n_282);
  nand g711 (n_909, A[10], n_283);
  nand g712 (n_300, n_907, n_908, n_909);
  xor g713 (n_910, n_284, A[13]);
  xor g714 (n_287, n_910, n_285);
  nand g715 (n_911, n_284, A[13]);
  nand g716 (n_912, n_285, A[13]);
  nand g717 (n_913, n_284, n_285);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, A[14], n_286);
  xor g720 (n_289, n_914, n_287);
  nand g721 (n_915, A[14], n_286);
  nand g722 (n_916, n_287, n_286);
  nand g723 (n_917, A[14], n_287);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, n_288, A[17]);
  xor g726 (n_291, n_918, n_289);
  nand g727 (n_919, n_288, A[17]);
  nand g728 (n_920, n_289, A[17]);
  nand g729 (n_921, n_288, n_289);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, A[18], n_290);
  xor g732 (n_293, n_922, A[20]);
  nand g733 (n_923, A[18], n_290);
  nand g734 (n_924, A[20], n_290);
  nand g735 (n_925, A[18], A[20]);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g755 (n_938, n_183, A[10]);
  xor g756 (n_299, n_938, n_208);
  nand g757 (n_939, n_183, A[10]);
  nand g759 (n_941, n_183, n_208);
  nand g760 (n_315, n_939, n_724, n_941);
  xor g761 (n_942, A[11], n_298);
  xor g762 (n_301, n_942, n_299);
  nand g763 (n_943, A[11], n_298);
  nand g764 (n_944, n_299, n_298);
  nand g765 (n_945, A[11], n_299);
  nand g766 (n_317, n_943, n_944, n_945);
  xor g767 (n_946, n_300, A[14]);
  xor g768 (n_303, n_946, A[15]);
  nand g769 (n_947, n_300, A[14]);
  nand g770 (n_948, A[15], A[14]);
  nand g771 (n_949, n_300, A[15]);
  nand g772 (n_319, n_947, n_948, n_949);
  xor g773 (n_950, n_301, n_302);
  xor g774 (n_305, n_950, n_303);
  nand g775 (n_951, n_301, n_302);
  nand g776 (n_952, n_303, n_302);
  nand g777 (n_953, n_301, n_303);
  nand g778 (n_321, n_951, n_952, n_953);
  xor g779 (n_954, n_304, A[18]);
  xor g780 (n_307, n_954, n_305);
  nand g781 (n_955, n_304, A[18]);
  nand g782 (n_956, n_305, A[18]);
  nand g783 (n_957, n_304, n_305);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, A[19], n_306);
  xor g786 (n_309, n_958, A[21]);
  nand g787 (n_959, A[19], n_306);
  nand g788 (n_960, A[21], n_306);
  nand g789 (n_961, A[19], A[21]);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g806 (n_314, n_670, n_188);
  nand g808 (n_972, n_188, A[8]);
  nand g809 (n_973, n_67, n_188);
  nand g810 (n_332, n_671, n_972, n_973);
  xor g811 (n_974, n_187, A[11]);
  xor g812 (n_316, n_974, n_314);
  nand g814 (n_976, n_314, A[11]);
  nand g815 (n_977, n_187, n_314);
  nand g816 (n_334, n_745, n_976, n_977);
  xor g817 (n_978, A[12], n_315);
  xor g818 (n_318, n_978, n_316);
  nand g819 (n_979, A[12], n_315);
  nand g820 (n_980, n_316, n_315);
  nand g821 (n_981, A[12], n_316);
  nand g822 (n_336, n_979, n_980, n_981);
  xor g823 (n_982, n_317, A[15]);
  xor g824 (n_320, n_982, A[16]);
  nand g825 (n_983, n_317, A[15]);
  nand g826 (n_984, A[16], A[15]);
  nand g827 (n_985, n_317, A[16]);
  nand g828 (n_338, n_983, n_984, n_985);
  xor g829 (n_986, n_318, n_319);
  xor g830 (n_322, n_986, n_320);
  nand g831 (n_987, n_318, n_319);
  nand g832 (n_988, n_320, n_319);
  nand g833 (n_989, n_318, n_320);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, n_321, A[19]);
  xor g836 (n_324, n_990, A[20]);
  nand g837 (n_991, n_321, A[19]);
  nand g838 (n_992, A[20], A[19]);
  nand g839 (n_993, n_321, A[20]);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, n_322, n_323);
  xor g842 (n_326, n_994, A[22]);
  nand g843 (n_995, n_322, n_323);
  nand g844 (n_996, A[22], n_323);
  nand g845 (n_997, n_322, A[22]);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, n_324, n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, n_324, n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, n_324, n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g873 (n_1014, n_332, A[12]);
  xor g874 (n_335, n_1014, n_269);
  nand g875 (n_1015, n_332, A[12]);
  nand g876 (n_1016, n_269, A[12]);
  nand g877 (n_1017, n_332, n_269);
  nand g878 (n_356, n_1015, n_1016, n_1017);
  xor g879 (n_1018, A[13], n_334);
  xor g880 (n_337, n_1018, n_335);
  nand g881 (n_1019, A[13], n_334);
  nand g882 (n_1020, n_335, n_334);
  nand g883 (n_1021, A[13], n_335);
  nand g884 (n_358, n_1019, n_1020, n_1021);
  xor g885 (n_1022, A[16], n_336);
  xor g886 (n_339, n_1022, A[17]);
  nand g887 (n_1023, A[16], n_336);
  nand g888 (n_1024, A[17], n_336);
  nand g889 (n_1025, A[16], A[17]);
  nand g890 (n_360, n_1023, n_1024, n_1025);
  xor g891 (n_1026, n_337, n_338);
  xor g892 (n_341, n_1026, n_339);
  nand g893 (n_1027, n_337, n_338);
  nand g894 (n_1028, n_339, n_338);
  nand g895 (n_1029, n_337, n_339);
  nand g896 (n_362, n_1027, n_1028, n_1029);
  xor g897 (n_1030, A[20], n_340);
  xor g898 (n_343, n_1030, n_341);
  nand g899 (n_1031, A[20], n_340);
  nand g900 (n_1032, n_341, n_340);
  nand g901 (n_1033, A[20], n_341);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, A[21], n_342);
  xor g904 (n_345, n_1034, n_343);
  nand g905 (n_1035, A[21], n_342);
  nand g906 (n_1036, n_343, n_342);
  nand g907 (n_1037, A[21], n_343);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, A[23], n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, A[23], n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, A[23], n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  xor g917 (n_1042, A[2], n_171);
  nand g922 (n_371, n_624, n_1044, n_1045);
  xor g923 (n_1046, A[5], n_349);
  xor g924 (n_351, n_1046, n_179);
  nand g925 (n_1047, A[5], n_349);
  nand g926 (n_1048, n_179, n_349);
  nand g928 (n_373, n_1047, n_1048, n_701);
  xor g929 (n_1050, A[6], n_351);
  xor g930 (n_353, n_1050, A[9]);
  nand g931 (n_1051, A[6], n_351);
  nand g932 (n_1052, A[9], n_351);
  nand g934 (n_375, n_1051, n_1052, n_705);
  xor g936 (n_355, n_906, n_353);
  nand g938 (n_1056, n_353, n_282);
  nand g939 (n_1057, A[10], n_353);
  nand g940 (n_377, n_907, n_1056, n_1057);
  xor g942 (n_357, n_910, n_355);
  nand g944 (n_1060, n_355, A[13]);
  nand g945 (n_1061, n_284, n_355);
  nand g946 (n_379, n_911, n_1060, n_1061);
  xor g947 (n_1062, A[14], n_356);
  xor g948 (n_359, n_1062, n_357);
  nand g949 (n_1063, A[14], n_356);
  nand g950 (n_1064, n_357, n_356);
  nand g951 (n_1065, A[14], n_357);
  nand g952 (n_381, n_1063, n_1064, n_1065);
  xor g953 (n_1066, n_358, A[17]);
  xor g954 (n_361, n_1066, A[18]);
  nand g955 (n_1067, n_358, A[17]);
  nand g956 (n_1068, A[18], A[17]);
  nand g957 (n_1069, n_358, A[18]);
  nand g958 (n_383, n_1067, n_1068, n_1069);
  xor g959 (n_1070, n_359, n_360);
  xor g960 (n_363, n_1070, n_361);
  nand g961 (n_1071, n_359, n_360);
  nand g962 (n_1072, n_361, n_360);
  nand g963 (n_1073, n_359, n_361);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, A[21], n_362);
  xor g966 (n_365, n_1074, A[22]);
  nand g967 (n_1075, A[21], n_362);
  nand g968 (n_1076, A[22], n_362);
  nand g969 (n_1077, A[21], A[22]);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g971 (n_1078, n_363, n_364);
  nand g973 (n_1079, n_363, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  xor g985 (n_1086, A[3], A[1]);
  nand g987 (n_1087, A[3], A[1]);
  nand g990 (n_392, n_1087, n_1088, n_1089);
  xor g991 (n_1090, n_371, n_372);
  xor g992 (n_374, n_1090, A[6]);
  nand g993 (n_1091, n_371, n_372);
  nand g994 (n_1092, A[6], n_372);
  nand g995 (n_1093, n_371, A[6]);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, n_374);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, n_374, n_373);
  nand g1001 (n_1097, A[7], n_374);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, A[10], A[11]);
  xor g1004 (n_378, n_1098, n_375);
  nand g1005 (n_1099, A[10], A[11]);
  nand g1006 (n_1100, n_375, A[11]);
  nand g1007 (n_1101, A[10], n_375);
  nand g1008 (n_398, n_1099, n_1100, n_1101);
  xor g1009 (n_1102, n_376, n_377);
  xor g1010 (n_380, n_1102, n_378);
  nand g1011 (n_1103, n_376, n_377);
  nand g1012 (n_1104, n_378, n_377);
  nand g1013 (n_1105, n_376, n_378);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, A[14], A[15]);
  xor g1016 (n_382, n_1106, n_379);
  nand g1018 (n_1108, n_379, A[15]);
  nand g1019 (n_1109, A[14], n_379);
  nand g1020 (n_402, n_948, n_1108, n_1109);
  xor g1021 (n_1110, n_380, A[18]);
  xor g1022 (n_384, n_1110, n_381);
  nand g1023 (n_1111, n_380, A[18]);
  nand g1024 (n_1112, n_381, A[18]);
  nand g1025 (n_1113, n_380, n_381);
  nand g1026 (n_404, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, n_382, A[19]);
  xor g1028 (n_386, n_1114, n_383);
  nand g1029 (n_1115, n_382, A[19]);
  nand g1030 (n_1116, n_383, A[19]);
  nand g1031 (n_1117, n_382, n_383);
  nand g1032 (n_406, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_384, n_385);
  xor g1034 (n_388, n_1118, n_386);
  nand g1035 (n_1119, n_384, n_385);
  nand g1036 (n_1120, n_386, n_385);
  nand g1037 (n_1121, n_384, n_386);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, A[22], A[23]);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, A[22], A[23]);
  nand g1042 (n_1124, n_387, A[23]);
  nand g1043 (n_1125, A[22], n_387);
  nand g1044 (n_411, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1052 (n_393, n_626, A[4]);
  nand g1054 (n_1132, A[4], A[2]);
  nand g1055 (n_1133, A[3], A[4]);
  nand g1056 (n_412, n_627, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, n_396, A[11]);
  xor g1070 (n_399, n_1142, n_397);
  nand g1071 (n_1143, n_396, A[11]);
  nand g1072 (n_1144, n_397, A[11]);
  nand g1073 (n_1145, n_396, n_397);
  nand g1074 (n_417, n_1143, n_1144, n_1145);
  xor g1075 (n_1146, A[12], n_398);
  xor g1076 (n_401, n_1146, n_399);
  nand g1077 (n_1147, A[12], n_398);
  nand g1078 (n_1148, n_399, n_398);
  nand g1079 (n_1149, A[12], n_399);
  nand g1080 (n_420, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, A[15], n_400);
  xor g1082 (n_403, n_1150, A[16]);
  nand g1083 (n_1151, A[15], n_400);
  nand g1084 (n_1152, A[16], n_400);
  nand g1086 (n_421, n_1151, n_1152, n_984);
  xor g1087 (n_1154, n_401, n_402);
  xor g1088 (n_405, n_1154, A[19]);
  nand g1089 (n_1155, n_401, n_402);
  nand g1090 (n_1156, A[19], n_402);
  nand g1091 (n_1157, n_401, A[19]);
  nand g1092 (n_424, n_1155, n_1156, n_1157);
  xor g1093 (n_1158, n_403, n_404);
  xor g1094 (n_407, n_1158, A[20]);
  nand g1095 (n_1159, n_403, n_404);
  nand g1096 (n_1160, A[20], n_404);
  nand g1097 (n_1161, n_403, A[20]);
  nand g1098 (n_425, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_405, n_406);
  xor g1100 (n_409, n_1162, n_407);
  nand g1101 (n_1163, n_405, n_406);
  nand g1102 (n_1164, n_407, n_406);
  nand g1103 (n_1165, n_405, n_407);
  nand g1104 (n_428, n_1163, n_1164, n_1165);
  xor g1106 (n_410, n_1166, n_408);
  nand g1108 (n_1168, n_408, A[23]);
  nand g1110 (n_430, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1123 (n_1178, A[8], n_413);
  xor g1124 (n_415, n_1178, A[9]);
  nand g1125 (n_1179, A[8], n_413);
  nand g1126 (n_1180, A[9], n_413);
  nand g1127 (n_1181, A[8], A[9]);
  nand g1128 (n_435, n_1179, n_1180, n_1181);
  xor g1129 (n_1182, n_414, n_415);
  xor g1130 (n_418, n_1182, n_416);
  nand g1131 (n_1183, n_414, n_415);
  nand g1132 (n_1184, n_416, n_415);
  nand g1133 (n_1185, n_414, n_416);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, A[12], A[13]);
  xor g1136 (n_419, n_1186, n_417);
  nand g1138 (n_1188, n_417, A[13]);
  nand g1139 (n_1189, A[12], n_417);
  nand g1140 (n_439, n_876, n_1188, n_1189);
  xor g1141 (n_1190, n_418, n_419);
  xor g1142 (n_422, n_1190, n_420);
  nand g1143 (n_1191, n_418, n_419);
  nand g1144 (n_1192, n_420, n_419);
  nand g1145 (n_1193, n_418, n_420);
  nand g1146 (n_441, n_1191, n_1192, n_1193);
  xor g1147 (n_1194, A[16], A[17]);
  xor g1148 (n_423, n_1194, n_421);
  nand g1150 (n_1196, n_421, A[17]);
  nand g1151 (n_1197, A[16], n_421);
  nand g1152 (n_443, n_1025, n_1196, n_1197);
  xor g1153 (n_1198, n_422, A[20]);
  xor g1154 (n_426, n_1198, n_423);
  nand g1155 (n_1199, n_422, A[20]);
  nand g1156 (n_1200, n_423, A[20]);
  nand g1157 (n_1201, n_422, n_423);
  nand g1158 (n_445, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_424, A[21]);
  xor g1160 (n_427, n_1202, n_425);
  nand g1161 (n_1203, n_424, A[21]);
  nand g1162 (n_1204, n_425, A[21]);
  nand g1163 (n_1205, n_424, n_425);
  nand g1164 (n_446, n_1203, n_1204, n_1205);
  xor g1166 (n_429, n_1206, n_427);
  nand g1169 (n_1209, n_426, n_427);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, n_433);
  nand g1183 (n_1217, A[6], n_433);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, A[9], A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, A[9], A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, A[9], n_434);
  nand g1190 (n_456, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, n_435, n_436);
  xor g1192 (n_438, n_1222, A[13]);
  nand g1193 (n_1223, n_435, n_436);
  nand g1194 (n_1224, A[13], n_436);
  nand g1195 (n_1225, n_435, A[13]);
  nand g1196 (n_457, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, n_437, A[14]);
  xor g1198 (n_440, n_1226, n_438);
  nand g1199 (n_1227, n_437, A[14]);
  nand g1200 (n_1228, n_438, A[14]);
  nand g1201 (n_1229, n_437, n_438);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, n_439, A[17]);
  xor g1204 (n_442, n_1230, A[18]);
  nand g1205 (n_1231, n_439, A[17]);
  nand g1207 (n_1233, n_439, A[18]);
  nand g1208 (n_461, n_1231, n_1068, n_1233);
  xor g1209 (n_1234, n_440, n_441);
  xor g1210 (n_444, n_1234, n_442);
  nand g1211 (n_1235, n_440, n_441);
  nand g1212 (n_1236, n_442, n_441);
  nand g1213 (n_1237, n_440, n_442);
  nand g1214 (n_463, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_443, A[21]);
  xor g1216 (n_447, n_1238, A[22]);
  nand g1217 (n_1239, n_443, A[21]);
  nand g1219 (n_1241, n_443, A[22]);
  nand g1220 (n_465, n_1239, n_1077, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[5], A[7]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], n_453);
  xor g1242 (n_455, n_1254, n_454);
  nand g1243 (n_1255, A[10], n_453);
  nand g1244 (n_1256, n_454, n_453);
  nand g1245 (n_1257, A[10], n_454);
  nand g1246 (n_472, n_1255, n_1256, n_1257);
  xor g1247 (n_1258, A[11], n_455);
  xor g1248 (n_458, n_1258, n_456);
  nand g1249 (n_1259, A[11], n_455);
  nand g1250 (n_1260, n_456, n_455);
  nand g1251 (n_1261, A[11], n_456);
  nand g1252 (n_474, n_1259, n_1260, n_1261);
  xor g1253 (n_1262, A[14], n_457);
  xor g1254 (n_460, n_1262, A[15]);
  nand g1255 (n_1263, A[14], n_457);
  nand g1256 (n_1264, A[15], n_457);
  nand g1258 (n_476, n_1263, n_1264, n_948);
  xor g1259 (n_1266, n_458, A[18]);
  xor g1260 (n_462, n_1266, n_459);
  nand g1261 (n_1267, n_458, A[18]);
  nand g1262 (n_1268, n_459, A[18]);
  nand g1263 (n_1269, n_458, n_459);
  nand g1264 (n_479, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, n_460, A[19]);
  xor g1266 (n_464, n_1270, n_461);
  nand g1267 (n_1271, n_460, A[19]);
  nand g1268 (n_1272, n_461, A[19]);
  nand g1269 (n_1273, n_460, n_461);
  nand g1270 (n_480, n_1271, n_1272, n_1273);
  xor g1271 (n_1274, n_462, n_463);
  xor g1272 (n_466, n_1274, n_464);
  nand g1273 (n_1275, n_462, n_463);
  nand g1274 (n_1276, n_464, n_463);
  nand g1275 (n_1277, n_462, n_464);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1278 (n_467, n_1122, n_465);
  nand g1280 (n_1280, n_465, A[23]);
  nand g1281 (n_1281, A[22], n_465);
  nand g1282 (n_485, n_1123, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1290 (n_471, n_718, A[8]);
  nand g1292 (n_1288, A[8], A[6]);
  nand g1294 (n_486, n_661, n_1288, n_739);
  xor g1295 (n_1290, n_470, n_471);
  xor g1296 (n_473, n_1290, A[11]);
  nand g1297 (n_1291, n_470, n_471);
  nand g1298 (n_1292, A[11], n_471);
  nand g1299 (n_1293, n_470, A[11]);
  nand g1300 (n_488, n_1291, n_1292, n_1293);
  xor g1301 (n_1294, A[12], n_472);
  xor g1302 (n_475, n_1294, n_473);
  nand g1303 (n_1295, A[12], n_472);
  nand g1304 (n_1296, n_473, n_472);
  nand g1305 (n_1297, A[12], n_473);
  nand g1306 (n_489, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, A[15], n_474);
  xor g1308 (n_477, n_1298, n_475);
  nand g1309 (n_1299, A[15], n_474);
  nand g1310 (n_1300, n_475, n_474);
  nand g1311 (n_1301, A[15], n_475);
  nand g1312 (n_491, n_1299, n_1300, n_1301);
  xor g1313 (n_1302, A[16], n_476);
  xor g1314 (n_478, n_1302, n_477);
  nand g1315 (n_1303, A[16], n_476);
  nand g1316 (n_1304, n_477, n_476);
  nand g1317 (n_1305, A[16], n_477);
  nand g1318 (n_494, n_1303, n_1304, n_1305);
  xor g1319 (n_1306, A[19], n_478);
  xor g1320 (n_481, n_1306, n_479);
  nand g1321 (n_1307, A[19], n_478);
  nand g1322 (n_1308, n_479, n_478);
  nand g1323 (n_1309, A[19], n_479);
  nand g1324 (n_495, n_1307, n_1308, n_1309);
  xor g1325 (n_1310, A[20], n_480);
  xor g1326 (n_483, n_1310, n_481);
  nand g1327 (n_1311, A[20], n_480);
  nand g1328 (n_1312, n_481, n_480);
  nand g1329 (n_1313, A[20], n_481);
  nand g1330 (n_498, n_1311, n_1312, n_1313);
  xor g1332 (n_484, n_1166, n_482);
  nand g1335 (n_1317, A[23], n_482);
  nand g1336 (n_500, n_1167, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1343 (n_1322, A[8], A[9]);
  xor g1344 (n_487, n_1322, n_486);
  nand g1346 (n_1324, n_486, A[9]);
  nand g1347 (n_1325, A[8], n_486);
  nand g1348 (n_503, n_1181, n_1324, n_1325);
  xor g1349 (n_1326, A[12], n_487);
  xor g1350 (n_490, n_1326, A[13]);
  nand g1351 (n_1327, A[12], n_487);
  nand g1352 (n_1328, A[13], n_487);
  nand g1354 (n_504, n_1327, n_1328, n_876);
  xor g1355 (n_1330, n_488, n_489);
  xor g1356 (n_492, n_1330, n_490);
  nand g1357 (n_1331, n_488, n_489);
  nand g1358 (n_1332, n_490, n_489);
  nand g1359 (n_1333, n_488, n_490);
  nand g1360 (n_507, n_1331, n_1332, n_1333);
  xor g1362 (n_493, n_1194, n_491);
  nand g1364 (n_1336, n_491, A[17]);
  nand g1365 (n_1337, A[16], n_491);
  nand g1366 (n_508, n_1025, n_1336, n_1337);
  xor g1367 (n_1338, n_492, n_493);
  xor g1368 (n_496, n_1338, n_494);
  nand g1369 (n_1339, n_492, n_493);
  nand g1370 (n_1340, n_494, n_493);
  nand g1371 (n_1341, n_492, n_494);
  nand g1372 (n_511, n_1339, n_1340, n_1341);
  xor g1373 (n_1342, A[20], A[21]);
  xor g1374 (n_497, n_1342, n_495);
  nand g1375 (n_1343, A[20], A[21]);
  nand g1376 (n_1344, n_495, A[21]);
  nand g1377 (n_1345, A[20], n_495);
  nand g1378 (n_512, n_1343, n_1344, n_1345);
  xor g1380 (n_499, n_1346, n_497);
  nand g1383 (n_1349, n_496, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  nand g1397 (n_1357, A[10], n_503);
  nand g1398 (n_520, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], A[14]);
  xor g1400 (n_506, n_1358, n_504);
  nand g1401 (n_1359, A[13], A[14]);
  nand g1402 (n_1360, n_504, A[14]);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_521, n_1359, n_1360, n_1361);
  xor g1405 (n_1362, n_505, A[17]);
  xor g1406 (n_509, n_1362, n_506);
  nand g1407 (n_1363, n_505, A[17]);
  nand g1408 (n_1364, n_506, A[17]);
  nand g1409 (n_1365, n_505, n_506);
  nand g1410 (n_523, n_1363, n_1364, n_1365);
  xor g1411 (n_1366, A[18], n_507);
  xor g1412 (n_510, n_1366, n_508);
  nand g1413 (n_1367, A[18], n_507);
  nand g1414 (n_1368, n_508, n_507);
  nand g1415 (n_1369, A[18], n_508);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_509, A[21]);
  xor g1418 (n_513, n_1370, A[22]);
  nand g1419 (n_1371, n_509, A[21]);
  nand g1421 (n_1373, n_509, A[22]);
  nand g1422 (n_527, n_1371, n_1077, n_1373);
  xor g1423 (n_1374, n_510, n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, n_510, n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, n_510, n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1437 (n_1382, A[9], A[11]);
  nand g1439 (n_1383, A[9], A[11]);
  nand g1442 (n_532, n_1383, n_1384, n_1385);
  xor g1443 (n_1386, A[14], n_519);
  xor g1444 (n_522, n_1386, n_520);
  nand g1445 (n_1387, A[14], n_519);
  nand g1446 (n_1388, n_520, n_519);
  nand g1447 (n_1389, A[14], n_520);
  nand g1448 (n_534, n_1387, n_1388, n_1389);
  xor g1449 (n_1390, A[15], n_521);
  xor g1450 (n_524, n_1390, n_522);
  nand g1451 (n_1391, A[15], n_521);
  nand g1452 (n_1392, n_522, n_521);
  nand g1453 (n_1393, A[15], n_522);
  nand g1454 (n_536, n_1391, n_1392, n_1393);
  xor g1455 (n_1394, A[18], n_523);
  xor g1456 (n_525, n_1394, A[19]);
  nand g1457 (n_1395, A[18], n_523);
  nand g1458 (n_1396, A[19], n_523);
  nand g1459 (n_1397, A[18], A[19]);
  nand g1460 (n_538, n_1395, n_1396, n_1397);
  xor g1461 (n_1398, n_524, n_525);
  xor g1462 (n_528, n_1398, n_526);
  nand g1463 (n_1399, n_524, n_525);
  nand g1464 (n_1400, n_526, n_525);
  nand g1465 (n_1401, n_524, n_526);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1468 (n_529, n_1122, n_527);
  nand g1470 (n_1404, n_527, A[23]);
  nand g1471 (n_1405, A[22], n_527);
  nand g1472 (n_543, n_1123, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1480 (n_533, n_1098, A[12]);
  nand g1482 (n_1412, A[12], A[10]);
  nand g1483 (n_1413, A[11], A[12]);
  nand g1484 (n_544, n_1099, n_1412, n_1413);
  xor g1485 (n_1414, n_532, n_533);
  xor g1486 (n_535, n_1414, A[15]);
  nand g1487 (n_1415, n_532, n_533);
  nand g1488 (n_1416, A[15], n_533);
  nand g1489 (n_1417, n_532, A[15]);
  nand g1490 (n_546, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, A[16], n_534);
  xor g1492 (n_537, n_1418, n_535);
  nand g1493 (n_1419, A[16], n_534);
  nand g1494 (n_1420, n_535, n_534);
  nand g1495 (n_1421, A[16], n_535);
  nand g1496 (n_547, n_1419, n_1420, n_1421);
  xor g1497 (n_1422, A[19], n_536);
  xor g1498 (n_539, n_1422, A[20]);
  nand g1499 (n_1423, A[19], n_536);
  nand g1500 (n_1424, A[20], n_536);
  nand g1502 (n_549, n_1423, n_1424, n_992);
  xor g1503 (n_1426, n_537, n_538);
  xor g1504 (n_541, n_1426, n_539);
  nand g1505 (n_1427, n_537, n_538);
  nand g1506 (n_1428, n_539, n_538);
  nand g1507 (n_1429, n_537, n_539);
  nand g1508 (n_551, n_1427, n_1428, n_1429);
  xor g1510 (n_542, n_1166, n_540);
  nand g1513 (n_1433, A[23], n_540);
  nand g1514 (n_554, n_1167, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1522 (n_545, n_1186, n_544);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_876, n_1440, n_1441);
  xor g1527 (n_1442, A[16], n_545);
  xor g1528 (n_548, n_1442, A[17]);
  nand g1529 (n_1443, A[16], n_545);
  nand g1530 (n_1444, A[17], n_545);
  nand g1532 (n_559, n_1443, n_1444, n_1025);
  xor g1533 (n_1446, n_546, n_547);
  xor g1534 (n_550, n_1446, n_548);
  nand g1535 (n_1447, n_546, n_547);
  nand g1536 (n_1448, n_548, n_547);
  nand g1537 (n_1449, n_546, n_548);
  nand g1538 (n_561, n_1447, n_1448, n_1449);
  xor g1540 (n_552, n_1342, n_549);
  nand g1542 (n_1452, n_549, A[21]);
  nand g1543 (n_1453, A[20], n_549);
  nand g1544 (n_563, n_1343, n_1452, n_1453);
  xor g1546 (n_553, n_1454, n_551);
  nand g1549 (n_1457, n_550, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1563 (n_1465, A[14], n_557);
  nand g1564 (n_570, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, A[17], A[18]);
  xor g1566 (n_560, n_1466, n_558);
  nand g1568 (n_1468, n_558, A[18]);
  nand g1569 (n_1469, A[17], n_558);
  nand g1570 (n_571, n_1068, n_1468, n_1469);
  xor g1571 (n_1470, n_559, n_560);
  xor g1572 (n_562, n_1470, n_561);
  nand g1573 (n_1471, n_559, n_560);
  nand g1574 (n_1472, n_561, n_560);
  nand g1575 (n_1473, n_559, n_561);
  nand g1576 (n_574, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, A[21], A[22]);
  xor g1578 (n_564, n_1474, n_562);
  nand g1580 (n_1476, n_562, A[22]);
  nand g1581 (n_1477, A[21], n_562);
  nand g1582 (n_575, n_1077, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  nand g1596 (n_578, n_948, n_1484, n_1463);
  xor g1597 (n_1486, A[18], n_569);
  xor g1598 (n_572, n_1486, n_570);
  nand g1599 (n_1487, A[18], n_569);
  nand g1600 (n_1488, n_570, n_569);
  nand g1601 (n_1489, A[18], n_570);
  nand g1602 (n_580, n_1487, n_1488, n_1489);
  xor g1603 (n_1490, A[19], n_571);
  xor g1604 (n_573, n_1490, n_572);
  nand g1605 (n_1491, A[19], n_571);
  nand g1606 (n_1492, n_572, n_571);
  nand g1607 (n_1493, A[19], n_572);
  nand g1608 (n_582, n_1491, n_1492, n_1493);
  xor g1609 (n_1494, A[22], n_573);
  xor g1610 (n_576, n_1494, A[23]);
  nand g1611 (n_1495, A[22], n_573);
  nand g1612 (n_1496, A[23], n_573);
  nand g1614 (n_584, n_1495, n_1496, n_1123);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1621 (n_1502, A[15], A[13]);
  xor g1622 (n_579, n_1502, A[16]);
  nand g1624 (n_1504, A[16], A[13]);
  nand g1626 (n_586, n_773, n_1504, n_984);
  xor g1627 (n_1506, n_578, n_579);
  xor g1628 (n_581, n_1506, A[19]);
  nand g1629 (n_1507, n_578, n_579);
  nand g1630 (n_1508, A[19], n_579);
  nand g1631 (n_1509, n_578, A[19]);
  nand g1632 (n_588, n_1507, n_1508, n_1509);
  xor g1633 (n_1510, A[20], n_580);
  xor g1634 (n_583, n_1510, n_581);
  nand g1635 (n_1511, A[20], n_580);
  nand g1636 (n_1512, n_581, n_580);
  nand g1637 (n_1513, A[20], n_581);
  nand g1638 (n_589, n_1511, n_1512, n_1513);
  xor g1639 (n_1514, n_582, n_583);
  xor g1640 (n_585, n_1514, A[23]);
  nand g1641 (n_1515, n_582, n_583);
  nand g1642 (n_1516, A[23], n_583);
  nand g1643 (n_1517, n_582, A[23]);
  nand g1644 (n_591, n_1515, n_1516, n_1517);
  xor g1646 (n_83, n_1518, n_585);
  nand g1648 (n_1520, n_585, n_584);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1652 (n_587, n_1194, n_586);
  nand g1654 (n_1524, n_586, A[17]);
  nand g1655 (n_1525, A[16], n_586);
  nand g1656 (n_595, n_1025, n_1524, n_1525);
  xor g1657 (n_1526, A[20], n_587);
  xor g1658 (n_590, n_1526, n_588);
  nand g1659 (n_1527, A[20], n_587);
  nand g1660 (n_1528, n_588, n_587);
  nand g1661 (n_1529, A[20], n_588);
  nand g1662 (n_597, n_1527, n_1528, n_1529);
  xor g1664 (n_592, n_1530, n_589);
  nand g1667 (n_1533, A[21], n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_81, n_1535, n_1536, n_1537);
  nand g1681 (n_1541, A[18], n_595);
  nand g1682 (n_604, n_1539, n_1540, n_1541);
  xor g1684 (n_598, n_1474, n_596);
  nand g1686 (n_1544, n_596, A[22]);
  nand g1687 (n_1545, A[21], n_596);
  nand g1688 (n_606, n_1077, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_33, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[17], A[19]);
  nand g1702 (n_608, n_889, n_1552, n_1553);
  xor g1703 (n_1554, A[22], n_603);
  xor g1704 (n_605, n_1554, n_604);
  nand g1705 (n_1555, A[22], n_603);
  nand g1706 (n_1556, n_604, n_603);
  nand g1707 (n_1557, A[22], n_604);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, A[23], n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, A[23], n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, A[23], n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1715 (n_1562, A[19], A[18]);
  xor g1716 (n_609, n_1562, A[20]);
  nand g1720 (n_612, n_1397, n_925, n_992);
  xor g1721 (n_1566, n_608, n_609);
  xor g1722 (n_611, n_1566, A[23]);
  nand g1723 (n_1567, n_608, n_609);
  nand g1724 (n_1568, A[23], n_609);
  nand g1725 (n_1569, n_608, A[23]);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1728 (n_79, n_1570, n_611);
  nand g1730 (n_1572, n_611, n_610);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1734 (n_613, n_1342, n_612);
  nand g1736 (n_1576, n_612, A[21]);
  nand g1737 (n_1577, A[20], n_612);
  nand g1738 (n_617, n_1343, n_1576, n_1577);
  xor g1740 (n_78, n_1578, n_614);
  nand g1742 (n_1580, n_614, n_613);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_617);
  nand g1752 (n_28, n_1583, n_1584, n_1585);
  nand g1759 (n_1589, A[21], A[23]);
  nand g1760 (n_27, n_1587, n_1588, n_1589);
  xor g1762 (n_75, n_1166, A[22]);
  nand g1766 (n_74, n_1167, n_1123, n_1593);
  nand g16 (n_1606, A[0], A[2]);
  xor g20 (Z[2], A[0], A[2]);
  nand g22 (n_1611, A[3], n_68);
  nand g25 (n_1615, n_1611, n_1612, n_1613);
  xor g26 (n_1614, A[3], n_68);
  nand g28 (n_1616, A[4], n_117);
  nand g29 (n_1617, A[4], n_1615);
  nand g30 (n_1618, n_117, n_1615);
  nand g31 (n_1620, n_1616, n_1617, n_1618);
  xor g32 (n_1619, A[4], n_117);
  xor g33 (Z[4], n_1615, n_1619);
  nand g34 (n_1621, A[5], n_116);
  nand g35 (n_1622, A[5], n_1620);
  nand g36 (n_1623, n_116, n_1620);
  nand g37 (n_1625, n_1621, n_1622, n_1623);
  xor g38 (n_1624, A[5], n_116);
  xor g39 (Z[5], n_1620, n_1624);
  nand g40 (n_1626, n_67, n_115);
  nand g41 (n_1627, n_67, n_1625);
  nand g42 (n_1628, n_115, n_1625);
  nand g43 (n_1630, n_1626, n_1627, n_1628);
  xor g44 (n_1629, n_67, n_115);
  xor g45 (Z[6], n_1625, n_1629);
  nand g46 (n_1631, n_66, n_114);
  nand g47 (n_1632, n_66, n_1630);
  nand g48 (n_1633, n_114, n_1630);
  nand g49 (n_1635, n_1631, n_1632, n_1633);
  xor g50 (n_1634, n_66, n_114);
  xor g51 (Z[7], n_1630, n_1634);
  nand g52 (n_1636, n_65, n_113);
  nand g53 (n_1637, n_65, n_1635);
  nand g54 (n_1638, n_113, n_1635);
  nand g55 (n_1640, n_1636, n_1637, n_1638);
  xor g56 (n_1639, n_65, n_113);
  xor g57 (Z[8], n_1635, n_1639);
  nand g58 (n_1641, n_64, n_112);
  nand g59 (n_1642, n_64, n_1640);
  nand g60 (n_1643, n_112, n_1640);
  nand g61 (n_1645, n_1641, n_1642, n_1643);
  xor g62 (n_1644, n_64, n_112);
  xor g63 (Z[9], n_1640, n_1644);
  nand g64 (n_1646, n_63, n_111);
  nand g65 (n_1647, n_63, n_1645);
  nand g66 (n_1648, n_111, n_1645);
  nand g67 (n_1650, n_1646, n_1647, n_1648);
  xor g68 (n_1649, n_63, n_111);
  xor g69 (Z[10], n_1645, n_1649);
  nand g70 (n_1651, n_62, n_110);
  nand g71 (n_1652, n_62, n_1650);
  nand g72 (n_1653, n_110, n_1650);
  nand g73 (n_1655, n_1651, n_1652, n_1653);
  xor g74 (n_1654, n_62, n_110);
  xor g75 (Z[11], n_1650, n_1654);
  nand g76 (n_1656, n_61, n_109);
  nand g77 (n_1657, n_61, n_1655);
  nand g78 (n_1658, n_109, n_1655);
  nand g79 (n_1660, n_1656, n_1657, n_1658);
  xor g80 (n_1659, n_61, n_109);
  xor g81 (Z[12], n_1655, n_1659);
  nand g82 (n_1661, n_60, n_108);
  nand g83 (n_1662, n_60, n_1660);
  nand g84 (n_1663, n_108, n_1660);
  nand g85 (n_1665, n_1661, n_1662, n_1663);
  xor g86 (n_1664, n_60, n_108);
  xor g87 (Z[13], n_1660, n_1664);
  nand g88 (n_1666, n_59, n_107);
  nand g89 (n_1667, n_59, n_1665);
  nand g90 (n_1668, n_107, n_1665);
  nand g91 (n_1670, n_1666, n_1667, n_1668);
  xor g92 (n_1669, n_59, n_107);
  xor g93 (Z[14], n_1665, n_1669);
  nand g94 (n_1671, n_58, n_106);
  nand g95 (n_1672, n_58, n_1670);
  nand g96 (n_1673, n_106, n_1670);
  nand g97 (n_1675, n_1671, n_1672, n_1673);
  xor g98 (n_1674, n_58, n_106);
  xor g99 (Z[15], n_1670, n_1674);
  nand g100 (n_1676, n_57, n_105);
  nand g101 (n_1677, n_57, n_1675);
  nand g102 (n_1678, n_105, n_1675);
  nand g103 (n_1680, n_1676, n_1677, n_1678);
  xor g104 (n_1679, n_57, n_105);
  xor g105 (Z[16], n_1675, n_1679);
  nand g106 (n_1681, n_56, n_104);
  nand g107 (n_1682, n_56, n_1680);
  nand g108 (n_1683, n_104, n_1680);
  nand g109 (n_1685, n_1681, n_1682, n_1683);
  xor g110 (n_1684, n_56, n_104);
  xor g111 (Z[17], n_1680, n_1684);
  nand g112 (n_1686, n_55, n_103);
  nand g113 (n_1687, n_55, n_1685);
  nand g114 (n_1688, n_103, n_1685);
  nand g115 (n_1690, n_1686, n_1687, n_1688);
  xor g116 (n_1689, n_55, n_103);
  xor g117 (Z[18], n_1685, n_1689);
  nand g118 (n_1691, n_54, n_102);
  nand g119 (n_1692, n_54, n_1690);
  nand g120 (n_1693, n_102, n_1690);
  nand g121 (n_1695, n_1691, n_1692, n_1693);
  xor g122 (n_1694, n_54, n_102);
  xor g123 (Z[19], n_1690, n_1694);
  nand g124 (n_1696, n_53, n_101);
  nand g125 (n_1697, n_53, n_1695);
  nand g126 (n_1698, n_101, n_1695);
  nand g127 (n_1700, n_1696, n_1697, n_1698);
  xor g128 (n_1699, n_53, n_101);
  xor g129 (Z[20], n_1695, n_1699);
  nand g130 (n_1701, n_52, n_100);
  nand g131 (n_1702, n_52, n_1700);
  nand g132 (n_1703, n_100, n_1700);
  nand g133 (n_1705, n_1701, n_1702, n_1703);
  xor g134 (n_1704, n_52, n_100);
  xor g135 (Z[21], n_1700, n_1704);
  nand g136 (n_1706, n_51, n_99);
  nand g137 (n_1707, n_51, n_1705);
  nand g138 (n_1708, n_99, n_1705);
  nand g139 (n_1710, n_1706, n_1707, n_1708);
  xor g140 (n_1709, n_51, n_99);
  xor g141 (Z[22], n_1705, n_1709);
  nand g142 (n_1711, n_50, n_98);
  nand g143 (n_1712, n_50, n_1710);
  nand g144 (n_1713, n_98, n_1710);
  nand g145 (n_1715, n_1711, n_1712, n_1713);
  xor g146 (n_1714, n_50, n_98);
  xor g147 (Z[23], n_1710, n_1714);
  nand g148 (n_1716, n_49, n_97);
  nand g149 (n_1717, n_49, n_1715);
  nand g150 (n_1718, n_97, n_1715);
  nand g151 (n_1720, n_1716, n_1717, n_1718);
  xor g152 (n_1719, n_49, n_97);
  xor g153 (Z[24], n_1715, n_1719);
  nand g154 (n_1721, n_48, n_96);
  nand g155 (n_1722, n_48, n_1720);
  nand g156 (n_1723, n_96, n_1720);
  nand g157 (n_1725, n_1721, n_1722, n_1723);
  xor g158 (n_1724, n_48, n_96);
  xor g159 (Z[25], n_1720, n_1724);
  nand g160 (n_1726, n_47, n_95);
  nand g161 (n_1727, n_47, n_1725);
  nand g162 (n_1728, n_95, n_1725);
  nand g163 (n_1730, n_1726, n_1727, n_1728);
  xor g164 (n_1729, n_47, n_95);
  xor g165 (Z[26], n_1725, n_1729);
  nand g166 (n_1731, n_46, n_94);
  nand g167 (n_1732, n_46, n_1730);
  nand g168 (n_1733, n_94, n_1730);
  nand g169 (n_1735, n_1731, n_1732, n_1733);
  xor g170 (n_1734, n_46, n_94);
  xor g171 (Z[27], n_1730, n_1734);
  nand g172 (n_1736, n_45, n_93);
  nand g173 (n_1737, n_45, n_1735);
  nand g174 (n_1738, n_93, n_1735);
  nand g175 (n_1740, n_1736, n_1737, n_1738);
  xor g176 (n_1739, n_45, n_93);
  xor g177 (Z[28], n_1735, n_1739);
  nand g178 (n_1741, n_44, n_92);
  nand g179 (n_1742, n_44, n_1740);
  nand g180 (n_1743, n_92, n_1740);
  nand g181 (n_1745, n_1741, n_1742, n_1743);
  xor g182 (n_1744, n_44, n_92);
  xor g183 (Z[29], n_1740, n_1744);
  nand g184 (n_1746, n_43, n_91);
  nand g185 (n_1747, n_43, n_1745);
  nand g186 (n_1748, n_91, n_1745);
  nand g187 (n_1750, n_1746, n_1747, n_1748);
  xor g188 (n_1749, n_43, n_91);
  xor g189 (Z[30], n_1745, n_1749);
  nand g190 (n_1751, n_42, n_90);
  nand g191 (n_1752, n_42, n_1750);
  nand g192 (n_1753, n_90, n_1750);
  nand g193 (n_1755, n_1751, n_1752, n_1753);
  xor g194 (n_1754, n_42, n_90);
  xor g195 (Z[31], n_1750, n_1754);
  nand g196 (n_1756, n_41, n_89);
  nand g197 (n_1757, n_41, n_1755);
  nand g198 (n_1758, n_89, n_1755);
  nand g199 (n_1760, n_1756, n_1757, n_1758);
  xor g200 (n_1759, n_41, n_89);
  xor g201 (Z[32], n_1755, n_1759);
  nand g202 (n_1761, n_40, n_88);
  nand g203 (n_1762, n_40, n_1760);
  nand g204 (n_1763, n_88, n_1760);
  nand g205 (n_1765, n_1761, n_1762, n_1763);
  xor g206 (n_1764, n_40, n_88);
  xor g207 (Z[33], n_1760, n_1764);
  nand g208 (n_1766, n_39, n_87);
  nand g209 (n_1767, n_39, n_1765);
  nand g210 (n_1768, n_87, n_1765);
  nand g211 (n_1770, n_1766, n_1767, n_1768);
  xor g212 (n_1769, n_39, n_87);
  xor g213 (Z[34], n_1765, n_1769);
  nand g214 (n_1771, n_38, n_86);
  nand g215 (n_1772, n_38, n_1770);
  nand g216 (n_1773, n_86, n_1770);
  nand g217 (n_1775, n_1771, n_1772, n_1773);
  xor g218 (n_1774, n_38, n_86);
  xor g219 (Z[35], n_1770, n_1774);
  nand g220 (n_1776, n_37, n_85);
  nand g221 (n_1777, n_37, n_1775);
  nand g222 (n_1778, n_85, n_1775);
  nand g223 (n_1780, n_1776, n_1777, n_1778);
  xor g224 (n_1779, n_37, n_85);
  xor g225 (Z[36], n_1775, n_1779);
  nand g226 (n_1781, n_36, n_84);
  nand g227 (n_1782, n_36, n_1780);
  nand g228 (n_1783, n_84, n_1780);
  nand g229 (n_1785, n_1781, n_1782, n_1783);
  xor g230 (n_1784, n_36, n_84);
  xor g231 (Z[37], n_1780, n_1784);
  nand g232 (n_1786, n_35, n_83);
  nand g233 (n_1787, n_35, n_1785);
  nand g234 (n_1788, n_83, n_1785);
  nand g235 (n_1790, n_1786, n_1787, n_1788);
  xor g236 (n_1789, n_35, n_83);
  xor g237 (Z[38], n_1785, n_1789);
  nand g238 (n_1791, n_34, n_82);
  nand g239 (n_1792, n_34, n_1790);
  nand g240 (n_1793, n_82, n_1790);
  nand g241 (n_1795, n_1791, n_1792, n_1793);
  xor g242 (n_1794, n_34, n_82);
  xor g243 (Z[39], n_1790, n_1794);
  nand g244 (n_1796, n_33, n_81);
  nand g245 (n_1797, n_33, n_1795);
  nand g246 (n_1798, n_81, n_1795);
  nand g247 (n_1800, n_1796, n_1797, n_1798);
  xor g248 (n_1799, n_33, n_81);
  xor g249 (Z[40], n_1795, n_1799);
  nand g250 (n_1801, n_32, n_80);
  nand g251 (n_1802, n_32, n_1800);
  nand g252 (n_1803, n_80, n_1800);
  nand g253 (n_1805, n_1801, n_1802, n_1803);
  xor g254 (n_1804, n_32, n_80);
  xor g255 (Z[41], n_1800, n_1804);
  nand g256 (n_1806, n_31, n_79);
  nand g257 (n_1807, n_31, n_1805);
  nand g258 (n_1808, n_79, n_1805);
  nand g259 (n_1810, n_1806, n_1807, n_1808);
  xor g260 (n_1809, n_31, n_79);
  xor g261 (Z[42], n_1805, n_1809);
  nand g262 (n_1811, n_30, n_78);
  nand g263 (n_1812, n_30, n_1810);
  nand g264 (n_1813, n_78, n_1810);
  nand g265 (n_1815, n_1811, n_1812, n_1813);
  xor g266 (n_1814, n_30, n_78);
  xor g267 (Z[43], n_1810, n_1814);
  nand g1772 (n_1816, n_29, n_77);
  nand g1773 (n_1817, n_29, n_1815);
  nand g1774 (n_1818, n_77, n_1815);
  nand g1775 (n_1820, n_1816, n_1817, n_1818);
  xor g1776 (n_1819, n_29, n_77);
  xor g1777 (Z[44], n_1815, n_1819);
  nand g1778 (n_1821, n_28, n_76);
  nand g1779 (n_1822, n_28, n_1820);
  nand g1780 (n_1823, n_76, n_1820);
  nand g1781 (n_1825, n_1821, n_1822, n_1823);
  xor g1782 (n_1824, n_28, n_76);
  xor g1783 (Z[45], n_1820, n_1824);
  nand g1784 (n_1826, n_27, n_75);
  nand g1785 (n_1827, n_27, n_1825);
  nand g1786 (n_1828, n_75, n_1825);
  nand g1787 (n_1830, n_1826, n_1827, n_1828);
  xor g1788 (n_1829, n_27, n_75);
  xor g1789 (Z[46], n_1825, n_1829);
  xor g1791 (Z[47], n_1830, n_1831);
  or g1803 (n_1044, A[1], wc);
  not gc (wc, n_171);
  or g1804 (n_1045, A[1], wc0);
  not gc0 (wc0, A[2]);
  or g1805 (n_1088, wc1, A[2]);
  not gc1 (wc1, A[1]);
  or g1806 (n_1089, A[2], wc2);
  not gc2 (wc2, A[3]);
  xnor g1807 (n_1166, A[24], A[23]);
  or g1808 (n_1167, wc3, A[24]);
  not gc3 (wc3, A[23]);
  xnor g1809 (n_1214, A[6], A[5]);
  or g1810 (n_1215, A[5], wc4);
  not gc4 (wc4, A[6]);
  or g1811 (n_1252, A[6], wc5);
  not gc5 (wc5, A[7]);
  or g1812 (n_1253, wc6, A[6]);
  not gc6 (wc6, A[5]);
  or g1814 (n_1355, A[9], wc7);
  not gc7 (wc7, A[10]);
  or g1815 (n_1384, A[10], wc8);
  not gc8 (wc8, A[11]);
  or g1816 (n_1385, wc9, A[10]);
  not gc9 (wc9, A[9]);
  or g1818 (n_1463, A[13], wc10);
  not gc10 (wc10, A[14]);
  xnor g1819 (n_1530, A[24], A[21]);
  or g1820 (n_1531, wc11, A[24]);
  not gc11 (wc11, A[21]);
  or g1822 (n_1539, A[17], wc12);
  not gc12 (wc12, A[18]);
  or g1823 (n_1552, A[18], wc13);
  not gc13 (wc13, A[19]);
  or g1824 (n_1553, wc14, A[18]);
  not gc14 (wc14, A[17]);
  or g1826 (n_1583, A[21], wc15);
  not gc15 (wc15, A[22]);
  or g1827 (n_1587, wc16, A[22]);
  not gc16 (wc16, A[21]);
  or g1828 (n_1588, A[22], wc17);
  not gc17 (wc17, A[23]);
  or g1829 (n_1593, wc18, A[24]);
  not gc18 (wc18, A[22]);
  xnor g1830 (n_349, n_1042, A[1]);
  xnor g1831 (n_372, n_1086, A[2]);
  xnor g1832 (n_453, n_1250, A[6]);
  xnor g1833 (n_519, n_1382, A[10]);
  xnor g1834 (n_569, n_1106, A[13]);
  or g1835 (n_1484, A[13], wc19);
  not gc19 (wc19, A[15]);
  xnor g1836 (n_603, n_1550, A[18]);
  xnor g1837 (n_76, n_1474, A[23]);
  xnor g1838 (n_1578, n_613, A[24]);
  or g1839 (n_1579, A[24], wc20);
  not gc20 (wc20, n_613);
  xnor g1840 (n_1831, n_74, A[24]);
  or g1841 (n_1216, A[5], wc21);
  not gc21 (wc21, n_433);
  xnor g1842 (n_505, n_1218, n_503);
  or g1843 (n_1356, A[9], wc22);
  not gc22 (wc22, n_503);
  xnor g1844 (n_558, n_1358, n_557);
  or g1845 (n_1464, A[13], wc23);
  not gc23 (wc23, n_557);
  or g1846 (n_1573, A[24], wc24);
  not gc24 (wc24, n_611);
  or g1847 (n_1581, A[24], wc25);
  not gc25 (wc25, n_614);
  xnor g1848 (n_29, n_1474, n_617);
  or g1849 (n_1584, A[21], wc26);
  not gc26 (wc26, n_617);
  xnor g1851 (n_596, n_1466, n_595);
  or g1852 (n_1540, A[17], wc27);
  not gc27 (wc27, n_595);
  or g1853 (n_1612, wc28, n_1606);
  not gc28 (wc28, A[3]);
  or g1854 (n_1613, n_1606, wc29);
  not gc29 (wc29, n_68);
  xnor g1855 (Z[3], n_1606, n_1614);
  xnor g1856 (n_1570, n_610, A[24]);
  or g1857 (n_1571, A[24], wc30);
  not gc30 (wc30, n_610);
  or g1858 (n_1532, A[24], wc31);
  not gc31 (wc31, n_589);
  xnor g1859 (n_1518, n_584, A[24]);
  or g1860 (n_1519, A[24], wc32);
  not gc32 (wc32, n_584);
  xnor g1861 (n_1454, n_550, A[24]);
  or g1862 (n_1455, A[24], wc33);
  not gc33 (wc33, n_550);
  or g1863 (n_1521, A[24], wc34);
  not gc34 (wc34, n_585);
  or g1864 (n_1081, A[24], wc35);
  not gc35 (wc35, n_363);
  or g1865 (n_1456, A[24], wc36);
  not gc36 (wc36, n_551);
  or g1866 (n_1080, A[24], wc37);
  not gc37 (wc37, n_364);
  xnor g1867 (n_1206, n_426, A[24]);
  or g1868 (n_1207, A[24], wc38);
  not gc38 (wc38, n_426);
  xnor g1869 (n_367, n_1078, A[24]);
  or g1870 (n_1208, A[24], wc39);
  not gc39 (wc39, n_427);
  xnor g1871 (n_1346, n_496, A[24]);
  or g1872 (n_1347, A[24], wc40);
  not gc40 (wc40, n_496);
  or g1873 (n_1348, A[24], wc41);
  not gc41 (wc41, n_497);
  or g1874 (n_1169, A[24], wc42);
  not gc42 (wc42, n_408);
  or g1875 (n_1316, A[24], wc43);
  not gc43 (wc43, n_482);
  or g1876 (n_1432, A[24], wc44);
  not gc44 (wc44, n_540);
endmodule

module mult_signed_const_4953_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_4953_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_5220_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_176;
  wire n_179, n_180, n_183, n_184, n_187, n_188, n_189, n_196;
  wire n_201, n_202, n_203, n_204, n_209, n_210, n_211, n_212;
  wire n_217, n_218, n_219, n_220, n_221, n_223, n_224, n_225;
  wire n_226, n_227, n_234, n_236, n_237, n_238, n_239, n_248;
  wire n_249, n_250, n_251, n_258, n_260, n_261, n_262, n_267;
  wire n_269, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_282, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_300, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_333, n_335, n_337, n_338;
  wire n_340, n_341, n_342, n_343, n_344, n_345, n_354, n_356;
  wire n_357, n_358, n_359, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_449, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_470, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_498, n_499, n_500, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_519, n_520, n_521, n_522, n_523, n_524;
  wire n_525, n_526, n_527, n_528, n_529, n_530, n_532, n_533;
  wire n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541;
  wire n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_557, n_558, n_559;
  wire n_560, n_561, n_562, n_563, n_564, n_565, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_578, n_579;
  wire n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587;
  wire n_588, n_589, n_590, n_591, n_592, n_595, n_596, n_597;
  wire n_598, n_599, n_603, n_604, n_605, n_606, n_608, n_609;
  wire n_610, n_611, n_612, n_613, n_614, n_617, n_622, n_623;
  wire n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631;
  wire n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639;
  wire n_640, n_641, n_646, n_647, n_648, n_649, n_650, n_651;
  wire n_652, n_653, n_658, n_659, n_660, n_661, n_662, n_663;
  wire n_664, n_665, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_684, n_685, n_686, n_687;
  wire n_688, n_689, n_690, n_691, n_692, n_693, n_704, n_705;
  wire n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_722, n_724, n_725, n_726, n_727, n_728, n_729, n_730;
  wire n_731, n_732, n_733, n_738, n_742, n_743, n_744, n_745;
  wire n_746, n_747, n_748, n_749, n_750, n_751, n_752, n_753;
  wire n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771;
  wire n_772, n_773, n_774, n_775, n_776, n_777, n_794, n_795;
  wire n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803;
  wire n_804, n_805, n_822, n_823, n_824, n_826, n_827, n_828;
  wire n_829, n_830, n_831, n_832, n_833, n_842, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_868, n_869, n_870, n_871;
  wire n_872, n_873, n_876, n_877, n_880, n_881, n_882, n_883;
  wire n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891;
  wire n_892, n_893, n_906, n_907, n_908, n_910, n_911, n_912;
  wire n_913, n_914, n_915, n_916, n_917, n_918, n_919, n_920;
  wire n_921, n_922, n_923, n_924, n_925, n_926, n_927, n_928;
  wire n_929, n_946, n_947, n_949, n_950, n_951, n_952, n_953;
  wire n_954, n_955, n_956, n_957, n_958, n_959, n_960, n_961;
  wire n_962, n_963, n_964, n_965, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_996, n_997, n_998, n_999, n_1000, n_1001, n_1013, n_1014;
  wire n_1015, n_1016, n_1017, n_1020, n_1021, n_1026, n_1027, n_1028;
  wire n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036;
  wire n_1037, n_1038, n_1039, n_1040, n_1041, n_1043, n_1044, n_1047;
  wire n_1049, n_1051, n_1052, n_1056, n_1057, n_1058, n_1059, n_1060;
  wire n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068;
  wire n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076;
  wire n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084;
  wire n_1085, n_1086, n_1088, n_1090, n_1091, n_1092, n_1093, n_1094;
  wire n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102;
  wire n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110;
  wire n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118;
  wire n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126;
  wire n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134;
  wire n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142;
  wire n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150;
  wire n_1151, n_1152, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159;
  wire n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167;
  wire n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175;
  wire n_1176, n_1177, n_1178, n_1179, n_1180, n_1182, n_1183, n_1184;
  wire n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192;
  wire n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200;
  wire n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208;
  wire n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216;
  wire n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224;
  wire n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232;
  wire n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1241;
  wire n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249;
  wire n_1250, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258;
  wire n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1266, n_1267;
  wire n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275;
  wire n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283;
  wire n_1284, n_1285, n_1286, n_1288, n_1290, n_1291, n_1292, n_1293;
  wire n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301;
  wire n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309;
  wire n_1310, n_1311, n_1312, n_1313, n_1316, n_1317, n_1318, n_1319;
  wire n_1320, n_1321, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329;
  wire n_1330, n_1331, n_1332, n_1333, n_1334, n_1336, n_1337, n_1338;
  wire n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346;
  wire n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1355;
  wire n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363;
  wire n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371;
  wire n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379;
  wire n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387;
  wire n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395;
  wire n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403;
  wire n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1412, n_1413;
  wire n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421;
  wire n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429;
  wire n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1440, n_1441;
  wire n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451;
  wire n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459;
  wire n_1460, n_1461, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468;
  wire n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476;
  wire n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1484, n_1485;
  wire n_1486, n_1487, n_1488, n_1490, n_1491, n_1492, n_1493, n_1496;
  wire n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1506, n_1507;
  wire n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515;
  wire n_1516, n_1518, n_1519, n_1520, n_1521, n_1524, n_1525, n_1526;
  wire n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534;
  wire n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542;
  wire n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551;
  wire n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559;
  wire n_1560, n_1561, n_1562, n_1565, n_1566, n_1567, n_1568, n_1569;
  wire n_1570, n_1571, n_1572, n_1573, n_1576, n_1577, n_1578, n_1579;
  wire n_1580, n_1581, n_1583, n_1584, n_1585, n_1587, n_1588, n_1589;
  wire n_1593, n_1606, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616;
  wire n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624;
  wire n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632;
  wire n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640;
  wire n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648;
  wire n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656;
  wire n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664;
  wire n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672;
  wire n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680;
  wire n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688;
  wire n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696;
  wire n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704;
  wire n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712;
  wire n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720;
  wire n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728;
  wire n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736;
  wire n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744;
  wire n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752;
  wire n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760;
  wire n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768;
  wire n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776;
  wire n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784;
  wire n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792;
  wire n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800;
  wire n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], n_171);
  xor g270 (n_117, n_622, A[2]);
  nand g3 (n_623, A[1], n_171);
  nand g271 (n_624, A[2], n_171);
  nand g272 (n_625, A[1], A[2]);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, A[4]);
  xor g288 (n_176, n_634, n_69);
  nand g289 (n_635, n_68, A[4]);
  nand g290 (n_636, n_69, A[4]);
  nand g291 (n_637, n_68, n_69);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_176);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_176);
  nand g296 (n_640, A[7], n_176);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g305 (n_646, n_117, A[5]);
  xor g306 (n_180, n_646, A[6]);
  nand g307 (n_647, n_117, A[5]);
  nand g308 (n_648, A[6], A[5]);
  nand g309 (n_649, n_117, A[6]);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, n_179, n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, n_179, n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, n_179, A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_188, n_659, n_660, n_661);
  xor g329 (n_662, n_183, A[9]);
  xor g330 (n_112, n_662, n_184);
  nand g331 (n_663, n_183, A[9]);
  nand g332 (n_664, n_184, A[9]);
  nand g333 (n_665, n_183, n_184);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_187, n_630, n_67);
  nand g340 (n_668, n_67, n_173);
  nand g341 (n_669, A[4], n_67);
  nand g342 (n_71, n_631, n_668, n_669);
  xor g343 (n_670, A[7], n_187);
  xor g344 (n_189, n_670, A[8]);
  nand g345 (n_671, A[7], n_187);
  nand g346 (n_672, A[8], n_187);
  nand g347 (n_673, A[7], A[8]);
  nand g348 (n_73, n_671, n_672, n_673);
  xor g349 (n_674, n_188, A[10]);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, n_188, A[10]);
  nand g352 (n_676, n_189, A[10]);
  nand g353 (n_677, n_188, n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_72, n_638, n_71);
  nand g366 (n_684, n_71, n_176);
  nand g367 (n_685, A[5], n_71);
  nand g368 (n_201, n_639, n_684, n_685);
  xor g369 (n_686, A[8], A[9]);
  xor g370 (n_196, n_686, n_73);
  nand g371 (n_687, A[8], A[9]);
  nand g372 (n_688, n_73, A[9]);
  nand g373 (n_689, A[8], n_73);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, n_72, A[11]);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, n_72, A[11]);
  nand g378 (n_692, n_196, A[11]);
  nand g379 (n_693, n_72, n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g394 (n_202, n_650, A[9]);
  nand g396 (n_704, A[9], n_180);
  nand g397 (n_705, n_179, A[9]);
  nand g398 (n_209, n_651, n_704, n_705);
  xor g399 (n_706, A[10], n_201);
  xor g400 (n_204, n_706, n_202);
  nand g401 (n_707, A[10], n_201);
  nand g402 (n_708, n_202, n_201);
  nand g403 (n_709, A[10], n_202);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, A[12], n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, A[12], n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, A[12], n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g423 (n_722, n_183, n_184);
  xor g424 (n_210, n_722, A[10]);
  nand g426 (n_724, A[10], n_184);
  nand g427 (n_725, n_183, A[10]);
  nand g428 (n_218, n_665, n_724, n_725);
  xor g429 (n_726, A[11], n_209);
  xor g430 (n_212, n_726, n_210);
  nand g431 (n_727, A[11], n_209);
  nand g432 (n_728, n_210, n_209);
  nand g433 (n_729, A[11], n_210);
  nand g434 (n_220, n_727, n_728, n_729);
  xor g435 (n_730, n_211, A[13]);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, n_211, A[13]);
  nand g438 (n_732, n_212, A[13]);
  nand g439 (n_733, n_211, n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_217, n_738, n_187);
  xor g455 (n_742, n_188, n_217);
  xor g456 (n_219, n_742, A[11]);
  nand g457 (n_743, n_188, n_217);
  nand g458 (n_744, A[11], n_217);
  nand g459 (n_745, n_188, A[11]);
  nand g460 (n_224, n_743, n_744, n_745);
  xor g461 (n_746, n_218, A[12]);
  xor g462 (n_221, n_746, A[14]);
  nand g463 (n_747, n_218, A[12]);
  nand g464 (n_748, A[14], A[12]);
  nand g465 (n_749, n_218, A[14]);
  nand g466 (n_226, n_747, n_748, n_749);
  xor g467 (n_750, n_219, n_220);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, n_219, n_220);
  nand g470 (n_752, n_221, n_220);
  nand g471 (n_753, n_219, n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g488 (n_223, n_686, n_72);
  nand g490 (n_764, n_72, A[9]);
  nand g491 (n_765, A[8], n_72);
  nand g492 (n_234, n_687, n_764, n_765);
  xor g493 (n_766, n_73, A[12]);
  xor g494 (n_225, n_766, n_223);
  nand g495 (n_767, n_73, A[12]);
  nand g496 (n_768, n_223, A[12]);
  nand g497 (n_769, n_73, n_223);
  nand g498 (n_236, n_767, n_768, n_769);
  xor g499 (n_770, A[13], n_224);
  xor g500 (n_227, n_770, A[15]);
  nand g501 (n_771, A[13], n_224);
  nand g502 (n_772, A[15], n_224);
  nand g503 (n_773, A[13], A[15]);
  nand g504 (n_238, n_771, n_772, n_773);
  xor g505 (n_774, n_225, n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, n_225, n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, n_225, n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g535 (n_794, n_234, A[13]);
  xor g536 (n_237, n_794, n_204);
  nand g537 (n_795, n_234, A[13]);
  nand g538 (n_796, n_204, A[13]);
  nand g539 (n_797, n_234, n_204);
  nand g540 (n_248, n_795, n_796, n_797);
  xor g541 (n_798, A[14], n_236);
  xor g542 (n_239, n_798, A[16]);
  nand g543 (n_799, A[14], n_236);
  nand g544 (n_800, A[16], n_236);
  nand g545 (n_801, A[14], A[16]);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, n_237, n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, n_237, n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, n_237, n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g577 (n_822, n_211, A[14]);
  xor g578 (n_249, n_822, n_212);
  nand g579 (n_823, n_211, A[14]);
  nand g580 (n_824, n_212, A[14]);
  nand g582 (n_261, n_823, n_824, n_733);
  xor g583 (n_826, A[15], n_248);
  xor g584 (n_251, n_826, A[17]);
  nand g585 (n_827, A[15], n_248);
  nand g586 (n_828, A[17], n_248);
  nand g587 (n_829, A[15], A[17]);
  nand g588 (n_118, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g609 (n_842, n_188, A[11]);
  xor g610 (n_258, n_842, n_217);
  xor g616 (n_260, n_746, n_258);
  nand g618 (n_848, n_258, n_218);
  nand g619 (n_849, A[12], n_258);
  nand g620 (n_272, n_747, n_848, n_849);
  xor g621 (n_850, n_220, A[15]);
  xor g622 (n_262, n_850, n_260);
  nand g623 (n_851, n_220, A[15]);
  nand g624 (n_852, n_260, A[15]);
  nand g625 (n_853, n_220, n_260);
  nand g626 (n_274, n_851, n_852, n_853);
  xor g627 (n_854, A[16], n_261);
  xor g628 (n_119, n_854, A[18]);
  nand g629 (n_855, A[16], n_261);
  nand g630 (n_856, A[18], n_261);
  nand g631 (n_857, A[16], A[18]);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_262, n_118);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_262, n_118);
  nand g636 (n_860, n_119, n_118);
  nand g637 (n_861, n_262, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g648 (n_267, n_638, A[8]);
  nand g650 (n_868, A[8], n_176);
  nand g651 (n_869, A[5], A[8]);
  nand g652 (n_282, n_639, n_868, n_869);
  xor g653 (n_870, n_71, A[9]);
  xor g654 (n_269, n_870, n_267);
  nand g655 (n_871, n_71, A[9]);
  nand g656 (n_872, n_267, A[9]);
  nand g657 (n_873, n_71, n_267);
  nand g658 (n_284, n_871, n_872, n_873);
  xor g660 (n_271, n_766, n_269);
  nand g662 (n_876, n_269, A[12]);
  nand g663 (n_877, n_73, n_269);
  nand g664 (n_286, n_767, n_876, n_877);
  xor g666 (n_273, n_770, n_271);
  nand g668 (n_880, n_271, A[13]);
  nand g669 (n_881, n_224, n_271);
  nand g670 (n_288, n_771, n_880, n_881);
  xor g671 (n_882, n_272, A[16]);
  xor g672 (n_275, n_882, A[17]);
  nand g673 (n_883, n_272, A[16]);
  nand g674 (n_884, A[17], A[16]);
  nand g675 (n_885, n_272, A[17]);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, n_273, n_274);
  xor g678 (n_277, n_886, A[19]);
  nand g679 (n_887, n_273, n_274);
  nand g680 (n_888, A[19], n_274);
  nand g681 (n_889, n_273, A[19]);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g707 (n_906, A[10], n_282);
  xor g708 (n_285, n_906, n_202);
  nand g709 (n_907, A[10], n_282);
  nand g710 (n_908, n_202, n_282);
  nand g712 (n_300, n_907, n_908, n_709);
  xor g713 (n_910, n_284, A[13]);
  xor g714 (n_287, n_910, n_285);
  nand g715 (n_911, n_284, A[13]);
  nand g716 (n_912, n_285, A[13]);
  nand g717 (n_913, n_284, n_285);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, A[14], n_286);
  xor g720 (n_289, n_914, n_287);
  nand g721 (n_915, A[14], n_286);
  nand g722 (n_916, n_287, n_286);
  nand g723 (n_917, A[14], n_287);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, A[17], n_288);
  xor g726 (n_291, n_918, n_289);
  nand g727 (n_919, A[17], n_288);
  nand g728 (n_920, n_289, n_288);
  nand g729 (n_921, A[17], n_289);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, A[18], n_290);
  xor g732 (n_293, n_922, A[20]);
  nand g733 (n_923, A[18], n_290);
  nand g734 (n_924, A[20], n_290);
  nand g735 (n_925, A[18], A[20]);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g767 (n_946, n_300, A[14]);
  xor g768 (n_303, n_946, n_212);
  nand g769 (n_947, n_300, A[14]);
  nand g771 (n_949, n_300, n_212);
  nand g772 (n_319, n_947, n_824, n_949);
  xor g773 (n_950, n_302, A[15]);
  xor g774 (n_305, n_950, n_303);
  nand g775 (n_951, n_302, A[15]);
  nand g776 (n_952, n_303, A[15]);
  nand g777 (n_953, n_302, n_303);
  nand g778 (n_321, n_951, n_952, n_953);
  xor g779 (n_954, n_304, A[18]);
  xor g780 (n_307, n_954, n_305);
  nand g781 (n_955, n_304, A[18]);
  nand g782 (n_956, n_305, A[18]);
  nand g783 (n_957, n_304, n_305);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, A[19], n_306);
  xor g786 (n_309, n_958, A[21]);
  nand g787 (n_959, A[19], n_306);
  nand g788 (n_960, A[21], n_306);
  nand g789 (n_961, A[19], A[21]);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g824 (n_320, n_850, A[16]);
  nand g826 (n_984, A[16], A[15]);
  nand g827 (n_985, n_220, A[16]);
  nand g828 (n_338, n_851, n_984, n_985);
  xor g829 (n_986, n_260, n_319);
  xor g830 (n_322, n_986, n_320);
  nand g831 (n_987, n_260, n_319);
  nand g832 (n_988, n_320, n_319);
  nand g833 (n_989, n_260, n_320);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, n_321, A[19]);
  xor g836 (n_324, n_990, n_322);
  nand g837 (n_991, n_321, A[19]);
  nand g838 (n_992, n_322, A[19]);
  nand g839 (n_993, n_321, n_322);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, A[20], n_323);
  xor g842 (n_326, n_994, A[22]);
  nand g843 (n_995, A[20], n_323);
  nand g844 (n_996, A[22], n_323);
  nand g845 (n_997, A[20], A[22]);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, n_324, n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, n_324, n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, n_324, n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g868 (n_333, n_870, n_73);
  nand g871 (n_1013, n_71, n_73);
  nand g872 (n_354, n_871, n_688, n_1013);
  xor g873 (n_1014, n_267, A[12]);
  xor g874 (n_335, n_1014, n_333);
  nand g875 (n_1015, n_267, A[12]);
  nand g876 (n_1016, n_333, A[12]);
  nand g877 (n_1017, n_267, n_333);
  nand g878 (n_356, n_1015, n_1016, n_1017);
  xor g880 (n_337, n_770, n_335);
  nand g882 (n_1020, n_335, A[13]);
  nand g883 (n_1021, n_224, n_335);
  nand g884 (n_358, n_771, n_1020, n_1021);
  xor g891 (n_1026, n_337, n_338);
  xor g892 (n_341, n_1026, n_275);
  nand g893 (n_1027, n_337, n_338);
  nand g894 (n_1028, n_275, n_338);
  nand g895 (n_1029, n_337, n_275);
  nand g896 (n_362, n_1027, n_1028, n_1029);
  xor g897 (n_1030, A[20], n_340);
  xor g898 (n_343, n_1030, n_341);
  nand g899 (n_1031, A[20], n_340);
  nand g900 (n_1032, n_341, n_340);
  nand g901 (n_1033, A[20], n_341);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, A[21], n_342);
  xor g904 (n_345, n_1034, n_343);
  nand g905 (n_1035, A[21], n_342);
  nand g906 (n_1036, n_343, n_342);
  nand g907 (n_1037, A[21], n_343);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, A[23], n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, A[23], n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, A[23], n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  nand g922 (n_371, n_1043, n_1044, n_624);
  nand g928 (n_373, n_1047, n_648, n_1049);
  nand g934 (n_375, n_1051, n_1052, n_705);
  nand g940 (n_377, n_907, n_1056, n_1057);
  xor g941 (n_1058, n_354, A[13]);
  nand g943 (n_1059, n_354, A[13]);
  nand g946 (n_379, n_1059, n_1060, n_1061);
  xor g947 (n_1062, A[14], n_356);
  xor g948 (n_359, n_1062, n_357);
  nand g949 (n_1063, A[14], n_356);
  nand g950 (n_1064, n_357, n_356);
  nand g951 (n_1065, A[14], n_357);
  nand g952 (n_381, n_1063, n_1064, n_1065);
  xor g953 (n_1066, A[17], n_358);
  xor g954 (n_361, n_1066, A[18]);
  nand g955 (n_1067, A[17], n_358);
  nand g956 (n_1068, A[18], n_358);
  nand g957 (n_1069, A[17], A[18]);
  nand g958 (n_383, n_1067, n_1068, n_1069);
  xor g959 (n_1070, n_359, n_290);
  xor g960 (n_363, n_1070, n_361);
  nand g961 (n_1071, n_359, n_290);
  nand g962 (n_1072, n_361, n_290);
  nand g963 (n_1073, n_359, n_361);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, A[21], n_362);
  xor g966 (n_365, n_1074, A[22]);
  nand g967 (n_1075, A[21], n_362);
  nand g968 (n_1076, A[22], n_362);
  nand g969 (n_1077, A[21], A[22]);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g972 (n_367, n_1078, n_364);
  nand g975 (n_1081, n_363, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  xor g986 (n_372, n_1086, A[3]);
  nand g990 (n_392, n_1044, n_1088, n_627);
  xor g991 (n_1090, n_371, n_372);
  xor g992 (n_374, n_1090, A[6]);
  nand g993 (n_1091, n_371, n_372);
  nand g994 (n_1092, A[6], n_372);
  nand g995 (n_1093, n_371, A[6]);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, n_374);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, n_374, n_373);
  nand g1001 (n_1097, A[7], n_374);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, A[10], A[11]);
  xor g1004 (n_378, n_1098, n_375);
  nand g1005 (n_1099, A[10], A[11]);
  nand g1006 (n_1100, n_375, A[11]);
  nand g1007 (n_1101, A[10], n_375);
  nand g1008 (n_398, n_1099, n_1100, n_1101);
  xor g1009 (n_1102, n_376, n_377);
  xor g1010 (n_380, n_1102, n_378);
  nand g1011 (n_1103, n_376, n_377);
  nand g1012 (n_1104, n_378, n_377);
  nand g1013 (n_1105, n_376, n_378);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, A[14], n_379);
  xor g1016 (n_382, n_1106, A[15]);
  nand g1017 (n_1107, A[14], n_379);
  nand g1018 (n_1108, A[15], n_379);
  nand g1019 (n_1109, A[14], A[15]);
  nand g1020 (n_402, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, n_380, A[18]);
  xor g1022 (n_384, n_1110, n_381);
  nand g1023 (n_1111, n_380, A[18]);
  nand g1024 (n_1112, n_381, A[18]);
  nand g1025 (n_1113, n_380, n_381);
  nand g1026 (n_404, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, n_382, A[19]);
  xor g1028 (n_386, n_1114, n_383);
  nand g1029 (n_1115, n_382, A[19]);
  nand g1030 (n_1116, n_383, A[19]);
  nand g1031 (n_1117, n_382, n_383);
  nand g1032 (n_406, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_384, A[22]);
  xor g1034 (n_388, n_1118, n_385);
  nand g1035 (n_1119, n_384, A[22]);
  nand g1036 (n_1120, n_385, A[22]);
  nand g1037 (n_1121, n_384, n_385);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, n_386, A[23]);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, n_386, A[23]);
  nand g1042 (n_1124, n_387, A[23]);
  nand g1043 (n_1125, n_386, n_387);
  nand g1044 (n_410, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1051 (n_1130, A[1], A[3]);
  xor g1052 (n_393, n_1130, A[4]);
  nand g1053 (n_1131, A[1], A[3]);
  nand g1054 (n_1132, A[4], A[3]);
  nand g1055 (n_1133, A[1], A[4]);
  nand g1056 (n_412, n_1131, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, n_396, A[11]);
  xor g1070 (n_399, n_1142, n_397);
  nand g1071 (n_1143, n_396, A[11]);
  nand g1072 (n_1144, n_397, A[11]);
  nand g1073 (n_1145, n_396, n_397);
  nand g1074 (n_418, n_1143, n_1144, n_1145);
  xor g1075 (n_1146, A[12], n_398);
  xor g1076 (n_401, n_1146, n_399);
  nand g1077 (n_1147, A[12], n_398);
  nand g1078 (n_1148, n_399, n_398);
  nand g1079 (n_1149, A[12], n_399);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, A[15], n_400);
  xor g1082 (n_403, n_1150, A[16]);
  nand g1083 (n_1151, A[15], n_400);
  nand g1084 (n_1152, A[16], n_400);
  nand g1086 (n_421, n_1151, n_1152, n_984);
  xor g1087 (n_1154, n_401, n_402);
  xor g1088 (n_405, n_1154, A[19]);
  nand g1089 (n_1155, n_401, n_402);
  nand g1090 (n_1156, A[19], n_402);
  nand g1091 (n_1157, n_401, A[19]);
  nand g1092 (n_424, n_1155, n_1156, n_1157);
  xor g1093 (n_1158, n_403, n_404);
  xor g1094 (n_407, n_1158, A[20]);
  nand g1095 (n_1159, n_403, n_404);
  nand g1096 (n_1160, A[20], n_404);
  nand g1097 (n_1161, n_403, A[20]);
  nand g1098 (n_425, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_405, n_406);
  xor g1100 (n_409, n_1162, n_407);
  nand g1101 (n_1163, n_405, n_406);
  nand g1102 (n_1164, n_407, n_406);
  nand g1103 (n_1165, n_405, n_407);
  nand g1104 (n_428, n_1163, n_1164, n_1165);
  xor g1106 (n_411, n_1166, n_408);
  nand g1108 (n_1168, n_408, A[23]);
  nand g1110 (n_430, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1123 (n_1178, A[8], n_413);
  xor g1124 (n_415, n_1178, A[9]);
  nand g1125 (n_1179, A[8], n_413);
  nand g1126 (n_1180, A[9], n_413);
  nand g1128 (n_435, n_1179, n_1180, n_687);
  xor g1129 (n_1182, n_414, n_415);
  xor g1130 (n_417, n_1182, n_416);
  nand g1131 (n_1183, n_414, n_415);
  nand g1132 (n_1184, n_416, n_415);
  nand g1133 (n_1185, n_414, n_416);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, A[12], A[13]);
  xor g1136 (n_420, n_1186, n_417);
  nand g1137 (n_1187, A[12], A[13]);
  nand g1138 (n_1188, n_417, A[13]);
  nand g1139 (n_1189, A[12], n_417);
  nand g1140 (n_439, n_1187, n_1188, n_1189);
  xor g1141 (n_1190, n_418, n_419);
  xor g1142 (n_422, n_1190, A[16]);
  nand g1143 (n_1191, n_418, n_419);
  nand g1144 (n_1192, A[16], n_419);
  nand g1145 (n_1193, n_418, A[16]);
  nand g1146 (n_440, n_1191, n_1192, n_1193);
  xor g1147 (n_1194, n_420, A[17]);
  xor g1148 (n_423, n_1194, n_421);
  nand g1149 (n_1195, n_420, A[17]);
  nand g1150 (n_1196, n_421, A[17]);
  nand g1151 (n_1197, n_420, n_421);
  nand g1152 (n_442, n_1195, n_1196, n_1197);
  xor g1153 (n_1198, n_422, A[20]);
  xor g1154 (n_426, n_1198, n_423);
  nand g1155 (n_1199, n_422, A[20]);
  nand g1156 (n_1200, n_423, A[20]);
  nand g1157 (n_1201, n_422, n_423);
  nand g1158 (n_445, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_424, A[21]);
  xor g1160 (n_427, n_1202, n_425);
  nand g1161 (n_1203, n_424, A[21]);
  nand g1162 (n_1204, n_425, A[21]);
  nand g1163 (n_1205, n_424, n_425);
  nand g1164 (n_447, n_1203, n_1204, n_1205);
  xor g1166 (n_429, n_1206, n_427);
  nand g1168 (n_1208, n_427, n_426);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, n_433);
  nand g1183 (n_1217, A[6], n_433);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, A[9], A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, A[9], A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, A[9], n_434);
  nand g1190 (n_455, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, n_435, n_436);
  xor g1192 (n_438, n_1222, A[13]);
  nand g1193 (n_1223, n_435, n_436);
  nand g1194 (n_1224, A[13], n_436);
  nand g1195 (n_1225, n_435, A[13]);
  nand g1196 (n_457, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, A[14], n_437);
  xor g1198 (n_441, n_1226, n_438);
  nand g1199 (n_1227, A[14], n_437);
  nand g1200 (n_1228, n_438, n_437);
  nand g1201 (n_1229, A[14], n_438);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, n_439, A[17]);
  xor g1204 (n_443, n_1230, n_440);
  nand g1205 (n_1231, n_439, A[17]);
  nand g1206 (n_1232, n_440, A[17]);
  nand g1207 (n_1233, n_439, n_440);
  nand g1208 (n_461, n_1231, n_1232, n_1233);
  xor g1209 (n_1234, A[18], n_441);
  xor g1210 (n_444, n_1234, n_442);
  nand g1211 (n_1235, A[18], n_441);
  nand g1212 (n_1236, n_442, n_441);
  nand g1213 (n_1237, A[18], n_442);
  nand g1214 (n_464, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_443, A[21]);
  xor g1216 (n_446, n_1238, A[22]);
  nand g1217 (n_1239, n_443, A[21]);
  nand g1219 (n_1241, n_443, A[22]);
  nand g1220 (n_465, n_1239, n_1077, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[5], A[7]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], n_453);
  xor g1242 (n_456, n_1254, n_454);
  nand g1243 (n_1255, A[10], n_453);
  nand g1244 (n_1256, n_454, n_453);
  nand g1245 (n_1257, A[10], n_454);
  nand g1246 (n_472, n_1255, n_1256, n_1257);
  xor g1247 (n_1258, A[11], n_455);
  xor g1248 (n_458, n_1258, n_456);
  nand g1249 (n_1259, A[11], n_455);
  nand g1250 (n_1260, n_456, n_455);
  nand g1251 (n_1261, A[11], n_456);
  nand g1252 (n_474, n_1259, n_1260, n_1261);
  xor g1253 (n_1262, A[14], n_457);
  xor g1254 (n_460, n_1262, A[15]);
  nand g1255 (n_1263, A[14], n_457);
  nand g1256 (n_1264, A[15], n_457);
  nand g1258 (n_476, n_1263, n_1264, n_1109);
  xor g1259 (n_1266, n_458, A[18]);
  xor g1260 (n_462, n_1266, n_459);
  nand g1261 (n_1267, n_458, A[18]);
  nand g1262 (n_1268, n_459, A[18]);
  nand g1263 (n_1269, n_458, n_459);
  nand g1264 (n_479, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, n_460, A[19]);
  xor g1266 (n_463, n_1270, n_461);
  nand g1267 (n_1271, n_460, A[19]);
  nand g1268 (n_1272, n_461, A[19]);
  nand g1269 (n_1273, n_460, n_461);
  nand g1270 (n_480, n_1271, n_1272, n_1273);
  xor g1271 (n_1274, n_462, A[22]);
  xor g1272 (n_466, n_1274, n_463);
  nand g1273 (n_1275, n_462, A[22]);
  nand g1274 (n_1276, n_463, A[22]);
  nand g1275 (n_1277, n_462, n_463);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1277 (n_1278, n_464, A[23]);
  xor g1278 (n_467, n_1278, n_465);
  nand g1279 (n_1279, n_464, A[23]);
  nand g1280 (n_1280, n_465, A[23]);
  nand g1281 (n_1281, n_464, n_465);
  nand g1282 (n_484, n_1279, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1289 (n_1286, A[7], A[6]);
  xor g1290 (n_471, n_1286, A[8]);
  nand g1292 (n_1288, A[8], A[6]);
  nand g1294 (n_486, n_661, n_1288, n_673);
  xor g1295 (n_1290, n_470, n_471);
  xor g1296 (n_473, n_1290, A[11]);
  nand g1297 (n_1291, n_470, n_471);
  nand g1298 (n_1292, A[11], n_471);
  nand g1299 (n_1293, n_470, A[11]);
  nand g1300 (n_488, n_1291, n_1292, n_1293);
  xor g1301 (n_1294, A[12], n_472);
  xor g1302 (n_475, n_1294, n_473);
  nand g1303 (n_1295, A[12], n_472);
  nand g1304 (n_1296, n_473, n_472);
  nand g1305 (n_1297, A[12], n_473);
  nand g1306 (n_489, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, A[15], n_474);
  xor g1308 (n_477, n_1298, n_475);
  nand g1309 (n_1299, A[15], n_474);
  nand g1310 (n_1300, n_475, n_474);
  nand g1311 (n_1301, A[15], n_475);
  nand g1312 (n_491, n_1299, n_1300, n_1301);
  xor g1313 (n_1302, A[16], n_476);
  xor g1314 (n_478, n_1302, n_477);
  nand g1315 (n_1303, A[16], n_476);
  nand g1316 (n_1304, n_477, n_476);
  nand g1317 (n_1305, A[16], n_477);
  nand g1318 (n_494, n_1303, n_1304, n_1305);
  xor g1319 (n_1306, A[19], n_478);
  xor g1320 (n_481, n_1306, n_479);
  nand g1321 (n_1307, A[19], n_478);
  nand g1322 (n_1308, n_479, n_478);
  nand g1323 (n_1309, A[19], n_479);
  nand g1324 (n_496, n_1307, n_1308, n_1309);
  xor g1325 (n_1310, A[20], n_480);
  xor g1326 (n_483, n_1310, n_481);
  nand g1327 (n_1311, A[20], n_480);
  nand g1328 (n_1312, n_481, n_480);
  nand g1329 (n_1313, A[20], n_481);
  nand g1330 (n_498, n_1311, n_1312, n_1313);
  xor g1332 (n_485, n_1166, n_482);
  nand g1335 (n_1317, A[23], n_482);
  nand g1336 (n_500, n_1167, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1344 (n_487, n_686, n_486);
  nand g1346 (n_1324, n_486, A[9]);
  nand g1347 (n_1325, A[8], n_486);
  nand g1348 (n_503, n_687, n_1324, n_1325);
  xor g1349 (n_1326, A[12], n_487);
  xor g1350 (n_490, n_1326, n_488);
  nand g1351 (n_1327, A[12], n_487);
  nand g1352 (n_1328, n_488, n_487);
  nand g1353 (n_1329, A[12], n_488);
  nand g1354 (n_505, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, A[13], n_489);
  xor g1356 (n_492, n_1330, n_490);
  nand g1357 (n_1331, A[13], n_489);
  nand g1358 (n_1332, n_490, n_489);
  nand g1359 (n_1333, A[13], n_490);
  nand g1360 (n_507, n_1331, n_1332, n_1333);
  xor g1361 (n_1334, A[16], A[17]);
  xor g1362 (n_493, n_1334, n_491);
  nand g1364 (n_1336, n_491, A[17]);
  nand g1365 (n_1337, A[16], n_491);
  nand g1366 (n_509, n_884, n_1336, n_1337);
  xor g1367 (n_1338, n_492, n_493);
  xor g1368 (n_495, n_1338, A[20]);
  nand g1369 (n_1339, n_492, n_493);
  nand g1370 (n_1340, A[20], n_493);
  nand g1371 (n_1341, n_492, A[20]);
  nand g1372 (n_511, n_1339, n_1340, n_1341);
  xor g1373 (n_1342, n_494, A[21]);
  xor g1374 (n_497, n_1342, n_495);
  nand g1375 (n_1343, n_494, A[21]);
  nand g1376 (n_1344, n_495, A[21]);
  nand g1377 (n_1345, n_494, n_495);
  nand g1378 (n_513, n_1343, n_1344, n_1345);
  xor g1380 (n_499, n_1346, n_497);
  nand g1383 (n_1349, n_496, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  nand g1397 (n_1357, A[10], n_503);
  nand g1398 (n_520, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], A[14]);
  xor g1400 (n_506, n_1358, n_504);
  nand g1401 (n_1359, A[13], A[14]);
  nand g1402 (n_1360, n_504, A[14]);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_521, n_1359, n_1360, n_1361);
  xor g1405 (n_1362, n_505, A[17]);
  xor g1406 (n_508, n_1362, n_506);
  nand g1407 (n_1363, n_505, A[17]);
  nand g1408 (n_1364, n_506, A[17]);
  nand g1409 (n_1365, n_505, n_506);
  nand g1410 (n_523, n_1363, n_1364, n_1365);
  xor g1411 (n_1366, n_507, A[18]);
  xor g1412 (n_510, n_1366, n_508);
  nand g1413 (n_1367, n_507, A[18]);
  nand g1414 (n_1368, n_508, A[18]);
  nand g1415 (n_1369, n_507, n_508);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_509, A[21]);
  xor g1418 (n_512, n_1370, n_510);
  nand g1419 (n_1371, n_509, A[21]);
  nand g1420 (n_1372, n_510, A[21]);
  nand g1421 (n_1373, n_509, n_510);
  nand g1422 (n_527, n_1371, n_1372, n_1373);
  xor g1423 (n_1374, A[22], n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, A[22], n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, A[22], n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1437 (n_1382, A[9], A[11]);
  nand g1439 (n_1383, A[9], A[11]);
  nand g1442 (n_532, n_1383, n_1384, n_1385);
  xor g1443 (n_1386, A[14], n_519);
  xor g1444 (n_522, n_1386, n_520);
  nand g1445 (n_1387, A[14], n_519);
  nand g1446 (n_1388, n_520, n_519);
  nand g1447 (n_1389, A[14], n_520);
  nand g1448 (n_534, n_1387, n_1388, n_1389);
  xor g1449 (n_1390, A[15], n_521);
  xor g1450 (n_524, n_1390, n_522);
  nand g1451 (n_1391, A[15], n_521);
  nand g1452 (n_1392, n_522, n_521);
  nand g1453 (n_1393, A[15], n_522);
  nand g1454 (n_536, n_1391, n_1392, n_1393);
  xor g1455 (n_1394, A[18], n_523);
  xor g1456 (n_525, n_1394, A[19]);
  nand g1457 (n_1395, A[18], n_523);
  nand g1458 (n_1396, A[19], n_523);
  nand g1459 (n_1397, A[18], A[19]);
  nand g1460 (n_538, n_1395, n_1396, n_1397);
  xor g1461 (n_1398, n_524, n_525);
  xor g1462 (n_528, n_1398, n_526);
  nand g1463 (n_1399, n_524, n_525);
  nand g1464 (n_1400, n_526, n_525);
  nand g1465 (n_1401, n_524, n_526);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1467 (n_1402, A[22], A[23]);
  xor g1468 (n_529, n_1402, n_527);
  nand g1469 (n_1403, A[22], A[23]);
  nand g1470 (n_1404, n_527, A[23]);
  nand g1471 (n_1405, A[22], n_527);
  nand g1472 (n_543, n_1403, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1480 (n_533, n_1098, A[12]);
  nand g1482 (n_1412, A[12], A[10]);
  nand g1483 (n_1413, A[11], A[12]);
  nand g1484 (n_544, n_1099, n_1412, n_1413);
  xor g1485 (n_1414, n_532, n_533);
  xor g1486 (n_535, n_1414, A[15]);
  nand g1487 (n_1415, n_532, n_533);
  nand g1488 (n_1416, A[15], n_533);
  nand g1489 (n_1417, n_532, A[15]);
  nand g1490 (n_546, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, A[16], n_534);
  xor g1492 (n_537, n_1418, n_535);
  nand g1493 (n_1419, A[16], n_534);
  nand g1494 (n_1420, n_535, n_534);
  nand g1495 (n_1421, A[16], n_535);
  nand g1496 (n_547, n_1419, n_1420, n_1421);
  xor g1497 (n_1422, A[19], n_536);
  xor g1498 (n_539, n_1422, n_537);
  nand g1499 (n_1423, A[19], n_536);
  nand g1500 (n_1424, n_537, n_536);
  nand g1501 (n_1425, A[19], n_537);
  nand g1502 (n_549, n_1423, n_1424, n_1425);
  xor g1503 (n_1426, A[20], n_538);
  xor g1504 (n_541, n_1426, n_539);
  nand g1505 (n_1427, A[20], n_538);
  nand g1506 (n_1428, n_539, n_538);
  nand g1507 (n_1429, A[20], n_539);
  nand g1508 (n_552, n_1427, n_1428, n_1429);
  xor g1510 (n_542, n_1166, n_540);
  nand g1513 (n_1433, A[23], n_540);
  nand g1514 (n_554, n_1167, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1522 (n_545, n_1186, n_544);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_1187, n_1440, n_1441);
  xor g1528 (n_548, n_1334, n_545);
  nand g1530 (n_1444, n_545, A[17]);
  nand g1531 (n_1445, A[16], n_545);
  nand g1532 (n_558, n_884, n_1444, n_1445);
  xor g1533 (n_1446, n_546, n_547);
  xor g1534 (n_550, n_1446, n_548);
  nand g1535 (n_1447, n_546, n_547);
  nand g1536 (n_1448, n_548, n_547);
  nand g1537 (n_1449, n_546, n_548);
  nand g1538 (n_561, n_1447, n_1448, n_1449);
  xor g1539 (n_1450, A[20], A[21]);
  xor g1540 (n_551, n_1450, n_549);
  nand g1541 (n_1451, A[20], A[21]);
  nand g1542 (n_1452, n_549, A[21]);
  nand g1543 (n_1453, A[20], n_549);
  nand g1544 (n_562, n_1451, n_1452, n_1453);
  xor g1546 (n_553, n_1454, n_551);
  nand g1549 (n_1457, n_550, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1563 (n_1465, A[14], A[17]);
  nand g1564 (n_570, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, n_557, A[18]);
  xor g1566 (n_560, n_1466, n_558);
  nand g1567 (n_1467, n_557, A[18]);
  nand g1568 (n_1468, n_558, A[18]);
  nand g1569 (n_1469, n_557, n_558);
  nand g1570 (n_571, n_1467, n_1468, n_1469);
  xor g1571 (n_1470, n_559, n_560);
  xor g1572 (n_563, n_1470, A[21]);
  nand g1573 (n_1471, n_559, n_560);
  nand g1574 (n_1472, A[21], n_560);
  nand g1575 (n_1473, n_559, A[21]);
  nand g1576 (n_573, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, n_561, A[22]);
  xor g1578 (n_564, n_1474, n_562);
  nand g1579 (n_1475, n_561, A[22]);
  nand g1580 (n_1476, n_562, A[22]);
  nand g1581 (n_1477, n_561, n_562);
  nand g1582 (n_576, n_1475, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  xor g1591 (n_1482, A[13], A[15]);
  nand g1596 (n_578, n_773, n_1484, n_1485);
  xor g1597 (n_1486, A[18], n_569);
  xor g1598 (n_572, n_1486, A[19]);
  nand g1599 (n_1487, A[18], n_569);
  nand g1600 (n_1488, A[19], n_569);
  nand g1602 (n_580, n_1487, n_1488, n_1397);
  xor g1603 (n_1490, n_570, n_571);
  xor g1604 (n_574, n_1490, n_572);
  nand g1605 (n_1491, n_570, n_571);
  nand g1606 (n_1492, n_572, n_571);
  nand g1607 (n_1493, n_570, n_572);
  nand g1608 (n_582, n_1491, n_1492, n_1493);
  xor g1610 (n_575, n_1402, n_573);
  nand g1612 (n_1496, n_573, A[23]);
  nand g1613 (n_1497, A[22], n_573);
  nand g1614 (n_584, n_1403, n_1496, n_1497);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1621 (n_1502, A[15], A[14]);
  xor g1622 (n_579, n_1502, A[16]);
  nand g1626 (n_586, n_1109, n_801, n_984);
  xor g1627 (n_1506, n_578, n_579);
  xor g1628 (n_581, n_1506, A[19]);
  nand g1629 (n_1507, n_578, n_579);
  nand g1630 (n_1508, A[19], n_579);
  nand g1631 (n_1509, n_578, A[19]);
  nand g1632 (n_588, n_1507, n_1508, n_1509);
  xor g1633 (n_1510, A[20], n_580);
  xor g1634 (n_583, n_1510, n_581);
  nand g1635 (n_1511, A[20], n_580);
  nand g1636 (n_1512, n_581, n_580);
  nand g1637 (n_1513, A[20], n_581);
  nand g1638 (n_589, n_1511, n_1512, n_1513);
  xor g1639 (n_1514, A[23], n_582);
  nand g1641 (n_1515, A[23], n_582);
  nand g1644 (n_591, n_1515, n_1516, n_1167);
  xor g1645 (n_1518, n_583, n_584);
  xor g1646 (n_83, n_1518, n_585);
  nand g1647 (n_1519, n_583, n_584);
  nand g1648 (n_1520, n_585, n_584);
  nand g1649 (n_1521, n_583, n_585);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1652 (n_587, n_1334, n_586);
  nand g1654 (n_1524, n_586, A[17]);
  nand g1655 (n_1525, A[16], n_586);
  nand g1656 (n_595, n_884, n_1524, n_1525);
  xor g1657 (n_1526, A[20], n_587);
  xor g1658 (n_590, n_1526, n_588);
  nand g1659 (n_1527, A[20], n_587);
  nand g1660 (n_1528, n_588, n_587);
  nand g1661 (n_1529, A[20], n_588);
  nand g1662 (n_597, n_1527, n_1528, n_1529);
  xor g1664 (n_592, n_1530, n_589);
  nand g1667 (n_1533, A[21], n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_81, n_1535, n_1536, n_1537);
  xor g1678 (n_596, n_1538, n_595);
  nand g1681 (n_1541, A[18], n_595);
  nand g1682 (n_604, n_1539, n_1540, n_1541);
  xor g1683 (n_1542, A[21], A[22]);
  xor g1684 (n_598, n_1542, n_596);
  nand g1686 (n_1544, n_596, A[22]);
  nand g1687 (n_1545, A[21], n_596);
  nand g1688 (n_606, n_1077, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_33, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[17], A[19]);
  nand g1699 (n_1551, A[17], A[19]);
  nand g1702 (n_608, n_1551, n_1552, n_1553);
  xor g1703 (n_1554, A[22], n_603);
  xor g1704 (n_605, n_1554, n_604);
  nand g1705 (n_1555, A[22], n_603);
  nand g1706 (n_1556, n_604, n_603);
  nand g1707 (n_1557, A[22], n_604);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, A[23], n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, A[23], n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, A[23], n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1715 (n_1562, A[19], A[18]);
  xor g1716 (n_609, n_1562, A[20]);
  nand g1719 (n_1565, A[19], A[20]);
  nand g1720 (n_612, n_1397, n_925, n_1565);
  xor g1721 (n_1566, n_608, n_609);
  xor g1722 (n_611, n_1566, A[23]);
  nand g1723 (n_1567, n_608, n_609);
  nand g1724 (n_1568, A[23], n_609);
  nand g1725 (n_1569, n_608, A[23]);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1728 (n_79, n_1570, n_611);
  nand g1730 (n_1572, n_611, n_610);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1734 (n_613, n_1450, n_612);
  nand g1736 (n_1576, n_612, A[21]);
  nand g1737 (n_1577, A[20], n_612);
  nand g1738 (n_617, n_1451, n_1576, n_1577);
  xor g1740 (n_78, n_1578, n_614);
  nand g1742 (n_1580, n_614, n_613);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_617);
  nand g1752 (n_76, n_1583, n_1584, n_1585);
  nand g1759 (n_1589, A[21], A[23]);
  nand g1760 (n_27, n_1587, n_1588, n_1589);
  xor g1762 (n_75, n_1166, A[22]);
  nand g1766 (n_74, n_1167, n_1403, n_1593);
  nand g16 (n_1606, A[0], A[2]);
  xor g20 (Z[2], A[0], A[2]);
  nand g22 (n_1611, n_68, A[3]);
  nand g25 (n_1615, n_1611, n_1612, n_1613);
  xor g26 (n_1614, n_68, A[3]);
  nand g28 (n_1616, A[4], n_117);
  nand g29 (n_1617, A[4], n_1615);
  nand g30 (n_1618, n_117, n_1615);
  nand g31 (n_1620, n_1616, n_1617, n_1618);
  xor g32 (n_1619, A[4], n_117);
  xor g33 (Z[4], n_1615, n_1619);
  nand g34 (n_1621, A[5], n_116);
  nand g35 (n_1622, A[5], n_1620);
  nand g36 (n_1623, n_116, n_1620);
  nand g37 (n_1625, n_1621, n_1622, n_1623);
  xor g38 (n_1624, A[5], n_116);
  xor g39 (Z[5], n_1620, n_1624);
  nand g40 (n_1626, n_67, n_115);
  nand g41 (n_1627, n_67, n_1625);
  nand g42 (n_1628, n_115, n_1625);
  nand g43 (n_1630, n_1626, n_1627, n_1628);
  xor g44 (n_1629, n_67, n_115);
  xor g45 (Z[6], n_1625, n_1629);
  nand g46 (n_1631, n_66, n_114);
  nand g47 (n_1632, n_66, n_1630);
  nand g48 (n_1633, n_114, n_1630);
  nand g49 (n_1635, n_1631, n_1632, n_1633);
  xor g50 (n_1634, n_66, n_114);
  xor g51 (Z[7], n_1630, n_1634);
  nand g52 (n_1636, n_65, n_113);
  nand g53 (n_1637, n_65, n_1635);
  nand g54 (n_1638, n_113, n_1635);
  nand g55 (n_1640, n_1636, n_1637, n_1638);
  xor g56 (n_1639, n_65, n_113);
  xor g57 (Z[8], n_1635, n_1639);
  nand g58 (n_1641, n_64, n_112);
  nand g59 (n_1642, n_64, n_1640);
  nand g60 (n_1643, n_112, n_1640);
  nand g61 (n_1645, n_1641, n_1642, n_1643);
  xor g62 (n_1644, n_64, n_112);
  xor g63 (Z[9], n_1640, n_1644);
  nand g64 (n_1646, n_63, n_111);
  nand g65 (n_1647, n_63, n_1645);
  nand g66 (n_1648, n_111, n_1645);
  nand g67 (n_1650, n_1646, n_1647, n_1648);
  xor g68 (n_1649, n_63, n_111);
  xor g69 (Z[10], n_1645, n_1649);
  nand g70 (n_1651, n_62, n_110);
  nand g71 (n_1652, n_62, n_1650);
  nand g72 (n_1653, n_110, n_1650);
  nand g73 (n_1655, n_1651, n_1652, n_1653);
  xor g74 (n_1654, n_62, n_110);
  xor g75 (Z[11], n_1650, n_1654);
  nand g76 (n_1656, n_61, n_109);
  nand g77 (n_1657, n_61, n_1655);
  nand g78 (n_1658, n_109, n_1655);
  nand g79 (n_1660, n_1656, n_1657, n_1658);
  xor g80 (n_1659, n_61, n_109);
  xor g81 (Z[12], n_1655, n_1659);
  nand g82 (n_1661, n_60, n_108);
  nand g83 (n_1662, n_60, n_1660);
  nand g84 (n_1663, n_108, n_1660);
  nand g85 (n_1665, n_1661, n_1662, n_1663);
  xor g86 (n_1664, n_60, n_108);
  xor g87 (Z[13], n_1660, n_1664);
  nand g88 (n_1666, n_59, n_107);
  nand g89 (n_1667, n_59, n_1665);
  nand g90 (n_1668, n_107, n_1665);
  nand g91 (n_1670, n_1666, n_1667, n_1668);
  xor g92 (n_1669, n_59, n_107);
  xor g93 (Z[14], n_1665, n_1669);
  nand g94 (n_1671, n_58, n_106);
  nand g95 (n_1672, n_58, n_1670);
  nand g96 (n_1673, n_106, n_1670);
  nand g97 (n_1675, n_1671, n_1672, n_1673);
  xor g98 (n_1674, n_58, n_106);
  xor g99 (Z[15], n_1670, n_1674);
  nand g100 (n_1676, n_57, n_105);
  nand g101 (n_1677, n_57, n_1675);
  nand g102 (n_1678, n_105, n_1675);
  nand g103 (n_1680, n_1676, n_1677, n_1678);
  xor g104 (n_1679, n_57, n_105);
  xor g105 (Z[16], n_1675, n_1679);
  nand g106 (n_1681, n_56, n_104);
  nand g107 (n_1682, n_56, n_1680);
  nand g108 (n_1683, n_104, n_1680);
  nand g109 (n_1685, n_1681, n_1682, n_1683);
  xor g110 (n_1684, n_56, n_104);
  xor g111 (Z[17], n_1680, n_1684);
  nand g112 (n_1686, n_55, n_103);
  nand g113 (n_1687, n_55, n_1685);
  nand g114 (n_1688, n_103, n_1685);
  nand g115 (n_1690, n_1686, n_1687, n_1688);
  xor g116 (n_1689, n_55, n_103);
  xor g117 (Z[18], n_1685, n_1689);
  nand g118 (n_1691, n_54, n_102);
  nand g119 (n_1692, n_54, n_1690);
  nand g120 (n_1693, n_102, n_1690);
  nand g121 (n_1695, n_1691, n_1692, n_1693);
  xor g122 (n_1694, n_54, n_102);
  xor g123 (Z[19], n_1690, n_1694);
  nand g124 (n_1696, n_53, n_101);
  nand g125 (n_1697, n_53, n_1695);
  nand g126 (n_1698, n_101, n_1695);
  nand g127 (n_1700, n_1696, n_1697, n_1698);
  xor g128 (n_1699, n_53, n_101);
  xor g129 (Z[20], n_1695, n_1699);
  nand g130 (n_1701, n_52, n_100);
  nand g131 (n_1702, n_52, n_1700);
  nand g132 (n_1703, n_100, n_1700);
  nand g133 (n_1705, n_1701, n_1702, n_1703);
  xor g134 (n_1704, n_52, n_100);
  xor g135 (Z[21], n_1700, n_1704);
  nand g136 (n_1706, n_51, n_99);
  nand g137 (n_1707, n_51, n_1705);
  nand g138 (n_1708, n_99, n_1705);
  nand g139 (n_1710, n_1706, n_1707, n_1708);
  xor g140 (n_1709, n_51, n_99);
  xor g141 (Z[22], n_1705, n_1709);
  nand g142 (n_1711, n_50, n_98);
  nand g143 (n_1712, n_50, n_1710);
  nand g144 (n_1713, n_98, n_1710);
  nand g145 (n_1715, n_1711, n_1712, n_1713);
  xor g146 (n_1714, n_50, n_98);
  xor g147 (Z[23], n_1710, n_1714);
  nand g148 (n_1716, n_49, n_97);
  nand g149 (n_1717, n_49, n_1715);
  nand g150 (n_1718, n_97, n_1715);
  nand g151 (n_1720, n_1716, n_1717, n_1718);
  xor g152 (n_1719, n_49, n_97);
  xor g153 (Z[24], n_1715, n_1719);
  nand g154 (n_1721, n_48, n_96);
  nand g155 (n_1722, n_48, n_1720);
  nand g156 (n_1723, n_96, n_1720);
  nand g157 (n_1725, n_1721, n_1722, n_1723);
  xor g158 (n_1724, n_48, n_96);
  xor g159 (Z[25], n_1720, n_1724);
  nand g160 (n_1726, n_47, n_95);
  nand g161 (n_1727, n_47, n_1725);
  nand g162 (n_1728, n_95, n_1725);
  nand g163 (n_1730, n_1726, n_1727, n_1728);
  xor g164 (n_1729, n_47, n_95);
  xor g165 (Z[26], n_1725, n_1729);
  nand g166 (n_1731, n_46, n_94);
  nand g167 (n_1732, n_46, n_1730);
  nand g168 (n_1733, n_94, n_1730);
  nand g169 (n_1735, n_1731, n_1732, n_1733);
  xor g170 (n_1734, n_46, n_94);
  xor g171 (Z[27], n_1730, n_1734);
  nand g172 (n_1736, n_45, n_93);
  nand g173 (n_1737, n_45, n_1735);
  nand g174 (n_1738, n_93, n_1735);
  nand g175 (n_1740, n_1736, n_1737, n_1738);
  xor g176 (n_1739, n_45, n_93);
  xor g177 (Z[28], n_1735, n_1739);
  nand g178 (n_1741, n_44, n_92);
  nand g179 (n_1742, n_44, n_1740);
  nand g180 (n_1743, n_92, n_1740);
  nand g181 (n_1745, n_1741, n_1742, n_1743);
  xor g182 (n_1744, n_44, n_92);
  xor g183 (Z[29], n_1740, n_1744);
  nand g184 (n_1746, n_43, n_91);
  nand g185 (n_1747, n_43, n_1745);
  nand g186 (n_1748, n_91, n_1745);
  nand g187 (n_1750, n_1746, n_1747, n_1748);
  xor g188 (n_1749, n_43, n_91);
  xor g189 (Z[30], n_1745, n_1749);
  nand g190 (n_1751, n_42, n_90);
  nand g191 (n_1752, n_42, n_1750);
  nand g192 (n_1753, n_90, n_1750);
  nand g193 (n_1755, n_1751, n_1752, n_1753);
  xor g194 (n_1754, n_42, n_90);
  xor g195 (Z[31], n_1750, n_1754);
  nand g196 (n_1756, n_41, n_89);
  nand g197 (n_1757, n_41, n_1755);
  nand g198 (n_1758, n_89, n_1755);
  nand g199 (n_1760, n_1756, n_1757, n_1758);
  xor g200 (n_1759, n_41, n_89);
  xor g201 (Z[32], n_1755, n_1759);
  nand g202 (n_1761, n_40, n_88);
  nand g203 (n_1762, n_40, n_1760);
  nand g204 (n_1763, n_88, n_1760);
  nand g205 (n_1765, n_1761, n_1762, n_1763);
  xor g206 (n_1764, n_40, n_88);
  xor g207 (Z[33], n_1760, n_1764);
  nand g208 (n_1766, n_39, n_87);
  nand g209 (n_1767, n_39, n_1765);
  nand g210 (n_1768, n_87, n_1765);
  nand g211 (n_1770, n_1766, n_1767, n_1768);
  xor g212 (n_1769, n_39, n_87);
  xor g213 (Z[34], n_1765, n_1769);
  nand g214 (n_1771, n_38, n_86);
  nand g215 (n_1772, n_38, n_1770);
  nand g216 (n_1773, n_86, n_1770);
  nand g217 (n_1775, n_1771, n_1772, n_1773);
  xor g218 (n_1774, n_38, n_86);
  xor g219 (Z[35], n_1770, n_1774);
  nand g220 (n_1776, n_37, n_85);
  nand g221 (n_1777, n_37, n_1775);
  nand g222 (n_1778, n_85, n_1775);
  nand g223 (n_1780, n_1776, n_1777, n_1778);
  xor g224 (n_1779, n_37, n_85);
  xor g225 (Z[36], n_1775, n_1779);
  nand g226 (n_1781, n_36, n_84);
  nand g227 (n_1782, n_36, n_1780);
  nand g228 (n_1783, n_84, n_1780);
  nand g229 (n_1785, n_1781, n_1782, n_1783);
  xor g230 (n_1784, n_36, n_84);
  xor g231 (Z[37], n_1780, n_1784);
  nand g232 (n_1786, n_35, n_83);
  nand g233 (n_1787, n_35, n_1785);
  nand g234 (n_1788, n_83, n_1785);
  nand g235 (n_1790, n_1786, n_1787, n_1788);
  xor g236 (n_1789, n_35, n_83);
  xor g237 (Z[38], n_1785, n_1789);
  nand g238 (n_1791, n_34, n_82);
  nand g239 (n_1792, n_34, n_1790);
  nand g240 (n_1793, n_82, n_1790);
  nand g241 (n_1795, n_1791, n_1792, n_1793);
  xor g242 (n_1794, n_34, n_82);
  xor g243 (Z[39], n_1790, n_1794);
  nand g244 (n_1796, n_33, n_81);
  nand g245 (n_1797, n_33, n_1795);
  nand g246 (n_1798, n_81, n_1795);
  nand g247 (n_1800, n_1796, n_1797, n_1798);
  xor g248 (n_1799, n_33, n_81);
  xor g249 (Z[40], n_1795, n_1799);
  nand g250 (n_1801, n_32, n_80);
  nand g251 (n_1802, n_32, n_1800);
  nand g252 (n_1803, n_80, n_1800);
  nand g253 (n_1805, n_1801, n_1802, n_1803);
  xor g254 (n_1804, n_32, n_80);
  xor g255 (Z[41], n_1800, n_1804);
  nand g256 (n_1806, n_31, n_79);
  nand g257 (n_1807, n_31, n_1805);
  nand g258 (n_1808, n_79, n_1805);
  nand g259 (n_1810, n_1806, n_1807, n_1808);
  xor g260 (n_1809, n_31, n_79);
  xor g261 (Z[42], n_1805, n_1809);
  nand g262 (n_1811, n_30, n_78);
  nand g263 (n_1812, n_30, n_1810);
  nand g264 (n_1813, n_78, n_1810);
  nand g265 (n_1815, n_1811, n_1812, n_1813);
  xor g266 (n_1814, n_30, n_78);
  xor g267 (Z[43], n_1810, n_1814);
  nand g1772 (n_1816, n_29, n_77);
  nand g1773 (n_1817, n_29, n_1815);
  nand g1774 (n_1818, n_77, n_1815);
  nand g1775 (n_1820, n_1816, n_1817, n_1818);
  xor g1776 (n_1819, n_29, n_77);
  xor g1777 (Z[44], n_1815, n_1819);
  nand g1778 (n_1821, n_28, n_76);
  nand g1779 (n_1822, n_28, n_1820);
  nand g1780 (n_1823, n_76, n_1820);
  nand g1781 (n_1825, n_1821, n_1822, n_1823);
  xor g1782 (n_1824, n_28, n_76);
  xor g1783 (Z[45], n_1820, n_1824);
  nand g1784 (n_1826, n_27, n_75);
  nand g1785 (n_1827, n_27, n_1825);
  nand g1786 (n_1828, n_75, n_1825);
  nand g1787 (n_1830, n_1826, n_1827, n_1828);
  xor g1788 (n_1829, n_27, n_75);
  xor g1789 (Z[46], n_1825, n_1829);
  xor g1791 (Z[47], n_1830, n_1831);
  or g1804 (n_1043, A[1], wc);
  not gc (wc, n_171);
  or g1805 (n_1044, A[1], wc0);
  not gc0 (wc0, A[2]);
  xnor g1807 (n_1166, A[24], A[23]);
  or g1808 (n_1167, wc1, A[24]);
  not gc1 (wc1, A[23]);
  xnor g1809 (n_1214, A[6], A[5]);
  or g1810 (n_1215, A[5], wc2);
  not gc2 (wc2, A[6]);
  or g1811 (n_1252, A[6], wc3);
  not gc3 (wc3, A[7]);
  or g1812 (n_1253, wc4, A[6]);
  not gc4 (wc4, A[5]);
  or g1814 (n_1355, A[9], wc5);
  not gc5 (wc5, A[10]);
  or g1815 (n_1384, A[10], wc6);
  not gc6 (wc6, A[11]);
  or g1816 (n_1385, wc7, A[10]);
  not gc7 (wc7, A[9]);
  or g1818 (n_1463, A[13], wc8);
  not gc8 (wc8, A[14]);
  or g1819 (n_1464, A[13], wc9);
  not gc9 (wc9, A[17]);
  or g1820 (n_1484, A[14], wc10);
  not gc10 (wc10, A[15]);
  or g1821 (n_1485, wc11, A[14]);
  not gc11 (wc11, A[13]);
  xnor g1822 (n_1530, A[24], A[21]);
  or g1823 (n_1531, wc12, A[24]);
  not gc12 (wc12, A[21]);
  xnor g1824 (n_1538, A[18], A[17]);
  or g1825 (n_1539, A[17], wc13);
  not gc13 (wc13, A[18]);
  or g1826 (n_1552, A[18], wc14);
  not gc14 (wc14, A[19]);
  or g1827 (n_1553, wc15, A[18]);
  not gc15 (wc15, A[17]);
  or g1829 (n_1583, A[21], wc16);
  not gc16 (wc16, A[22]);
  or g1830 (n_1587, wc17, A[22]);
  not gc17 (wc17, A[21]);
  or g1831 (n_1588, A[22], wc18);
  not gc18 (wc18, A[23]);
  or g1832 (n_1593, wc19, A[24]);
  not gc19 (wc19, A[22]);
  xnor g1834 (n_1086, A[2], A[1]);
  or g1835 (n_1088, A[1], wc20);
  not gc20 (wc20, A[3]);
  xnor g1836 (n_453, n_1250, A[6]);
  xnor g1837 (n_519, n_1382, A[10]);
  xnor g1838 (n_559, n_1358, A[17]);
  xnor g1839 (n_569, n_1482, A[14]);
  xnor g1840 (n_603, n_1550, A[18]);
  xnor g1841 (n_28, n_1542, A[23]);
  or g1843 (n_1047, wc21, n_117);
  not gc21 (wc21, A[5]);
  or g1844 (n_1049, wc22, n_117);
  not gc22 (wc22, A[6]);
  xnor g1846 (n_1578, n_613, A[24]);
  or g1847 (n_1579, A[24], wc23);
  not gc23 (wc23, n_613);
  xnor g1848 (n_1831, n_74, A[24]);
  or g1850 (n_1051, n_180, wc24);
  not gc24 (wc24, n_179);
  or g1851 (n_1052, wc25, n_180);
  not gc25 (wc25, A[9]);
  xnor g1852 (n_504, n_1218, n_503);
  or g1853 (n_1356, A[9], wc26);
  not gc26 (wc26, n_503);
  or g1854 (n_1540, A[17], wc27);
  not gc27 (wc27, n_595);
  or g1855 (n_1573, A[24], wc28);
  not gc28 (wc28, n_611);
  or g1856 (n_1581, A[24], wc29);
  not gc29 (wc29, n_614);
  xnor g1857 (n_29, n_1542, n_617);
  or g1858 (n_1584, A[21], wc30);
  not gc30 (wc30, n_617);
  or g1861 (n_1216, A[5], wc31);
  not gc31 (wc31, n_433);
  or g1862 (n_1612, n_1606, wc32);
  not gc32 (wc32, n_68);
  or g1863 (n_1613, wc33, n_1606);
  not gc33 (wc33, A[3]);
  xnor g1864 (Z[3], n_1606, n_1614);
  or g1866 (n_1056, wc34, n_202);
  not gc34 (wc34, A[10]);
  or g1867 (n_1057, wc35, n_202);
  not gc35 (wc35, n_282);
  or g1868 (n_1532, A[24], wc36);
  not gc36 (wc36, n_589);
  or g1869 (n_1060, wc37, n_285);
  not gc37 (wc37, A[13]);
  xnor g1870 (n_1570, n_610, A[24]);
  or g1871 (n_1571, A[24], wc38);
  not gc38 (wc38, n_610);
  or g1872 (n_1061, wc39, n_285);
  not gc39 (wc39, n_354);
  or g1873 (n_1516, A[24], wc40);
  not gc40 (wc40, n_582);
  xnor g1874 (n_357, n_285, n_1058);
  xnor g1875 (n_585, n_1514, A[24]);
  xnor g1876 (n_1454, n_550, A[24]);
  or g1877 (n_1455, A[24], wc41);
  not gc41 (wc41, n_550);
  or g1878 (n_1456, A[24], wc42);
  not gc42 (wc42, n_551);
  xnor g1879 (n_1078, n_363, A[24]);
  or g1880 (n_1079, A[24], wc43);
  not gc43 (wc43, n_363);
  or g1881 (n_1080, A[24], wc44);
  not gc44 (wc44, n_364);
  xnor g1882 (n_1206, n_426, A[24]);
  or g1883 (n_1207, A[24], wc45);
  not gc45 (wc45, n_426);
  xnor g1884 (n_1346, n_496, A[24]);
  or g1885 (n_1347, A[24], wc46);
  not gc46 (wc46, n_496);
  or g1886 (n_1169, A[24], wc47);
  not gc47 (wc47, n_408);
  or g1887 (n_1348, A[24], wc48);
  not gc48 (wc48, n_497);
  or g1888 (n_1432, A[24], wc49);
  not gc49 (wc49, n_540);
  or g1889 (n_1209, A[24], wc50);
  not gc50 (wc50, n_427);
  or g1890 (n_1316, A[24], wc51);
  not gc51 (wc51, n_482);
endmodule

module mult_signed_const_5220_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_5220_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_5487_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_176;
  wire n_179, n_180, n_183, n_184, n_187, n_188, n_189, n_195;
  wire n_196, n_201, n_202, n_203, n_204, n_209, n_210, n_211;
  wire n_212, n_217, n_218, n_219, n_220, n_221, n_223, n_224;
  wire n_225, n_226, n_227, n_232, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_246, n_248, n_249, n_250, n_251, n_261;
  wire n_262, n_265, n_267, n_269, n_271, n_273, n_274, n_275;
  wire n_276, n_277, n_281, n_282, n_283, n_284, n_285, n_286;
  wire n_287, n_288, n_289, n_290, n_291, n_292, n_293, n_296;
  wire n_298, n_299, n_300, n_301, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_315, n_317, n_318, n_319;
  wire n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_333;
  wire n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342;
  wire n_343, n_344, n_345, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_371, n_372, n_373, n_374, n_375, n_376, n_377;
  wire n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385;
  wire n_386, n_387, n_388, n_389, n_390, n_392, n_393, n_394;
  wire n_395, n_396, n_397, n_398, n_399, n_400, n_401, n_402;
  wire n_403, n_404, n_405, n_406, n_407, n_408, n_409, n_410;
  wire n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418;
  wire n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426;
  wire n_427, n_428, n_429, n_430, n_433, n_434, n_435, n_436;
  wire n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444;
  wire n_445, n_446, n_447, n_448, n_449, n_453, n_454, n_455;
  wire n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463;
  wire n_464, n_465, n_466, n_467, n_468, n_470, n_471, n_472;
  wire n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480;
  wire n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488;
  wire n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496;
  wire n_497, n_498, n_499, n_500, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_519, n_520, n_521, n_522, n_523, n_524, n_525;
  wire n_526, n_527, n_528, n_529, n_530, n_532, n_533, n_534;
  wire n_535, n_536, n_537, n_538, n_539, n_540, n_541, n_542;
  wire n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550;
  wire n_551, n_552, n_553, n_554, n_557, n_558, n_559, n_560;
  wire n_561, n_562, n_563, n_564, n_565, n_569, n_570, n_571;
  wire n_572, n_573, n_574, n_575, n_576, n_578, n_579, n_580;
  wire n_581, n_582, n_583, n_584, n_585, n_586, n_587, n_588;
  wire n_589, n_590, n_591, n_592, n_595, n_596, n_597, n_598;
  wire n_599, n_603, n_604, n_605, n_606, n_608, n_609, n_610;
  wire n_611, n_612, n_613, n_614, n_617, n_622, n_623, n_624;
  wire n_625, n_626, n_627, n_628, n_629, n_630, n_631, n_632;
  wire n_633, n_634, n_635, n_636, n_637, n_638, n_639, n_640;
  wire n_641, n_646, n_647, n_648, n_649, n_650, n_651, n_652;
  wire n_653, n_658, n_659, n_660, n_661, n_662, n_663, n_664;
  wire n_665, n_668, n_669, n_670, n_671, n_672, n_673, n_674;
  wire n_675, n_676, n_677, n_684, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_691, n_692, n_693, n_704, n_705, n_706;
  wire n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_724;
  wire n_725, n_726, n_727, n_728, n_729, n_730, n_731, n_732;
  wire n_733, n_738, n_742, n_743, n_744, n_745, n_746, n_747;
  wire n_748, n_749, n_750, n_751, n_752, n_753, n_760, n_761;
  wire n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769;
  wire n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777;
  wire n_790, n_791, n_792, n_794, n_795, n_796, n_797, n_798;
  wire n_799, n_800, n_801, n_802, n_803, n_804, n_805, n_822;
  wire n_823, n_824, n_825, n_826, n_827, n_828, n_829, n_830;
  wire n_831, n_832, n_833, n_850, n_851, n_852, n_854, n_855;
  wire n_856, n_857, n_858, n_859, n_860, n_861, n_862, n_866;
  wire n_867, n_868, n_872, n_873, n_876, n_877, n_878, n_879;
  wire n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887;
  wire n_888, n_889, n_890, n_891, n_892, n_893, n_900, n_901;
  wire n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909;
  wire n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917;
  wire n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925;
  wire n_926, n_927, n_928, n_929, n_938, n_939, n_941, n_942;
  wire n_943, n_944, n_945, n_946, n_947, n_948, n_949, n_950;
  wire n_951, n_952, n_953, n_954, n_955, n_956, n_957, n_958;
  wire n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_978;
  wire n_979, n_980, n_982, n_983, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_996, n_997, n_998, n_999, n_1000, n_1001, n_1013, n_1014;
  wire n_1015, n_1016, n_1017, n_1020, n_1021, n_1022, n_1023, n_1024;
  wire n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040;
  wire n_1041, n_1043, n_1044, n_1047, n_1049, n_1051, n_1052, n_1056;
  wire n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064;
  wire n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072;
  wire n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080;
  wire n_1081, n_1082, n_1083, n_1084, n_1085, n_1088, n_1090, n_1091;
  wire n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099;
  wire n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107;
  wire n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115;
  wire n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123;
  wire n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131;
  wire n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139;
  wire n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147;
  wire n_1148, n_1149, n_1150, n_1151, n_1152, n_1154, n_1155, n_1156;
  wire n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164;
  wire n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172;
  wire n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180;
  wire n_1182, n_1183, n_1184, n_1185, n_1186, n_1188, n_1189, n_1190;
  wire n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198;
  wire n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206;
  wire n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214;
  wire n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222;
  wire n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230;
  wire n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238;
  wire n_1239, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247;
  wire n_1248, n_1249, n_1250, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1266;
  wire n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274;
  wire n_1275, n_1276, n_1277, n_1280, n_1281, n_1282, n_1283, n_1284;
  wire n_1285, n_1286, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295;
  wire n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303;
  wire n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311;
  wire n_1312, n_1313, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321;
  wire n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331;
  wire n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339;
  wire n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347;
  wire n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1355, n_1356;
  wire n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364;
  wire n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381;
  wire n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
  wire n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397;
  wire n_1398, n_1399, n_1400, n_1401, n_1404, n_1405, n_1406, n_1407;
  wire n_1408, n_1409, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417;
  wire n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1426;
  wire n_1427, n_1428, n_1429, n_1432, n_1433, n_1434, n_1435, n_1436;
  wire n_1437, n_1440, n_1441, n_1442, n_1443, n_1444, n_1446, n_1447;
  wire n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455;
  wire n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1463, n_1464;
  wire n_1465, n_1466, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473;
  wire n_1474, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1484;
  wire n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493;
  wire n_1494, n_1495, n_1496, n_1498, n_1499, n_1500, n_1501, n_1502;
  wire n_1504, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512;
  wire n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520;
  wire n_1521, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530;
  wire n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1539;
  wire n_1540, n_1541, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558;
  wire n_1559, n_1560, n_1561, n_1562, n_1566, n_1567, n_1568, n_1569;
  wire n_1570, n_1571, n_1572, n_1573, n_1576, n_1577, n_1578, n_1579;
  wire n_1580, n_1581, n_1583, n_1584, n_1585, n_1587, n_1588, n_1589;
  wire n_1593, n_1606, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616;
  wire n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624;
  wire n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632;
  wire n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640;
  wire n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648;
  wire n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656;
  wire n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664;
  wire n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672;
  wire n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680;
  wire n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688;
  wire n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696;
  wire n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704;
  wire n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712;
  wire n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720;
  wire n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728;
  wire n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736;
  wire n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744;
  wire n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752;
  wire n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760;
  wire n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768;
  wire n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776;
  wire n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784;
  wire n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792;
  wire n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800;
  wire n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], n_171);
  xor g270 (n_117, n_622, A[2]);
  nand g3 (n_623, A[1], n_171);
  nand g271 (n_624, A[2], n_171);
  nand g272 (n_625, A[1], A[2]);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, n_69);
  xor g288 (n_176, n_634, A[4]);
  nand g289 (n_635, n_68, n_69);
  nand g290 (n_636, A[4], n_69);
  nand g291 (n_637, n_68, A[4]);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_176);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_176);
  nand g296 (n_640, A[7], n_176);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g305 (n_646, n_117, A[5]);
  xor g306 (n_180, n_646, n_179);
  nand g307 (n_647, n_117, A[5]);
  nand g308 (n_648, n_179, A[5]);
  nand g309 (n_649, n_117, n_179);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, A[6], n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, A[6], n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, A[6], A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_188, n_659, n_660, n_661);
  xor g329 (n_662, n_183, n_184);
  xor g330 (n_112, n_662, A[9]);
  nand g331 (n_663, n_183, n_184);
  nand g332 (n_664, A[9], n_184);
  nand g333 (n_665, n_183, A[9]);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_187, n_630, n_67);
  nand g340 (n_668, n_67, n_173);
  nand g341 (n_669, A[4], n_67);
  nand g342 (n_71, n_631, n_668, n_669);
  xor g343 (n_670, A[7], n_187);
  xor g344 (n_189, n_670, A[8]);
  nand g345 (n_671, A[7], n_187);
  nand g346 (n_672, A[8], n_187);
  nand g347 (n_673, A[7], A[8]);
  nand g348 (n_73, n_671, n_672, n_673);
  xor g349 (n_674, n_188, A[10]);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, n_188, A[10]);
  nand g352 (n_676, n_189, A[10]);
  nand g353 (n_677, n_188, n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_195, n_638, n_71);
  nand g366 (n_684, n_71, n_176);
  nand g367 (n_685, A[5], n_71);
  nand g368 (n_201, n_639, n_684, n_685);
  xor g369 (n_686, A[8], A[9]);
  xor g370 (n_196, n_686, n_73);
  nand g371 (n_687, A[8], A[9]);
  nand g372 (n_688, n_73, A[9]);
  nand g373 (n_689, A[8], n_73);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, A[11], n_195);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, A[11], n_195);
  nand g378 (n_692, n_196, n_195);
  nand g379 (n_693, A[11], n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g394 (n_202, n_650, A[9]);
  nand g396 (n_704, A[9], n_180);
  nand g397 (n_705, A[6], A[9]);
  nand g398 (n_209, n_651, n_704, n_705);
  xor g399 (n_706, A[10], n_201);
  xor g400 (n_204, n_706, n_202);
  nand g401 (n_707, A[10], n_201);
  nand g402 (n_708, n_202, n_201);
  nand g403 (n_709, A[10], n_202);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, A[12], n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, A[12], n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, A[12], n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g424 (n_210, n_662, A[10]);
  nand g426 (n_724, A[10], n_184);
  nand g427 (n_725, n_183, A[10]);
  nand g428 (n_218, n_663, n_724, n_725);
  xor g429 (n_726, A[11], n_209);
  xor g430 (n_212, n_726, n_210);
  nand g431 (n_727, A[11], n_209);
  nand g432 (n_728, n_210, n_209);
  nand g433 (n_729, A[11], n_210);
  nand g434 (n_220, n_727, n_728, n_729);
  xor g435 (n_730, A[13], n_211);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, A[13], n_211);
  nand g438 (n_732, n_212, n_211);
  nand g439 (n_733, A[13], n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_217, n_738, n_187);
  xor g455 (n_742, n_188, A[11]);
  xor g456 (n_219, n_742, n_217);
  nand g457 (n_743, n_188, A[11]);
  nand g458 (n_744, n_217, A[11]);
  nand g459 (n_745, n_188, n_217);
  nand g460 (n_224, n_743, n_744, n_745);
  xor g461 (n_746, n_218, A[12]);
  xor g462 (n_221, n_746, n_219);
  nand g463 (n_747, n_218, A[12]);
  nand g464 (n_748, n_219, A[12]);
  nand g465 (n_749, n_218, n_219);
  nand g466 (n_226, n_747, n_748, n_749);
  xor g467 (n_750, n_220, A[14]);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, n_220, A[14]);
  nand g470 (n_752, n_221, A[14]);
  nand g471 (n_753, n_220, n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g482 (n_72, n_638, A[8]);
  nand g484 (n_760, A[8], n_176);
  nand g485 (n_761, A[5], A[8]);
  nand g486 (n_232, n_639, n_760, n_761);
  xor g487 (n_762, n_71, A[9]);
  xor g488 (n_223, n_762, n_72);
  nand g489 (n_763, n_71, A[9]);
  nand g490 (n_764, n_72, A[9]);
  nand g491 (n_765, n_71, n_72);
  nand g492 (n_234, n_763, n_764, n_765);
  xor g493 (n_766, n_73, A[12]);
  xor g494 (n_225, n_766, n_223);
  nand g495 (n_767, n_73, A[12]);
  nand g496 (n_768, n_223, A[12]);
  nand g497 (n_769, n_73, n_223);
  nand g498 (n_236, n_767, n_768, n_769);
  xor g499 (n_770, A[13], n_224);
  xor g500 (n_227, n_770, A[15]);
  nand g501 (n_771, A[13], n_224);
  nand g502 (n_772, A[15], n_224);
  nand g503 (n_773, A[13], A[15]);
  nand g504 (n_238, n_771, n_772, n_773);
  xor g505 (n_774, n_225, n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, n_225, n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, n_225, n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g529 (n_790, A[10], n_232);
  xor g530 (n_235, n_790, n_202);
  nand g531 (n_791, A[10], n_232);
  nand g532 (n_792, n_202, n_232);
  nand g534 (n_246, n_791, n_792, n_709);
  xor g535 (n_794, n_234, A[13]);
  xor g536 (n_237, n_794, n_235);
  nand g537 (n_795, n_234, A[13]);
  nand g538 (n_796, n_235, A[13]);
  nand g539 (n_797, n_234, n_235);
  nand g540 (n_248, n_795, n_796, n_797);
  xor g541 (n_798, A[14], n_236);
  xor g542 (n_239, n_798, A[16]);
  nand g543 (n_799, A[14], n_236);
  nand g544 (n_800, A[16], n_236);
  nand g545 (n_801, A[14], A[16]);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, n_237, n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, n_237, n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, n_237, n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g577 (n_822, n_246, A[14]);
  xor g578 (n_249, n_822, n_212);
  nand g579 (n_823, n_246, A[14]);
  nand g580 (n_824, n_212, A[14]);
  nand g581 (n_825, n_246, n_212);
  nand g582 (n_261, n_823, n_824, n_825);
  xor g583 (n_826, A[15], n_248);
  xor g584 (n_251, n_826, A[17]);
  nand g585 (n_827, A[15], n_248);
  nand g586 (n_828, A[17], n_248);
  nand g587 (n_829, A[15], A[17]);
  nand g588 (n_118, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g621 (n_850, n_220, A[15]);
  xor g622 (n_262, n_850, n_221);
  nand g623 (n_851, n_220, A[15]);
  nand g624 (n_852, n_221, A[15]);
  nand g626 (n_274, n_851, n_852, n_753);
  xor g627 (n_854, A[16], n_261);
  xor g628 (n_119, n_854, A[18]);
  nand g629 (n_855, A[16], n_261);
  nand g630 (n_856, A[18], n_261);
  nand g631 (n_857, A[16], A[18]);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_262, n_118);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_262, n_118);
  nand g636 (n_860, n_119, n_118);
  nand g637 (n_861, n_262, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g641 (n_862, n_68, A[4]);
  xor g642 (n_265, n_862, n_69);
  xor g647 (n_866, A[5], n_265);
  xor g648 (n_267, n_866, A[8]);
  nand g649 (n_867, A[5], n_265);
  nand g650 (n_868, A[8], n_265);
  nand g652 (n_282, n_867, n_868, n_761);
  xor g654 (n_269, n_762, n_267);
  nand g656 (n_872, n_267, A[9]);
  nand g657 (n_873, n_71, n_267);
  nand g658 (n_284, n_763, n_872, n_873);
  xor g660 (n_271, n_766, A[13]);
  nand g662 (n_876, A[13], A[12]);
  nand g663 (n_877, n_73, A[13]);
  nand g664 (n_286, n_767, n_876, n_877);
  xor g665 (n_878, n_269, n_224);
  xor g666 (n_273, n_878, n_271);
  nand g667 (n_879, n_269, n_224);
  nand g668 (n_880, n_271, n_224);
  nand g669 (n_881, n_269, n_271);
  nand g670 (n_288, n_879, n_880, n_881);
  xor g671 (n_882, n_226, A[16]);
  xor g672 (n_275, n_882, n_273);
  nand g673 (n_883, n_226, A[16]);
  nand g674 (n_884, n_273, A[16]);
  nand g675 (n_885, n_226, n_273);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, A[17], n_274);
  xor g678 (n_277, n_886, A[19]);
  nand g679 (n_887, A[17], n_274);
  nand g680 (n_888, A[19], n_274);
  nand g681 (n_889, A[17], A[19]);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g696 (n_281, n_646, A[6]);
  nand g698 (n_900, A[6], A[5]);
  nand g699 (n_901, n_117, A[6]);
  nand g700 (n_296, n_647, n_900, n_901);
  xor g701 (n_902, n_179, n_281);
  xor g702 (n_283, n_902, A[9]);
  nand g703 (n_903, n_179, n_281);
  nand g704 (n_904, A[9], n_281);
  nand g705 (n_905, n_179, A[9]);
  nand g706 (n_298, n_903, n_904, n_905);
  xor g707 (n_906, A[10], n_282);
  xor g708 (n_285, n_906, n_283);
  nand g709 (n_907, A[10], n_282);
  nand g710 (n_908, n_283, n_282);
  nand g711 (n_909, A[10], n_283);
  nand g712 (n_300, n_907, n_908, n_909);
  xor g713 (n_910, n_284, A[13]);
  xor g714 (n_287, n_910, n_285);
  nand g715 (n_911, n_284, A[13]);
  nand g716 (n_912, n_285, A[13]);
  nand g717 (n_913, n_284, n_285);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, A[14], n_286);
  xor g720 (n_289, n_914, n_287);
  nand g721 (n_915, A[14], n_286);
  nand g722 (n_916, n_287, n_286);
  nand g723 (n_917, A[14], n_287);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, n_288, A[17]);
  xor g726 (n_291, n_918, n_289);
  nand g727 (n_919, n_288, A[17]);
  nand g728 (n_920, n_289, A[17]);
  nand g729 (n_921, n_288, n_289);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, A[18], n_290);
  xor g732 (n_293, n_922, A[20]);
  nand g733 (n_923, A[18], n_290);
  nand g734 (n_924, A[20], n_290);
  nand g735 (n_925, A[18], A[20]);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g755 (n_938, n_296, n_184);
  xor g756 (n_299, n_938, A[10]);
  nand g757 (n_939, n_296, n_184);
  nand g759 (n_941, n_296, A[10]);
  nand g760 (n_315, n_939, n_724, n_941);
  xor g761 (n_942, A[11], n_298);
  xor g762 (n_301, n_942, n_299);
  nand g763 (n_943, A[11], n_298);
  nand g764 (n_944, n_299, n_298);
  nand g765 (n_945, A[11], n_299);
  nand g766 (n_317, n_943, n_944, n_945);
  xor g767 (n_946, n_300, A[14]);
  xor g768 (n_303, n_946, n_301);
  nand g769 (n_947, n_300, A[14]);
  nand g770 (n_948, n_301, A[14]);
  nand g771 (n_949, n_300, n_301);
  nand g772 (n_319, n_947, n_948, n_949);
  xor g773 (n_950, A[15], n_302);
  xor g774 (n_305, n_950, n_303);
  nand g775 (n_951, A[15], n_302);
  nand g776 (n_952, n_303, n_302);
  nand g777 (n_953, A[15], n_303);
  nand g778 (n_321, n_951, n_952, n_953);
  xor g779 (n_954, n_304, A[18]);
  xor g780 (n_307, n_954, n_305);
  nand g781 (n_955, n_304, A[18]);
  nand g782 (n_956, n_305, A[18]);
  nand g783 (n_957, n_304, n_305);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, A[19], n_306);
  xor g786 (n_309, n_958, A[21]);
  nand g787 (n_959, A[19], n_306);
  nand g788 (n_960, A[21], n_306);
  nand g789 (n_961, A[19], A[21]);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g817 (n_978, A[12], n_315);
  xor g818 (n_318, n_978, n_219);
  nand g819 (n_979, A[12], n_315);
  nand g820 (n_980, n_219, n_315);
  nand g822 (n_336, n_979, n_980, n_748);
  xor g823 (n_982, n_317, A[15]);
  xor g824 (n_320, n_982, A[16]);
  nand g825 (n_983, n_317, A[15]);
  nand g826 (n_984, A[16], A[15]);
  nand g827 (n_985, n_317, A[16]);
  nand g828 (n_338, n_983, n_984, n_985);
  xor g829 (n_986, n_318, n_319);
  xor g830 (n_322, n_986, n_320);
  nand g831 (n_987, n_318, n_319);
  nand g832 (n_988, n_320, n_319);
  nand g833 (n_989, n_318, n_320);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, n_321, A[19]);
  xor g836 (n_324, n_990, n_322);
  nand g837 (n_991, n_321, A[19]);
  nand g838 (n_992, n_322, A[19]);
  nand g839 (n_993, n_321, n_322);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, A[20], n_323);
  xor g842 (n_326, n_994, n_324);
  nand g843 (n_995, A[20], n_323);
  nand g844 (n_996, n_324, n_323);
  nand g845 (n_997, A[20], n_324);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, A[22], n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, A[22], n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, A[22], n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g868 (n_333, n_762, n_73);
  nand g871 (n_1013, n_71, n_73);
  nand g872 (n_354, n_763, n_688, n_1013);
  xor g873 (n_1014, n_267, A[12]);
  xor g874 (n_335, n_1014, n_333);
  nand g875 (n_1015, n_267, A[12]);
  nand g876 (n_1016, n_333, A[12]);
  nand g877 (n_1017, n_267, n_333);
  nand g878 (n_356, n_1015, n_1016, n_1017);
  xor g880 (n_337, n_770, n_335);
  nand g882 (n_1020, n_335, n_224);
  nand g883 (n_1021, A[13], n_335);
  nand g884 (n_358, n_771, n_1020, n_1021);
  xor g885 (n_1022, n_336, A[16]);
  xor g886 (n_339, n_1022, n_337);
  nand g887 (n_1023, n_336, A[16]);
  nand g888 (n_1024, n_337, A[16]);
  nand g889 (n_1025, n_336, n_337);
  nand g890 (n_360, n_1023, n_1024, n_1025);
  xor g891 (n_1026, A[17], n_338);
  xor g892 (n_341, n_1026, n_339);
  nand g893 (n_1027, A[17], n_338);
  nand g894 (n_1028, n_339, n_338);
  nand g895 (n_1029, A[17], n_339);
  nand g896 (n_362, n_1027, n_1028, n_1029);
  xor g897 (n_1030, A[20], n_340);
  xor g898 (n_343, n_1030, n_341);
  nand g899 (n_1031, A[20], n_340);
  nand g900 (n_1032, n_341, n_340);
  nand g901 (n_1033, A[20], n_341);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, A[21], n_342);
  xor g904 (n_345, n_1034, n_343);
  nand g905 (n_1035, A[21], n_342);
  nand g906 (n_1036, n_343, n_342);
  nand g907 (n_1037, A[21], n_343);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, A[23], n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, A[23], n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, A[23], n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  nand g922 (n_371, n_1043, n_1044, n_624);
  nand g928 (n_373, n_1047, n_648, n_1049);
  nand g934 (n_375, n_1051, n_1052, n_705);
  nand g940 (n_377, n_907, n_1056, n_1057);
  xor g941 (n_1058, n_354, A[13]);
  xor g942 (n_357, n_1058, n_355);
  nand g943 (n_1059, n_354, A[13]);
  nand g944 (n_1060, n_355, A[13]);
  nand g945 (n_1061, n_354, n_355);
  nand g946 (n_379, n_1059, n_1060, n_1061);
  xor g947 (n_1062, A[14], n_356);
  xor g948 (n_359, n_1062, n_357);
  nand g949 (n_1063, A[14], n_356);
  nand g950 (n_1064, n_357, n_356);
  nand g951 (n_1065, A[14], n_357);
  nand g952 (n_381, n_1063, n_1064, n_1065);
  xor g953 (n_1066, n_358, A[17]);
  xor g954 (n_361, n_1066, A[18]);
  nand g955 (n_1067, n_358, A[17]);
  nand g956 (n_1068, A[18], A[17]);
  nand g957 (n_1069, n_358, A[18]);
  nand g958 (n_383, n_1067, n_1068, n_1069);
  xor g959 (n_1070, n_359, n_360);
  xor g960 (n_363, n_1070, n_361);
  nand g961 (n_1071, n_359, n_360);
  nand g962 (n_1072, n_361, n_360);
  nand g963 (n_1073, n_359, n_361);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, A[21], n_362);
  xor g966 (n_365, n_1074, A[22]);
  nand g967 (n_1075, A[21], n_362);
  nand g968 (n_1076, A[22], n_362);
  nand g969 (n_1077, A[21], A[22]);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g971 (n_1078, n_363, n_364);
  nand g973 (n_1079, n_363, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  nand g990 (n_392, n_627, n_1088, n_1044);
  xor g991 (n_1090, n_371, n_372);
  xor g992 (n_374, n_1090, A[6]);
  nand g993 (n_1091, n_371, n_372);
  nand g994 (n_1092, A[6], n_372);
  nand g995 (n_1093, n_371, A[6]);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, n_374);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, n_374, n_373);
  nand g1001 (n_1097, A[7], n_374);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, A[10], A[11]);
  xor g1004 (n_378, n_1098, n_375);
  nand g1005 (n_1099, A[10], A[11]);
  nand g1006 (n_1100, n_375, A[11]);
  nand g1007 (n_1101, A[10], n_375);
  nand g1008 (n_398, n_1099, n_1100, n_1101);
  xor g1009 (n_1102, n_376, n_377);
  xor g1010 (n_380, n_1102, n_378);
  nand g1011 (n_1103, n_376, n_377);
  nand g1012 (n_1104, n_378, n_377);
  nand g1013 (n_1105, n_376, n_378);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, A[14], A[15]);
  xor g1016 (n_382, n_1106, n_379);
  nand g1017 (n_1107, A[14], A[15]);
  nand g1018 (n_1108, n_379, A[15]);
  nand g1019 (n_1109, A[14], n_379);
  nand g1020 (n_402, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, n_380, A[18]);
  xor g1022 (n_384, n_1110, n_381);
  nand g1023 (n_1111, n_380, A[18]);
  nand g1024 (n_1112, n_381, A[18]);
  nand g1025 (n_1113, n_380, n_381);
  nand g1026 (n_404, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, n_382, A[19]);
  xor g1028 (n_386, n_1114, n_383);
  nand g1029 (n_1115, n_382, A[19]);
  nand g1030 (n_1116, n_383, A[19]);
  nand g1031 (n_1117, n_382, n_383);
  nand g1032 (n_406, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_384, n_385);
  xor g1034 (n_388, n_1118, n_386);
  nand g1035 (n_1119, n_384, n_385);
  nand g1036 (n_1120, n_386, n_385);
  nand g1037 (n_1121, n_384, n_386);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, A[22], A[23]);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, A[22], A[23]);
  nand g1042 (n_1124, n_387, A[23]);
  nand g1043 (n_1125, A[22], n_387);
  nand g1044 (n_411, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1051 (n_1130, A[3], A[1]);
  xor g1052 (n_393, n_1130, A[4]);
  nand g1053 (n_1131, A[3], A[1]);
  nand g1054 (n_1132, A[4], A[1]);
  nand g1055 (n_1133, A[3], A[4]);
  nand g1056 (n_412, n_1131, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, n_396, A[11]);
  xor g1070 (n_399, n_1142, n_397);
  nand g1071 (n_1143, n_396, A[11]);
  nand g1072 (n_1144, n_397, A[11]);
  nand g1073 (n_1145, n_396, n_397);
  nand g1074 (n_417, n_1143, n_1144, n_1145);
  xor g1075 (n_1146, A[12], n_398);
  xor g1076 (n_401, n_1146, n_399);
  nand g1077 (n_1147, A[12], n_398);
  nand g1078 (n_1148, n_399, n_398);
  nand g1079 (n_1149, A[12], n_399);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, A[15], n_400);
  xor g1082 (n_403, n_1150, A[16]);
  nand g1083 (n_1151, A[15], n_400);
  nand g1084 (n_1152, A[16], n_400);
  nand g1086 (n_421, n_1151, n_1152, n_984);
  xor g1087 (n_1154, n_401, n_402);
  xor g1088 (n_405, n_1154, n_403);
  nand g1089 (n_1155, n_401, n_402);
  nand g1090 (n_1156, n_403, n_402);
  nand g1091 (n_1157, n_401, n_403);
  nand g1092 (n_424, n_1155, n_1156, n_1157);
  xor g1093 (n_1158, A[19], n_404);
  xor g1094 (n_407, n_1158, A[20]);
  nand g1095 (n_1159, A[19], n_404);
  nand g1096 (n_1160, A[20], n_404);
  nand g1097 (n_1161, A[19], A[20]);
  nand g1098 (n_425, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_405, n_406);
  xor g1100 (n_409, n_1162, n_407);
  nand g1101 (n_1163, n_405, n_406);
  nand g1102 (n_1164, n_407, n_406);
  nand g1103 (n_1165, n_405, n_407);
  nand g1104 (n_428, n_1163, n_1164, n_1165);
  xor g1106 (n_410, n_1166, n_408);
  nand g1109 (n_1169, A[23], n_408);
  nand g1110 (n_430, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1123 (n_1178, A[8], n_413);
  xor g1124 (n_415, n_1178, A[9]);
  nand g1125 (n_1179, A[8], n_413);
  nand g1126 (n_1180, A[9], n_413);
  nand g1128 (n_435, n_1179, n_1180, n_687);
  xor g1129 (n_1182, n_414, n_415);
  xor g1130 (n_418, n_1182, n_416);
  nand g1131 (n_1183, n_414, n_415);
  nand g1132 (n_1184, n_416, n_415);
  nand g1133 (n_1185, n_414, n_416);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, A[12], A[13]);
  xor g1136 (n_420, n_1186, n_417);
  nand g1138 (n_1188, n_417, A[13]);
  nand g1139 (n_1189, A[12], n_417);
  nand g1140 (n_439, n_876, n_1188, n_1189);
  xor g1141 (n_1190, n_418, n_419);
  xor g1142 (n_422, n_1190, A[16]);
  nand g1143 (n_1191, n_418, n_419);
  nand g1144 (n_1192, A[16], n_419);
  nand g1145 (n_1193, n_418, A[16]);
  nand g1146 (n_440, n_1191, n_1192, n_1193);
  xor g1147 (n_1194, n_420, A[17]);
  xor g1148 (n_423, n_1194, n_421);
  nand g1149 (n_1195, n_420, A[17]);
  nand g1150 (n_1196, n_421, A[17]);
  nand g1151 (n_1197, n_420, n_421);
  nand g1152 (n_442, n_1195, n_1196, n_1197);
  xor g1153 (n_1198, n_422, A[20]);
  xor g1154 (n_426, n_1198, n_423);
  nand g1155 (n_1199, n_422, A[20]);
  nand g1156 (n_1200, n_423, A[20]);
  nand g1157 (n_1201, n_422, n_423);
  nand g1158 (n_445, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_424, A[21]);
  xor g1160 (n_427, n_1202, n_425);
  nand g1161 (n_1203, n_424, A[21]);
  nand g1162 (n_1204, n_425, A[21]);
  nand g1163 (n_1205, n_424, n_425);
  nand g1164 (n_447, n_1203, n_1204, n_1205);
  xor g1166 (n_429, n_1206, n_427);
  nand g1169 (n_1209, n_426, n_427);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, n_433);
  nand g1183 (n_1217, A[6], n_433);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, A[9], A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, A[9], A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, A[9], n_434);
  nand g1190 (n_456, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, n_435, n_436);
  xor g1192 (n_438, n_1222, A[13]);
  nand g1193 (n_1223, n_435, n_436);
  nand g1194 (n_1224, A[13], n_436);
  nand g1195 (n_1225, n_435, A[13]);
  nand g1196 (n_457, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, n_437, A[14]);
  xor g1198 (n_441, n_1226, n_438);
  nand g1199 (n_1227, n_437, A[14]);
  nand g1200 (n_1228, n_438, A[14]);
  nand g1201 (n_1229, n_437, n_438);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, n_439, A[17]);
  xor g1204 (n_443, n_1230, n_440);
  nand g1205 (n_1231, n_439, A[17]);
  nand g1206 (n_1232, n_440, A[17]);
  nand g1207 (n_1233, n_439, n_440);
  nand g1208 (n_461, n_1231, n_1232, n_1233);
  xor g1209 (n_1234, A[18], n_441);
  xor g1210 (n_444, n_1234, n_442);
  nand g1211 (n_1235, A[18], n_441);
  nand g1212 (n_1236, n_442, n_441);
  nand g1213 (n_1237, A[18], n_442);
  nand g1214 (n_463, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_443, A[21]);
  xor g1216 (n_446, n_1238, A[22]);
  nand g1217 (n_1239, n_443, A[21]);
  nand g1219 (n_1241, n_443, A[22]);
  nand g1220 (n_465, n_1239, n_1077, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[5], A[7]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], n_453);
  xor g1242 (n_455, n_1254, A[11]);
  nand g1243 (n_1255, A[10], n_453);
  nand g1244 (n_1256, A[11], n_453);
  nand g1246 (n_472, n_1255, n_1256, n_1099);
  xor g1247 (n_1258, n_454, n_455);
  xor g1248 (n_458, n_1258, n_456);
  nand g1249 (n_1259, n_454, n_455);
  nand g1250 (n_1260, n_456, n_455);
  nand g1251 (n_1261, n_454, n_456);
  nand g1252 (n_474, n_1259, n_1260, n_1261);
  xor g1253 (n_1262, A[14], n_457);
  xor g1254 (n_460, n_1262, A[15]);
  nand g1255 (n_1263, A[14], n_457);
  nand g1256 (n_1264, A[15], n_457);
  nand g1258 (n_476, n_1263, n_1264, n_1107);
  xor g1259 (n_1266, n_458, A[18]);
  xor g1260 (n_462, n_1266, n_459);
  nand g1261 (n_1267, n_458, A[18]);
  nand g1262 (n_1268, n_459, A[18]);
  nand g1263 (n_1269, n_458, n_459);
  nand g1264 (n_479, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, n_460, A[19]);
  xor g1266 (n_464, n_1270, n_461);
  nand g1267 (n_1271, n_460, A[19]);
  nand g1268 (n_1272, n_461, A[19]);
  nand g1269 (n_1273, n_460, n_461);
  nand g1270 (n_480, n_1271, n_1272, n_1273);
  xor g1271 (n_1274, n_462, n_463);
  xor g1272 (n_466, n_1274, n_464);
  nand g1273 (n_1275, n_462, n_463);
  nand g1274 (n_1276, n_464, n_463);
  nand g1275 (n_1277, n_462, n_464);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1278 (n_467, n_1122, n_465);
  nand g1280 (n_1280, n_465, A[23]);
  nand g1281 (n_1281, A[22], n_465);
  nand g1282 (n_485, n_1123, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1289 (n_1286, A[7], A[6]);
  xor g1290 (n_471, n_1286, A[8]);
  nand g1294 (n_486, n_661, n_653, n_673);
  xor g1295 (n_1290, n_470, A[11]);
  xor g1296 (n_473, n_1290, n_471);
  nand g1297 (n_1291, n_470, A[11]);
  nand g1298 (n_1292, n_471, A[11]);
  nand g1299 (n_1293, n_470, n_471);
  nand g1300 (n_487, n_1291, n_1292, n_1293);
  xor g1301 (n_1294, A[12], n_472);
  xor g1302 (n_475, n_1294, n_473);
  nand g1303 (n_1295, A[12], n_472);
  nand g1304 (n_1296, n_473, n_472);
  nand g1305 (n_1297, A[12], n_473);
  nand g1306 (n_490, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, A[15], n_474);
  xor g1308 (n_477, n_1298, n_475);
  nand g1309 (n_1299, A[15], n_474);
  nand g1310 (n_1300, n_475, n_474);
  nand g1311 (n_1301, A[15], n_475);
  nand g1312 (n_491, n_1299, n_1300, n_1301);
  xor g1313 (n_1302, A[16], n_476);
  xor g1314 (n_478, n_1302, n_477);
  nand g1315 (n_1303, A[16], n_476);
  nand g1316 (n_1304, n_477, n_476);
  nand g1317 (n_1305, A[16], n_477);
  nand g1318 (n_494, n_1303, n_1304, n_1305);
  xor g1319 (n_1306, A[19], n_478);
  xor g1320 (n_481, n_1306, n_479);
  nand g1321 (n_1307, A[19], n_478);
  nand g1322 (n_1308, n_479, n_478);
  nand g1323 (n_1309, A[19], n_479);
  nand g1324 (n_495, n_1307, n_1308, n_1309);
  xor g1325 (n_1310, A[20], n_480);
  xor g1326 (n_483, n_1310, n_481);
  nand g1327 (n_1311, A[20], n_480);
  nand g1328 (n_1312, n_481, n_480);
  nand g1329 (n_1313, A[20], n_481);
  nand g1330 (n_498, n_1311, n_1312, n_1313);
  xor g1332 (n_484, n_1166, n_482);
  nand g1335 (n_1317, A[23], n_482);
  nand g1336 (n_500, n_1167, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1344 (n_488, n_686, n_486);
  nand g1346 (n_1324, n_486, A[9]);
  nand g1347 (n_1325, A[8], n_486);
  nand g1348 (n_503, n_687, n_1324, n_1325);
  xor g1349 (n_1326, A[12], n_487);
  xor g1350 (n_489, n_1326, n_488);
  nand g1351 (n_1327, A[12], n_487);
  nand g1352 (n_1328, n_488, n_487);
  nand g1353 (n_1329, A[12], n_488);
  nand g1354 (n_504, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, A[13], n_489);
  xor g1356 (n_492, n_1330, n_490);
  nand g1357 (n_1331, A[13], n_489);
  nand g1358 (n_1332, n_490, n_489);
  nand g1359 (n_1333, A[13], n_490);
  nand g1360 (n_507, n_1331, n_1332, n_1333);
  xor g1361 (n_1334, A[16], A[17]);
  xor g1362 (n_493, n_1334, n_491);
  nand g1363 (n_1335, A[16], A[17]);
  nand g1364 (n_1336, n_491, A[17]);
  nand g1365 (n_1337, A[16], n_491);
  nand g1366 (n_508, n_1335, n_1336, n_1337);
  xor g1367 (n_1338, n_492, A[20]);
  xor g1368 (n_496, n_1338, n_493);
  nand g1369 (n_1339, n_492, A[20]);
  nand g1370 (n_1340, n_493, A[20]);
  nand g1371 (n_1341, n_492, n_493);
  nand g1372 (n_511, n_1339, n_1340, n_1341);
  xor g1373 (n_1342, n_494, A[21]);
  xor g1374 (n_497, n_1342, n_495);
  nand g1375 (n_1343, n_494, A[21]);
  nand g1376 (n_1344, n_495, A[21]);
  nand g1377 (n_1345, n_494, n_495);
  nand g1378 (n_512, n_1343, n_1344, n_1345);
  xor g1380 (n_499, n_1346, n_497);
  nand g1383 (n_1349, n_496, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  nand g1397 (n_1357, A[10], n_503);
  nand g1398 (n_520, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], A[14]);
  xor g1400 (n_506, n_1358, n_504);
  nand g1401 (n_1359, A[13], A[14]);
  nand g1402 (n_1360, n_504, A[14]);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_521, n_1359, n_1360, n_1361);
  xor g1405 (n_1362, n_505, A[17]);
  xor g1406 (n_509, n_1362, n_506);
  nand g1407 (n_1363, n_505, A[17]);
  nand g1408 (n_1364, n_506, A[17]);
  nand g1409 (n_1365, n_505, n_506);
  nand g1410 (n_523, n_1363, n_1364, n_1365);
  xor g1411 (n_1366, A[18], n_507);
  xor g1412 (n_510, n_1366, n_508);
  nand g1413 (n_1367, A[18], n_507);
  nand g1414 (n_1368, n_508, n_507);
  nand g1415 (n_1369, A[18], n_508);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_509, A[21]);
  xor g1418 (n_513, n_1370, A[22]);
  nand g1419 (n_1371, n_509, A[21]);
  nand g1421 (n_1373, n_509, A[22]);
  nand g1422 (n_527, n_1371, n_1077, n_1373);
  xor g1423 (n_1374, n_510, n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, n_510, n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, n_510, n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1437 (n_1382, A[11], A[9]);
  nand g1439 (n_1383, A[11], A[9]);
  nand g1442 (n_532, n_1383, n_1384, n_1385);
  xor g1443 (n_1386, n_519, A[14]);
  xor g1444 (n_522, n_1386, n_520);
  nand g1445 (n_1387, n_519, A[14]);
  nand g1446 (n_1388, n_520, A[14]);
  nand g1447 (n_1389, n_519, n_520);
  nand g1448 (n_534, n_1387, n_1388, n_1389);
  xor g1449 (n_1390, A[15], n_521);
  xor g1450 (n_524, n_1390, n_522);
  nand g1451 (n_1391, A[15], n_521);
  nand g1452 (n_1392, n_522, n_521);
  nand g1453 (n_1393, A[15], n_522);
  nand g1454 (n_536, n_1391, n_1392, n_1393);
  xor g1455 (n_1394, A[18], n_523);
  xor g1456 (n_525, n_1394, A[19]);
  nand g1457 (n_1395, A[18], n_523);
  nand g1458 (n_1396, A[19], n_523);
  nand g1459 (n_1397, A[18], A[19]);
  nand g1460 (n_538, n_1395, n_1396, n_1397);
  xor g1461 (n_1398, n_524, n_525);
  xor g1462 (n_528, n_1398, n_526);
  nand g1463 (n_1399, n_524, n_525);
  nand g1464 (n_1400, n_526, n_525);
  nand g1465 (n_1401, n_524, n_526);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1468 (n_529, n_1122, n_527);
  nand g1470 (n_1404, n_527, A[23]);
  nand g1471 (n_1405, A[22], n_527);
  nand g1472 (n_543, n_1123, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1480 (n_533, n_1098, A[12]);
  nand g1482 (n_1412, A[12], A[10]);
  nand g1483 (n_1413, A[11], A[12]);
  nand g1484 (n_544, n_1099, n_1412, n_1413);
  xor g1485 (n_1414, n_532, n_533);
  xor g1486 (n_535, n_1414, A[15]);
  nand g1487 (n_1415, n_532, n_533);
  nand g1488 (n_1416, A[15], n_533);
  nand g1489 (n_1417, n_532, A[15]);
  nand g1490 (n_546, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, A[16], n_534);
  xor g1492 (n_537, n_1418, n_535);
  nand g1493 (n_1419, A[16], n_534);
  nand g1494 (n_1420, n_535, n_534);
  nand g1495 (n_1421, A[16], n_535);
  nand g1496 (n_547, n_1419, n_1420, n_1421);
  xor g1497 (n_1422, A[19], n_536);
  xor g1498 (n_539, n_1422, A[20]);
  nand g1499 (n_1423, A[19], n_536);
  nand g1500 (n_1424, A[20], n_536);
  nand g1502 (n_549, n_1423, n_1424, n_1161);
  xor g1503 (n_1426, n_537, n_538);
  xor g1504 (n_541, n_1426, n_539);
  nand g1505 (n_1427, n_537, n_538);
  nand g1506 (n_1428, n_539, n_538);
  nand g1507 (n_1429, n_537, n_539);
  nand g1508 (n_551, n_1427, n_1428, n_1429);
  xor g1510 (n_542, n_1166, n_540);
  nand g1513 (n_1433, A[23], n_540);
  nand g1514 (n_554, n_1167, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1522 (n_545, n_1186, n_544);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_876, n_1440, n_1441);
  xor g1527 (n_1442, A[16], n_545);
  xor g1528 (n_548, n_1442, A[17]);
  nand g1529 (n_1443, A[16], n_545);
  nand g1530 (n_1444, A[17], n_545);
  nand g1532 (n_559, n_1443, n_1444, n_1335);
  xor g1533 (n_1446, n_546, n_547);
  xor g1534 (n_550, n_1446, n_548);
  nand g1535 (n_1447, n_546, n_547);
  nand g1536 (n_1448, n_548, n_547);
  nand g1537 (n_1449, n_546, n_548);
  nand g1538 (n_561, n_1447, n_1448, n_1449);
  xor g1539 (n_1450, A[20], A[21]);
  xor g1540 (n_552, n_1450, n_549);
  nand g1541 (n_1451, A[20], A[21]);
  nand g1542 (n_1452, n_549, A[21]);
  nand g1543 (n_1453, A[20], n_549);
  nand g1544 (n_563, n_1451, n_1452, n_1453);
  xor g1546 (n_553, n_1454, n_551);
  nand g1549 (n_1457, n_550, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1563 (n_1465, A[14], n_557);
  nand g1564 (n_570, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, A[17], A[18]);
  xor g1566 (n_560, n_1466, n_558);
  nand g1568 (n_1468, n_558, A[18]);
  nand g1569 (n_1469, A[17], n_558);
  nand g1570 (n_571, n_1068, n_1468, n_1469);
  xor g1571 (n_1470, n_559, n_560);
  xor g1572 (n_562, n_1470, n_561);
  nand g1573 (n_1471, n_559, n_560);
  nand g1574 (n_1472, n_561, n_560);
  nand g1575 (n_1473, n_559, n_561);
  nand g1576 (n_574, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, A[21], A[22]);
  xor g1578 (n_564, n_1474, n_562);
  nand g1580 (n_1476, n_562, A[22]);
  nand g1581 (n_1477, A[21], n_562);
  nand g1582 (n_575, n_1077, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  nand g1596 (n_578, n_1107, n_1484, n_1463);
  xor g1597 (n_1486, A[18], n_569);
  xor g1598 (n_572, n_1486, n_570);
  nand g1599 (n_1487, A[18], n_569);
  nand g1600 (n_1488, n_570, n_569);
  nand g1601 (n_1489, A[18], n_570);
  nand g1602 (n_580, n_1487, n_1488, n_1489);
  xor g1603 (n_1490, A[19], n_571);
  xor g1604 (n_573, n_1490, n_572);
  nand g1605 (n_1491, A[19], n_571);
  nand g1606 (n_1492, n_572, n_571);
  nand g1607 (n_1493, A[19], n_572);
  nand g1608 (n_582, n_1491, n_1492, n_1493);
  xor g1609 (n_1494, A[22], n_573);
  xor g1610 (n_576, n_1494, A[23]);
  nand g1611 (n_1495, A[22], n_573);
  nand g1612 (n_1496, A[23], n_573);
  nand g1614 (n_584, n_1495, n_1496, n_1123);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1621 (n_1502, A[15], A[16]);
  xor g1622 (n_579, n_1502, A[13]);
  nand g1624 (n_1504, A[13], A[16]);
  nand g1626 (n_586, n_984, n_1504, n_773);
  xor g1627 (n_1506, n_578, n_579);
  xor g1628 (n_581, n_1506, A[19]);
  nand g1629 (n_1507, n_578, n_579);
  nand g1630 (n_1508, A[19], n_579);
  nand g1631 (n_1509, n_578, A[19]);
  nand g1632 (n_588, n_1507, n_1508, n_1509);
  xor g1633 (n_1510, A[20], n_580);
  xor g1634 (n_583, n_1510, n_581);
  nand g1635 (n_1511, A[20], n_580);
  nand g1636 (n_1512, n_581, n_580);
  nand g1637 (n_1513, A[20], n_581);
  nand g1638 (n_589, n_1511, n_1512, n_1513);
  xor g1639 (n_1514, n_582, n_583);
  xor g1640 (n_585, n_1514, A[23]);
  nand g1641 (n_1515, n_582, n_583);
  nand g1642 (n_1516, A[23], n_583);
  nand g1643 (n_1517, n_582, A[23]);
  nand g1644 (n_591, n_1515, n_1516, n_1517);
  xor g1646 (n_83, n_1518, n_585);
  nand g1648 (n_1520, n_585, n_584);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1652 (n_587, n_1334, n_586);
  nand g1654 (n_1524, n_586, A[17]);
  nand g1655 (n_1525, A[16], n_586);
  nand g1656 (n_595, n_1335, n_1524, n_1525);
  xor g1657 (n_1526, A[20], n_587);
  xor g1658 (n_590, n_1526, n_588);
  nand g1659 (n_1527, A[20], n_587);
  nand g1660 (n_1528, n_588, n_587);
  nand g1661 (n_1529, A[20], n_588);
  nand g1662 (n_597, n_1527, n_1528, n_1529);
  xor g1664 (n_592, n_1530, n_589);
  nand g1667 (n_1533, A[21], n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_81, n_1535, n_1536, n_1537);
  nand g1681 (n_1541, A[18], n_595);
  nand g1682 (n_603, n_1539, n_1540, n_1541);
  xor g1684 (n_598, n_1474, n_596);
  nand g1686 (n_1544, n_596, A[22]);
  nand g1687 (n_1545, A[21], n_596);
  nand g1688 (n_605, n_1077, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_33, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_80, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[17], A[19]);
  nand g1702 (n_608, n_889, n_1552, n_1553);
  xor g1703 (n_1554, n_603, n_604);
  xor g1704 (n_606, n_1554, A[22]);
  nand g1705 (n_1555, n_603, n_604);
  nand g1706 (n_1556, A[22], n_604);
  nand g1707 (n_1557, n_603, A[22]);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, A[23], n_605);
  xor g1710 (n_32, n_1558, n_606);
  nand g1711 (n_1559, A[23], n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, A[23], n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1715 (n_1562, A[19], A[18]);
  xor g1716 (n_609, n_1562, A[20]);
  nand g1720 (n_612, n_1397, n_925, n_1161);
  xor g1721 (n_1566, n_608, n_609);
  xor g1722 (n_611, n_1566, A[23]);
  nand g1723 (n_1567, n_608, n_609);
  nand g1724 (n_1568, A[23], n_609);
  nand g1725 (n_1569, n_608, A[23]);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1728 (n_79, n_1570, n_611);
  nand g1730 (n_1572, n_611, n_610);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1734 (n_613, n_1450, n_612);
  nand g1736 (n_1576, n_612, A[21]);
  nand g1737 (n_1577, A[20], n_612);
  nand g1738 (n_617, n_1451, n_1576, n_1577);
  xor g1740 (n_78, n_1578, n_614);
  nand g1742 (n_1580, n_614, n_613);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_617);
  nand g1752 (n_28, n_1583, n_1584, n_1585);
  nand g1759 (n_1589, A[21], A[23]);
  nand g1760 (n_27, n_1587, n_1588, n_1589);
  xor g1762 (n_75, n_1166, A[22]);
  nand g1766 (n_74, n_1167, n_1123, n_1593);
  nand g16 (n_1606, A[0], A[2]);
  xor g20 (Z[2], A[0], A[2]);
  nand g22 (n_1611, n_68, A[3]);
  nand g25 (n_1615, n_1611, n_1612, n_1613);
  xor g26 (n_1614, n_68, A[3]);
  nand g28 (n_1616, A[4], n_117);
  nand g29 (n_1617, A[4], n_1615);
  nand g30 (n_1618, n_117, n_1615);
  nand g31 (n_1620, n_1616, n_1617, n_1618);
  xor g32 (n_1619, A[4], n_117);
  xor g33 (Z[4], n_1615, n_1619);
  nand g34 (n_1621, A[5], n_116);
  nand g35 (n_1622, A[5], n_1620);
  nand g36 (n_1623, n_116, n_1620);
  nand g37 (n_1625, n_1621, n_1622, n_1623);
  xor g38 (n_1624, A[5], n_116);
  xor g39 (Z[5], n_1620, n_1624);
  nand g40 (n_1626, n_67, n_115);
  nand g41 (n_1627, n_67, n_1625);
  nand g42 (n_1628, n_115, n_1625);
  nand g43 (n_1630, n_1626, n_1627, n_1628);
  xor g44 (n_1629, n_67, n_115);
  xor g45 (Z[6], n_1625, n_1629);
  nand g46 (n_1631, n_66, n_114);
  nand g47 (n_1632, n_66, n_1630);
  nand g48 (n_1633, n_114, n_1630);
  nand g49 (n_1635, n_1631, n_1632, n_1633);
  xor g50 (n_1634, n_66, n_114);
  xor g51 (Z[7], n_1630, n_1634);
  nand g52 (n_1636, n_65, n_113);
  nand g53 (n_1637, n_65, n_1635);
  nand g54 (n_1638, n_113, n_1635);
  nand g55 (n_1640, n_1636, n_1637, n_1638);
  xor g56 (n_1639, n_65, n_113);
  xor g57 (Z[8], n_1635, n_1639);
  nand g58 (n_1641, n_64, n_112);
  nand g59 (n_1642, n_64, n_1640);
  nand g60 (n_1643, n_112, n_1640);
  nand g61 (n_1645, n_1641, n_1642, n_1643);
  xor g62 (n_1644, n_64, n_112);
  xor g63 (Z[9], n_1640, n_1644);
  nand g64 (n_1646, n_63, n_111);
  nand g65 (n_1647, n_63, n_1645);
  nand g66 (n_1648, n_111, n_1645);
  nand g67 (n_1650, n_1646, n_1647, n_1648);
  xor g68 (n_1649, n_63, n_111);
  xor g69 (Z[10], n_1645, n_1649);
  nand g70 (n_1651, n_62, n_110);
  nand g71 (n_1652, n_62, n_1650);
  nand g72 (n_1653, n_110, n_1650);
  nand g73 (n_1655, n_1651, n_1652, n_1653);
  xor g74 (n_1654, n_62, n_110);
  xor g75 (Z[11], n_1650, n_1654);
  nand g76 (n_1656, n_61, n_109);
  nand g77 (n_1657, n_61, n_1655);
  nand g78 (n_1658, n_109, n_1655);
  nand g79 (n_1660, n_1656, n_1657, n_1658);
  xor g80 (n_1659, n_61, n_109);
  xor g81 (Z[12], n_1655, n_1659);
  nand g82 (n_1661, n_60, n_108);
  nand g83 (n_1662, n_60, n_1660);
  nand g84 (n_1663, n_108, n_1660);
  nand g85 (n_1665, n_1661, n_1662, n_1663);
  xor g86 (n_1664, n_60, n_108);
  xor g87 (Z[13], n_1660, n_1664);
  nand g88 (n_1666, n_59, n_107);
  nand g89 (n_1667, n_59, n_1665);
  nand g90 (n_1668, n_107, n_1665);
  nand g91 (n_1670, n_1666, n_1667, n_1668);
  xor g92 (n_1669, n_59, n_107);
  xor g93 (Z[14], n_1665, n_1669);
  nand g94 (n_1671, n_58, n_106);
  nand g95 (n_1672, n_58, n_1670);
  nand g96 (n_1673, n_106, n_1670);
  nand g97 (n_1675, n_1671, n_1672, n_1673);
  xor g98 (n_1674, n_58, n_106);
  xor g99 (Z[15], n_1670, n_1674);
  nand g100 (n_1676, n_57, n_105);
  nand g101 (n_1677, n_57, n_1675);
  nand g102 (n_1678, n_105, n_1675);
  nand g103 (n_1680, n_1676, n_1677, n_1678);
  xor g104 (n_1679, n_57, n_105);
  xor g105 (Z[16], n_1675, n_1679);
  nand g106 (n_1681, n_56, n_104);
  nand g107 (n_1682, n_56, n_1680);
  nand g108 (n_1683, n_104, n_1680);
  nand g109 (n_1685, n_1681, n_1682, n_1683);
  xor g110 (n_1684, n_56, n_104);
  xor g111 (Z[17], n_1680, n_1684);
  nand g112 (n_1686, n_55, n_103);
  nand g113 (n_1687, n_55, n_1685);
  nand g114 (n_1688, n_103, n_1685);
  nand g115 (n_1690, n_1686, n_1687, n_1688);
  xor g116 (n_1689, n_55, n_103);
  xor g117 (Z[18], n_1685, n_1689);
  nand g118 (n_1691, n_54, n_102);
  nand g119 (n_1692, n_54, n_1690);
  nand g120 (n_1693, n_102, n_1690);
  nand g121 (n_1695, n_1691, n_1692, n_1693);
  xor g122 (n_1694, n_54, n_102);
  xor g123 (Z[19], n_1690, n_1694);
  nand g124 (n_1696, n_53, n_101);
  nand g125 (n_1697, n_53, n_1695);
  nand g126 (n_1698, n_101, n_1695);
  nand g127 (n_1700, n_1696, n_1697, n_1698);
  xor g128 (n_1699, n_53, n_101);
  xor g129 (Z[20], n_1695, n_1699);
  nand g130 (n_1701, n_52, n_100);
  nand g131 (n_1702, n_52, n_1700);
  nand g132 (n_1703, n_100, n_1700);
  nand g133 (n_1705, n_1701, n_1702, n_1703);
  xor g134 (n_1704, n_52, n_100);
  xor g135 (Z[21], n_1700, n_1704);
  nand g136 (n_1706, n_51, n_99);
  nand g137 (n_1707, n_51, n_1705);
  nand g138 (n_1708, n_99, n_1705);
  nand g139 (n_1710, n_1706, n_1707, n_1708);
  xor g140 (n_1709, n_51, n_99);
  xor g141 (Z[22], n_1705, n_1709);
  nand g142 (n_1711, n_50, n_98);
  nand g143 (n_1712, n_50, n_1710);
  nand g144 (n_1713, n_98, n_1710);
  nand g145 (n_1715, n_1711, n_1712, n_1713);
  xor g146 (n_1714, n_50, n_98);
  xor g147 (Z[23], n_1710, n_1714);
  nand g148 (n_1716, n_49, n_97);
  nand g149 (n_1717, n_49, n_1715);
  nand g150 (n_1718, n_97, n_1715);
  nand g151 (n_1720, n_1716, n_1717, n_1718);
  xor g152 (n_1719, n_49, n_97);
  xor g153 (Z[24], n_1715, n_1719);
  nand g154 (n_1721, n_48, n_96);
  nand g155 (n_1722, n_48, n_1720);
  nand g156 (n_1723, n_96, n_1720);
  nand g157 (n_1725, n_1721, n_1722, n_1723);
  xor g158 (n_1724, n_48, n_96);
  xor g159 (Z[25], n_1720, n_1724);
  nand g160 (n_1726, n_47, n_95);
  nand g161 (n_1727, n_47, n_1725);
  nand g162 (n_1728, n_95, n_1725);
  nand g163 (n_1730, n_1726, n_1727, n_1728);
  xor g164 (n_1729, n_47, n_95);
  xor g165 (Z[26], n_1725, n_1729);
  nand g166 (n_1731, n_46, n_94);
  nand g167 (n_1732, n_46, n_1730);
  nand g168 (n_1733, n_94, n_1730);
  nand g169 (n_1735, n_1731, n_1732, n_1733);
  xor g170 (n_1734, n_46, n_94);
  xor g171 (Z[27], n_1730, n_1734);
  nand g172 (n_1736, n_45, n_93);
  nand g173 (n_1737, n_45, n_1735);
  nand g174 (n_1738, n_93, n_1735);
  nand g175 (n_1740, n_1736, n_1737, n_1738);
  xor g176 (n_1739, n_45, n_93);
  xor g177 (Z[28], n_1735, n_1739);
  nand g178 (n_1741, n_44, n_92);
  nand g179 (n_1742, n_44, n_1740);
  nand g180 (n_1743, n_92, n_1740);
  nand g181 (n_1745, n_1741, n_1742, n_1743);
  xor g182 (n_1744, n_44, n_92);
  xor g183 (Z[29], n_1740, n_1744);
  nand g184 (n_1746, n_43, n_91);
  nand g185 (n_1747, n_43, n_1745);
  nand g186 (n_1748, n_91, n_1745);
  nand g187 (n_1750, n_1746, n_1747, n_1748);
  xor g188 (n_1749, n_43, n_91);
  xor g189 (Z[30], n_1745, n_1749);
  nand g190 (n_1751, n_42, n_90);
  nand g191 (n_1752, n_42, n_1750);
  nand g192 (n_1753, n_90, n_1750);
  nand g193 (n_1755, n_1751, n_1752, n_1753);
  xor g194 (n_1754, n_42, n_90);
  xor g195 (Z[31], n_1750, n_1754);
  nand g196 (n_1756, n_41, n_89);
  nand g197 (n_1757, n_41, n_1755);
  nand g198 (n_1758, n_89, n_1755);
  nand g199 (n_1760, n_1756, n_1757, n_1758);
  xor g200 (n_1759, n_41, n_89);
  xor g201 (Z[32], n_1755, n_1759);
  nand g202 (n_1761, n_40, n_88);
  nand g203 (n_1762, n_40, n_1760);
  nand g204 (n_1763, n_88, n_1760);
  nand g205 (n_1765, n_1761, n_1762, n_1763);
  xor g206 (n_1764, n_40, n_88);
  xor g207 (Z[33], n_1760, n_1764);
  nand g208 (n_1766, n_39, n_87);
  nand g209 (n_1767, n_39, n_1765);
  nand g210 (n_1768, n_87, n_1765);
  nand g211 (n_1770, n_1766, n_1767, n_1768);
  xor g212 (n_1769, n_39, n_87);
  xor g213 (Z[34], n_1765, n_1769);
  nand g214 (n_1771, n_38, n_86);
  nand g215 (n_1772, n_38, n_1770);
  nand g216 (n_1773, n_86, n_1770);
  nand g217 (n_1775, n_1771, n_1772, n_1773);
  xor g218 (n_1774, n_38, n_86);
  xor g219 (Z[35], n_1770, n_1774);
  nand g220 (n_1776, n_37, n_85);
  nand g221 (n_1777, n_37, n_1775);
  nand g222 (n_1778, n_85, n_1775);
  nand g223 (n_1780, n_1776, n_1777, n_1778);
  xor g224 (n_1779, n_37, n_85);
  xor g225 (Z[36], n_1775, n_1779);
  nand g226 (n_1781, n_36, n_84);
  nand g227 (n_1782, n_36, n_1780);
  nand g228 (n_1783, n_84, n_1780);
  nand g229 (n_1785, n_1781, n_1782, n_1783);
  xor g230 (n_1784, n_36, n_84);
  xor g231 (Z[37], n_1780, n_1784);
  nand g232 (n_1786, n_35, n_83);
  nand g233 (n_1787, n_35, n_1785);
  nand g234 (n_1788, n_83, n_1785);
  nand g235 (n_1790, n_1786, n_1787, n_1788);
  xor g236 (n_1789, n_35, n_83);
  xor g237 (Z[38], n_1785, n_1789);
  nand g238 (n_1791, n_34, n_82);
  nand g239 (n_1792, n_34, n_1790);
  nand g240 (n_1793, n_82, n_1790);
  nand g241 (n_1795, n_1791, n_1792, n_1793);
  xor g242 (n_1794, n_34, n_82);
  xor g243 (Z[39], n_1790, n_1794);
  nand g244 (n_1796, n_33, n_81);
  nand g245 (n_1797, n_33, n_1795);
  nand g246 (n_1798, n_81, n_1795);
  nand g247 (n_1800, n_1796, n_1797, n_1798);
  xor g248 (n_1799, n_33, n_81);
  xor g249 (Z[40], n_1795, n_1799);
  nand g250 (n_1801, n_32, n_80);
  nand g251 (n_1802, n_32, n_1800);
  nand g252 (n_1803, n_80, n_1800);
  nand g253 (n_1805, n_1801, n_1802, n_1803);
  xor g254 (n_1804, n_32, n_80);
  xor g255 (Z[41], n_1800, n_1804);
  nand g256 (n_1806, n_31, n_79);
  nand g257 (n_1807, n_31, n_1805);
  nand g258 (n_1808, n_79, n_1805);
  nand g259 (n_1810, n_1806, n_1807, n_1808);
  xor g260 (n_1809, n_31, n_79);
  xor g261 (Z[42], n_1805, n_1809);
  nand g262 (n_1811, n_30, n_78);
  nand g263 (n_1812, n_30, n_1810);
  nand g264 (n_1813, n_78, n_1810);
  nand g265 (n_1815, n_1811, n_1812, n_1813);
  xor g266 (n_1814, n_30, n_78);
  xor g267 (Z[43], n_1810, n_1814);
  nand g1772 (n_1816, n_29, n_77);
  nand g1773 (n_1817, n_29, n_1815);
  nand g1774 (n_1818, n_77, n_1815);
  nand g1775 (n_1820, n_1816, n_1817, n_1818);
  xor g1776 (n_1819, n_29, n_77);
  xor g1777 (Z[44], n_1815, n_1819);
  nand g1778 (n_1821, n_28, n_76);
  nand g1779 (n_1822, n_28, n_1820);
  nand g1780 (n_1823, n_76, n_1820);
  nand g1781 (n_1825, n_1821, n_1822, n_1823);
  xor g1782 (n_1824, n_28, n_76);
  xor g1783 (Z[45], n_1820, n_1824);
  nand g1784 (n_1826, n_27, n_75);
  nand g1785 (n_1827, n_27, n_1825);
  nand g1786 (n_1828, n_75, n_1825);
  nand g1787 (n_1830, n_1826, n_1827, n_1828);
  xor g1788 (n_1829, n_27, n_75);
  xor g1789 (Z[46], n_1825, n_1829);
  xor g1791 (Z[47], n_1830, n_1831);
  or g1803 (n_1043, A[1], wc);
  not gc (wc, n_171);
  or g1804 (n_1044, A[1], wc0);
  not gc0 (wc0, A[2]);
  xnor g1806 (n_1166, A[24], A[23]);
  or g1807 (n_1167, wc1, A[24]);
  not gc1 (wc1, A[23]);
  xnor g1808 (n_1214, A[6], A[5]);
  or g1809 (n_1215, A[5], wc2);
  not gc2 (wc2, A[6]);
  or g1810 (n_1252, A[6], wc3);
  not gc3 (wc3, A[7]);
  or g1811 (n_1253, wc4, A[6]);
  not gc4 (wc4, A[5]);
  or g1813 (n_1355, A[9], wc5);
  not gc5 (wc5, A[10]);
  or g1814 (n_1384, wc6, A[10]);
  not gc6 (wc6, A[9]);
  or g1815 (n_1385, A[10], wc7);
  not gc7 (wc7, A[11]);
  or g1817 (n_1463, A[13], wc8);
  not gc8 (wc8, A[14]);
  xnor g1818 (n_1530, A[24], A[21]);
  or g1819 (n_1531, wc9, A[24]);
  not gc9 (wc9, A[21]);
  or g1821 (n_1539, A[17], wc10);
  not gc10 (wc10, A[18]);
  or g1822 (n_1552, A[18], wc11);
  not gc11 (wc11, A[19]);
  or g1823 (n_1553, wc12, A[18]);
  not gc12 (wc12, A[17]);
  or g1825 (n_1583, A[21], wc13);
  not gc13 (wc13, A[22]);
  or g1826 (n_1587, wc14, A[22]);
  not gc14 (wc14, A[21]);
  or g1827 (n_1588, A[22], wc15);
  not gc15 (wc15, A[23]);
  or g1828 (n_1593, wc16, A[24]);
  not gc16 (wc16, A[22]);
  xnor g1830 (n_372, n_626, A[1]);
  or g1831 (n_1088, A[1], wc17);
  not gc17 (wc17, A[3]);
  xnor g1832 (n_453, n_1250, A[6]);
  xnor g1833 (n_519, n_1382, A[10]);
  xnor g1834 (n_569, n_1106, A[13]);
  or g1835 (n_1484, A[13], wc18);
  not gc18 (wc18, A[15]);
  xnor g1836 (n_604, n_1550, A[18]);
  xnor g1837 (n_76, n_1474, A[23]);
  or g1839 (n_1047, wc19, n_117);
  not gc19 (wc19, A[5]);
  or g1840 (n_1049, wc20, n_117);
  not gc20 (wc20, n_179);
  xnor g1842 (n_1578, n_613, A[24]);
  or g1843 (n_1579, A[24], wc21);
  not gc21 (wc21, n_613);
  xnor g1844 (n_1831, n_74, A[24]);
  or g1846 (n_1051, wc22, n_180);
  not gc22 (wc22, A[6]);
  or g1847 (n_1052, wc23, n_180);
  not gc23 (wc23, A[9]);
  xnor g1848 (n_505, n_1218, n_503);
  or g1849 (n_1356, A[9], wc24);
  not gc24 (wc24, n_503);
  xnor g1850 (n_558, n_1358, n_557);
  or g1851 (n_1464, A[13], wc25);
  not gc25 (wc25, n_557);
  or g1852 (n_1573, A[24], wc26);
  not gc26 (wc26, n_611);
  or g1853 (n_1581, A[24], wc27);
  not gc27 (wc27, n_614);
  xnor g1854 (n_29, n_1474, n_617);
  or g1855 (n_1584, A[21], wc28);
  not gc28 (wc28, n_617);
  or g1858 (n_1216, A[5], wc29);
  not gc29 (wc29, n_433);
  xnor g1859 (n_596, n_1466, n_595);
  or g1860 (n_1540, A[17], wc30);
  not gc30 (wc30, n_595);
  or g1861 (n_1612, n_1606, wc31);
  not gc31 (wc31, n_68);
  or g1862 (n_1613, wc32, n_1606);
  not gc32 (wc32, A[3]);
  xnor g1863 (Z[3], n_1606, n_1614);
  xnor g1864 (n_355, n_202, n_906);
  or g1865 (n_1056, wc33, n_202);
  not gc33 (wc33, n_282);
  or g1866 (n_1057, wc34, n_202);
  not gc34 (wc34, A[10]);
  xnor g1867 (n_1570, n_610, A[24]);
  or g1868 (n_1571, A[24], wc35);
  not gc35 (wc35, n_610);
  or g1869 (n_1532, A[24], wc36);
  not gc36 (wc36, n_589);
  xnor g1870 (n_1518, n_584, A[24]);
  or g1871 (n_1519, A[24], wc37);
  not gc37 (wc37, n_584);
  xnor g1872 (n_1454, n_550, A[24]);
  or g1873 (n_1455, A[24], wc38);
  not gc38 (wc38, n_550);
  or g1874 (n_1521, A[24], wc39);
  not gc39 (wc39, n_585);
  or g1875 (n_1081, A[24], wc40);
  not gc40 (wc40, n_363);
  xnor g1876 (n_1206, n_426, A[24]);
  or g1877 (n_1207, A[24], wc41);
  not gc41 (wc41, n_426);
  xnor g1878 (n_1346, n_496, A[24]);
  or g1879 (n_1347, A[24], wc42);
  not gc42 (wc42, n_496);
  or g1880 (n_1456, A[24], wc43);
  not gc43 (wc43, n_551);
  or g1881 (n_1080, A[24], wc44);
  not gc44 (wc44, n_364);
  xnor g1882 (n_367, n_1078, A[24]);
  or g1883 (n_1348, A[24], wc45);
  not gc45 (wc45, n_497);
  or g1884 (n_1168, A[24], wc46);
  not gc46 (wc46, n_408);
  or g1885 (n_1208, A[24], wc47);
  not gc47 (wc47, n_427);
  or g1886 (n_1316, A[24], wc48);
  not gc48 (wc48, n_482);
  or g1887 (n_1432, A[24], wc49);
  not gc49 (wc49, n_540);
endmodule

module mult_signed_const_5487_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_5487_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_5754_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_176;
  wire n_179, n_180, n_183, n_184, n_187, n_188, n_189, n_196;
  wire n_201, n_202, n_203, n_204, n_209, n_210, n_211, n_212;
  wire n_217, n_218, n_219, n_220, n_221, n_223, n_224, n_225;
  wire n_226, n_227, n_234, n_236, n_237, n_238, n_239, n_248;
  wire n_249, n_250, n_251, n_258, n_260, n_261, n_262, n_267;
  wire n_269, n_271, n_272, n_273, n_274, n_275, n_276, n_277;
  wire n_282, n_284, n_285, n_286, n_287, n_288, n_289, n_290;
  wire n_291, n_292, n_293, n_300, n_302, n_303, n_304, n_305;
  wire n_306, n_307, n_308, n_309, n_319, n_320, n_321, n_322;
  wire n_323, n_324, n_325, n_326, n_333, n_335, n_337, n_338;
  wire n_339, n_340, n_341, n_342, n_343, n_344, n_345, n_354;
  wire n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363;
  wire n_364, n_365, n_366, n_367, n_371, n_372, n_373, n_374;
  wire n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382;
  wire n_383, n_384, n_385, n_386, n_387, n_388, n_389, n_390;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407;
  wire n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415;
  wire n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423;
  wire n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_433;
  wire n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441;
  wire n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449;
  wire n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460;
  wire n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468;
  wire n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477;
  wire n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485;
  wire n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493;
  wire n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_503;
  wire n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511;
  wire n_512, n_513, n_514, n_515, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539;
  wire n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547;
  wire n_548, n_549, n_550, n_551, n_552, n_553, n_554, n_557;
  wire n_558, n_559, n_560, n_561, n_562, n_563, n_564, n_565;
  wire n_569, n_570, n_571, n_572, n_573, n_574, n_575, n_576;
  wire n_578, n_579, n_580, n_581, n_582, n_583, n_584, n_585;
  wire n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_595;
  wire n_596, n_597, n_598, n_599, n_603, n_604, n_605, n_606;
  wire n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_617;
  wire n_622, n_623, n_624, n_625, n_626, n_627, n_628, n_629;
  wire n_630, n_631, n_632, n_633, n_634, n_635, n_636, n_637;
  wire n_638, n_639, n_640, n_641, n_646, n_647, n_648, n_649;
  wire n_650, n_651, n_652, n_653, n_658, n_659, n_660, n_661;
  wire n_662, n_663, n_664, n_665, n_668, n_669, n_670, n_671;
  wire n_672, n_673, n_674, n_675, n_676, n_677, n_684, n_685;
  wire n_686, n_687, n_688, n_689, n_690, n_691, n_692, n_693;
  wire n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711;
  wire n_712, n_713, n_722, n_724, n_725, n_726, n_727, n_728;
  wire n_729, n_730, n_731, n_732, n_733, n_738, n_742, n_743;
  wire n_744, n_745, n_746, n_747, n_748, n_749, n_750, n_751;
  wire n_752, n_753, n_764, n_765, n_766, n_767, n_768, n_769;
  wire n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777;
  wire n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801;
  wire n_802, n_803, n_804, n_805, n_822, n_823, n_824, n_826;
  wire n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_842;
  wire n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855;
  wire n_856, n_857, n_858, n_859, n_860, n_861, n_868, n_869;
  wire n_870, n_871, n_872, n_873, n_876, n_877, n_880, n_881;
  wire n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889;
  wire n_890, n_891, n_892, n_893, n_906, n_907, n_908, n_910;
  wire n_911, n_912, n_913, n_914, n_915, n_916, n_917, n_918;
  wire n_919, n_920, n_921, n_922, n_923, n_924, n_925, n_926;
  wire n_927, n_928, n_929, n_946, n_947, n_949, n_950, n_951;
  wire n_952, n_953, n_954, n_955, n_956, n_957, n_958, n_959;
  wire n_960, n_961, n_962, n_963, n_964, n_965, n_984, n_985;
  wire n_986, n_987, n_988, n_989, n_990, n_991, n_992, n_993;
  wire n_994, n_995, n_996, n_997, n_998, n_999, n_1000, n_1001;
  wire n_1013, n_1014, n_1015, n_1016, n_1017, n_1020, n_1021, n_1024;
  wire n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040;
  wire n_1041, n_1043, n_1044, n_1047, n_1049, n_1051, n_1052, n_1056;
  wire n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064;
  wire n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072;
  wire n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080;
  wire n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1088, n_1090;
  wire n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098;
  wire n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106;
  wire n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114;
  wire n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122;
  wire n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130;
  wire n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138;
  wire n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146;
  wire n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1154, n_1155;
  wire n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163;
  wire n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171;
  wire n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179;
  wire n_1180, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188;
  wire n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196;
  wire n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204;
  wire n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212;
  wire n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220;
  wire n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228;
  wire n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236;
  wire n_1237, n_1238, n_1239, n_1241, n_1242, n_1243, n_1244, n_1245;
  wire n_1246, n_1247, n_1248, n_1249, n_1250, n_1252, n_1253, n_1254;
  wire n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262;
  wire n_1263, n_1264, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271;
  wire n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279;
  wire n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1288;
  wire n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297;
  wire n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305;
  wire n_1306, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1316;
  wire n_1317, n_1318, n_1319, n_1320, n_1321, n_1324, n_1325, n_1326;
  wire n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334;
  wire n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342;
  wire n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350;
  wire n_1351, n_1352, n_1353, n_1355, n_1356, n_1357, n_1358, n_1359;
  wire n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367;
  wire n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375;
  wire n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383;
  wire n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391;
  wire n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399;
  wire n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407;
  wire n_1408, n_1409, n_1410, n_1412, n_1414, n_1415, n_1416, n_1417;
  wire n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1426;
  wire n_1427, n_1428, n_1429, n_1432, n_1433, n_1434, n_1435, n_1436;
  wire n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444;
  wire n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453;
  wire n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461;
  wire n_1463, n_1464, n_1465, n_1466, n_1468, n_1469, n_1470, n_1471;
  wire n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479;
  wire n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487;
  wire n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495;
  wire n_1496, n_1498, n_1499, n_1500, n_1501, n_1502, n_1506, n_1507;
  wire n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515;
  wire n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1524, n_1525;
  wire n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533;
  wire n_1534, n_1535, n_1536, n_1537, n_1539, n_1540, n_1541, n_1542;
  wire n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1552;
  wire n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560;
  wire n_1561, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572;
  wire n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580;
  wire n_1581, n_1583, n_1584, n_1585, n_1587, n_1588, n_1589, n_1593;
  wire n_1606, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617;
  wire n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625;
  wire n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633;
  wire n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641;
  wire n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649;
  wire n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657;
  wire n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665;
  wire n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673;
  wire n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681;
  wire n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689;
  wire n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697;
  wire n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705;
  wire n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713;
  wire n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721;
  wire n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729;
  wire n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737;
  wire n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745;
  wire n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753;
  wire n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761;
  wire n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769;
  wire n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777;
  wire n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785;
  wire n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793;
  wire n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801;
  wire n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809;
  wire n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817;
  wire n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825;
  wire n_1826, n_1827, n_1828, n_1829, n_1830, n_1831;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], n_171);
  xor g270 (n_117, n_622, A[2]);
  nand g3 (n_623, A[1], n_171);
  nand g271 (n_624, A[2], n_171);
  nand g272 (n_625, A[1], A[2]);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, A[4]);
  xor g288 (n_176, n_634, n_69);
  nand g289 (n_635, n_68, A[4]);
  nand g290 (n_636, n_69, A[4]);
  nand g291 (n_637, n_68, n_69);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_176);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_176);
  nand g296 (n_640, A[7], n_176);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g305 (n_646, n_117, A[5]);
  xor g306 (n_180, n_646, A[6]);
  nand g307 (n_647, n_117, A[5]);
  nand g308 (n_648, A[6], A[5]);
  nand g309 (n_649, n_117, A[6]);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, n_179, n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, n_179, n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, n_179, A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_188, n_659, n_660, n_661);
  xor g329 (n_662, n_183, A[9]);
  xor g330 (n_112, n_662, n_184);
  nand g331 (n_663, n_183, A[9]);
  nand g332 (n_664, n_184, A[9]);
  nand g333 (n_665, n_183, n_184);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_187, n_630, n_67);
  nand g340 (n_668, n_67, n_173);
  nand g341 (n_669, A[4], n_67);
  nand g342 (n_71, n_631, n_668, n_669);
  xor g343 (n_670, A[7], n_187);
  xor g344 (n_189, n_670, A[8]);
  nand g345 (n_671, A[7], n_187);
  nand g346 (n_672, A[8], n_187);
  nand g347 (n_673, A[7], A[8]);
  nand g348 (n_73, n_671, n_672, n_673);
  xor g349 (n_674, n_188, A[10]);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, n_188, A[10]);
  nand g352 (n_676, n_189, A[10]);
  nand g353 (n_677, n_188, n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_72, n_638, n_71);
  nand g366 (n_684, n_71, n_176);
  nand g367 (n_685, A[5], n_71);
  nand g368 (n_201, n_639, n_684, n_685);
  xor g369 (n_686, A[8], A[9]);
  xor g370 (n_196, n_686, n_73);
  nand g371 (n_687, A[8], A[9]);
  nand g372 (n_688, n_73, A[9]);
  nand g373 (n_689, A[8], n_73);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, n_72, A[11]);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, n_72, A[11]);
  nand g378 (n_692, n_196, A[11]);
  nand g379 (n_693, n_72, n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g394 (n_202, n_650, A[9]);
  nand g396 (n_704, A[9], n_180);
  nand g397 (n_705, n_179, A[9]);
  nand g398 (n_209, n_651, n_704, n_705);
  xor g399 (n_706, A[10], n_201);
  xor g400 (n_204, n_706, n_202);
  nand g401 (n_707, A[10], n_201);
  nand g402 (n_708, n_202, n_201);
  nand g403 (n_709, A[10], n_202);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, A[12], n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, A[12], n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, A[12], n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g423 (n_722, n_183, n_184);
  xor g424 (n_210, n_722, A[10]);
  nand g426 (n_724, A[10], n_184);
  nand g427 (n_725, n_183, A[10]);
  nand g428 (n_218, n_665, n_724, n_725);
  xor g429 (n_726, A[11], n_209);
  xor g430 (n_212, n_726, n_210);
  nand g431 (n_727, A[11], n_209);
  nand g432 (n_728, n_210, n_209);
  nand g433 (n_729, A[11], n_210);
  nand g434 (n_220, n_727, n_728, n_729);
  xor g435 (n_730, n_211, A[13]);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, n_211, A[13]);
  nand g438 (n_732, n_212, A[13]);
  nand g439 (n_733, n_211, n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_217, n_738, n_187);
  xor g455 (n_742, n_188, n_217);
  xor g456 (n_219, n_742, A[11]);
  nand g457 (n_743, n_188, n_217);
  nand g458 (n_744, A[11], n_217);
  nand g459 (n_745, n_188, A[11]);
  nand g460 (n_224, n_743, n_744, n_745);
  xor g461 (n_746, A[12], n_218);
  xor g462 (n_221, n_746, A[14]);
  nand g463 (n_747, A[12], n_218);
  nand g464 (n_748, A[14], n_218);
  nand g465 (n_749, A[12], A[14]);
  nand g466 (n_226, n_747, n_748, n_749);
  xor g467 (n_750, n_219, n_220);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, n_219, n_220);
  nand g470 (n_752, n_221, n_220);
  nand g471 (n_753, n_219, n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g488 (n_223, n_686, n_72);
  nand g490 (n_764, n_72, A[9]);
  nand g491 (n_765, A[8], n_72);
  nand g492 (n_234, n_687, n_764, n_765);
  xor g493 (n_766, n_73, A[12]);
  xor g494 (n_225, n_766, n_223);
  nand g495 (n_767, n_73, A[12]);
  nand g496 (n_768, n_223, A[12]);
  nand g497 (n_769, n_73, n_223);
  nand g498 (n_236, n_767, n_768, n_769);
  xor g499 (n_770, A[13], n_224);
  xor g500 (n_227, n_770, n_225);
  nand g501 (n_771, A[13], n_224);
  nand g502 (n_772, n_225, n_224);
  nand g503 (n_773, A[13], n_225);
  nand g504 (n_238, n_771, n_772, n_773);
  xor g505 (n_774, A[15], n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, A[15], n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, A[15], n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g535 (n_794, n_234, A[13]);
  xor g536 (n_237, n_794, n_204);
  nand g537 (n_795, n_234, A[13]);
  nand g538 (n_796, n_204, A[13]);
  nand g539 (n_797, n_234, n_204);
  nand g540 (n_248, n_795, n_796, n_797);
  xor g541 (n_798, A[14], n_236);
  xor g542 (n_239, n_798, A[16]);
  nand g543 (n_799, A[14], n_236);
  nand g544 (n_800, A[16], n_236);
  nand g545 (n_801, A[14], A[16]);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, n_237, n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, n_237, n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, n_237, n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g577 (n_822, n_211, A[14]);
  xor g578 (n_249, n_822, n_212);
  nand g579 (n_823, n_211, A[14]);
  nand g580 (n_824, n_212, A[14]);
  nand g582 (n_261, n_823, n_824, n_733);
  xor g583 (n_826, A[15], n_248);
  xor g584 (n_251, n_826, A[17]);
  nand g585 (n_827, A[15], n_248);
  nand g586 (n_828, A[17], n_248);
  nand g587 (n_829, A[15], A[17]);
  nand g588 (n_118, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g609 (n_842, n_188, A[11]);
  xor g610 (n_258, n_842, n_217);
  xor g616 (n_260, n_746, n_258);
  nand g618 (n_848, n_258, n_218);
  nand g619 (n_849, A[12], n_258);
  nand g620 (n_272, n_747, n_848, n_849);
  xor g621 (n_850, n_220, A[15]);
  xor g622 (n_262, n_850, n_260);
  nand g623 (n_851, n_220, A[15]);
  nand g624 (n_852, n_260, A[15]);
  nand g625 (n_853, n_220, n_260);
  nand g626 (n_274, n_851, n_852, n_853);
  xor g627 (n_854, A[16], n_261);
  xor g628 (n_119, n_854, A[18]);
  nand g629 (n_855, A[16], n_261);
  nand g630 (n_856, A[18], n_261);
  nand g631 (n_857, A[16], A[18]);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_262, n_118);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_262, n_118);
  nand g636 (n_860, n_119, n_118);
  nand g637 (n_861, n_262, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g648 (n_267, n_638, A[8]);
  nand g650 (n_868, A[8], n_176);
  nand g651 (n_869, A[5], A[8]);
  nand g652 (n_282, n_639, n_868, n_869);
  xor g653 (n_870, n_71, A[9]);
  xor g654 (n_269, n_870, n_267);
  nand g655 (n_871, n_71, A[9]);
  nand g656 (n_872, n_267, A[9]);
  nand g657 (n_873, n_71, n_267);
  nand g658 (n_284, n_871, n_872, n_873);
  xor g660 (n_271, n_766, n_269);
  nand g662 (n_876, n_269, A[12]);
  nand g663 (n_877, n_73, n_269);
  nand g664 (n_286, n_767, n_876, n_877);
  xor g666 (n_273, n_770, n_271);
  nand g668 (n_880, n_271, A[13]);
  nand g669 (n_881, n_224, n_271);
  nand g670 (n_288, n_771, n_880, n_881);
  xor g671 (n_882, n_272, A[16]);
  xor g672 (n_275, n_882, n_273);
  nand g673 (n_883, n_272, A[16]);
  nand g674 (n_884, n_273, A[16]);
  nand g675 (n_885, n_272, n_273);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, A[17], n_274);
  xor g678 (n_277, n_886, A[19]);
  nand g679 (n_887, A[17], n_274);
  nand g680 (n_888, A[19], n_274);
  nand g681 (n_889, A[17], A[19]);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g707 (n_906, A[10], n_282);
  xor g708 (n_285, n_906, n_202);
  nand g709 (n_907, A[10], n_282);
  nand g710 (n_908, n_202, n_282);
  nand g712 (n_300, n_907, n_908, n_709);
  xor g713 (n_910, n_284, A[13]);
  xor g714 (n_287, n_910, n_285);
  nand g715 (n_911, n_284, A[13]);
  nand g716 (n_912, n_285, A[13]);
  nand g717 (n_913, n_284, n_285);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, A[14], n_286);
  xor g720 (n_289, n_914, n_287);
  nand g721 (n_915, A[14], n_286);
  nand g722 (n_916, n_287, n_286);
  nand g723 (n_917, A[14], n_287);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, n_288, A[17]);
  xor g726 (n_291, n_918, n_289);
  nand g727 (n_919, n_288, A[17]);
  nand g728 (n_920, n_289, A[17]);
  nand g729 (n_921, n_288, n_289);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, A[18], n_290);
  xor g732 (n_293, n_922, A[20]);
  nand g733 (n_923, A[18], n_290);
  nand g734 (n_924, A[20], n_290);
  nand g735 (n_925, A[18], A[20]);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g767 (n_946, n_300, A[14]);
  xor g768 (n_303, n_946, n_212);
  nand g769 (n_947, n_300, A[14]);
  nand g771 (n_949, n_300, n_212);
  nand g772 (n_319, n_947, n_824, n_949);
  xor g773 (n_950, n_302, A[15]);
  xor g774 (n_305, n_950, n_303);
  nand g775 (n_951, n_302, A[15]);
  nand g776 (n_952, n_303, A[15]);
  nand g777 (n_953, n_302, n_303);
  nand g778 (n_321, n_951, n_952, n_953);
  xor g779 (n_954, n_304, A[18]);
  xor g780 (n_307, n_954, n_305);
  nand g781 (n_955, n_304, A[18]);
  nand g782 (n_956, n_305, A[18]);
  nand g783 (n_957, n_304, n_305);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, A[19], n_306);
  xor g786 (n_309, n_958, A[21]);
  nand g787 (n_959, A[19], n_306);
  nand g788 (n_960, A[21], n_306);
  nand g789 (n_961, A[19], A[21]);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g824 (n_320, n_850, A[16]);
  nand g826 (n_984, A[16], A[15]);
  nand g827 (n_985, n_220, A[16]);
  nand g828 (n_338, n_851, n_984, n_985);
  xor g829 (n_986, n_260, n_319);
  xor g830 (n_322, n_986, n_320);
  nand g831 (n_987, n_260, n_319);
  nand g832 (n_988, n_320, n_319);
  nand g833 (n_989, n_260, n_320);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, n_321, A[19]);
  xor g836 (n_324, n_990, A[20]);
  nand g837 (n_991, n_321, A[19]);
  nand g838 (n_992, A[20], A[19]);
  nand g839 (n_993, n_321, A[20]);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, n_322, n_323);
  xor g842 (n_326, n_994, n_324);
  nand g843 (n_995, n_322, n_323);
  nand g844 (n_996, n_324, n_323);
  nand g845 (n_997, n_322, n_324);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, A[22], n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, A[22], n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, A[22], n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g868 (n_333, n_870, n_73);
  nand g871 (n_1013, n_71, n_73);
  nand g872 (n_354, n_871, n_688, n_1013);
  xor g873 (n_1014, n_267, A[12]);
  xor g874 (n_335, n_1014, n_333);
  nand g875 (n_1015, n_267, A[12]);
  nand g876 (n_1016, n_333, A[12]);
  nand g877 (n_1017, n_267, n_333);
  nand g878 (n_356, n_1015, n_1016, n_1017);
  xor g880 (n_337, n_770, n_335);
  nand g882 (n_1020, n_335, A[13]);
  nand g883 (n_1021, n_224, n_335);
  nand g884 (n_358, n_771, n_1020, n_1021);
  xor g886 (n_339, n_882, n_337);
  nand g888 (n_1024, n_337, A[16]);
  nand g889 (n_1025, n_272, n_337);
  nand g890 (n_360, n_883, n_1024, n_1025);
  xor g891 (n_1026, A[17], n_338);
  xor g892 (n_341, n_1026, n_339);
  nand g893 (n_1027, A[17], n_338);
  nand g894 (n_1028, n_339, n_338);
  nand g895 (n_1029, A[17], n_339);
  nand g896 (n_362, n_1027, n_1028, n_1029);
  xor g897 (n_1030, A[20], n_340);
  xor g898 (n_343, n_1030, n_341);
  nand g899 (n_1031, A[20], n_340);
  nand g900 (n_1032, n_341, n_340);
  nand g901 (n_1033, A[20], n_341);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, A[21], n_342);
  xor g904 (n_345, n_1034, n_343);
  nand g905 (n_1035, A[21], n_342);
  nand g906 (n_1036, n_343, n_342);
  nand g907 (n_1037, A[21], n_343);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, A[23], n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, A[23], n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, A[23], n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  nand g922 (n_371, n_1043, n_1044, n_624);
  nand g928 (n_373, n_1047, n_648, n_1049);
  nand g934 (n_375, n_1051, n_1052, n_705);
  nand g940 (n_377, n_907, n_1056, n_1057);
  xor g941 (n_1058, n_354, A[13]);
  nand g943 (n_1059, n_354, A[13]);
  nand g946 (n_379, n_1059, n_1060, n_1061);
  xor g947 (n_1062, A[14], n_356);
  xor g948 (n_359, n_1062, n_357);
  nand g949 (n_1063, A[14], n_356);
  nand g950 (n_1064, n_357, n_356);
  nand g951 (n_1065, A[14], n_357);
  nand g952 (n_381, n_1063, n_1064, n_1065);
  xor g953 (n_1066, n_358, A[17]);
  xor g954 (n_361, n_1066, A[18]);
  nand g955 (n_1067, n_358, A[17]);
  nand g956 (n_1068, A[18], A[17]);
  nand g957 (n_1069, n_358, A[18]);
  nand g958 (n_383, n_1067, n_1068, n_1069);
  xor g959 (n_1070, n_359, n_360);
  xor g960 (n_363, n_1070, n_361);
  nand g961 (n_1071, n_359, n_360);
  nand g962 (n_1072, n_361, n_360);
  nand g963 (n_1073, n_359, n_361);
  nand g964 (n_385, n_1071, n_1072, n_1073);
  xor g965 (n_1074, A[21], n_362);
  xor g966 (n_365, n_1074, A[22]);
  nand g967 (n_1075, A[21], n_362);
  nand g968 (n_1076, A[22], n_362);
  nand g969 (n_1077, A[21], A[22]);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g972 (n_367, n_1078, n_364);
  nand g975 (n_1081, n_363, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  xor g986 (n_372, n_1086, A[3]);
  nand g990 (n_392, n_1044, n_1088, n_627);
  xor g991 (n_1090, n_371, n_372);
  xor g992 (n_374, n_1090, A[6]);
  nand g993 (n_1091, n_371, n_372);
  nand g994 (n_1092, A[6], n_372);
  nand g995 (n_1093, n_371, A[6]);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, n_374);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, n_374, n_373);
  nand g1001 (n_1097, A[7], n_374);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, A[10], A[11]);
  xor g1004 (n_378, n_1098, n_375);
  nand g1005 (n_1099, A[10], A[11]);
  nand g1006 (n_1100, n_375, A[11]);
  nand g1007 (n_1101, A[10], n_375);
  nand g1008 (n_398, n_1099, n_1100, n_1101);
  xor g1009 (n_1102, n_376, n_377);
  xor g1010 (n_380, n_1102, n_378);
  nand g1011 (n_1103, n_376, n_377);
  nand g1012 (n_1104, n_378, n_377);
  nand g1013 (n_1105, n_376, n_378);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, A[14], n_379);
  xor g1016 (n_382, n_1106, A[15]);
  nand g1017 (n_1107, A[14], n_379);
  nand g1018 (n_1108, A[15], n_379);
  nand g1019 (n_1109, A[14], A[15]);
  nand g1020 (n_402, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, n_380, A[18]);
  xor g1022 (n_384, n_1110, n_381);
  nand g1023 (n_1111, n_380, A[18]);
  nand g1024 (n_1112, n_381, A[18]);
  nand g1025 (n_1113, n_380, n_381);
  nand g1026 (n_404, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, n_382, A[19]);
  xor g1028 (n_386, n_1114, n_383);
  nand g1029 (n_1115, n_382, A[19]);
  nand g1030 (n_1116, n_383, A[19]);
  nand g1031 (n_1117, n_382, n_383);
  nand g1032 (n_407, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_384, A[22]);
  xor g1034 (n_388, n_1118, n_385);
  nand g1035 (n_1119, n_384, A[22]);
  nand g1036 (n_1120, n_385, A[22]);
  nand g1037 (n_1121, n_384, n_385);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, n_386, A[23]);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, n_386, A[23]);
  nand g1042 (n_1124, n_387, A[23]);
  nand g1043 (n_1125, n_386, n_387);
  nand g1044 (n_410, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1051 (n_1130, A[1], A[3]);
  xor g1052 (n_393, n_1130, A[4]);
  nand g1053 (n_1131, A[1], A[3]);
  nand g1054 (n_1132, A[4], A[3]);
  nand g1055 (n_1133, A[1], A[4]);
  nand g1056 (n_412, n_1131, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, n_396, A[11]);
  xor g1070 (n_399, n_1142, A[12]);
  nand g1071 (n_1143, n_396, A[11]);
  nand g1072 (n_1144, A[12], A[11]);
  nand g1073 (n_1145, n_396, A[12]);
  nand g1074 (n_418, n_1143, n_1144, n_1145);
  xor g1075 (n_1146, n_397, n_398);
  xor g1076 (n_401, n_1146, n_399);
  nand g1077 (n_1147, n_397, n_398);
  nand g1078 (n_1148, n_399, n_398);
  nand g1079 (n_1149, n_397, n_399);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, A[15], n_400);
  xor g1082 (n_403, n_1150, A[16]);
  nand g1083 (n_1151, A[15], n_400);
  nand g1084 (n_1152, A[16], n_400);
  nand g1086 (n_421, n_1151, n_1152, n_984);
  xor g1087 (n_1154, n_401, n_402);
  xor g1088 (n_405, n_1154, A[19]);
  nand g1089 (n_1155, n_401, n_402);
  nand g1090 (n_1156, A[19], n_402);
  nand g1091 (n_1157, n_401, A[19]);
  nand g1092 (n_424, n_1155, n_1156, n_1157);
  xor g1093 (n_1158, n_403, A[20]);
  xor g1094 (n_406, n_1158, n_404);
  nand g1095 (n_1159, n_403, A[20]);
  nand g1096 (n_1160, n_404, A[20]);
  nand g1097 (n_1161, n_403, n_404);
  nand g1098 (n_425, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_405, n_406);
  xor g1100 (n_409, n_1162, n_407);
  nand g1101 (n_1163, n_405, n_406);
  nand g1102 (n_1164, n_407, n_406);
  nand g1103 (n_1165, n_405, n_407);
  nand g1104 (n_427, n_1163, n_1164, n_1165);
  xor g1106 (n_411, n_1166, n_408);
  nand g1108 (n_1168, n_408, A[23]);
  nand g1110 (n_430, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1123 (n_1178, A[8], n_413);
  xor g1124 (n_415, n_1178, A[9]);
  nand g1125 (n_1179, A[8], n_413);
  nand g1126 (n_1180, A[9], n_413);
  nand g1128 (n_435, n_1179, n_1180, n_687);
  xor g1129 (n_1182, n_414, n_415);
  xor g1130 (n_417, n_1182, A[12]);
  nand g1131 (n_1183, n_414, n_415);
  nand g1132 (n_1184, A[12], n_415);
  nand g1133 (n_1185, n_414, A[12]);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, n_416, A[13]);
  xor g1136 (n_420, n_1186, n_417);
  nand g1137 (n_1187, n_416, A[13]);
  nand g1138 (n_1188, n_417, A[13]);
  nand g1139 (n_1189, n_416, n_417);
  nand g1140 (n_439, n_1187, n_1188, n_1189);
  xor g1141 (n_1190, n_418, n_419);
  xor g1142 (n_422, n_1190, A[16]);
  nand g1143 (n_1191, n_418, n_419);
  nand g1144 (n_1192, A[16], n_419);
  nand g1145 (n_1193, n_418, A[16]);
  nand g1146 (n_440, n_1191, n_1192, n_1193);
  xor g1147 (n_1194, n_420, A[17]);
  xor g1148 (n_423, n_1194, n_421);
  nand g1149 (n_1195, n_420, A[17]);
  nand g1150 (n_1196, n_421, A[17]);
  nand g1151 (n_1197, n_420, n_421);
  nand g1152 (n_442, n_1195, n_1196, n_1197);
  xor g1153 (n_1198, n_422, A[20]);
  xor g1154 (n_426, n_1198, n_423);
  nand g1155 (n_1199, n_422, A[20]);
  nand g1156 (n_1200, n_423, A[20]);
  nand g1157 (n_1201, n_422, n_423);
  nand g1158 (n_445, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_424, A[21]);
  xor g1160 (n_428, n_1202, n_425);
  nand g1161 (n_1203, n_424, A[21]);
  nand g1162 (n_1204, n_425, A[21]);
  nand g1163 (n_1205, n_424, n_425);
  nand g1164 (n_447, n_1203, n_1204, n_1205);
  xor g1166 (n_429, n_1206, n_427);
  nand g1169 (n_1209, n_426, n_427);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, n_433);
  nand g1183 (n_1217, A[6], n_433);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, A[9], A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, A[9], A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, A[9], n_434);
  nand g1190 (n_455, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, n_435, n_436);
  xor g1192 (n_438, n_1222, A[13]);
  nand g1193 (n_1223, n_435, n_436);
  nand g1194 (n_1224, A[13], n_436);
  nand g1195 (n_1225, n_435, A[13]);
  nand g1196 (n_457, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, A[14], n_437);
  xor g1198 (n_441, n_1226, n_438);
  nand g1199 (n_1227, A[14], n_437);
  nand g1200 (n_1228, n_438, n_437);
  nand g1201 (n_1229, A[14], n_438);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, n_439, A[17]);
  xor g1204 (n_443, n_1230, n_440);
  nand g1205 (n_1231, n_439, A[17]);
  nand g1206 (n_1232, n_440, A[17]);
  nand g1207 (n_1233, n_439, n_440);
  nand g1208 (n_461, n_1231, n_1232, n_1233);
  xor g1209 (n_1234, A[18], n_441);
  xor g1210 (n_444, n_1234, n_442);
  nand g1211 (n_1235, A[18], n_441);
  nand g1212 (n_1236, n_442, n_441);
  nand g1213 (n_1237, A[18], n_442);
  nand g1214 (n_464, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_443, A[21]);
  xor g1216 (n_446, n_1238, A[22]);
  nand g1217 (n_1239, n_443, A[21]);
  nand g1219 (n_1241, n_443, A[22]);
  nand g1220 (n_465, n_1239, n_1077, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[5], A[7]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], n_453);
  xor g1242 (n_456, n_1254, n_454);
  nand g1243 (n_1255, A[10], n_453);
  nand g1244 (n_1256, n_454, n_453);
  nand g1245 (n_1257, A[10], n_454);
  nand g1246 (n_472, n_1255, n_1256, n_1257);
  xor g1247 (n_1258, A[11], n_455);
  xor g1248 (n_458, n_1258, n_456);
  nand g1249 (n_1259, A[11], n_455);
  nand g1250 (n_1260, n_456, n_455);
  nand g1251 (n_1261, A[11], n_456);
  nand g1252 (n_474, n_1259, n_1260, n_1261);
  xor g1253 (n_1262, A[14], n_457);
  xor g1254 (n_460, n_1262, A[15]);
  nand g1255 (n_1263, A[14], n_457);
  nand g1256 (n_1264, A[15], n_457);
  nand g1258 (n_476, n_1263, n_1264, n_1109);
  xor g1259 (n_1266, n_458, A[18]);
  xor g1260 (n_462, n_1266, n_459);
  nand g1261 (n_1267, n_458, A[18]);
  nand g1262 (n_1268, n_459, A[18]);
  nand g1263 (n_1269, n_458, n_459);
  nand g1264 (n_478, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, n_460, A[19]);
  xor g1266 (n_463, n_1270, n_461);
  nand g1267 (n_1271, n_460, A[19]);
  nand g1268 (n_1272, n_461, A[19]);
  nand g1269 (n_1273, n_460, n_461);
  nand g1270 (n_480, n_1271, n_1272, n_1273);
  xor g1271 (n_1274, n_462, A[22]);
  xor g1272 (n_466, n_1274, n_463);
  nand g1273 (n_1275, n_462, A[22]);
  nand g1274 (n_1276, n_463, A[22]);
  nand g1275 (n_1277, n_462, n_463);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1277 (n_1278, n_464, A[23]);
  xor g1278 (n_467, n_1278, n_465);
  nand g1279 (n_1279, n_464, A[23]);
  nand g1280 (n_1280, n_465, A[23]);
  nand g1281 (n_1281, n_464, n_465);
  nand g1282 (n_484, n_1279, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1289 (n_1286, A[7], A[6]);
  xor g1290 (n_471, n_1286, A[8]);
  nand g1292 (n_1288, A[8], A[6]);
  nand g1294 (n_486, n_661, n_1288, n_673);
  xor g1295 (n_1290, n_470, n_471);
  xor g1296 (n_473, n_1290, A[11]);
  nand g1297 (n_1291, n_470, n_471);
  nand g1298 (n_1292, A[11], n_471);
  nand g1299 (n_1293, n_470, A[11]);
  nand g1300 (n_488, n_1291, n_1292, n_1293);
  xor g1301 (n_1294, A[12], n_472);
  xor g1302 (n_475, n_1294, n_473);
  nand g1303 (n_1295, A[12], n_472);
  nand g1304 (n_1296, n_473, n_472);
  nand g1305 (n_1297, A[12], n_473);
  nand g1306 (n_489, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, A[15], n_474);
  xor g1308 (n_477, n_1298, n_475);
  nand g1309 (n_1299, A[15], n_474);
  nand g1310 (n_1300, n_475, n_474);
  nand g1311 (n_1301, A[15], n_475);
  nand g1312 (n_491, n_1299, n_1300, n_1301);
  xor g1313 (n_1302, A[16], n_476);
  xor g1314 (n_479, n_1302, n_477);
  nand g1315 (n_1303, A[16], n_476);
  nand g1316 (n_1304, n_477, n_476);
  nand g1317 (n_1305, A[16], n_477);
  nand g1318 (n_494, n_1303, n_1304, n_1305);
  xor g1319 (n_1306, A[19], A[20]);
  xor g1320 (n_481, n_1306, n_478);
  nand g1322 (n_1308, n_478, A[20]);
  nand g1323 (n_1309, A[19], n_478);
  nand g1324 (n_496, n_992, n_1308, n_1309);
  xor g1325 (n_1310, n_479, n_480);
  xor g1326 (n_483, n_1310, n_481);
  nand g1327 (n_1311, n_479, n_480);
  nand g1328 (n_1312, n_481, n_480);
  nand g1329 (n_1313, n_479, n_481);
  nand g1330 (n_497, n_1311, n_1312, n_1313);
  xor g1332 (n_485, n_1166, n_482);
  nand g1335 (n_1317, A[23], n_482);
  nand g1336 (n_500, n_1167, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1344 (n_487, n_686, n_486);
  nand g1346 (n_1324, n_486, A[9]);
  nand g1347 (n_1325, A[8], n_486);
  nand g1348 (n_503, n_687, n_1324, n_1325);
  xor g1349 (n_1326, A[12], n_487);
  xor g1350 (n_490, n_1326, n_488);
  nand g1351 (n_1327, A[12], n_487);
  nand g1352 (n_1328, n_488, n_487);
  nand g1353 (n_1329, A[12], n_488);
  nand g1354 (n_505, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, A[13], n_489);
  xor g1356 (n_492, n_1330, n_490);
  nand g1357 (n_1331, A[13], n_489);
  nand g1358 (n_1332, n_490, n_489);
  nand g1359 (n_1333, A[13], n_490);
  nand g1360 (n_507, n_1331, n_1332, n_1333);
  xor g1361 (n_1334, A[16], A[17]);
  xor g1362 (n_493, n_1334, n_491);
  nand g1363 (n_1335, A[16], A[17]);
  nand g1364 (n_1336, n_491, A[17]);
  nand g1365 (n_1337, A[16], n_491);
  nand g1366 (n_509, n_1335, n_1336, n_1337);
  xor g1367 (n_1338, n_492, A[20]);
  xor g1368 (n_495, n_1338, n_493);
  nand g1369 (n_1339, n_492, A[20]);
  nand g1370 (n_1340, n_493, A[20]);
  nand g1371 (n_1341, n_492, n_493);
  nand g1372 (n_511, n_1339, n_1340, n_1341);
  xor g1373 (n_1342, n_494, A[21]);
  xor g1374 (n_498, n_1342, n_495);
  nand g1375 (n_1343, n_494, A[21]);
  nand g1376 (n_1344, n_495, A[21]);
  nand g1377 (n_1345, n_494, n_495);
  nand g1378 (n_513, n_1343, n_1344, n_1345);
  xor g1380 (n_499, n_1346, n_497);
  nand g1383 (n_1349, n_496, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  nand g1397 (n_1357, A[10], n_503);
  nand g1398 (n_520, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], A[14]);
  xor g1400 (n_506, n_1358, n_504);
  nand g1401 (n_1359, A[13], A[14]);
  nand g1402 (n_1360, n_504, A[14]);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_521, n_1359, n_1360, n_1361);
  xor g1405 (n_1362, n_505, A[17]);
  xor g1406 (n_508, n_1362, n_506);
  nand g1407 (n_1363, n_505, A[17]);
  nand g1408 (n_1364, n_506, A[17]);
  nand g1409 (n_1365, n_505, n_506);
  nand g1410 (n_523, n_1363, n_1364, n_1365);
  xor g1411 (n_1366, n_507, A[18]);
  xor g1412 (n_510, n_1366, n_508);
  nand g1413 (n_1367, n_507, A[18]);
  nand g1414 (n_1368, n_508, A[18]);
  nand g1415 (n_1369, n_507, n_508);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_509, A[21]);
  xor g1418 (n_512, n_1370, n_510);
  nand g1419 (n_1371, n_509, A[21]);
  nand g1420 (n_1372, n_510, A[21]);
  nand g1421 (n_1373, n_509, n_510);
  nand g1422 (n_527, n_1371, n_1372, n_1373);
  xor g1423 (n_1374, A[22], n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, A[22], n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, A[22], n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1437 (n_1382, A[9], A[11]);
  nand g1439 (n_1383, A[9], A[11]);
  nand g1442 (n_532, n_1383, n_1384, n_1385);
  xor g1443 (n_1386, A[14], n_519);
  xor g1444 (n_522, n_1386, n_520);
  nand g1445 (n_1387, A[14], n_519);
  nand g1446 (n_1388, n_520, n_519);
  nand g1447 (n_1389, A[14], n_520);
  nand g1448 (n_534, n_1387, n_1388, n_1389);
  xor g1449 (n_1390, A[15], n_521);
  xor g1450 (n_524, n_1390, n_522);
  nand g1451 (n_1391, A[15], n_521);
  nand g1452 (n_1392, n_522, n_521);
  nand g1453 (n_1393, A[15], n_522);
  nand g1454 (n_536, n_1391, n_1392, n_1393);
  xor g1455 (n_1394, A[18], n_523);
  xor g1456 (n_525, n_1394, A[19]);
  nand g1457 (n_1395, A[18], n_523);
  nand g1458 (n_1396, A[19], n_523);
  nand g1459 (n_1397, A[18], A[19]);
  nand g1460 (n_538, n_1395, n_1396, n_1397);
  xor g1461 (n_1398, n_524, n_525);
  xor g1462 (n_528, n_1398, n_526);
  nand g1463 (n_1399, n_524, n_525);
  nand g1464 (n_1400, n_526, n_525);
  nand g1465 (n_1401, n_524, n_526);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1467 (n_1402, A[22], A[23]);
  xor g1468 (n_529, n_1402, n_527);
  nand g1469 (n_1403, A[22], A[23]);
  nand g1470 (n_1404, n_527, A[23]);
  nand g1471 (n_1405, A[22], n_527);
  nand g1472 (n_543, n_1403, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1479 (n_1410, A[11], A[12]);
  xor g1480 (n_533, n_1410, A[10]);
  nand g1482 (n_1412, A[10], A[12]);
  nand g1484 (n_544, n_1144, n_1412, n_1099);
  xor g1485 (n_1414, n_532, n_533);
  xor g1486 (n_535, n_1414, A[15]);
  nand g1487 (n_1415, n_532, n_533);
  nand g1488 (n_1416, A[15], n_533);
  nand g1489 (n_1417, n_532, A[15]);
  nand g1490 (n_546, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, A[16], n_534);
  xor g1492 (n_537, n_1418, n_535);
  nand g1493 (n_1419, A[16], n_534);
  nand g1494 (n_1420, n_535, n_534);
  nand g1495 (n_1421, A[16], n_535);
  nand g1496 (n_548, n_1419, n_1420, n_1421);
  xor g1497 (n_1422, A[19], n_536);
  xor g1498 (n_539, n_1422, A[20]);
  nand g1499 (n_1423, A[19], n_536);
  nand g1500 (n_1424, A[20], n_536);
  nand g1502 (n_549, n_1423, n_1424, n_992);
  xor g1503 (n_1426, n_537, n_538);
  xor g1504 (n_541, n_1426, n_539);
  nand g1505 (n_1427, n_537, n_538);
  nand g1506 (n_1428, n_539, n_538);
  nand g1507 (n_1429, n_537, n_539);
  nand g1508 (n_551, n_1427, n_1428, n_1429);
  xor g1510 (n_542, n_1166, n_540);
  nand g1513 (n_1433, A[23], n_540);
  nand g1514 (n_554, n_1167, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1521 (n_1438, A[12], A[13]);
  xor g1522 (n_545, n_1438, n_544);
  nand g1523 (n_1439, A[12], A[13]);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_1439, n_1440, n_1441);
  xor g1527 (n_1442, A[16], n_545);
  xor g1528 (n_547, n_1442, A[17]);
  nand g1529 (n_1443, A[16], n_545);
  nand g1530 (n_1444, A[17], n_545);
  nand g1532 (n_559, n_1443, n_1444, n_1335);
  xor g1533 (n_1446, n_546, n_547);
  xor g1534 (n_550, n_1446, A[20]);
  nand g1535 (n_1447, n_546, n_547);
  nand g1536 (n_1448, A[20], n_547);
  nand g1537 (n_1449, n_546, A[20]);
  nand g1538 (n_561, n_1447, n_1448, n_1449);
  xor g1539 (n_1450, n_548, A[21]);
  xor g1540 (n_552, n_1450, n_549);
  nand g1541 (n_1451, n_548, A[21]);
  nand g1542 (n_1452, n_549, A[21]);
  nand g1543 (n_1453, n_548, n_549);
  nand g1544 (n_562, n_1451, n_1452, n_1453);
  xor g1546 (n_553, n_1454, n_551);
  nand g1549 (n_1457, n_550, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1563 (n_1465, A[14], n_557);
  nand g1564 (n_569, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, A[17], A[18]);
  xor g1566 (n_560, n_1466, n_558);
  nand g1568 (n_1468, n_558, A[18]);
  nand g1569 (n_1469, A[17], n_558);
  nand g1570 (n_571, n_1068, n_1468, n_1469);
  xor g1571 (n_1470, n_559, n_560);
  xor g1572 (n_563, n_1470, A[21]);
  nand g1573 (n_1471, n_559, n_560);
  nand g1574 (n_1472, A[21], n_560);
  nand g1575 (n_1473, n_559, A[21]);
  nand g1576 (n_574, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, A[22], n_561);
  xor g1578 (n_564, n_1474, n_562);
  nand g1579 (n_1475, A[22], n_561);
  nand g1580 (n_1476, n_562, n_561);
  nand g1581 (n_1477, A[22], n_562);
  nand g1582 (n_576, n_1475, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  xor g1591 (n_1482, A[13], A[15]);
  nand g1593 (n_1483, A[13], A[15]);
  nand g1596 (n_578, n_1483, n_1484, n_1485);
  xor g1597 (n_1486, A[18], n_569);
  xor g1598 (n_572, n_1486, n_570);
  nand g1599 (n_1487, A[18], n_569);
  nand g1600 (n_1488, n_570, n_569);
  nand g1601 (n_1489, A[18], n_570);
  nand g1602 (n_580, n_1487, n_1488, n_1489);
  xor g1603 (n_1490, A[19], n_571);
  xor g1604 (n_573, n_1490, n_572);
  nand g1605 (n_1491, A[19], n_571);
  nand g1606 (n_1492, n_572, n_571);
  nand g1607 (n_1493, A[19], n_572);
  nand g1608 (n_583, n_1491, n_1492, n_1493);
  xor g1609 (n_1494, A[22], n_573);
  xor g1610 (n_575, n_1494, A[23]);
  nand g1611 (n_1495, A[22], n_573);
  nand g1612 (n_1496, A[23], n_573);
  nand g1614 (n_584, n_1495, n_1496, n_1403);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1621 (n_1502, A[15], A[14]);
  xor g1622 (n_579, n_1502, A[16]);
  nand g1626 (n_586, n_1109, n_801, n_984);
  xor g1627 (n_1506, n_578, n_579);
  xor g1628 (n_581, n_1506, A[19]);
  nand g1629 (n_1507, n_578, n_579);
  nand g1630 (n_1508, A[19], n_579);
  nand g1631 (n_1509, n_578, A[19]);
  nand g1632 (n_588, n_1507, n_1508, n_1509);
  xor g1633 (n_1510, A[20], n_580);
  xor g1634 (n_582, n_1510, n_581);
  nand g1635 (n_1511, A[20], n_580);
  nand g1636 (n_1512, n_581, n_580);
  nand g1637 (n_1513, A[20], n_581);
  nand g1638 (n_589, n_1511, n_1512, n_1513);
  xor g1639 (n_1514, A[23], n_582);
  xor g1640 (n_585, n_1514, n_583);
  nand g1641 (n_1515, A[23], n_582);
  nand g1642 (n_1516, n_583, n_582);
  nand g1643 (n_1517, A[23], n_583);
  nand g1644 (n_591, n_1515, n_1516, n_1517);
  xor g1646 (n_83, n_1518, n_585);
  nand g1648 (n_1520, n_585, n_584);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1652 (n_587, n_1334, n_586);
  nand g1654 (n_1524, n_586, A[17]);
  nand g1655 (n_1525, A[16], n_586);
  nand g1656 (n_595, n_1335, n_1524, n_1525);
  xor g1657 (n_1526, A[20], n_587);
  xor g1658 (n_590, n_1526, n_588);
  nand g1659 (n_1527, A[20], n_587);
  nand g1660 (n_1528, n_588, n_587);
  nand g1661 (n_1529, A[20], n_588);
  nand g1662 (n_597, n_1527, n_1528, n_1529);
  xor g1664 (n_592, n_1530, n_589);
  nand g1667 (n_1533, A[21], n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_81, n_1535, n_1536, n_1537);
  nand g1681 (n_1541, A[18], n_595);
  nand g1682 (n_604, n_1539, n_1540, n_1541);
  xor g1683 (n_1542, A[21], A[22]);
  xor g1684 (n_598, n_1542, n_596);
  nand g1686 (n_1544, n_596, A[22]);
  nand g1687 (n_1545, A[21], n_596);
  nand g1688 (n_606, n_1077, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_33, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[17], A[19]);
  nand g1702 (n_608, n_889, n_1552, n_1553);
  xor g1703 (n_1554, A[22], n_603);
  xor g1704 (n_605, n_1554, n_604);
  nand g1705 (n_1555, A[22], n_603);
  nand g1706 (n_1556, n_604, n_603);
  nand g1707 (n_1557, A[22], n_604);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, A[23], n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, A[23], n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, A[23], n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1716 (n_609, n_1306, A[18]);
  nand g1720 (n_612, n_992, n_925, n_1397);
  xor g1721 (n_1566, n_608, n_609);
  xor g1722 (n_611, n_1566, A[23]);
  nand g1723 (n_1567, n_608, n_609);
  nand g1724 (n_1568, A[23], n_609);
  nand g1725 (n_1569, n_608, A[23]);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1728 (n_79, n_1570, n_611);
  nand g1730 (n_1572, n_611, n_610);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1733 (n_1574, A[20], A[21]);
  xor g1734 (n_613, n_1574, n_612);
  nand g1735 (n_1575, A[20], A[21]);
  nand g1736 (n_1576, n_612, A[21]);
  nand g1737 (n_1577, A[20], n_612);
  nand g1738 (n_617, n_1575, n_1576, n_1577);
  xor g1740 (n_78, n_1578, n_614);
  nand g1742 (n_1580, n_614, n_613);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_617);
  nand g1752 (n_28, n_1583, n_1584, n_1585);
  nand g1759 (n_1589, A[21], A[23]);
  nand g1760 (n_27, n_1587, n_1588, n_1589);
  xor g1762 (n_75, n_1166, A[22]);
  nand g1766 (n_74, n_1167, n_1403, n_1593);
  nand g16 (n_1606, A[0], A[2]);
  xor g20 (Z[2], A[0], A[2]);
  nand g22 (n_1611, n_68, A[3]);
  nand g25 (n_1615, n_1611, n_1612, n_1613);
  xor g26 (n_1614, n_68, A[3]);
  nand g28 (n_1616, A[4], n_117);
  nand g29 (n_1617, A[4], n_1615);
  nand g30 (n_1618, n_117, n_1615);
  nand g31 (n_1620, n_1616, n_1617, n_1618);
  xor g32 (n_1619, A[4], n_117);
  xor g33 (Z[4], n_1615, n_1619);
  nand g34 (n_1621, A[5], n_116);
  nand g35 (n_1622, A[5], n_1620);
  nand g36 (n_1623, n_116, n_1620);
  nand g37 (n_1625, n_1621, n_1622, n_1623);
  xor g38 (n_1624, A[5], n_116);
  xor g39 (Z[5], n_1620, n_1624);
  nand g40 (n_1626, n_67, n_115);
  nand g41 (n_1627, n_67, n_1625);
  nand g42 (n_1628, n_115, n_1625);
  nand g43 (n_1630, n_1626, n_1627, n_1628);
  xor g44 (n_1629, n_67, n_115);
  xor g45 (Z[6], n_1625, n_1629);
  nand g46 (n_1631, n_66, n_114);
  nand g47 (n_1632, n_66, n_1630);
  nand g48 (n_1633, n_114, n_1630);
  nand g49 (n_1635, n_1631, n_1632, n_1633);
  xor g50 (n_1634, n_66, n_114);
  xor g51 (Z[7], n_1630, n_1634);
  nand g52 (n_1636, n_65, n_113);
  nand g53 (n_1637, n_65, n_1635);
  nand g54 (n_1638, n_113, n_1635);
  nand g55 (n_1640, n_1636, n_1637, n_1638);
  xor g56 (n_1639, n_65, n_113);
  xor g57 (Z[8], n_1635, n_1639);
  nand g58 (n_1641, n_64, n_112);
  nand g59 (n_1642, n_64, n_1640);
  nand g60 (n_1643, n_112, n_1640);
  nand g61 (n_1645, n_1641, n_1642, n_1643);
  xor g62 (n_1644, n_64, n_112);
  xor g63 (Z[9], n_1640, n_1644);
  nand g64 (n_1646, n_63, n_111);
  nand g65 (n_1647, n_63, n_1645);
  nand g66 (n_1648, n_111, n_1645);
  nand g67 (n_1650, n_1646, n_1647, n_1648);
  xor g68 (n_1649, n_63, n_111);
  xor g69 (Z[10], n_1645, n_1649);
  nand g70 (n_1651, n_62, n_110);
  nand g71 (n_1652, n_62, n_1650);
  nand g72 (n_1653, n_110, n_1650);
  nand g73 (n_1655, n_1651, n_1652, n_1653);
  xor g74 (n_1654, n_62, n_110);
  xor g75 (Z[11], n_1650, n_1654);
  nand g76 (n_1656, n_61, n_109);
  nand g77 (n_1657, n_61, n_1655);
  nand g78 (n_1658, n_109, n_1655);
  nand g79 (n_1660, n_1656, n_1657, n_1658);
  xor g80 (n_1659, n_61, n_109);
  xor g81 (Z[12], n_1655, n_1659);
  nand g82 (n_1661, n_60, n_108);
  nand g83 (n_1662, n_60, n_1660);
  nand g84 (n_1663, n_108, n_1660);
  nand g85 (n_1665, n_1661, n_1662, n_1663);
  xor g86 (n_1664, n_60, n_108);
  xor g87 (Z[13], n_1660, n_1664);
  nand g88 (n_1666, n_59, n_107);
  nand g89 (n_1667, n_59, n_1665);
  nand g90 (n_1668, n_107, n_1665);
  nand g91 (n_1670, n_1666, n_1667, n_1668);
  xor g92 (n_1669, n_59, n_107);
  xor g93 (Z[14], n_1665, n_1669);
  nand g94 (n_1671, n_58, n_106);
  nand g95 (n_1672, n_58, n_1670);
  nand g96 (n_1673, n_106, n_1670);
  nand g97 (n_1675, n_1671, n_1672, n_1673);
  xor g98 (n_1674, n_58, n_106);
  xor g99 (Z[15], n_1670, n_1674);
  nand g100 (n_1676, n_57, n_105);
  nand g101 (n_1677, n_57, n_1675);
  nand g102 (n_1678, n_105, n_1675);
  nand g103 (n_1680, n_1676, n_1677, n_1678);
  xor g104 (n_1679, n_57, n_105);
  xor g105 (Z[16], n_1675, n_1679);
  nand g106 (n_1681, n_56, n_104);
  nand g107 (n_1682, n_56, n_1680);
  nand g108 (n_1683, n_104, n_1680);
  nand g109 (n_1685, n_1681, n_1682, n_1683);
  xor g110 (n_1684, n_56, n_104);
  xor g111 (Z[17], n_1680, n_1684);
  nand g112 (n_1686, n_55, n_103);
  nand g113 (n_1687, n_55, n_1685);
  nand g114 (n_1688, n_103, n_1685);
  nand g115 (n_1690, n_1686, n_1687, n_1688);
  xor g116 (n_1689, n_55, n_103);
  xor g117 (Z[18], n_1685, n_1689);
  nand g118 (n_1691, n_54, n_102);
  nand g119 (n_1692, n_54, n_1690);
  nand g120 (n_1693, n_102, n_1690);
  nand g121 (n_1695, n_1691, n_1692, n_1693);
  xor g122 (n_1694, n_54, n_102);
  xor g123 (Z[19], n_1690, n_1694);
  nand g124 (n_1696, n_53, n_101);
  nand g125 (n_1697, n_53, n_1695);
  nand g126 (n_1698, n_101, n_1695);
  nand g127 (n_1700, n_1696, n_1697, n_1698);
  xor g128 (n_1699, n_53, n_101);
  xor g129 (Z[20], n_1695, n_1699);
  nand g130 (n_1701, n_52, n_100);
  nand g131 (n_1702, n_52, n_1700);
  nand g132 (n_1703, n_100, n_1700);
  nand g133 (n_1705, n_1701, n_1702, n_1703);
  xor g134 (n_1704, n_52, n_100);
  xor g135 (Z[21], n_1700, n_1704);
  nand g136 (n_1706, n_51, n_99);
  nand g137 (n_1707, n_51, n_1705);
  nand g138 (n_1708, n_99, n_1705);
  nand g139 (n_1710, n_1706, n_1707, n_1708);
  xor g140 (n_1709, n_51, n_99);
  xor g141 (Z[22], n_1705, n_1709);
  nand g142 (n_1711, n_50, n_98);
  nand g143 (n_1712, n_50, n_1710);
  nand g144 (n_1713, n_98, n_1710);
  nand g145 (n_1715, n_1711, n_1712, n_1713);
  xor g146 (n_1714, n_50, n_98);
  xor g147 (Z[23], n_1710, n_1714);
  nand g148 (n_1716, n_49, n_97);
  nand g149 (n_1717, n_49, n_1715);
  nand g150 (n_1718, n_97, n_1715);
  nand g151 (n_1720, n_1716, n_1717, n_1718);
  xor g152 (n_1719, n_49, n_97);
  xor g153 (Z[24], n_1715, n_1719);
  nand g154 (n_1721, n_48, n_96);
  nand g155 (n_1722, n_48, n_1720);
  nand g156 (n_1723, n_96, n_1720);
  nand g157 (n_1725, n_1721, n_1722, n_1723);
  xor g158 (n_1724, n_48, n_96);
  xor g159 (Z[25], n_1720, n_1724);
  nand g160 (n_1726, n_47, n_95);
  nand g161 (n_1727, n_47, n_1725);
  nand g162 (n_1728, n_95, n_1725);
  nand g163 (n_1730, n_1726, n_1727, n_1728);
  xor g164 (n_1729, n_47, n_95);
  xor g165 (Z[26], n_1725, n_1729);
  nand g166 (n_1731, n_46, n_94);
  nand g167 (n_1732, n_46, n_1730);
  nand g168 (n_1733, n_94, n_1730);
  nand g169 (n_1735, n_1731, n_1732, n_1733);
  xor g170 (n_1734, n_46, n_94);
  xor g171 (Z[27], n_1730, n_1734);
  nand g172 (n_1736, n_45, n_93);
  nand g173 (n_1737, n_45, n_1735);
  nand g174 (n_1738, n_93, n_1735);
  nand g175 (n_1740, n_1736, n_1737, n_1738);
  xor g176 (n_1739, n_45, n_93);
  xor g177 (Z[28], n_1735, n_1739);
  nand g178 (n_1741, n_44, n_92);
  nand g179 (n_1742, n_44, n_1740);
  nand g180 (n_1743, n_92, n_1740);
  nand g181 (n_1745, n_1741, n_1742, n_1743);
  xor g182 (n_1744, n_44, n_92);
  xor g183 (Z[29], n_1740, n_1744);
  nand g184 (n_1746, n_43, n_91);
  nand g185 (n_1747, n_43, n_1745);
  nand g186 (n_1748, n_91, n_1745);
  nand g187 (n_1750, n_1746, n_1747, n_1748);
  xor g188 (n_1749, n_43, n_91);
  xor g189 (Z[30], n_1745, n_1749);
  nand g190 (n_1751, n_42, n_90);
  nand g191 (n_1752, n_42, n_1750);
  nand g192 (n_1753, n_90, n_1750);
  nand g193 (n_1755, n_1751, n_1752, n_1753);
  xor g194 (n_1754, n_42, n_90);
  xor g195 (Z[31], n_1750, n_1754);
  nand g196 (n_1756, n_41, n_89);
  nand g197 (n_1757, n_41, n_1755);
  nand g198 (n_1758, n_89, n_1755);
  nand g199 (n_1760, n_1756, n_1757, n_1758);
  xor g200 (n_1759, n_41, n_89);
  xor g201 (Z[32], n_1755, n_1759);
  nand g202 (n_1761, n_40, n_88);
  nand g203 (n_1762, n_40, n_1760);
  nand g204 (n_1763, n_88, n_1760);
  nand g205 (n_1765, n_1761, n_1762, n_1763);
  xor g206 (n_1764, n_40, n_88);
  xor g207 (Z[33], n_1760, n_1764);
  nand g208 (n_1766, n_39, n_87);
  nand g209 (n_1767, n_39, n_1765);
  nand g210 (n_1768, n_87, n_1765);
  nand g211 (n_1770, n_1766, n_1767, n_1768);
  xor g212 (n_1769, n_39, n_87);
  xor g213 (Z[34], n_1765, n_1769);
  nand g214 (n_1771, n_38, n_86);
  nand g215 (n_1772, n_38, n_1770);
  nand g216 (n_1773, n_86, n_1770);
  nand g217 (n_1775, n_1771, n_1772, n_1773);
  xor g218 (n_1774, n_38, n_86);
  xor g219 (Z[35], n_1770, n_1774);
  nand g220 (n_1776, n_37, n_85);
  nand g221 (n_1777, n_37, n_1775);
  nand g222 (n_1778, n_85, n_1775);
  nand g223 (n_1780, n_1776, n_1777, n_1778);
  xor g224 (n_1779, n_37, n_85);
  xor g225 (Z[36], n_1775, n_1779);
  nand g226 (n_1781, n_36, n_84);
  nand g227 (n_1782, n_36, n_1780);
  nand g228 (n_1783, n_84, n_1780);
  nand g229 (n_1785, n_1781, n_1782, n_1783);
  xor g230 (n_1784, n_36, n_84);
  xor g231 (Z[37], n_1780, n_1784);
  nand g232 (n_1786, n_35, n_83);
  nand g233 (n_1787, n_35, n_1785);
  nand g234 (n_1788, n_83, n_1785);
  nand g235 (n_1790, n_1786, n_1787, n_1788);
  xor g236 (n_1789, n_35, n_83);
  xor g237 (Z[38], n_1785, n_1789);
  nand g238 (n_1791, n_34, n_82);
  nand g239 (n_1792, n_34, n_1790);
  nand g240 (n_1793, n_82, n_1790);
  nand g241 (n_1795, n_1791, n_1792, n_1793);
  xor g242 (n_1794, n_34, n_82);
  xor g243 (Z[39], n_1790, n_1794);
  nand g244 (n_1796, n_33, n_81);
  nand g245 (n_1797, n_33, n_1795);
  nand g246 (n_1798, n_81, n_1795);
  nand g247 (n_1800, n_1796, n_1797, n_1798);
  xor g248 (n_1799, n_33, n_81);
  xor g249 (Z[40], n_1795, n_1799);
  nand g250 (n_1801, n_32, n_80);
  nand g251 (n_1802, n_32, n_1800);
  nand g252 (n_1803, n_80, n_1800);
  nand g253 (n_1805, n_1801, n_1802, n_1803);
  xor g254 (n_1804, n_32, n_80);
  xor g255 (Z[41], n_1800, n_1804);
  nand g256 (n_1806, n_31, n_79);
  nand g257 (n_1807, n_31, n_1805);
  nand g258 (n_1808, n_79, n_1805);
  nand g259 (n_1810, n_1806, n_1807, n_1808);
  xor g260 (n_1809, n_31, n_79);
  xor g261 (Z[42], n_1805, n_1809);
  nand g262 (n_1811, n_30, n_78);
  nand g263 (n_1812, n_30, n_1810);
  nand g264 (n_1813, n_78, n_1810);
  nand g265 (n_1815, n_1811, n_1812, n_1813);
  xor g266 (n_1814, n_30, n_78);
  xor g267 (Z[43], n_1810, n_1814);
  nand g1772 (n_1816, n_29, n_77);
  nand g1773 (n_1817, n_29, n_1815);
  nand g1774 (n_1818, n_77, n_1815);
  nand g1775 (n_1820, n_1816, n_1817, n_1818);
  xor g1776 (n_1819, n_29, n_77);
  xor g1777 (Z[44], n_1815, n_1819);
  nand g1778 (n_1821, n_28, n_76);
  nand g1779 (n_1822, n_28, n_1820);
  nand g1780 (n_1823, n_76, n_1820);
  nand g1781 (n_1825, n_1821, n_1822, n_1823);
  xor g1782 (n_1824, n_28, n_76);
  xor g1783 (Z[45], n_1820, n_1824);
  nand g1784 (n_1826, n_27, n_75);
  nand g1785 (n_1827, n_27, n_1825);
  nand g1786 (n_1828, n_75, n_1825);
  nand g1787 (n_1830, n_1826, n_1827, n_1828);
  xor g1788 (n_1829, n_27, n_75);
  xor g1789 (Z[46], n_1825, n_1829);
  xor g1791 (Z[47], n_1830, n_1831);
  or g1804 (n_1043, A[1], wc);
  not gc (wc, n_171);
  or g1805 (n_1044, A[1], wc0);
  not gc0 (wc0, A[2]);
  xnor g1807 (n_1166, A[24], A[23]);
  or g1808 (n_1167, wc1, A[24]);
  not gc1 (wc1, A[23]);
  xnor g1809 (n_1214, A[6], A[5]);
  or g1810 (n_1215, A[5], wc2);
  not gc2 (wc2, A[6]);
  or g1811 (n_1252, A[6], wc3);
  not gc3 (wc3, A[7]);
  or g1812 (n_1253, wc4, A[6]);
  not gc4 (wc4, A[5]);
  or g1814 (n_1355, A[9], wc5);
  not gc5 (wc5, A[10]);
  or g1815 (n_1384, A[10], wc6);
  not gc6 (wc6, A[11]);
  or g1816 (n_1385, wc7, A[10]);
  not gc7 (wc7, A[9]);
  or g1818 (n_1463, A[13], wc8);
  not gc8 (wc8, A[14]);
  or g1819 (n_1484, A[14], wc9);
  not gc9 (wc9, A[15]);
  or g1820 (n_1485, wc10, A[14]);
  not gc10 (wc10, A[13]);
  xnor g1821 (n_1530, A[24], A[21]);
  or g1822 (n_1531, wc11, A[24]);
  not gc11 (wc11, A[21]);
  or g1824 (n_1539, A[17], wc12);
  not gc12 (wc12, A[18]);
  or g1825 (n_1552, A[18], wc13);
  not gc13 (wc13, A[19]);
  or g1826 (n_1553, wc14, A[18]);
  not gc14 (wc14, A[17]);
  or g1828 (n_1583, A[21], wc15);
  not gc15 (wc15, A[22]);
  or g1829 (n_1587, wc16, A[22]);
  not gc16 (wc16, A[21]);
  or g1830 (n_1588, A[22], wc17);
  not gc17 (wc17, A[23]);
  or g1831 (n_1593, wc18, A[24]);
  not gc18 (wc18, A[22]);
  xnor g1833 (n_1086, A[2], A[1]);
  or g1834 (n_1088, A[1], wc19);
  not gc19 (wc19, A[3]);
  xnor g1835 (n_453, n_1250, A[6]);
  xnor g1836 (n_519, n_1382, A[10]);
  xnor g1837 (n_570, n_1482, A[14]);
  xnor g1838 (n_603, n_1550, A[18]);
  xnor g1839 (n_76, n_1542, A[23]);
  or g1841 (n_1047, wc20, n_117);
  not gc20 (wc20, A[5]);
  or g1842 (n_1049, wc21, n_117);
  not gc21 (wc21, A[6]);
  xnor g1844 (n_1578, n_613, A[24]);
  or g1845 (n_1579, A[24], wc22);
  not gc22 (wc22, n_613);
  xnor g1846 (n_1831, n_74, A[24]);
  or g1848 (n_1051, n_180, wc23);
  not gc23 (wc23, n_179);
  or g1849 (n_1052, wc24, n_180);
  not gc24 (wc24, A[9]);
  xnor g1850 (n_504, n_1218, n_503);
  or g1851 (n_1356, A[9], wc25);
  not gc25 (wc25, n_503);
  xnor g1852 (n_558, n_1358, n_557);
  or g1853 (n_1464, A[13], wc26);
  not gc26 (wc26, n_557);
  xnor g1854 (n_596, n_1466, n_595);
  or g1855 (n_1540, A[17], wc27);
  not gc27 (wc27, n_595);
  or g1856 (n_1573, A[24], wc28);
  not gc28 (wc28, n_611);
  or g1857 (n_1581, A[24], wc29);
  not gc29 (wc29, n_614);
  xnor g1858 (n_29, n_1542, n_617);
  or g1859 (n_1584, A[21], wc30);
  not gc30 (wc30, n_617);
  or g1862 (n_1216, A[5], wc31);
  not gc31 (wc31, n_433);
  or g1863 (n_1612, n_1606, wc32);
  not gc32 (wc32, n_68);
  or g1864 (n_1613, wc33, n_1606);
  not gc33 (wc33, A[3]);
  xnor g1865 (Z[3], n_1606, n_1614);
  or g1867 (n_1056, wc34, n_202);
  not gc34 (wc34, A[10]);
  or g1868 (n_1057, wc35, n_202);
  not gc35 (wc35, n_282);
  or g1869 (n_1060, wc36, n_285);
  not gc36 (wc36, A[13]);
  xnor g1870 (n_1454, n_550, A[24]);
  or g1871 (n_1455, A[24], wc37);
  not gc37 (wc37, n_550);
  xnor g1872 (n_1570, n_610, A[24]);
  or g1873 (n_1571, A[24], wc38);
  not gc38 (wc38, n_610);
  or g1874 (n_1061, wc39, n_285);
  not gc39 (wc39, n_354);
  xnor g1875 (n_357, n_285, n_1058);
  or g1876 (n_1532, A[24], wc40);
  not gc40 (wc40, n_589);
  xnor g1877 (n_1518, n_584, A[24]);
  or g1878 (n_1519, A[24], wc41);
  not gc41 (wc41, n_584);
  or g1879 (n_1521, A[24], wc42);
  not gc42 (wc42, n_585);
  or g1880 (n_1456, A[24], wc43);
  not gc43 (wc43, n_551);
  xnor g1881 (n_1078, n_363, A[24]);
  or g1882 (n_1079, A[24], wc44);
  not gc44 (wc44, n_363);
  or g1883 (n_1080, A[24], wc45);
  not gc45 (wc45, n_364);
  xnor g1884 (n_1206, n_426, A[24]);
  or g1885 (n_1207, A[24], wc46);
  not gc46 (wc46, n_426);
  xnor g1886 (n_1346, n_496, A[24]);
  or g1887 (n_1347, A[24], wc47);
  not gc47 (wc47, n_496);
  or g1888 (n_1169, A[24], wc48);
  not gc48 (wc48, n_408);
  or g1889 (n_1432, A[24], wc49);
  not gc49 (wc49, n_540);
  or g1890 (n_1208, A[24], wc50);
  not gc50 (wc50, n_427);
  or g1891 (n_1316, A[24], wc51);
  not gc51 (wc51, n_482);
  or g1892 (n_1348, A[24], wc52);
  not gc52 (wc52, n_497);
endmodule

module mult_signed_const_5754_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_5754_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

module mult_signed_const_6021_GENERIC_REAL(A, Z);
// synthesis_equation "assign Z = $signed(A) * 13421773;"
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  wire n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34;
  wire n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42;
  wire n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50;
  wire n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58;
  wire n_59, n_60, n_61, n_62, n_63, n_64, n_65, n_66;
  wire n_67, n_68, n_69, n_71, n_72, n_73, n_74, n_75;
  wire n_76, n_77, n_78, n_79, n_80, n_81, n_82, n_83;
  wire n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91;
  wire n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115;
  wire n_116, n_117, n_118, n_119, n_171, n_172, n_173, n_176;
  wire n_179, n_180, n_183, n_184, n_187, n_188, n_189, n_195;
  wire n_196, n_201, n_202, n_203, n_204, n_209, n_210, n_211;
  wire n_212, n_217, n_218, n_219, n_220, n_221, n_223, n_224;
  wire n_225, n_226, n_227, n_232, n_234, n_235, n_236, n_237;
  wire n_238, n_239, n_246, n_248, n_249, n_250, n_251, n_259;
  wire n_260, n_262, n_265, n_267, n_269, n_271, n_273, n_274;
  wire n_275, n_276, n_277, n_281, n_282, n_283, n_284, n_285;
  wire n_286, n_287, n_288, n_289, n_290, n_291, n_292, n_293;
  wire n_296, n_298, n_299, n_300, n_301, n_302, n_303, n_304;
  wire n_305, n_306, n_307, n_308, n_309, n_315, n_316, n_318;
  wire n_319, n_320, n_321, n_322, n_323, n_324, n_325, n_326;
  wire n_333, n_335, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_354, n_355, n_356, n_357;
  wire n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365;
  wire n_366, n_367, n_371, n_372, n_373, n_374, n_375, n_376;
  wire n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384;
  wire n_385, n_386, n_387, n_388, n_389, n_390, n_392, n_393;
  wire n_394, n_395, n_396, n_397, n_398, n_399, n_400, n_401;
  wire n_402, n_403, n_404, n_405, n_406, n_407, n_408, n_409;
  wire n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417;
  wire n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425;
  wire n_426, n_427, n_428, n_429, n_430, n_433, n_434, n_435;
  wire n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443;
  wire n_444, n_445, n_446, n_447, n_448, n_449, n_453, n_454;
  wire n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462;
  wire n_463, n_464, n_465, n_466, n_467, n_468, n_470, n_471;
  wire n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479;
  wire n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487;
  wire n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495;
  wire n_496, n_497, n_498, n_499, n_500, n_503, n_504, n_505;
  wire n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
  wire n_514, n_515, n_519, n_520, n_521, n_522, n_523, n_524;
  wire n_525, n_526, n_527, n_528, n_529, n_530, n_532, n_533;
  wire n_534, n_535, n_536, n_537, n_538, n_539, n_540, n_541;
  wire n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549;
  wire n_550, n_551, n_552, n_553, n_554, n_557, n_558, n_559;
  wire n_560, n_561, n_562, n_563, n_564, n_565, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_578, n_579;
  wire n_580, n_581, n_582, n_583, n_584, n_585, n_586, n_587;
  wire n_588, n_589, n_590, n_591, n_592, n_595, n_596, n_597;
  wire n_598, n_599, n_603, n_604, n_605, n_606, n_608, n_609;
  wire n_610, n_611, n_612, n_613, n_614, n_617, n_622, n_623;
  wire n_624, n_625, n_626, n_627, n_628, n_629, n_630, n_631;
  wire n_632, n_633, n_634, n_635, n_636, n_637, n_638, n_639;
  wire n_640, n_641, n_646, n_647, n_648, n_649, n_650, n_651;
  wire n_652, n_653, n_658, n_659, n_660, n_661, n_662, n_663;
  wire n_664, n_665, n_668, n_669, n_670, n_671, n_672, n_673;
  wire n_674, n_675, n_676, n_677, n_684, n_685, n_686, n_687;
  wire n_688, n_689, n_690, n_691, n_692, n_693, n_704, n_705;
  wire n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713;
  wire n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_738, n_742, n_743, n_744, n_745, n_746;
  wire n_747, n_748, n_749, n_750, n_751, n_752, n_753, n_760;
  wire n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768;
  wire n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776;
  wire n_777, n_790, n_791, n_792, n_794, n_795, n_796, n_797;
  wire n_798, n_799, n_800, n_801, n_802, n_803, n_804, n_805;
  wire n_822, n_823, n_824, n_825, n_826, n_827, n_828, n_829;
  wire n_830, n_831, n_832, n_833, n_842, n_850, n_851, n_852;
  wire n_853, n_854, n_855, n_856, n_857, n_858, n_859, n_860;
  wire n_861, n_862, n_866, n_867, n_868, n_872, n_873, n_876;
  wire n_877, n_880, n_881, n_882, n_883, n_884, n_885, n_886;
  wire n_887, n_888, n_889, n_890, n_891, n_892, n_893, n_900;
  wire n_901, n_902, n_903, n_904, n_905, n_906, n_907, n_908;
  wire n_909, n_910, n_911, n_912, n_913, n_914, n_915, n_916;
  wire n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924;
  wire n_925, n_926, n_927, n_928, n_929, n_938, n_939, n_941;
  wire n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949;
  wire n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957;
  wire n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965;
  wire n_978, n_979, n_980, n_981, n_984, n_985, n_986, n_987;
  wire n_988, n_989, n_990, n_991, n_992, n_993, n_994, n_995;
  wire n_996, n_997, n_998, n_999, n_1000, n_1001, n_1013, n_1014;
  wire n_1015, n_1016, n_1017, n_1020, n_1021, n_1022, n_1023, n_1024;
  wire n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032;
  wire n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040;
  wire n_1041, n_1043, n_1044, n_1047, n_1049, n_1051, n_1052, n_1056;
  wire n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064;
  wire n_1065, n_1066, n_1067, n_1069, n_1070, n_1071, n_1072, n_1073;
  wire n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081;
  wire n_1082, n_1083, n_1084, n_1085, n_1088, n_1090, n_1091, n_1092;
  wire n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100;
  wire n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108;
  wire n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116;
  wire n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124;
  wire n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132;
  wire n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140;
  wire n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148;
  wire n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156;
  wire n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164;
  wire n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172;
  wire n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180;
  wire n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189;
  wire n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197;
  wire n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205;
  wire n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213;
  wire n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221;
  wire n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229;
  wire n_1230, n_1231, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238;
  wire n_1239, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247;
  wire n_1248, n_1249, n_1250, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1257, n_1258, n_1259, n_1260, n_1261, n_1264, n_1265, n_1266;
  wire n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274;
  wire n_1275, n_1276, n_1277, n_1280, n_1281, n_1282, n_1283, n_1284;
  wire n_1285, n_1286, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295;
  wire n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303;
  wire n_1304, n_1305, n_1306, n_1307, n_1308, n_1310, n_1311, n_1312;
  wire n_1313, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1324;
  wire n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332;
  wire n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340;
  wire n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348;
  wire n_1349, n_1350, n_1351, n_1352, n_1353, n_1355, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373;
  wire n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381;
  wire n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
  wire n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397;
  wire n_1398, n_1399, n_1400, n_1401, n_1404, n_1405, n_1406, n_1407;
  wire n_1408, n_1409, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417;
  wire n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1426;
  wire n_1427, n_1428, n_1429, n_1432, n_1433, n_1434, n_1435, n_1436;
  wire n_1437, n_1440, n_1441, n_1442, n_1443, n_1444, n_1446, n_1447;
  wire n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455;
  wire n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1463, n_1464;
  wire n_1465, n_1466, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473;
  wire n_1474, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482;
  wire n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491;
  wire n_1492, n_1493, n_1494, n_1495, n_1496, n_1498, n_1499, n_1500;
  wire n_1501, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512;
  wire n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520;
  wire n_1521, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530;
  wire n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1539;
  wire n_1540, n_1541, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558;
  wire n_1559, n_1560, n_1561, n_1562, n_1564, n_1566, n_1567, n_1568;
  wire n_1569, n_1570, n_1571, n_1572, n_1573, n_1576, n_1577, n_1578;
  wire n_1579, n_1580, n_1581, n_1583, n_1584, n_1585, n_1587, n_1588;
  wire n_1589, n_1593, n_1606, n_1611, n_1612, n_1613, n_1614, n_1615;
  wire n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623;
  wire n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631;
  wire n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639;
  wire n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647;
  wire n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655;
  wire n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663;
  wire n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671;
  wire n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679;
  wire n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687;
  wire n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695;
  wire n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703;
  wire n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711;
  wire n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719;
  wire n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727;
  wire n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735;
  wire n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743;
  wire n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751;
  wire n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759;
  wire n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767;
  wire n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775;
  wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
  wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
  wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
  wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
  wire n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815;
  wire n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823;
  wire n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831;
  assign Z[0] = A[0];
  assign Z[1] = A[1];
  xor g268 (n_68, A[0], A[1]);
  and g2 (n_171, A[0], A[1]);
  xor g269 (n_622, A[1], n_171);
  xor g270 (n_117, n_622, A[2]);
  nand g3 (n_623, A[1], n_171);
  nand g271 (n_624, A[2], n_171);
  nand g272 (n_625, A[1], A[2]);
  nand g273 (n_172, n_623, n_624, n_625);
  xor g274 (n_626, A[2], A[3]);
  xor g275 (n_116, n_626, n_172);
  nand g276 (n_627, A[2], A[3]);
  nand g4 (n_628, n_172, A[3]);
  nand g277 (n_629, A[2], n_172);
  nand g278 (n_67, n_627, n_628, n_629);
  xor g279 (n_173, A[0], A[3]);
  and g280 (n_69, A[0], A[3]);
  xor g281 (n_630, A[4], n_173);
  xor g282 (n_115, n_630, A[6]);
  nand g283 (n_631, A[4], n_173);
  nand g284 (n_632, A[6], n_173);
  nand g5 (n_633, A[4], A[6]);
  nand g6 (n_66, n_631, n_632, n_633);
  xor g287 (n_634, n_68, n_69);
  xor g288 (n_176, n_634, A[4]);
  nand g289 (n_635, n_68, n_69);
  nand g290 (n_636, A[4], n_69);
  nand g291 (n_637, n_68, A[4]);
  nand g292 (n_179, n_635, n_636, n_637);
  xor g293 (n_638, A[5], n_176);
  xor g294 (n_114, n_638, A[7]);
  nand g295 (n_639, A[5], n_176);
  nand g296 (n_640, A[7], n_176);
  nand g297 (n_641, A[5], A[7]);
  nand g298 (n_65, n_639, n_640, n_641);
  xor g305 (n_646, n_117, A[5]);
  xor g306 (n_180, n_646, n_179);
  nand g307 (n_647, n_117, A[5]);
  nand g308 (n_648, n_179, A[5]);
  nand g309 (n_649, n_117, n_179);
  nand g310 (n_183, n_647, n_648, n_649);
  xor g311 (n_650, A[6], n_180);
  xor g312 (n_113, n_650, A[8]);
  nand g313 (n_651, A[6], n_180);
  nand g314 (n_652, A[8], n_180);
  nand g315 (n_653, A[6], A[8]);
  nand g316 (n_64, n_651, n_652, n_653);
  xor g323 (n_658, A[6], n_116);
  xor g324 (n_184, n_658, A[7]);
  nand g325 (n_659, A[6], n_116);
  nand g326 (n_660, A[7], n_116);
  nand g327 (n_661, A[6], A[7]);
  nand g328 (n_188, n_659, n_660, n_661);
  xor g329 (n_662, n_183, n_184);
  xor g330 (n_112, n_662, A[9]);
  nand g331 (n_663, n_183, n_184);
  nand g332 (n_664, A[9], n_184);
  nand g333 (n_665, n_183, A[9]);
  nand g334 (n_63, n_663, n_664, n_665);
  xor g338 (n_187, n_630, n_67);
  nand g340 (n_668, n_67, n_173);
  nand g341 (n_669, A[4], n_67);
  nand g342 (n_71, n_631, n_668, n_669);
  xor g343 (n_670, A[7], n_187);
  xor g344 (n_189, n_670, A[8]);
  nand g345 (n_671, A[7], n_187);
  nand g346 (n_672, A[8], n_187);
  nand g347 (n_673, A[7], A[8]);
  nand g348 (n_73, n_671, n_672, n_673);
  xor g349 (n_674, n_188, A[10]);
  xor g350 (n_111, n_674, n_189);
  nand g351 (n_675, n_188, A[10]);
  nand g352 (n_676, n_189, A[10]);
  nand g353 (n_677, n_188, n_189);
  nand g354 (n_62, n_675, n_676, n_677);
  xor g364 (n_195, n_638, n_71);
  nand g366 (n_684, n_71, n_176);
  nand g367 (n_685, A[5], n_71);
  nand g368 (n_201, n_639, n_684, n_685);
  xor g369 (n_686, A[8], A[9]);
  xor g370 (n_196, n_686, n_73);
  nand g371 (n_687, A[8], A[9]);
  nand g372 (n_688, n_73, A[9]);
  nand g373 (n_689, A[8], n_73);
  nand g374 (n_203, n_687, n_688, n_689);
  xor g375 (n_690, n_195, A[11]);
  xor g376 (n_110, n_690, n_196);
  nand g377 (n_691, n_195, A[11]);
  nand g378 (n_692, n_196, A[11]);
  nand g379 (n_693, n_195, n_196);
  nand g380 (n_61, n_691, n_692, n_693);
  xor g394 (n_202, n_650, A[9]);
  nand g396 (n_704, A[9], n_180);
  nand g397 (n_705, A[6], A[9]);
  nand g398 (n_209, n_651, n_704, n_705);
  xor g399 (n_706, A[10], n_201);
  xor g400 (n_204, n_706, n_202);
  nand g401 (n_707, A[10], n_201);
  nand g402 (n_708, n_202, n_201);
  nand g403 (n_709, A[10], n_202);
  nand g404 (n_211, n_707, n_708, n_709);
  xor g405 (n_710, A[12], n_203);
  xor g406 (n_109, n_710, n_204);
  nand g407 (n_711, A[12], n_203);
  nand g408 (n_712, n_204, n_203);
  nand g409 (n_713, A[12], n_204);
  nand g410 (n_60, n_711, n_712, n_713);
  xor g424 (n_210, n_662, A[10]);
  nand g426 (n_724, A[10], n_184);
  nand g427 (n_725, n_183, A[10]);
  nand g428 (n_218, n_663, n_724, n_725);
  xor g429 (n_726, A[11], n_209);
  xor g430 (n_212, n_726, n_210);
  nand g431 (n_727, A[11], n_209);
  nand g432 (n_728, n_210, n_209);
  nand g433 (n_729, A[11], n_210);
  nand g434 (n_219, n_727, n_728, n_729);
  xor g435 (n_730, n_211, A[13]);
  xor g436 (n_108, n_730, n_212);
  nand g437 (n_731, n_211, A[13]);
  nand g438 (n_732, n_212, A[13]);
  nand g439 (n_733, n_211, n_212);
  nand g440 (n_59, n_731, n_732, n_733);
  xor g449 (n_738, A[7], A[8]);
  xor g450 (n_217, n_738, n_187);
  xor g455 (n_742, n_188, n_217);
  xor g456 (n_220, n_742, A[11]);
  nand g457 (n_743, n_188, n_217);
  nand g458 (n_744, A[11], n_217);
  nand g459 (n_745, n_188, A[11]);
  nand g460 (n_224, n_743, n_744, n_745);
  xor g461 (n_746, n_218, A[12]);
  xor g462 (n_221, n_746, n_219);
  nand g463 (n_747, n_218, A[12]);
  nand g464 (n_748, n_219, A[12]);
  nand g465 (n_749, n_218, n_219);
  nand g466 (n_226, n_747, n_748, n_749);
  xor g467 (n_750, A[14], n_220);
  xor g468 (n_107, n_750, n_221);
  nand g469 (n_751, A[14], n_220);
  nand g470 (n_752, n_221, n_220);
  nand g471 (n_753, A[14], n_221);
  nand g472 (n_58, n_751, n_752, n_753);
  xor g482 (n_72, n_638, A[8]);
  nand g484 (n_760, A[8], n_176);
  nand g485 (n_761, A[5], A[8]);
  nand g486 (n_232, n_639, n_760, n_761);
  xor g487 (n_762, n_71, A[9]);
  xor g488 (n_223, n_762, n_72);
  nand g489 (n_763, n_71, A[9]);
  nand g490 (n_764, n_72, A[9]);
  nand g491 (n_765, n_71, n_72);
  nand g492 (n_234, n_763, n_764, n_765);
  xor g493 (n_766, n_73, A[12]);
  xor g494 (n_225, n_766, n_223);
  nand g495 (n_767, n_73, A[12]);
  nand g496 (n_768, n_223, A[12]);
  nand g497 (n_769, n_73, n_223);
  nand g498 (n_236, n_767, n_768, n_769);
  xor g499 (n_770, n_224, A[13]);
  xor g500 (n_227, n_770, A[15]);
  nand g501 (n_771, n_224, A[13]);
  nand g502 (n_772, A[15], A[13]);
  nand g503 (n_773, n_224, A[15]);
  nand g504 (n_238, n_771, n_772, n_773);
  xor g505 (n_774, n_225, n_226);
  xor g506 (n_106, n_774, n_227);
  nand g507 (n_775, n_225, n_226);
  nand g508 (n_776, n_227, n_226);
  nand g509 (n_777, n_225, n_227);
  nand g510 (n_57, n_775, n_776, n_777);
  xor g529 (n_790, A[10], n_232);
  xor g530 (n_235, n_790, n_202);
  nand g531 (n_791, A[10], n_232);
  nand g532 (n_792, n_202, n_232);
  nand g534 (n_246, n_791, n_792, n_709);
  xor g535 (n_794, n_234, n_235);
  xor g536 (n_237, n_794, A[13]);
  nand g537 (n_795, n_234, n_235);
  nand g538 (n_796, A[13], n_235);
  nand g539 (n_797, n_234, A[13]);
  nand g540 (n_248, n_795, n_796, n_797);
  xor g541 (n_798, A[14], n_236);
  xor g542 (n_239, n_798, A[16]);
  nand g543 (n_799, A[14], n_236);
  nand g544 (n_800, A[16], n_236);
  nand g545 (n_801, A[14], A[16]);
  nand g546 (n_250, n_799, n_800, n_801);
  xor g547 (n_802, n_237, n_238);
  xor g548 (n_105, n_802, n_239);
  nand g549 (n_803, n_237, n_238);
  nand g550 (n_804, n_239, n_238);
  nand g551 (n_805, n_237, n_239);
  nand g552 (n_56, n_803, n_804, n_805);
  xor g577 (n_822, n_246, A[14]);
  xor g578 (n_249, n_822, n_212);
  nand g579 (n_823, n_246, A[14]);
  nand g580 (n_824, n_212, A[14]);
  nand g581 (n_825, n_246, n_212);
  nand g582 (n_260, n_823, n_824, n_825);
  xor g583 (n_826, A[15], n_248);
  xor g584 (n_251, n_826, A[17]);
  nand g585 (n_827, A[15], n_248);
  nand g586 (n_828, A[17], n_248);
  nand g587 (n_829, A[15], A[17]);
  nand g588 (n_118, n_827, n_828, n_829);
  xor g589 (n_830, n_249, n_250);
  xor g590 (n_104, n_830, n_251);
  nand g591 (n_831, n_249, n_250);
  nand g592 (n_832, n_251, n_250);
  nand g593 (n_833, n_249, n_251);
  nand g594 (n_55, n_831, n_832, n_833);
  xor g609 (n_842, n_188, A[11]);
  xor g610 (n_259, n_842, n_217);
  xor g621 (n_850, n_259, A[15]);
  xor g622 (n_262, n_850, n_260);
  nand g623 (n_851, n_259, A[15]);
  nand g624 (n_852, n_260, A[15]);
  nand g625 (n_853, n_259, n_260);
  nand g626 (n_274, n_851, n_852, n_853);
  xor g627 (n_854, n_221, A[16]);
  xor g628 (n_119, n_854, A[18]);
  nand g629 (n_855, n_221, A[16]);
  nand g630 (n_856, A[18], A[16]);
  nand g631 (n_857, n_221, A[18]);
  nand g632 (n_276, n_855, n_856, n_857);
  xor g633 (n_858, n_262, n_118);
  xor g634 (n_103, n_858, n_119);
  nand g635 (n_859, n_262, n_118);
  nand g636 (n_860, n_119, n_118);
  nand g637 (n_861, n_262, n_119);
  nand g638 (n_54, n_859, n_860, n_861);
  xor g641 (n_862, n_68, A[4]);
  xor g642 (n_265, n_862, n_69);
  xor g647 (n_866, A[5], n_265);
  xor g648 (n_267, n_866, A[8]);
  nand g649 (n_867, A[5], n_265);
  nand g650 (n_868, A[8], n_265);
  nand g652 (n_282, n_867, n_868, n_761);
  xor g654 (n_269, n_762, n_267);
  nand g656 (n_872, n_267, A[9]);
  nand g657 (n_873, n_71, n_267);
  nand g658 (n_284, n_763, n_872, n_873);
  xor g660 (n_271, n_766, n_269);
  nand g662 (n_876, n_269, A[12]);
  nand g663 (n_877, n_73, n_269);
  nand g664 (n_286, n_767, n_876, n_877);
  xor g666 (n_273, n_770, n_271);
  nand g668 (n_880, n_271, A[13]);
  nand g669 (n_881, n_224, n_271);
  nand g670 (n_288, n_771, n_880, n_881);
  xor g671 (n_882, n_226, A[16]);
  xor g672 (n_275, n_882, n_273);
  nand g673 (n_883, n_226, A[16]);
  nand g674 (n_884, n_273, A[16]);
  nand g675 (n_885, n_226, n_273);
  nand g676 (n_290, n_883, n_884, n_885);
  xor g677 (n_886, A[17], n_274);
  xor g678 (n_277, n_886, A[19]);
  nand g679 (n_887, A[17], n_274);
  nand g680 (n_888, A[19], n_274);
  nand g681 (n_889, A[17], A[19]);
  nand g682 (n_292, n_887, n_888, n_889);
  xor g683 (n_890, n_275, n_276);
  xor g684 (n_102, n_890, n_277);
  nand g685 (n_891, n_275, n_276);
  nand g686 (n_892, n_277, n_276);
  nand g687 (n_893, n_275, n_277);
  nand g688 (n_53, n_891, n_892, n_893);
  xor g696 (n_281, n_646, A[6]);
  nand g698 (n_900, A[6], A[5]);
  nand g699 (n_901, n_117, A[6]);
  nand g700 (n_296, n_647, n_900, n_901);
  xor g701 (n_902, n_179, n_281);
  xor g702 (n_283, n_902, A[9]);
  nand g703 (n_903, n_179, n_281);
  nand g704 (n_904, A[9], n_281);
  nand g705 (n_905, n_179, A[9]);
  nand g706 (n_298, n_903, n_904, n_905);
  xor g707 (n_906, A[10], n_282);
  xor g708 (n_285, n_906, n_283);
  nand g709 (n_907, A[10], n_282);
  nand g710 (n_908, n_283, n_282);
  nand g711 (n_909, A[10], n_283);
  nand g712 (n_300, n_907, n_908, n_909);
  xor g713 (n_910, n_284, A[13]);
  xor g714 (n_287, n_910, n_285);
  nand g715 (n_911, n_284, A[13]);
  nand g716 (n_912, n_285, A[13]);
  nand g717 (n_913, n_284, n_285);
  nand g718 (n_302, n_911, n_912, n_913);
  xor g719 (n_914, A[14], n_286);
  xor g720 (n_289, n_914, n_287);
  nand g721 (n_915, A[14], n_286);
  nand g722 (n_916, n_287, n_286);
  nand g723 (n_917, A[14], n_287);
  nand g724 (n_304, n_915, n_916, n_917);
  xor g725 (n_918, n_288, A[17]);
  xor g726 (n_291, n_918, A[18]);
  nand g727 (n_919, n_288, A[17]);
  nand g728 (n_920, A[18], A[17]);
  nand g729 (n_921, n_288, A[18]);
  nand g730 (n_306, n_919, n_920, n_921);
  xor g731 (n_922, n_289, n_290);
  xor g732 (n_293, n_922, A[20]);
  nand g733 (n_923, n_289, n_290);
  nand g734 (n_924, A[20], n_290);
  nand g735 (n_925, n_289, A[20]);
  nand g736 (n_308, n_923, n_924, n_925);
  xor g737 (n_926, n_291, n_292);
  xor g738 (n_101, n_926, n_293);
  nand g739 (n_927, n_291, n_292);
  nand g740 (n_928, n_293, n_292);
  nand g741 (n_929, n_291, n_293);
  nand g742 (n_52, n_927, n_928, n_929);
  xor g755 (n_938, n_296, n_184);
  xor g756 (n_299, n_938, A[10]);
  nand g757 (n_939, n_296, n_184);
  nand g759 (n_941, n_296, A[10]);
  nand g760 (n_315, n_939, n_724, n_941);
  xor g761 (n_942, A[11], n_298);
  xor g762 (n_301, n_942, n_299);
  nand g763 (n_943, A[11], n_298);
  nand g764 (n_944, n_299, n_298);
  nand g765 (n_945, A[11], n_299);
  nand g766 (n_316, n_943, n_944, n_945);
  xor g767 (n_946, n_300, A[14]);
  xor g768 (n_303, n_946, n_301);
  nand g769 (n_947, n_300, A[14]);
  nand g770 (n_948, n_301, A[14]);
  nand g771 (n_949, n_300, n_301);
  nand g772 (n_318, n_947, n_948, n_949);
  xor g773 (n_950, A[15], n_302);
  xor g774 (n_305, n_950, n_303);
  nand g775 (n_951, A[15], n_302);
  nand g776 (n_952, n_303, n_302);
  nand g777 (n_953, A[15], n_303);
  nand g778 (n_321, n_951, n_952, n_953);
  xor g779 (n_954, A[18], n_304);
  xor g780 (n_307, n_954, n_305);
  nand g781 (n_955, A[18], n_304);
  nand g782 (n_956, n_305, n_304);
  nand g783 (n_957, A[18], n_305);
  nand g784 (n_323, n_955, n_956, n_957);
  xor g785 (n_958, A[19], n_306);
  xor g786 (n_309, n_958, A[21]);
  nand g787 (n_959, A[19], n_306);
  nand g788 (n_960, A[21], n_306);
  nand g789 (n_961, A[19], A[21]);
  nand g790 (n_325, n_959, n_960, n_961);
  xor g791 (n_962, n_307, n_308);
  xor g792 (n_100, n_962, n_309);
  nand g793 (n_963, n_307, n_308);
  nand g794 (n_964, n_309, n_308);
  nand g795 (n_965, n_307, n_309);
  nand g796 (n_51, n_963, n_964, n_965);
  xor g817 (n_978, A[12], n_315);
  xor g818 (n_319, n_978, n_316);
  nand g819 (n_979, A[12], n_315);
  nand g820 (n_980, n_316, n_315);
  nand g821 (n_981, A[12], n_316);
  nand g822 (n_336, n_979, n_980, n_981);
  xor g824 (n_320, n_850, n_318);
  nand g826 (n_984, n_318, A[15]);
  nand g827 (n_985, n_259, n_318);
  nand g828 (n_338, n_851, n_984, n_985);
  xor g829 (n_986, A[16], n_319);
  xor g830 (n_322, n_986, n_320);
  nand g831 (n_987, A[16], n_319);
  nand g832 (n_988, n_320, n_319);
  nand g833 (n_989, A[16], n_320);
  nand g834 (n_340, n_987, n_988, n_989);
  xor g835 (n_990, A[19], n_321);
  xor g836 (n_324, n_990, A[20]);
  nand g837 (n_991, A[19], n_321);
  nand g838 (n_992, A[20], n_321);
  nand g839 (n_993, A[19], A[20]);
  nand g840 (n_342, n_991, n_992, n_993);
  xor g841 (n_994, n_322, n_323);
  xor g842 (n_326, n_994, n_324);
  nand g843 (n_995, n_322, n_323);
  nand g844 (n_996, n_324, n_323);
  nand g845 (n_997, n_322, n_324);
  nand g846 (n_344, n_995, n_996, n_997);
  xor g847 (n_998, A[22], n_325);
  xor g848 (n_99, n_998, n_326);
  nand g849 (n_999, A[22], n_325);
  nand g850 (n_1000, n_326, n_325);
  nand g851 (n_1001, A[22], n_326);
  nand g852 (n_50, n_999, n_1000, n_1001);
  xor g868 (n_333, n_762, n_73);
  nand g871 (n_1013, n_71, n_73);
  nand g872 (n_354, n_763, n_688, n_1013);
  xor g873 (n_1014, n_267, A[12]);
  xor g874 (n_335, n_1014, n_333);
  nand g875 (n_1015, n_267, A[12]);
  nand g876 (n_1016, n_333, A[12]);
  nand g877 (n_1017, n_267, n_333);
  nand g878 (n_356, n_1015, n_1016, n_1017);
  xor g880 (n_337, n_770, n_335);
  nand g882 (n_1020, n_335, A[13]);
  nand g883 (n_1021, n_224, n_335);
  nand g884 (n_358, n_771, n_1020, n_1021);
  xor g885 (n_1022, n_336, A[16]);
  xor g886 (n_339, n_1022, n_337);
  nand g887 (n_1023, n_336, A[16]);
  nand g888 (n_1024, n_337, A[16]);
  nand g889 (n_1025, n_336, n_337);
  nand g890 (n_360, n_1023, n_1024, n_1025);
  xor g891 (n_1026, A[17], n_338);
  xor g892 (n_341, n_1026, n_339);
  nand g893 (n_1027, A[17], n_338);
  nand g894 (n_1028, n_339, n_338);
  nand g895 (n_1029, A[17], n_339);
  nand g896 (n_362, n_1027, n_1028, n_1029);
  xor g897 (n_1030, A[20], n_340);
  xor g898 (n_343, n_1030, n_341);
  nand g899 (n_1031, A[20], n_340);
  nand g900 (n_1032, n_341, n_340);
  nand g901 (n_1033, A[20], n_341);
  nand g902 (n_364, n_1031, n_1032, n_1033);
  xor g903 (n_1034, A[21], n_342);
  xor g904 (n_345, n_1034, n_343);
  nand g905 (n_1035, A[21], n_342);
  nand g906 (n_1036, n_343, n_342);
  nand g907 (n_1037, A[21], n_343);
  nand g908 (n_366, n_1035, n_1036, n_1037);
  xor g909 (n_1038, A[23], n_344);
  xor g910 (n_98, n_1038, n_345);
  nand g911 (n_1039, A[23], n_344);
  nand g912 (n_1040, n_345, n_344);
  nand g913 (n_1041, A[23], n_345);
  nand g914 (n_49, n_1039, n_1040, n_1041);
  nand g922 (n_371, n_1043, n_1044, n_624);
  nand g928 (n_373, n_1047, n_648, n_1049);
  nand g934 (n_375, n_1051, n_1052, n_705);
  nand g940 (n_377, n_907, n_1056, n_1057);
  xor g941 (n_1058, n_354, A[13]);
  xor g942 (n_357, n_1058, n_355);
  nand g943 (n_1059, n_354, A[13]);
  nand g944 (n_1060, n_355, A[13]);
  nand g945 (n_1061, n_354, n_355);
  nand g946 (n_379, n_1059, n_1060, n_1061);
  xor g947 (n_1062, A[14], n_356);
  xor g948 (n_359, n_1062, n_357);
  nand g949 (n_1063, A[14], n_356);
  nand g950 (n_1064, n_357, n_356);
  nand g951 (n_1065, A[14], n_357);
  nand g952 (n_382, n_1063, n_1064, n_1065);
  xor g953 (n_1066, n_358, A[17]);
  xor g954 (n_361, n_1066, A[18]);
  nand g955 (n_1067, n_358, A[17]);
  nand g957 (n_1069, n_358, A[18]);
  nand g958 (n_383, n_1067, n_920, n_1069);
  xor g959 (n_1070, n_359, n_360);
  xor g960 (n_363, n_1070, n_361);
  nand g961 (n_1071, n_359, n_360);
  nand g962 (n_1072, n_361, n_360);
  nand g963 (n_1073, n_359, n_361);
  nand g964 (n_386, n_1071, n_1072, n_1073);
  xor g965 (n_1074, A[21], n_362);
  xor g966 (n_365, n_1074, A[22]);
  nand g967 (n_1075, A[21], n_362);
  nand g968 (n_1076, A[22], n_362);
  nand g969 (n_1077, A[21], A[22]);
  nand g970 (n_387, n_1075, n_1076, n_1077);
  xor g971 (n_1078, n_363, n_364);
  nand g973 (n_1079, n_363, n_364);
  nand g976 (n_389, n_1079, n_1080, n_1081);
  xor g977 (n_1082, n_365, n_366);
  xor g978 (n_97, n_1082, n_367);
  nand g979 (n_1083, n_365, n_366);
  nand g980 (n_1084, n_367, n_366);
  nand g981 (n_1085, n_365, n_367);
  nand g982 (n_48, n_1083, n_1084, n_1085);
  nand g990 (n_392, n_627, n_1088, n_1044);
  xor g991 (n_1090, n_371, n_372);
  xor g992 (n_374, n_1090, A[6]);
  nand g993 (n_1091, n_371, n_372);
  nand g994 (n_1092, A[6], n_372);
  nand g995 (n_1093, n_371, A[6]);
  nand g996 (n_394, n_1091, n_1092, n_1093);
  xor g997 (n_1094, A[7], n_373);
  xor g998 (n_376, n_1094, n_374);
  nand g999 (n_1095, A[7], n_373);
  nand g1000 (n_1096, n_374, n_373);
  nand g1001 (n_1097, A[7], n_374);
  nand g1002 (n_396, n_1095, n_1096, n_1097);
  xor g1003 (n_1098, A[10], A[11]);
  xor g1004 (n_378, n_1098, n_375);
  nand g1005 (n_1099, A[10], A[11]);
  nand g1006 (n_1100, n_375, A[11]);
  nand g1007 (n_1101, A[10], n_375);
  nand g1008 (n_398, n_1099, n_1100, n_1101);
  xor g1009 (n_1102, n_376, n_377);
  xor g1010 (n_380, n_1102, n_378);
  nand g1011 (n_1103, n_376, n_377);
  nand g1012 (n_1104, n_378, n_377);
  nand g1013 (n_1105, n_376, n_378);
  nand g1014 (n_400, n_1103, n_1104, n_1105);
  xor g1015 (n_1106, A[14], A[15]);
  xor g1016 (n_381, n_1106, n_379);
  nand g1017 (n_1107, A[14], A[15]);
  nand g1018 (n_1108, n_379, A[15]);
  nand g1019 (n_1109, A[14], n_379);
  nand g1020 (n_402, n_1107, n_1108, n_1109);
  xor g1021 (n_1110, n_380, A[18]);
  xor g1022 (n_384, n_1110, n_381);
  nand g1023 (n_1111, n_380, A[18]);
  nand g1024 (n_1112, n_381, A[18]);
  nand g1025 (n_1113, n_380, n_381);
  nand g1026 (n_404, n_1111, n_1112, n_1113);
  xor g1027 (n_1114, n_382, A[19]);
  xor g1028 (n_385, n_1114, n_383);
  nand g1029 (n_1115, n_382, A[19]);
  nand g1030 (n_1116, n_383, A[19]);
  nand g1031 (n_1117, n_382, n_383);
  nand g1032 (n_406, n_1115, n_1116, n_1117);
  xor g1033 (n_1118, n_384, n_385);
  xor g1034 (n_388, n_1118, n_386);
  nand g1035 (n_1119, n_384, n_385);
  nand g1036 (n_1120, n_386, n_385);
  nand g1037 (n_1121, n_384, n_386);
  nand g1038 (n_408, n_1119, n_1120, n_1121);
  xor g1039 (n_1122, A[22], A[23]);
  xor g1040 (n_390, n_1122, n_387);
  nand g1041 (n_1123, A[22], A[23]);
  nand g1042 (n_1124, n_387, A[23]);
  nand g1043 (n_1125, A[22], n_387);
  nand g1044 (n_411, n_1123, n_1124, n_1125);
  xor g1045 (n_1126, n_388, n_389);
  xor g1046 (n_96, n_1126, n_390);
  nand g1047 (n_1127, n_388, n_389);
  nand g1048 (n_1128, n_390, n_389);
  nand g1049 (n_1129, n_388, n_390);
  nand g1050 (n_47, n_1127, n_1128, n_1129);
  xor g1051 (n_1130, A[3], A[1]);
  xor g1052 (n_393, n_1130, A[4]);
  nand g1053 (n_1131, A[3], A[1]);
  nand g1054 (n_1132, A[4], A[1]);
  nand g1055 (n_1133, A[3], A[4]);
  nand g1056 (n_412, n_1131, n_1132, n_1133);
  xor g1057 (n_1134, n_392, n_393);
  xor g1058 (n_395, n_1134, A[7]);
  nand g1059 (n_1135, n_392, n_393);
  nand g1060 (n_1136, A[7], n_393);
  nand g1061 (n_1137, n_392, A[7]);
  nand g1062 (n_414, n_1135, n_1136, n_1137);
  xor g1063 (n_1138, A[8], n_394);
  xor g1064 (n_397, n_1138, n_395);
  nand g1065 (n_1139, A[8], n_394);
  nand g1066 (n_1140, n_395, n_394);
  nand g1067 (n_1141, A[8], n_395);
  nand g1068 (n_416, n_1139, n_1140, n_1141);
  xor g1069 (n_1142, n_396, A[11]);
  xor g1070 (n_399, n_1142, n_397);
  nand g1071 (n_1143, n_396, A[11]);
  nand g1072 (n_1144, n_397, A[11]);
  nand g1073 (n_1145, n_396, n_397);
  nand g1074 (n_417, n_1143, n_1144, n_1145);
  xor g1075 (n_1146, A[12], n_398);
  xor g1076 (n_401, n_1146, n_399);
  nand g1077 (n_1147, A[12], n_398);
  nand g1078 (n_1148, n_399, n_398);
  nand g1079 (n_1149, A[12], n_399);
  nand g1080 (n_419, n_1147, n_1148, n_1149);
  xor g1081 (n_1150, A[15], n_400);
  xor g1082 (n_403, n_1150, A[16]);
  nand g1083 (n_1151, A[15], n_400);
  nand g1084 (n_1152, A[16], n_400);
  nand g1085 (n_1153, A[15], A[16]);
  nand g1086 (n_421, n_1151, n_1152, n_1153);
  xor g1087 (n_1154, n_401, n_402);
  xor g1088 (n_405, n_1154, A[19]);
  nand g1089 (n_1155, n_401, n_402);
  nand g1090 (n_1156, A[19], n_402);
  nand g1091 (n_1157, n_401, A[19]);
  nand g1092 (n_424, n_1155, n_1156, n_1157);
  xor g1093 (n_1158, n_403, n_404);
  xor g1094 (n_407, n_1158, A[20]);
  nand g1095 (n_1159, n_403, n_404);
  nand g1096 (n_1160, A[20], n_404);
  nand g1097 (n_1161, n_403, A[20]);
  nand g1098 (n_425, n_1159, n_1160, n_1161);
  xor g1099 (n_1162, n_405, n_406);
  xor g1100 (n_409, n_1162, n_407);
  nand g1101 (n_1163, n_405, n_406);
  nand g1102 (n_1164, n_407, n_406);
  nand g1103 (n_1165, n_405, n_407);
  nand g1104 (n_428, n_1163, n_1164, n_1165);
  xor g1106 (n_410, n_1166, n_408);
  nand g1108 (n_1168, n_408, A[23]);
  nand g1110 (n_430, n_1167, n_1168, n_1169);
  xor g1111 (n_1170, n_409, n_410);
  xor g1112 (n_95, n_1170, n_411);
  nand g1113 (n_1171, n_409, n_410);
  nand g1114 (n_1172, n_411, n_410);
  nand g1115 (n_1173, n_409, n_411);
  nand g1116 (n_46, n_1171, n_1172, n_1173);
  xor g1117 (n_1174, A[4], A[5]);
  xor g1118 (n_413, n_1174, n_412);
  nand g1119 (n_1175, A[4], A[5]);
  nand g1120 (n_1176, n_412, A[5]);
  nand g1121 (n_1177, A[4], n_412);
  nand g1122 (n_433, n_1175, n_1176, n_1177);
  xor g1123 (n_1178, A[8], n_413);
  xor g1124 (n_415, n_1178, A[9]);
  nand g1125 (n_1179, A[8], n_413);
  nand g1126 (n_1180, A[9], n_413);
  nand g1128 (n_435, n_1179, n_1180, n_687);
  xor g1129 (n_1182, n_414, n_415);
  xor g1130 (n_418, n_1182, n_416);
  nand g1131 (n_1183, n_414, n_415);
  nand g1132 (n_1184, n_416, n_415);
  nand g1133 (n_1185, n_414, n_416);
  nand g1134 (n_437, n_1183, n_1184, n_1185);
  xor g1135 (n_1186, A[12], A[13]);
  xor g1136 (n_420, n_1186, n_417);
  nand g1137 (n_1187, A[12], A[13]);
  nand g1138 (n_1188, n_417, A[13]);
  nand g1139 (n_1189, A[12], n_417);
  nand g1140 (n_439, n_1187, n_1188, n_1189);
  xor g1141 (n_1190, n_418, n_419);
  xor g1142 (n_422, n_1190, A[16]);
  nand g1143 (n_1191, n_418, n_419);
  nand g1144 (n_1192, A[16], n_419);
  nand g1145 (n_1193, n_418, A[16]);
  nand g1146 (n_441, n_1191, n_1192, n_1193);
  xor g1147 (n_1194, n_420, A[17]);
  xor g1148 (n_423, n_1194, n_421);
  nand g1149 (n_1195, n_420, A[17]);
  nand g1150 (n_1196, n_421, A[17]);
  nand g1151 (n_1197, n_420, n_421);
  nand g1152 (n_443, n_1195, n_1196, n_1197);
  xor g1153 (n_1198, n_422, A[20]);
  xor g1154 (n_426, n_1198, n_423);
  nand g1155 (n_1199, n_422, A[20]);
  nand g1156 (n_1200, n_423, A[20]);
  nand g1157 (n_1201, n_422, n_423);
  nand g1158 (n_445, n_1199, n_1200, n_1201);
  xor g1159 (n_1202, n_424, A[21]);
  xor g1160 (n_427, n_1202, n_425);
  nand g1161 (n_1203, n_424, A[21]);
  nand g1162 (n_1204, n_425, A[21]);
  nand g1163 (n_1205, n_424, n_425);
  nand g1164 (n_446, n_1203, n_1204, n_1205);
  xor g1166 (n_429, n_1206, n_427);
  nand g1169 (n_1209, n_426, n_427);
  nand g1170 (n_449, n_1207, n_1208, n_1209);
  xor g1171 (n_1210, n_428, n_429);
  xor g1172 (n_94, n_1210, n_430);
  nand g1173 (n_1211, n_428, n_429);
  nand g1174 (n_1212, n_430, n_429);
  nand g1175 (n_1213, n_428, n_430);
  nand g1176 (n_45, n_1211, n_1212, n_1213);
  xor g1180 (n_434, n_1214, n_433);
  nand g1183 (n_1217, A[6], n_433);
  nand g1184 (n_454, n_1215, n_1216, n_1217);
  xor g1185 (n_1218, A[9], A[10]);
  xor g1186 (n_436, n_1218, n_434);
  nand g1187 (n_1219, A[9], A[10]);
  nand g1188 (n_1220, n_434, A[10]);
  nand g1189 (n_1221, A[9], n_434);
  nand g1190 (n_456, n_1219, n_1220, n_1221);
  xor g1191 (n_1222, n_435, n_436);
  xor g1192 (n_438, n_1222, A[13]);
  nand g1193 (n_1223, n_435, n_436);
  nand g1194 (n_1224, A[13], n_436);
  nand g1195 (n_1225, n_435, A[13]);
  nand g1196 (n_457, n_1223, n_1224, n_1225);
  xor g1197 (n_1226, n_437, A[14]);
  xor g1198 (n_440, n_1226, n_438);
  nand g1199 (n_1227, n_437, A[14]);
  nand g1200 (n_1228, n_438, A[14]);
  nand g1201 (n_1229, n_437, n_438);
  nand g1202 (n_459, n_1227, n_1228, n_1229);
  xor g1203 (n_1230, n_439, A[17]);
  xor g1204 (n_442, n_1230, A[18]);
  nand g1205 (n_1231, n_439, A[17]);
  nand g1207 (n_1233, n_439, A[18]);
  nand g1208 (n_461, n_1231, n_920, n_1233);
  xor g1209 (n_1234, n_440, n_441);
  xor g1210 (n_444, n_1234, n_442);
  nand g1211 (n_1235, n_440, n_441);
  nand g1212 (n_1236, n_442, n_441);
  nand g1213 (n_1237, n_440, n_442);
  nand g1214 (n_463, n_1235, n_1236, n_1237);
  xor g1215 (n_1238, n_443, A[21]);
  xor g1216 (n_447, n_1238, A[22]);
  nand g1217 (n_1239, n_443, A[21]);
  nand g1219 (n_1241, n_443, A[22]);
  nand g1220 (n_465, n_1239, n_1077, n_1241);
  xor g1221 (n_1242, n_444, n_445);
  xor g1222 (n_448, n_1242, n_446);
  nand g1223 (n_1243, n_444, n_445);
  nand g1224 (n_1244, n_446, n_445);
  nand g1225 (n_1245, n_444, n_446);
  nand g1226 (n_468, n_1243, n_1244, n_1245);
  xor g1227 (n_1246, n_447, n_448);
  xor g1228 (n_93, n_1246, n_449);
  nand g1229 (n_1247, n_447, n_448);
  nand g1230 (n_1248, n_449, n_448);
  nand g1231 (n_1249, n_447, n_449);
  nand g1232 (n_44, n_1247, n_1248, n_1249);
  xor g1235 (n_1250, A[7], A[5]);
  nand g1240 (n_470, n_641, n_1252, n_1253);
  xor g1241 (n_1254, A[10], n_453);
  xor g1242 (n_455, n_1254, n_454);
  nand g1243 (n_1255, A[10], n_453);
  nand g1244 (n_1256, n_454, n_453);
  nand g1245 (n_1257, A[10], n_454);
  nand g1246 (n_472, n_1255, n_1256, n_1257);
  xor g1247 (n_1258, A[11], n_455);
  xor g1248 (n_458, n_1258, n_456);
  nand g1249 (n_1259, A[11], n_455);
  nand g1250 (n_1260, n_456, n_455);
  nand g1251 (n_1261, A[11], n_456);
  nand g1252 (n_474, n_1259, n_1260, n_1261);
  xor g1254 (n_460, n_1106, n_457);
  nand g1256 (n_1264, n_457, A[15]);
  nand g1257 (n_1265, A[14], n_457);
  nand g1258 (n_476, n_1107, n_1264, n_1265);
  xor g1259 (n_1266, n_458, A[18]);
  xor g1260 (n_462, n_1266, n_459);
  nand g1261 (n_1267, n_458, A[18]);
  nand g1262 (n_1268, n_459, A[18]);
  nand g1263 (n_1269, n_458, n_459);
  nand g1264 (n_478, n_1267, n_1268, n_1269);
  xor g1265 (n_1270, n_460, A[19]);
  xor g1266 (n_464, n_1270, n_461);
  nand g1267 (n_1271, n_460, A[19]);
  nand g1268 (n_1272, n_461, A[19]);
  nand g1269 (n_1273, n_460, n_461);
  nand g1270 (n_480, n_1271, n_1272, n_1273);
  xor g1271 (n_1274, n_462, n_463);
  xor g1272 (n_466, n_1274, n_464);
  nand g1273 (n_1275, n_462, n_463);
  nand g1274 (n_1276, n_464, n_463);
  nand g1275 (n_1277, n_462, n_464);
  nand g1276 (n_482, n_1275, n_1276, n_1277);
  xor g1278 (n_467, n_1122, n_465);
  nand g1280 (n_1280, n_465, A[23]);
  nand g1281 (n_1281, A[22], n_465);
  nand g1282 (n_485, n_1123, n_1280, n_1281);
  xor g1283 (n_1282, n_466, n_467);
  xor g1284 (n_92, n_1282, n_468);
  nand g1285 (n_1283, n_466, n_467);
  nand g1286 (n_1284, n_468, n_467);
  nand g1287 (n_1285, n_466, n_468);
  nand g1288 (n_43, n_1283, n_1284, n_1285);
  xor g1289 (n_1286, A[7], A[6]);
  xor g1290 (n_471, n_1286, A[8]);
  nand g1294 (n_486, n_661, n_653, n_673);
  xor g1295 (n_1290, n_470, n_471);
  xor g1296 (n_473, n_1290, A[11]);
  nand g1297 (n_1291, n_470, n_471);
  nand g1298 (n_1292, A[11], n_471);
  nand g1299 (n_1293, n_470, A[11]);
  nand g1300 (n_488, n_1291, n_1292, n_1293);
  xor g1301 (n_1294, A[12], n_472);
  xor g1302 (n_475, n_1294, n_473);
  nand g1303 (n_1295, A[12], n_472);
  nand g1304 (n_1296, n_473, n_472);
  nand g1305 (n_1297, A[12], n_473);
  nand g1306 (n_489, n_1295, n_1296, n_1297);
  xor g1307 (n_1298, A[15], n_474);
  xor g1308 (n_477, n_1298, n_475);
  nand g1309 (n_1299, A[15], n_474);
  nand g1310 (n_1300, n_475, n_474);
  nand g1311 (n_1301, A[15], n_475);
  nand g1312 (n_491, n_1299, n_1300, n_1301);
  xor g1313 (n_1302, A[16], n_476);
  xor g1314 (n_479, n_1302, n_477);
  nand g1315 (n_1303, A[16], n_476);
  nand g1316 (n_1304, n_477, n_476);
  nand g1317 (n_1305, A[16], n_477);
  nand g1318 (n_494, n_1303, n_1304, n_1305);
  xor g1319 (n_1306, A[19], n_478);
  xor g1320 (n_481, n_1306, A[20]);
  nand g1321 (n_1307, A[19], n_478);
  nand g1322 (n_1308, A[20], n_478);
  nand g1324 (n_495, n_1307, n_1308, n_993);
  xor g1325 (n_1310, n_479, n_480);
  xor g1326 (n_483, n_1310, n_481);
  nand g1327 (n_1311, n_479, n_480);
  nand g1328 (n_1312, n_481, n_480);
  nand g1329 (n_1313, n_479, n_481);
  nand g1330 (n_498, n_1311, n_1312, n_1313);
  xor g1332 (n_484, n_1166, n_482);
  nand g1335 (n_1317, A[23], n_482);
  nand g1336 (n_500, n_1167, n_1316, n_1317);
  xor g1337 (n_1318, n_483, n_484);
  xor g1338 (n_91, n_1318, n_485);
  nand g1339 (n_1319, n_483, n_484);
  nand g1340 (n_1320, n_485, n_484);
  nand g1341 (n_1321, n_483, n_485);
  nand g1342 (n_42, n_1319, n_1320, n_1321);
  xor g1344 (n_487, n_686, n_486);
  nand g1346 (n_1324, n_486, A[9]);
  nand g1347 (n_1325, A[8], n_486);
  nand g1348 (n_503, n_687, n_1324, n_1325);
  xor g1349 (n_1326, A[12], n_487);
  xor g1350 (n_490, n_1326, n_488);
  nand g1351 (n_1327, A[12], n_487);
  nand g1352 (n_1328, n_488, n_487);
  nand g1353 (n_1329, A[12], n_488);
  nand g1354 (n_505, n_1327, n_1328, n_1329);
  xor g1355 (n_1330, A[13], n_489);
  xor g1356 (n_492, n_1330, n_490);
  nand g1357 (n_1331, A[13], n_489);
  nand g1358 (n_1332, n_490, n_489);
  nand g1359 (n_1333, A[13], n_490);
  nand g1360 (n_507, n_1331, n_1332, n_1333);
  xor g1361 (n_1334, A[16], A[17]);
  xor g1362 (n_493, n_1334, n_491);
  nand g1363 (n_1335, A[16], A[17]);
  nand g1364 (n_1336, n_491, A[17]);
  nand g1365 (n_1337, A[16], n_491);
  nand g1366 (n_508, n_1335, n_1336, n_1337);
  xor g1367 (n_1338, n_492, A[20]);
  xor g1368 (n_496, n_1338, n_493);
  nand g1369 (n_1339, n_492, A[20]);
  nand g1370 (n_1340, n_493, A[20]);
  nand g1371 (n_1341, n_492, n_493);
  nand g1372 (n_511, n_1339, n_1340, n_1341);
  xor g1373 (n_1342, n_494, A[21]);
  xor g1374 (n_497, n_1342, n_495);
  nand g1375 (n_1343, n_494, A[21]);
  nand g1376 (n_1344, n_495, A[21]);
  nand g1377 (n_1345, n_494, n_495);
  nand g1378 (n_512, n_1343, n_1344, n_1345);
  xor g1380 (n_499, n_1346, n_497);
  nand g1383 (n_1349, n_496, n_497);
  nand g1384 (n_515, n_1347, n_1348, n_1349);
  xor g1385 (n_1350, n_498, n_499);
  xor g1386 (n_90, n_1350, n_500);
  nand g1387 (n_1351, n_498, n_499);
  nand g1388 (n_1352, n_500, n_499);
  nand g1389 (n_1353, n_498, n_500);
  nand g1390 (n_41, n_1351, n_1352, n_1353);
  nand g1397 (n_1357, A[10], n_503);
  nand g1398 (n_520, n_1355, n_1356, n_1357);
  xor g1399 (n_1358, A[13], A[14]);
  xor g1400 (n_506, n_1358, n_504);
  nand g1401 (n_1359, A[13], A[14]);
  nand g1402 (n_1360, n_504, A[14]);
  nand g1403 (n_1361, A[13], n_504);
  nand g1404 (n_521, n_1359, n_1360, n_1361);
  xor g1405 (n_1362, n_505, A[17]);
  xor g1406 (n_509, n_1362, n_506);
  nand g1407 (n_1363, n_505, A[17]);
  nand g1408 (n_1364, n_506, A[17]);
  nand g1409 (n_1365, n_505, n_506);
  nand g1410 (n_523, n_1363, n_1364, n_1365);
  xor g1411 (n_1366, A[18], n_507);
  xor g1412 (n_510, n_1366, n_508);
  nand g1413 (n_1367, A[18], n_507);
  nand g1414 (n_1368, n_508, n_507);
  nand g1415 (n_1369, A[18], n_508);
  nand g1416 (n_526, n_1367, n_1368, n_1369);
  xor g1417 (n_1370, n_509, A[21]);
  xor g1418 (n_513, n_1370, n_510);
  nand g1419 (n_1371, n_509, A[21]);
  nand g1420 (n_1372, n_510, A[21]);
  nand g1421 (n_1373, n_509, n_510);
  nand g1422 (n_527, n_1371, n_1372, n_1373);
  xor g1423 (n_1374, A[22], n_511);
  xor g1424 (n_514, n_1374, n_512);
  nand g1425 (n_1375, A[22], n_511);
  nand g1426 (n_1376, n_512, n_511);
  nand g1427 (n_1377, A[22], n_512);
  nand g1428 (n_530, n_1375, n_1376, n_1377);
  xor g1429 (n_1378, n_513, n_514);
  xor g1430 (n_89, n_1378, n_515);
  nand g1431 (n_1379, n_513, n_514);
  nand g1432 (n_1380, n_515, n_514);
  nand g1433 (n_1381, n_513, n_515);
  nand g1434 (n_40, n_1379, n_1380, n_1381);
  xor g1437 (n_1382, A[9], A[11]);
  nand g1439 (n_1383, A[9], A[11]);
  nand g1442 (n_532, n_1383, n_1384, n_1385);
  xor g1443 (n_1386, A[14], n_519);
  xor g1444 (n_522, n_1386, n_520);
  nand g1445 (n_1387, A[14], n_519);
  nand g1446 (n_1388, n_520, n_519);
  nand g1447 (n_1389, A[14], n_520);
  nand g1448 (n_534, n_1387, n_1388, n_1389);
  xor g1449 (n_1390, A[15], n_521);
  xor g1450 (n_524, n_1390, n_522);
  nand g1451 (n_1391, A[15], n_521);
  nand g1452 (n_1392, n_522, n_521);
  nand g1453 (n_1393, A[15], n_522);
  nand g1454 (n_536, n_1391, n_1392, n_1393);
  xor g1455 (n_1394, A[18], n_523);
  xor g1456 (n_525, n_1394, A[19]);
  nand g1457 (n_1395, A[18], n_523);
  nand g1458 (n_1396, A[19], n_523);
  nand g1459 (n_1397, A[18], A[19]);
  nand g1460 (n_538, n_1395, n_1396, n_1397);
  xor g1461 (n_1398, n_524, n_525);
  xor g1462 (n_528, n_1398, n_526);
  nand g1463 (n_1399, n_524, n_525);
  nand g1464 (n_1400, n_526, n_525);
  nand g1465 (n_1401, n_524, n_526);
  nand g1466 (n_540, n_1399, n_1400, n_1401);
  xor g1468 (n_529, n_1122, n_527);
  nand g1470 (n_1404, n_527, A[23]);
  nand g1471 (n_1405, A[22], n_527);
  nand g1472 (n_543, n_1123, n_1404, n_1405);
  xor g1473 (n_1406, n_528, n_529);
  xor g1474 (n_88, n_1406, n_530);
  nand g1475 (n_1407, n_528, n_529);
  nand g1476 (n_1408, n_530, n_529);
  nand g1477 (n_1409, n_528, n_530);
  nand g1478 (n_39, n_1407, n_1408, n_1409);
  xor g1480 (n_533, n_1098, A[12]);
  nand g1482 (n_1412, A[12], A[10]);
  nand g1483 (n_1413, A[11], A[12]);
  nand g1484 (n_544, n_1099, n_1412, n_1413);
  xor g1485 (n_1414, n_532, n_533);
  xor g1486 (n_535, n_1414, A[15]);
  nand g1487 (n_1415, n_532, n_533);
  nand g1488 (n_1416, A[15], n_533);
  nand g1489 (n_1417, n_532, A[15]);
  nand g1490 (n_546, n_1415, n_1416, n_1417);
  xor g1491 (n_1418, A[16], n_534);
  xor g1492 (n_537, n_1418, n_535);
  nand g1493 (n_1419, A[16], n_534);
  nand g1494 (n_1420, n_535, n_534);
  nand g1495 (n_1421, A[16], n_535);
  nand g1496 (n_547, n_1419, n_1420, n_1421);
  xor g1497 (n_1422, A[19], n_536);
  xor g1498 (n_539, n_1422, A[20]);
  nand g1499 (n_1423, A[19], n_536);
  nand g1500 (n_1424, A[20], n_536);
  nand g1502 (n_549, n_1423, n_1424, n_993);
  xor g1503 (n_1426, n_537, n_538);
  xor g1504 (n_541, n_1426, n_539);
  nand g1505 (n_1427, n_537, n_538);
  nand g1506 (n_1428, n_539, n_538);
  nand g1507 (n_1429, n_537, n_539);
  nand g1508 (n_551, n_1427, n_1428, n_1429);
  xor g1510 (n_542, n_1166, n_540);
  nand g1513 (n_1433, A[23], n_540);
  nand g1514 (n_554, n_1167, n_1432, n_1433);
  xor g1515 (n_1434, n_541, n_542);
  xor g1516 (n_87, n_1434, n_543);
  nand g1517 (n_1435, n_541, n_542);
  nand g1518 (n_1436, n_543, n_542);
  nand g1519 (n_1437, n_541, n_543);
  nand g1520 (n_38, n_1435, n_1436, n_1437);
  xor g1522 (n_545, n_1186, n_544);
  nand g1524 (n_1440, n_544, A[13]);
  nand g1525 (n_1441, A[12], n_544);
  nand g1526 (n_557, n_1187, n_1440, n_1441);
  xor g1527 (n_1442, A[16], n_545);
  xor g1528 (n_548, n_1442, A[17]);
  nand g1529 (n_1443, A[16], n_545);
  nand g1530 (n_1444, A[17], n_545);
  nand g1532 (n_559, n_1443, n_1444, n_1335);
  xor g1533 (n_1446, n_546, n_547);
  xor g1534 (n_550, n_1446, n_548);
  nand g1535 (n_1447, n_546, n_547);
  nand g1536 (n_1448, n_548, n_547);
  nand g1537 (n_1449, n_546, n_548);
  nand g1538 (n_561, n_1447, n_1448, n_1449);
  xor g1539 (n_1450, A[20], A[21]);
  xor g1540 (n_552, n_1450, n_549);
  nand g1541 (n_1451, A[20], A[21]);
  nand g1542 (n_1452, n_549, A[21]);
  nand g1543 (n_1453, A[20], n_549);
  nand g1544 (n_563, n_1451, n_1452, n_1453);
  xor g1546 (n_553, n_1454, n_551);
  nand g1549 (n_1457, n_550, n_551);
  nand g1550 (n_565, n_1455, n_1456, n_1457);
  xor g1551 (n_1458, n_552, n_553);
  xor g1552 (n_86, n_1458, n_554);
  nand g1553 (n_1459, n_552, n_553);
  nand g1554 (n_1460, n_554, n_553);
  nand g1555 (n_1461, n_552, n_554);
  nand g1556 (n_37, n_1459, n_1460, n_1461);
  nand g1563 (n_1465, A[14], n_557);
  nand g1564 (n_570, n_1463, n_1464, n_1465);
  xor g1565 (n_1466, A[17], A[18]);
  xor g1566 (n_560, n_1466, n_558);
  nand g1568 (n_1468, n_558, A[18]);
  nand g1569 (n_1469, A[17], n_558);
  nand g1570 (n_571, n_920, n_1468, n_1469);
  xor g1571 (n_1470, n_559, n_560);
  xor g1572 (n_562, n_1470, n_561);
  nand g1573 (n_1471, n_559, n_560);
  nand g1574 (n_1472, n_561, n_560);
  nand g1575 (n_1473, n_559, n_561);
  nand g1576 (n_574, n_1471, n_1472, n_1473);
  xor g1577 (n_1474, A[21], A[22]);
  xor g1578 (n_564, n_1474, n_562);
  nand g1580 (n_1476, n_562, A[22]);
  nand g1581 (n_1477, A[21], n_562);
  nand g1582 (n_575, n_1077, n_1476, n_1477);
  xor g1583 (n_1478, n_563, n_564);
  xor g1584 (n_85, n_1478, n_565);
  nand g1585 (n_1479, n_563, n_564);
  nand g1586 (n_1480, n_565, n_564);
  nand g1587 (n_1481, n_563, n_565);
  nand g1588 (n_36, n_1479, n_1480, n_1481);
  xor g1591 (n_1482, A[13], A[15]);
  nand g1596 (n_578, n_772, n_1484, n_1485);
  xor g1597 (n_1486, A[18], n_569);
  xor g1598 (n_572, n_1486, n_570);
  nand g1599 (n_1487, A[18], n_569);
  nand g1600 (n_1488, n_570, n_569);
  nand g1601 (n_1489, A[18], n_570);
  nand g1602 (n_580, n_1487, n_1488, n_1489);
  xor g1603 (n_1490, A[19], n_571);
  xor g1604 (n_573, n_1490, n_572);
  nand g1605 (n_1491, A[19], n_571);
  nand g1606 (n_1492, n_572, n_571);
  nand g1607 (n_1493, A[19], n_572);
  nand g1608 (n_582, n_1491, n_1492, n_1493);
  xor g1609 (n_1494, A[22], n_573);
  xor g1610 (n_576, n_1494, A[23]);
  nand g1611 (n_1495, A[22], n_573);
  nand g1612 (n_1496, A[23], n_573);
  nand g1614 (n_584, n_1495, n_1496, n_1123);
  xor g1615 (n_1498, n_574, n_575);
  xor g1616 (n_84, n_1498, n_576);
  nand g1617 (n_1499, n_574, n_575);
  nand g1618 (n_1500, n_576, n_575);
  nand g1619 (n_1501, n_574, n_576);
  nand g1620 (n_35, n_1499, n_1500, n_1501);
  xor g1622 (n_579, n_1106, A[16]);
  nand g1626 (n_586, n_1107, n_801, n_1153);
  xor g1627 (n_1506, n_578, n_579);
  xor g1628 (n_581, n_1506, A[19]);
  nand g1629 (n_1507, n_578, n_579);
  nand g1630 (n_1508, A[19], n_579);
  nand g1631 (n_1509, n_578, A[19]);
  nand g1632 (n_588, n_1507, n_1508, n_1509);
  xor g1633 (n_1510, A[20], n_580);
  xor g1634 (n_583, n_1510, n_581);
  nand g1635 (n_1511, A[20], n_580);
  nand g1636 (n_1512, n_581, n_580);
  nand g1637 (n_1513, A[20], n_581);
  nand g1638 (n_589, n_1511, n_1512, n_1513);
  xor g1639 (n_1514, n_582, n_583);
  xor g1640 (n_585, n_1514, A[23]);
  nand g1641 (n_1515, n_582, n_583);
  nand g1642 (n_1516, A[23], n_583);
  nand g1643 (n_1517, n_582, A[23]);
  nand g1644 (n_591, n_1515, n_1516, n_1517);
  xor g1646 (n_83, n_1518, n_585);
  nand g1648 (n_1520, n_585, n_584);
  nand g1650 (n_34, n_1519, n_1520, n_1521);
  xor g1652 (n_587, n_1334, n_586);
  nand g1654 (n_1524, n_586, A[17]);
  nand g1655 (n_1525, A[16], n_586);
  nand g1656 (n_595, n_1335, n_1524, n_1525);
  xor g1657 (n_1526, A[20], n_587);
  xor g1658 (n_590, n_1526, n_588);
  nand g1659 (n_1527, A[20], n_587);
  nand g1660 (n_1528, n_588, n_587);
  nand g1661 (n_1529, A[20], n_588);
  nand g1662 (n_597, n_1527, n_1528, n_1529);
  xor g1664 (n_592, n_1530, n_589);
  nand g1667 (n_1533, A[21], n_589);
  nand g1668 (n_599, n_1531, n_1532, n_1533);
  xor g1669 (n_1534, n_590, n_591);
  xor g1670 (n_82, n_1534, n_592);
  nand g1671 (n_1535, n_590, n_591);
  nand g1672 (n_1536, n_592, n_591);
  nand g1673 (n_1537, n_590, n_592);
  nand g1674 (n_81, n_1535, n_1536, n_1537);
  nand g1681 (n_1541, A[18], n_595);
  nand g1682 (n_604, n_1539, n_1540, n_1541);
  xor g1684 (n_598, n_1474, n_596);
  nand g1686 (n_1544, n_596, A[22]);
  nand g1687 (n_1545, A[21], n_596);
  nand g1688 (n_606, n_1077, n_1544, n_1545);
  xor g1689 (n_1546, n_597, n_598);
  xor g1690 (n_33, n_1546, n_599);
  nand g1691 (n_1547, n_597, n_598);
  nand g1692 (n_1548, n_599, n_598);
  nand g1693 (n_1549, n_597, n_599);
  nand g1694 (n_32, n_1547, n_1548, n_1549);
  xor g1697 (n_1550, A[17], A[19]);
  nand g1702 (n_608, n_889, n_1552, n_1553);
  xor g1703 (n_1554, A[22], n_603);
  xor g1704 (n_605, n_1554, n_604);
  nand g1705 (n_1555, A[22], n_603);
  nand g1706 (n_1556, n_604, n_603);
  nand g1707 (n_1557, A[22], n_604);
  nand g1708 (n_610, n_1555, n_1556, n_1557);
  xor g1709 (n_1558, A[23], n_605);
  xor g1710 (n_80, n_1558, n_606);
  nand g1711 (n_1559, A[23], n_605);
  nand g1712 (n_1560, n_606, n_605);
  nand g1713 (n_1561, A[23], n_606);
  nand g1714 (n_31, n_1559, n_1560, n_1561);
  xor g1715 (n_1562, A[19], A[18]);
  xor g1716 (n_609, n_1562, A[20]);
  nand g1718 (n_1564, A[20], A[18]);
  nand g1720 (n_612, n_1397, n_1564, n_993);
  xor g1721 (n_1566, n_608, n_609);
  xor g1722 (n_611, n_1566, A[23]);
  nand g1723 (n_1567, n_608, n_609);
  nand g1724 (n_1568, A[23], n_609);
  nand g1725 (n_1569, n_608, A[23]);
  nand g1726 (n_614, n_1567, n_1568, n_1569);
  xor g1728 (n_79, n_1570, n_611);
  nand g1730 (n_1572, n_611, n_610);
  nand g1732 (n_30, n_1571, n_1572, n_1573);
  xor g1734 (n_613, n_1450, n_612);
  nand g1736 (n_1576, n_612, A[21]);
  nand g1737 (n_1577, A[20], n_612);
  nand g1738 (n_617, n_1451, n_1576, n_1577);
  xor g1740 (n_78, n_1578, n_614);
  nand g1742 (n_1580, n_614, n_613);
  nand g1744 (n_77, n_1579, n_1580, n_1581);
  nand g1751 (n_1585, A[22], n_617);
  nand g1752 (n_28, n_1583, n_1584, n_1585);
  nand g1759 (n_1589, A[21], A[23]);
  nand g1760 (n_27, n_1587, n_1588, n_1589);
  xor g1762 (n_75, n_1166, A[22]);
  nand g1766 (n_74, n_1167, n_1123, n_1593);
  nand g16 (n_1606, A[0], A[2]);
  xor g20 (Z[2], A[0], A[2]);
  nand g22 (n_1611, n_68, A[3]);
  nand g25 (n_1615, n_1611, n_1612, n_1613);
  xor g26 (n_1614, n_68, A[3]);
  nand g28 (n_1616, A[4], n_117);
  nand g29 (n_1617, A[4], n_1615);
  nand g30 (n_1618, n_117, n_1615);
  nand g31 (n_1620, n_1616, n_1617, n_1618);
  xor g32 (n_1619, A[4], n_117);
  xor g33 (Z[4], n_1615, n_1619);
  nand g34 (n_1621, A[5], n_116);
  nand g35 (n_1622, A[5], n_1620);
  nand g36 (n_1623, n_116, n_1620);
  nand g37 (n_1625, n_1621, n_1622, n_1623);
  xor g38 (n_1624, A[5], n_116);
  xor g39 (Z[5], n_1620, n_1624);
  nand g40 (n_1626, n_67, n_115);
  nand g41 (n_1627, n_67, n_1625);
  nand g42 (n_1628, n_115, n_1625);
  nand g43 (n_1630, n_1626, n_1627, n_1628);
  xor g44 (n_1629, n_67, n_115);
  xor g45 (Z[6], n_1625, n_1629);
  nand g46 (n_1631, n_66, n_114);
  nand g47 (n_1632, n_66, n_1630);
  nand g48 (n_1633, n_114, n_1630);
  nand g49 (n_1635, n_1631, n_1632, n_1633);
  xor g50 (n_1634, n_66, n_114);
  xor g51 (Z[7], n_1630, n_1634);
  nand g52 (n_1636, n_65, n_113);
  nand g53 (n_1637, n_65, n_1635);
  nand g54 (n_1638, n_113, n_1635);
  nand g55 (n_1640, n_1636, n_1637, n_1638);
  xor g56 (n_1639, n_65, n_113);
  xor g57 (Z[8], n_1635, n_1639);
  nand g58 (n_1641, n_64, n_112);
  nand g59 (n_1642, n_64, n_1640);
  nand g60 (n_1643, n_112, n_1640);
  nand g61 (n_1645, n_1641, n_1642, n_1643);
  xor g62 (n_1644, n_64, n_112);
  xor g63 (Z[9], n_1640, n_1644);
  nand g64 (n_1646, n_63, n_111);
  nand g65 (n_1647, n_63, n_1645);
  nand g66 (n_1648, n_111, n_1645);
  nand g67 (n_1650, n_1646, n_1647, n_1648);
  xor g68 (n_1649, n_63, n_111);
  xor g69 (Z[10], n_1645, n_1649);
  nand g70 (n_1651, n_62, n_110);
  nand g71 (n_1652, n_62, n_1650);
  nand g72 (n_1653, n_110, n_1650);
  nand g73 (n_1655, n_1651, n_1652, n_1653);
  xor g74 (n_1654, n_62, n_110);
  xor g75 (Z[11], n_1650, n_1654);
  nand g76 (n_1656, n_61, n_109);
  nand g77 (n_1657, n_61, n_1655);
  nand g78 (n_1658, n_109, n_1655);
  nand g79 (n_1660, n_1656, n_1657, n_1658);
  xor g80 (n_1659, n_61, n_109);
  xor g81 (Z[12], n_1655, n_1659);
  nand g82 (n_1661, n_60, n_108);
  nand g83 (n_1662, n_60, n_1660);
  nand g84 (n_1663, n_108, n_1660);
  nand g85 (n_1665, n_1661, n_1662, n_1663);
  xor g86 (n_1664, n_60, n_108);
  xor g87 (Z[13], n_1660, n_1664);
  nand g88 (n_1666, n_59, n_107);
  nand g89 (n_1667, n_59, n_1665);
  nand g90 (n_1668, n_107, n_1665);
  nand g91 (n_1670, n_1666, n_1667, n_1668);
  xor g92 (n_1669, n_59, n_107);
  xor g93 (Z[14], n_1665, n_1669);
  nand g94 (n_1671, n_58, n_106);
  nand g95 (n_1672, n_58, n_1670);
  nand g96 (n_1673, n_106, n_1670);
  nand g97 (n_1675, n_1671, n_1672, n_1673);
  xor g98 (n_1674, n_58, n_106);
  xor g99 (Z[15], n_1670, n_1674);
  nand g100 (n_1676, n_57, n_105);
  nand g101 (n_1677, n_57, n_1675);
  nand g102 (n_1678, n_105, n_1675);
  nand g103 (n_1680, n_1676, n_1677, n_1678);
  xor g104 (n_1679, n_57, n_105);
  xor g105 (Z[16], n_1675, n_1679);
  nand g106 (n_1681, n_56, n_104);
  nand g107 (n_1682, n_56, n_1680);
  nand g108 (n_1683, n_104, n_1680);
  nand g109 (n_1685, n_1681, n_1682, n_1683);
  xor g110 (n_1684, n_56, n_104);
  xor g111 (Z[17], n_1680, n_1684);
  nand g112 (n_1686, n_55, n_103);
  nand g113 (n_1687, n_55, n_1685);
  nand g114 (n_1688, n_103, n_1685);
  nand g115 (n_1690, n_1686, n_1687, n_1688);
  xor g116 (n_1689, n_55, n_103);
  xor g117 (Z[18], n_1685, n_1689);
  nand g118 (n_1691, n_54, n_102);
  nand g119 (n_1692, n_54, n_1690);
  nand g120 (n_1693, n_102, n_1690);
  nand g121 (n_1695, n_1691, n_1692, n_1693);
  xor g122 (n_1694, n_54, n_102);
  xor g123 (Z[19], n_1690, n_1694);
  nand g124 (n_1696, n_53, n_101);
  nand g125 (n_1697, n_53, n_1695);
  nand g126 (n_1698, n_101, n_1695);
  nand g127 (n_1700, n_1696, n_1697, n_1698);
  xor g128 (n_1699, n_53, n_101);
  xor g129 (Z[20], n_1695, n_1699);
  nand g130 (n_1701, n_52, n_100);
  nand g131 (n_1702, n_52, n_1700);
  nand g132 (n_1703, n_100, n_1700);
  nand g133 (n_1705, n_1701, n_1702, n_1703);
  xor g134 (n_1704, n_52, n_100);
  xor g135 (Z[21], n_1700, n_1704);
  nand g136 (n_1706, n_51, n_99);
  nand g137 (n_1707, n_51, n_1705);
  nand g138 (n_1708, n_99, n_1705);
  nand g139 (n_1710, n_1706, n_1707, n_1708);
  xor g140 (n_1709, n_51, n_99);
  xor g141 (Z[22], n_1705, n_1709);
  nand g142 (n_1711, n_50, n_98);
  nand g143 (n_1712, n_50, n_1710);
  nand g144 (n_1713, n_98, n_1710);
  nand g145 (n_1715, n_1711, n_1712, n_1713);
  xor g146 (n_1714, n_50, n_98);
  xor g147 (Z[23], n_1710, n_1714);
  nand g148 (n_1716, n_49, n_97);
  nand g149 (n_1717, n_49, n_1715);
  nand g150 (n_1718, n_97, n_1715);
  nand g151 (n_1720, n_1716, n_1717, n_1718);
  xor g152 (n_1719, n_49, n_97);
  xor g153 (Z[24], n_1715, n_1719);
  nand g154 (n_1721, n_48, n_96);
  nand g155 (n_1722, n_48, n_1720);
  nand g156 (n_1723, n_96, n_1720);
  nand g157 (n_1725, n_1721, n_1722, n_1723);
  xor g158 (n_1724, n_48, n_96);
  xor g159 (Z[25], n_1720, n_1724);
  nand g160 (n_1726, n_47, n_95);
  nand g161 (n_1727, n_47, n_1725);
  nand g162 (n_1728, n_95, n_1725);
  nand g163 (n_1730, n_1726, n_1727, n_1728);
  xor g164 (n_1729, n_47, n_95);
  xor g165 (Z[26], n_1725, n_1729);
  nand g166 (n_1731, n_46, n_94);
  nand g167 (n_1732, n_46, n_1730);
  nand g168 (n_1733, n_94, n_1730);
  nand g169 (n_1735, n_1731, n_1732, n_1733);
  xor g170 (n_1734, n_46, n_94);
  xor g171 (Z[27], n_1730, n_1734);
  nand g172 (n_1736, n_45, n_93);
  nand g173 (n_1737, n_45, n_1735);
  nand g174 (n_1738, n_93, n_1735);
  nand g175 (n_1740, n_1736, n_1737, n_1738);
  xor g176 (n_1739, n_45, n_93);
  xor g177 (Z[28], n_1735, n_1739);
  nand g178 (n_1741, n_44, n_92);
  nand g179 (n_1742, n_44, n_1740);
  nand g180 (n_1743, n_92, n_1740);
  nand g181 (n_1745, n_1741, n_1742, n_1743);
  xor g182 (n_1744, n_44, n_92);
  xor g183 (Z[29], n_1740, n_1744);
  nand g184 (n_1746, n_43, n_91);
  nand g185 (n_1747, n_43, n_1745);
  nand g186 (n_1748, n_91, n_1745);
  nand g187 (n_1750, n_1746, n_1747, n_1748);
  xor g188 (n_1749, n_43, n_91);
  xor g189 (Z[30], n_1745, n_1749);
  nand g190 (n_1751, n_42, n_90);
  nand g191 (n_1752, n_42, n_1750);
  nand g192 (n_1753, n_90, n_1750);
  nand g193 (n_1755, n_1751, n_1752, n_1753);
  xor g194 (n_1754, n_42, n_90);
  xor g195 (Z[31], n_1750, n_1754);
  nand g196 (n_1756, n_41, n_89);
  nand g197 (n_1757, n_41, n_1755);
  nand g198 (n_1758, n_89, n_1755);
  nand g199 (n_1760, n_1756, n_1757, n_1758);
  xor g200 (n_1759, n_41, n_89);
  xor g201 (Z[32], n_1755, n_1759);
  nand g202 (n_1761, n_40, n_88);
  nand g203 (n_1762, n_40, n_1760);
  nand g204 (n_1763, n_88, n_1760);
  nand g205 (n_1765, n_1761, n_1762, n_1763);
  xor g206 (n_1764, n_40, n_88);
  xor g207 (Z[33], n_1760, n_1764);
  nand g208 (n_1766, n_39, n_87);
  nand g209 (n_1767, n_39, n_1765);
  nand g210 (n_1768, n_87, n_1765);
  nand g211 (n_1770, n_1766, n_1767, n_1768);
  xor g212 (n_1769, n_39, n_87);
  xor g213 (Z[34], n_1765, n_1769);
  nand g214 (n_1771, n_38, n_86);
  nand g215 (n_1772, n_38, n_1770);
  nand g216 (n_1773, n_86, n_1770);
  nand g217 (n_1775, n_1771, n_1772, n_1773);
  xor g218 (n_1774, n_38, n_86);
  xor g219 (Z[35], n_1770, n_1774);
  nand g220 (n_1776, n_37, n_85);
  nand g221 (n_1777, n_37, n_1775);
  nand g222 (n_1778, n_85, n_1775);
  nand g223 (n_1780, n_1776, n_1777, n_1778);
  xor g224 (n_1779, n_37, n_85);
  xor g225 (Z[36], n_1775, n_1779);
  nand g226 (n_1781, n_36, n_84);
  nand g227 (n_1782, n_36, n_1780);
  nand g228 (n_1783, n_84, n_1780);
  nand g229 (n_1785, n_1781, n_1782, n_1783);
  xor g230 (n_1784, n_36, n_84);
  xor g231 (Z[37], n_1780, n_1784);
  nand g232 (n_1786, n_35, n_83);
  nand g233 (n_1787, n_35, n_1785);
  nand g234 (n_1788, n_83, n_1785);
  nand g235 (n_1790, n_1786, n_1787, n_1788);
  xor g236 (n_1789, n_35, n_83);
  xor g237 (Z[38], n_1785, n_1789);
  nand g238 (n_1791, n_34, n_82);
  nand g239 (n_1792, n_34, n_1790);
  nand g240 (n_1793, n_82, n_1790);
  nand g241 (n_1795, n_1791, n_1792, n_1793);
  xor g242 (n_1794, n_34, n_82);
  xor g243 (Z[39], n_1790, n_1794);
  nand g244 (n_1796, n_33, n_81);
  nand g245 (n_1797, n_33, n_1795);
  nand g246 (n_1798, n_81, n_1795);
  nand g247 (n_1800, n_1796, n_1797, n_1798);
  xor g248 (n_1799, n_33, n_81);
  xor g249 (Z[40], n_1795, n_1799);
  nand g250 (n_1801, n_32, n_80);
  nand g251 (n_1802, n_32, n_1800);
  nand g252 (n_1803, n_80, n_1800);
  nand g253 (n_1805, n_1801, n_1802, n_1803);
  xor g254 (n_1804, n_32, n_80);
  xor g255 (Z[41], n_1800, n_1804);
  nand g256 (n_1806, n_31, n_79);
  nand g257 (n_1807, n_31, n_1805);
  nand g258 (n_1808, n_79, n_1805);
  nand g259 (n_1810, n_1806, n_1807, n_1808);
  xor g260 (n_1809, n_31, n_79);
  xor g261 (Z[42], n_1805, n_1809);
  nand g262 (n_1811, n_30, n_78);
  nand g263 (n_1812, n_30, n_1810);
  nand g264 (n_1813, n_78, n_1810);
  nand g265 (n_1815, n_1811, n_1812, n_1813);
  xor g266 (n_1814, n_30, n_78);
  xor g267 (Z[43], n_1810, n_1814);
  nand g1772 (n_1816, n_29, n_77);
  nand g1773 (n_1817, n_29, n_1815);
  nand g1774 (n_1818, n_77, n_1815);
  nand g1775 (n_1820, n_1816, n_1817, n_1818);
  xor g1776 (n_1819, n_29, n_77);
  xor g1777 (Z[44], n_1815, n_1819);
  nand g1778 (n_1821, n_28, n_76);
  nand g1779 (n_1822, n_28, n_1820);
  nand g1780 (n_1823, n_76, n_1820);
  nand g1781 (n_1825, n_1821, n_1822, n_1823);
  xor g1782 (n_1824, n_28, n_76);
  xor g1783 (Z[45], n_1820, n_1824);
  nand g1784 (n_1826, n_27, n_75);
  nand g1785 (n_1827, n_27, n_1825);
  nand g1786 (n_1828, n_75, n_1825);
  nand g1787 (n_1830, n_1826, n_1827, n_1828);
  xor g1788 (n_1829, n_27, n_75);
  xor g1789 (Z[46], n_1825, n_1829);
  xor g1791 (Z[47], n_1830, n_1831);
  or g1804 (n_1043, A[1], wc);
  not gc (wc, n_171);
  or g1805 (n_1044, A[1], wc0);
  not gc0 (wc0, A[2]);
  xnor g1807 (n_1166, A[24], A[23]);
  or g1808 (n_1167, wc1, A[24]);
  not gc1 (wc1, A[23]);
  xnor g1809 (n_1214, A[6], A[5]);
  or g1810 (n_1215, A[5], wc2);
  not gc2 (wc2, A[6]);
  or g1811 (n_1252, wc3, A[6]);
  not gc3 (wc3, A[5]);
  or g1812 (n_1253, A[6], wc4);
  not gc4 (wc4, A[7]);
  or g1814 (n_1355, A[9], wc5);
  not gc5 (wc5, A[10]);
  or g1815 (n_1384, A[10], wc6);
  not gc6 (wc6, A[11]);
  or g1816 (n_1385, wc7, A[10]);
  not gc7 (wc7, A[9]);
  or g1818 (n_1463, A[13], wc8);
  not gc8 (wc8, A[14]);
  or g1819 (n_1484, A[14], wc9);
  not gc9 (wc9, A[15]);
  or g1820 (n_1485, wc10, A[14]);
  not gc10 (wc10, A[13]);
  xnor g1821 (n_1530, A[24], A[21]);
  or g1822 (n_1531, wc11, A[24]);
  not gc11 (wc11, A[21]);
  or g1824 (n_1539, A[17], wc12);
  not gc12 (wc12, A[18]);
  or g1825 (n_1552, A[18], wc13);
  not gc13 (wc13, A[19]);
  or g1826 (n_1553, wc14, A[18]);
  not gc14 (wc14, A[17]);
  or g1828 (n_1583, A[21], wc15);
  not gc15 (wc15, A[22]);
  or g1829 (n_1587, wc16, A[22]);
  not gc16 (wc16, A[21]);
  or g1830 (n_1588, A[22], wc17);
  not gc17 (wc17, A[23]);
  or g1831 (n_1593, wc18, A[24]);
  not gc18 (wc18, A[22]);
  xnor g1833 (n_372, n_626, A[1]);
  or g1834 (n_1088, A[1], wc19);
  not gc19 (wc19, A[3]);
  xnor g1835 (n_453, n_1250, A[6]);
  xnor g1836 (n_519, n_1382, A[10]);
  xnor g1837 (n_569, n_1482, A[14]);
  xnor g1838 (n_603, n_1550, A[18]);
  xnor g1839 (n_76, n_1474, A[23]);
  or g1841 (n_1047, wc20, n_117);
  not gc20 (wc20, A[5]);
  or g1842 (n_1049, wc21, n_117);
  not gc21 (wc21, n_179);
  xnor g1844 (n_1578, n_613, A[24]);
  or g1845 (n_1579, A[24], wc22);
  not gc22 (wc22, n_613);
  xnor g1846 (n_1831, n_74, A[24]);
  or g1848 (n_1051, wc23, n_180);
  not gc23 (wc23, A[6]);
  or g1849 (n_1052, wc24, n_180);
  not gc24 (wc24, A[9]);
  xnor g1850 (n_504, n_1218, n_503);
  or g1851 (n_1356, A[9], wc25);
  not gc25 (wc25, n_503);
  xnor g1852 (n_558, n_1358, n_557);
  or g1853 (n_1464, A[13], wc26);
  not gc26 (wc26, n_557);
  xnor g1854 (n_596, n_1466, n_595);
  or g1855 (n_1540, A[17], wc27);
  not gc27 (wc27, n_595);
  or g1856 (n_1573, A[24], wc28);
  not gc28 (wc28, n_611);
  or g1857 (n_1581, A[24], wc29);
  not gc29 (wc29, n_614);
  xnor g1858 (n_29, n_1474, n_617);
  or g1859 (n_1584, A[21], wc30);
  not gc30 (wc30, n_617);
  or g1862 (n_1216, A[5], wc31);
  not gc31 (wc31, n_433);
  or g1863 (n_1612, n_1606, wc32);
  not gc32 (wc32, n_68);
  or g1864 (n_1613, wc33, n_1606);
  not gc33 (wc33, A[3]);
  xnor g1865 (Z[3], n_1606, n_1614);
  xnor g1866 (n_355, n_202, n_906);
  or g1867 (n_1056, wc34, n_202);
  not gc34 (wc34, n_282);
  or g1868 (n_1057, wc35, n_202);
  not gc35 (wc35, A[10]);
  xnor g1869 (n_1570, n_610, A[24]);
  or g1870 (n_1571, A[24], wc36);
  not gc36 (wc36, n_610);
  or g1871 (n_1532, A[24], wc37);
  not gc37 (wc37, n_589);
  xnor g1872 (n_1518, n_584, A[24]);
  or g1873 (n_1519, A[24], wc38);
  not gc38 (wc38, n_584);
  xnor g1874 (n_1454, n_550, A[24]);
  or g1875 (n_1455, A[24], wc39);
  not gc39 (wc39, n_550);
  or g1876 (n_1521, A[24], wc40);
  not gc40 (wc40, n_585);
  or g1877 (n_1456, A[24], wc41);
  not gc41 (wc41, n_551);
  xnor g1878 (n_1206, n_426, A[24]);
  or g1879 (n_1207, A[24], wc42);
  not gc42 (wc42, n_426);
  or g1880 (n_1081, A[24], wc43);
  not gc43 (wc43, n_363);
  xnor g1881 (n_1346, n_496, A[24]);
  or g1882 (n_1347, A[24], wc44);
  not gc44 (wc44, n_496);
  or g1883 (n_1080, A[24], wc45);
  not gc45 (wc45, n_364);
  or g1884 (n_1316, A[24], wc46);
  not gc46 (wc46, n_482);
  or g1885 (n_1348, A[24], wc47);
  not gc47 (wc47, n_497);
  xnor g1886 (n_367, n_1078, A[24]);
  or g1887 (n_1169, A[24], wc48);
  not gc48 (wc48, n_408);
  or g1888 (n_1208, A[24], wc49);
  not gc49 (wc49, n_427);
  or g1889 (n_1432, A[24], wc50);
  not gc50 (wc50, n_540);
endmodule

module mult_signed_const_6021_GENERIC(A, Z);
  input [24:0] A;
  output [47:0] Z;
  wire [24:0] A;
  wire [47:0] Z;
  mult_signed_const_6021_GENERIC_REAL g1(.A (A), .Z (Z));
endmodule

